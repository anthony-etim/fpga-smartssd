`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
JOAFmN7MhR6w3yBSOfBKDeSsI5hm6ums6qxgGZ8dnYQ2KD9dpZfQcC2zI83GILRR5vF3Yyq1yTiZ
k8r5qKL0uA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
jfvg1X38SbMYNN3yqF1i56s2Du98wF9u+BpGnrlsJynaGFN+D7yBh09EZ4+vHQc22UKR7xPzubjt
tj8t0s0PTnYjaZGAUphNfxY5QAmJdeTodeJdjyG4yZXqDlBEWeObrITMlZHFvGuNhHV57mKM+oHB
UwuR26DLm74t7mYp+fA=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
qJKCED1BAc7BGYsTgK6P2gdbdfAkiAslu5vohHfYNzojGSIQGhjlwE/wVhz9WCndRinkmwH/yd5Y
HrPt4uwaIzSFHzQaUBW4ek51ZUJ9wXL600fEqP6Q7Etv27Kd+SW/8RaW+vssyWrmZYBeI1je1mmD
+JZAZ9xU6psu6F+V/SeWeC5tdoHAKBEe5m7ZMfxIRCq1wwD4Grp/NXldfGuwtv0tiD83nDrhRQnB
drW8D73Sno1zKHnhDnCQbZy6Wf5c9y6IneWmdGSYgDW0aazGTdYxLXBlA3VJGzT6kIvQL9bHuHa3
MLoi90a+FkZ4iF2HpnXRLghgvDITXtpMlrKEMg==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
rpUdZetpZGd19xednZhbjWa7Fe94yM5ATNaRDWPdBPH+YjfXelIOcjImIfDRWKdcp03BKtRNBjuo
sdecWhcDV8T7FqXhwhJWXzbkx+PSGGtS1PkVCZb1H0kvuuWUI5gClnMy1c9pPBVNEPTwRGl5xNQw
c6ghD/zlWY2ko6nb1DIsXwTB0QKig1Z6PB8M2JsLKwPhHvIA9VR5QcdJRU5MLdZqySwyhT6RRreF
QmorwwRgEfQOEEPZhRArkgp8SaGKHihpFlfZWNAEWuFlY2eK3SIGwI1fmNqMDGiocFyzVNlOmGsz
hnGeGLIHw0mWQjUB8DdCXyle8L6HjhL+1ya2mA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
WdFhWA8JPPIE3+vs5HNDO41Z7vDL0NLOxrwrbAIIWrsx8CAxfd6jJ4SrnOy/jA0ejbfhPSE6jhUo
qUn4G4Qgk2QMqPdOst9YPp45DQxeivdqK3ijLZih0OysQXcaXz05S2T2ywIw3ioLdpX+1mazlOnM
yOw7k+qbqAwgSLfNrj+Qh0POY2U8nJUX7qUQLHoeSe+crdjrxB3hkAZlJtcaPkc3mIMeQCIMHL9u
lQIhJlapNVct5bEdY+cUdxiOaFXGdY5kO3xH2KvLf16Wv+ERdf9HT1Lw9P4b4wbe6KtEbENEF6B+
2Non0bg02+XOiM4SbNSGAQDDCpUVHOicXs+TPQ==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
FcoOn31iKFNo5Blj0fbygoxDk2yIVUalIHnWjkQIJdCsC/wxJYTB0y1N0OdYfPv/FmQOpvJdIRMo
laqcbfB4joJWq4Tblp2GIT0MJy+KTUOku+lh6I921yHvrSP1ZuCzaYaRiVCWP9g7aKTAdT2EtSBa
KOa6YTx2Y08yDyOrXOs=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
mrJi2aNDh25xn/wLvAIO7Xn+RYfyQHLKtygjGCGYnuUYjNqwXoRJYOtJMRH9rIqR6kI+4IBsSCY7
raqLA4o5bAPMcvABO1If1Zxl1yIuVTrmIsNWKOFMbFFAw+XjS3j/8Aa6JrZp+J4QKfxeFuroUh52
nYZhmHxXzpQaBzqcKIWPjj/1k/RvsGEahMZbv/eyxd0DD0aihTFCXo1ToOFm3B2Lvt723n3IgmZi
rQRAP00JdTUdlYaDhuukqWgVKOdAZxhkL9HVWyQtq52r/Fwt+ZvQ6BYpknrcIqVRlo8v1GBpqQ6l
6ESIwWaF3jxRSHcx1qjCWt3oUGQVt4jVaT8xJA==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
0qNDA3WYKpLQi5qdid5aF9mZYXXU2AsTwZEDHibFK8R8ffUsdBZlLYdgIlx5DLUQG0OWmmxDi7GQ
jWOM0I311IFsTVjc1OmUHTTmtl4esgt+nOJtuLRK1Dmf7rndcQNFWHD1NcGFoiFe+jBB2LHH9NbY
lzxY1XdSXhVSF91DOa6GCbgX389gghvRCLL3zwoc573XpgRtodzwDsZPXlR5zJoPcgjZsz6srrax
wYChKVhvpHpmcbG++j457QcN5rggxRL4ArMyLHoE3ddTucB5EoQB+tQKJLZkxZ88CYVklAkRYYUU
dpyovSEzJbkdzmMFjdD5LC2++P/6XOKpddvLcw==

`pragma protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
lV2NyLkwq5JeziokX596vuUemekm72ZxBOIvSxbzoPY6BwLazKj2YXOuQqM+tFuI8C9ymBtG1pcT
c0bRNGkiJpIUrodPo4iB52+nW0uQ5SMph+h0UgERMmPpGtu1kKSh+nOTpIl3+aeGK5plW/G7iS7O
rogx62/4AngbIA7A4+wiDkWzquxhgzJ9Ty4WxLFzPfoqLCIzw+X2+6TmAQN0auU/szFZyAXQ1O7Z
3Ess0bL20n3cQKqX8vwPIL0AFCZlIDgRA3b5Xe+ZpBZT9HDMCNZdDlW5YhmMa1QipRomfAiEXSUt
sO1eqOabJ0NrRPbysuPsXf6P4j0nTHr0LIZ//g==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_11", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
CWg3E8yxKvbp1snsyLPAb5eOklquGqYQyi+yYlmkyLFHONLsQaSBafeT5XhzZS87C7uAnybQRIJp
Ik6AlzdsbqIeIxgXFRjq0keNc6GrtGr08UbrOTHbXR5VASSQcUh907Y5kqsD10Q/RbYSD+rPCfNg
YM8+zT8zHciB82Q4ArdxGOR7CXHohCpIEPqE+BW7ZNWz4ZqBR0nSuZ3pRP5QOKseGUaU/anfGLbv
cdf1+yG/avc31Y+9MAdsDpluxd0Hu3VkjGuYhY0AvL/GoDxR6bVd30CjbiUpf/+XGsz4rWh+5VQj
rV1nIXmHVdyCxbMOem9/i97kRWcGCtsTLtWYCw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2331584)
`pragma protect data_block
Du50BQgXza6URIW61t/+++Izc85FrC22yR3GcKJ8Z3Mxi0iQN6BQWkzDLgt+oOctB3TdAmcTcXo4
gSP4LU1Yl+Z7sofUCYrcnMt54brygi8b6zmM3hvZ4eHktmh37SDjgpKItVH22pgj89fO3J+ETrPy
82wGnkwYdX4FKZaKeYDk83Z+DzCU1N/KfhC2GIO4uKbQHxGAliwqry95FBfNsovO/rNJMu/+MxjL
bTEMc7gnGhXJ7PjjaaQ+KNSh3yPeuZGaK6WRi84xkOhKSTWDsy+h6EWCRMdSWBjaJ8vQh6z6lOds
XfmGx0jYFG6irpyiwg18dRzjuAylZZDUwN8cGzZWwbvbEKuxEFZDOJTv9dsAkIeAs69dLlBy1ULU
NoBu/r4sgrGTmC4UNvcb1yrHHqpKj1N34jRUXg8XVvzTFb8qla9wkztqhv6OtLkm3LyUkzyJPjpf
0ahBqFWECas+3pT+09pWJbx5ap/pLZwDnL31INwPVPwJ2qNC+0FocBYhtukY4+4l1h9UyUCah9dD
NSwvwBlKUNmOk4Ib6oS9M2TQs9GVdpmMRY2Z5DjT5HqOTQP/1fSubSjdq0eORc6RrxOuCQkd5Xjr
LPwVHiVCDdXtctpnViI2XAyu7nsGHQCWeQKbeST+pvCauHx0CgAqSw028/OsYIsfKUpmY19ZXWHv
/FQ/NF41+gNXCYjzUAroaLy4PX8cp7NNkVR4XKID9TkIgg92gWJYck82os1ArjtdRsJY1/otsSKV
15rMjK4nCsrCV4SCzw5HkXp0RIZ0wtMN5kLXE3tDjz96o/frvlrH5meo8DlL9n9PjKORMQU+IF3Z
3K1eqbAUh2LuZF01HvSBsKWlcOTS1D5Ux6AyfTzlFHIDolZjuxg6e/POhfIKjfaGxr3yjMee1HrR
vjR3yHEa446xpAdOAuwrOQnbRazAoTGSo2zzES1XoI2JpzoqnURiVMQNYbDpL7U/We+DZ76lpG7v
z0YxZ+HqZrA5wKFJbtyt7whqIPdm/MR8pVpA+Zd0U3UeEn3X9QanTxg1GWdygKaxTrWoLz/8sumt
2XZM15l/1ssms/U8QPTpUUlryEb9TDQ9p/c5FnSyYpd27rOjURz+iqabxq00zwSRDc+QFyQUrVK2
SYm7E3FVKoDkSWnAeGFxMUJIAgBw/M8sagyUbz+JFi2fQm4I9/l2M+5DOpRiSPJO1QWbK7MSq5Fh
ThD/bt4C692LBryjOewosn9oyw4Rsc65/LXz3xDVVfsh2dED8nSIP6pdMr5WedIyhLZOIAKmFXOM
JBWlxy2qKXWz0nm+iYYpk+z61Kaoqniq5qB8+Y3kbWnYWIqBxGC5GvDrc6Pcln33QpezJcXm2LA8
O6+mNFa49wOcNxkAFvQu/XEOSshkTgic5oH8yiRvgxYX1gV5x7oqmNYjMib+FoxiBeQyI6E3mqm3
3MNV2baeElpcJRToZXHXR0zQjnKk7YEka+XXq/oCYdEEOjitAFD0skfqCxRcFy/Kejb4H4Gp6q8h
aC5WKDKAO8PDkYdIld0TJdvgMf6yuuQYTbqiwwWR+fSdbXKvGQ4LRr7vk6TGWG13aIZDwl7sVxTM
U4Q62lsEMeFg5B0ZnXRCsNYtvRrPw91xquPwsj3A/lc9mmyGR+iy9X1jmA/4m0Kwmi9OKYGclRYX
PfUTpY25G5qqa+rfXJjwnCqI/6byw+IzoucYab9b0MPqZ224BFDJy2obmwUhu0+4ZLKPQDhAmE6g
L2Th1C7ihxlhTMxaih0cqEhqxz+f0hV6LuoVlWjfVj/ZegCD9EJIe0089doUcxVkxR2TixSzTI4E
5bDPzQ6TrbDdGUnu7SEOREHT2fI+AO9bCo8pytTozZcp8zpvCpETVhsE2hvj/YAQJXgDhgpjbzpW
4Nf78URlDB13QDwHmAI4bJxMc+ep/N3fC7Djnhv7Oucnpbk1O5KGR205Xk8F0euAQSJIPTUHNZi/
Py3tBE0vP6c3pTFI3oBJDYI4hOztgoMsQAsh4JWSTw0uE6QdO46a5mIapfpOj0tV+2YORN3kFlJD
r5KKGHBVy4C42a7Xa06TqypAI/imZMMAgFxaMXnPppQTgSzbZ2ws11lXvP/DpZPIqHFgfaCUL2LY
ZVo9XDFk6Ts9YP2MOQZacGtyCtRyuEY6P01+jm2cH4gfYWnObuUBcdyYn5cozOnKnuqMT4bdRcim
MhbeWWeiLQow6ng2iGpsrYQXURLtbw0eQwd1N3WwMxCFXFW7HEQWOg8NGumACk705xFzSLVZIVyJ
S6DRY4Fssi8orKd8gYAmafswgN/DughQdkVwFxcW67ioTjNug/4MUmcAPB/iKGOk4rPori+FB8a6
kh5QaiwzzL2ktzN/ZqoErZPPCzc3MJlN+dPR95jwTkD4zmnPkhLbmDKMjfEZQlauurIn5TsxevDe
yxr/SQnEU7Un6uTHwBiXbvNnZjXc2kl7H9H3B6K/YGgWdGo68jsUIxEavm3/HUrFD7J2JzsqaTNG
rR3NmngOUAoddwgYrxbOHKbYrtFvfPVST862TqKCc8L4rW96rcBSAo7vi+cgkhW95Mk5dSgDQk8+
WTGDoylgnU5SWDv42XXuo19+rMTf59KBJNpSEx0UQI6EjLmtsu9IrVeEj2gBiGTSg8XyuZk4i02c
vRmSh0+xGtK4EshozbMhNAIOqZaGvq2H0iK4fcus5B3q5BUqnZFi1R7YZOjor7T/PXVJwYbPu6EV
lLLYr0ChCeqJU4jmREDZQmJtq4ZMINFn4d3Ys3y8rmJEyQKD6qhB54IRQRmGntrMJrsrHXLmWL1u
3kll1MJyTGo4cMf6AJboS/RRev5rRYyr5HoTwblbq2I45QkpzXuRA/0WLPF07bjjPqq39EQF5gV7
0G9Glt7E1+9eAN8Dqq0SdqMs/FXR5Ws7USyJf+6wXgK1ayXBT7c25/9uNzQmQ2tqhJl+dB85/T2A
LS167/UCx5aB7HzBdJMbCpvbwQRxS2cMtSuWUGV8bjzbJ5UpR+7/oaYW0gq/fa/QLzs4MLe/idlA
N1SlaIjaffEEw6bMdmhVjOa7ZGPrFQ9H4zKh9OtCwCsd0+fW+apL20OTYRNWlcjbHmgXuv06qsp4
DLZxvQiM2y/iFlVjzMUT/aOMTHeeHrnL34g11IbwY1+p93f03VYISFicmfcm9Itr0Ut81QTz/jN0
yoslSPmRpwJS4irdMUbeMmQegauzHlDENXl/7cuJd+y9zuLozOq4WQZiY2h2TkyN6WCabX5JGXZn
f1aMlhHuHxAUsSu8gTbfIMfERPUygUW1aKo/mFkFt77uUTuoV9TnKbEizUrU4zhnDswKYMDvARTs
8M+kTHtInwRDT5NjAI2VBG1P4aVwPLev9l/hv8GsO4Jbr+FvbetoTEZ800VN6DgB+jWewBDU3/hY
MeUlZck2XeR1gezU9+PD8VVQsg2V3najzbyejG+DN9Njm20ghH85q4Amu5Q3vwsMvNdPq/j6vw5g
o84TNT/mSyt4+coHMbYcy00PyC03K1QqM77zB5HuhE/dk0e0UfiY1lHQwu9nTgl5HLi6uZ0isJcV
JHgjTE1AehL0c1nDdTCIN3bF7rd7knwv0wgRy9RgA1MGxt44geRECPoaTXOUDqpSDwjj3vNffJGD
Z9V+NVNpiAWELkVACzJv9BNBEgiLMz6MhWKESG1/7GF7CY79g5Rlscbx9yKTKbmhjsmmOpXlIwvy
RE3bXN6PnRDz9Lws9KzoC1Ds+0POUF8hEbLV1x54cjX5VOSzgiKDdmAKWzAjQh5ZqVyq2goKBcx/
i0ggHGzqcYpMcPQ5fH5pAm3XzlajUc1mqA2SOlfgI2jLKbajWkPePRy4pSr1KIltW8E2OWhvdYmJ
bVSL2MUtKLsSBtp7WqHS4puYziqhZ9Uy2wMEgD6l7yzOd+JDjEgoFlvTA1Hf6T6f11fQ7Xd8IN7A
modRNlu6RPuoQoxadIHKTeuwmLyzg+BnChshiirHqrF+fM+ABqfd6NaKNiivnloqkxHoOuUvKIqH
aOOuYJ2lq5A6GuPfiAzCiodaZWtGBhVJdH2dmR6OwSZJ9zugccjnlBSnMf+C0JML3F6ald7cfItH
FO73KbA7FP0VzZCsOYBg16CLr6dWQk9fG2k3HF+DtnDBGE4Tot2y2n25gE8WD/ndCz//yP8wLaBu
MsUfBpHvPWLX7ij45/6Wjh//BVFLlxwuBysb3aZMh1nqJOORY8U4ABpnIGC72B8K9wCnv+7nxi5g
rLmJewH0WLv6a/NUFx+jq4opDdYcimxNMLI+1wUesv1OzOKy+skhnviHGCVmgWKX59vwZ6v3rE2y
0EFPDVVplgp5n1ZXyoBg1i3jcxQS3DyL2218dN1rVSD0G8XpUEuSjUeGlWBk+FlX92LMx3xgU+hw
riuumhM0atO3nf72wY7qwNjxwUxlQEEe8JGGtuZMMCwlSEomsVR0M10REEzaB4/Ah1YtkgwuPJ6H
6UGcsqkz1Sqvu7ycpAZGdvBAI2A8iugerZVrTrnhI1wd36SsxqkyFwbJgrVwNV8nd9HcXPQUkfq0
Wz+dVhWAXzUBxFeB+K/9b0/oarD3CivMeDthSYpaHD5wk8Uqpj1785xcYbwphZoB7xX+c9i7SItK
ho2Zjz26gr5evyBs0WTYxPeko5GujQaXS96IzQxmxLsX3xPcq4DaDzrINGtGGYqFeH/HNH6HUxEf
viQbHKlLifZuILi5yvniFy+p/MojJz9IhBh9o5lZfh2wo+Mv68tIXlsIagtSSckV6qC7qRKHBOAG
VUIJA/ngKE/n9TGyonDNSXYN7UQCn6ptrgIDPr9YAs65ZL5umMU7urAES3yhlbkECeIHMi8VyMpn
p3/BDwSZDfDy+L9t7oaNeIgERPiLCwwqFhz/cLAP8LPs1TVHu54+XX0ZLQ+Te6yIdmFBXK6p/qkb
fR6Et0DmC8VhwLCYP+G5na5yykf3OMvjABEDWTg3WWJqwezDEqgvORXw0XesJ8D01pYoOJVe3ekf
sFBe9SUFeQ6cxrOcf/ieimdZ10/4B/EjG2bWGlOzd28aOhHhNAz/XdjM5FwN1u1gPcX/hwLje3Pb
yRZm6FaHH1C44fh9XREOuc581F2DbkbPeU9ycy6yfYbdiy3W4PYwYCcFC0VOaIsh3H1KlwZ4PyPB
3Sg41OWKenS9zvudHS9MBjU68rP3WtBSIOzNTnfpq851Wt+ez9PUHtj+tJ3jPnhCH1TTz+pZ5TL+
30Z7muvaESx70UCp53+bohMLD3DWcjgcEjGBu+5EDnaKNG+VPIcZ8/UTUG0rEme/ZRsSzPfAxSeR
cune/9Fzz/T2PlsMt+ZAJsrPKAFcIxWtaBXbtkX+osBlJ4GlLSY32g6ZqEnV0yjYMgkDc4zfqPxA
dg2z2k8DMx9Yu3YCfdwQ08TkwD9NmflTdLL/zf+jyBjU4ss7ai96YHylEzT1jQ/kH+BWw1StQWFv
6h1i4hQTkWfCBlgev1K55ctSMDvjhzRYQ3aou1VCtGIlQsEDcaZDOcsR6jADXODjDMk3JfJ+5UsB
05iw4E/tmRROyTsHM8hFohRl6Cth4OWAqJON5RpO28A7XoDD3je09znmAwP8C4THz00zETyxruMS
q0IJhX991MvoB3wqRDUT732NLBpW+AzhRhNVZXGOXnhKYTRlsmKBS/IOWxke5M+LCSAI5rAbjeAD
8C5ZmQOevep3bQL9IzCcyaex7jGPX9wtt0vp2e8SkGqCad2Boe6aOWQQmAF43WnrZ6MHO1+PT5ZA
EV3ljlbWlleLd8dnFOpxvcVwLBLvFHWCDEK6BMQil9gaZ5hCU1n+XyugIWM2iH5cF90dfvB23wxw
vOY37HZGHDEtUt6eFJPfSLuh64fflcbaLvatjlkyTpSIlRiqohmR8jS7OJ5VHR5AgjQU8bxvJptO
FNldhWwfeNulFeSN9AkKrRFYhO6XP5efLzKJHTB3V6K65UOdazWIO0Uw+Ak8Hm61YdNnK1xIP4E7
VMl7ggTlN2yYjgRyfUxZzZPqIsw6UuoHgd7RADdEEY/NjrfU5dBMu0kKbKo/LAPo2hC7ASboUafo
bwWCF2LexffdW5//6QclY8gbexwryvB8NG8/gQQInX5GQwmY4nZaCQNDh4zIh8LfUMHjEFhHIaU9
UlxVGE/woeUC7ldB1ZMpRCd4l2J/QWH097J59QlaV9PtE2YD1N46fPGC010SPBb9lzT6Wibvcath
Mq5o5dwKDwLo93rl4kjfDER5zSdDjso3LK5boPXcqoPOIo1CBVZ66KQ1VUc4hYkAth+BUiQLpTt5
/U5jvobqtS0Tf0MC+5n0Dhx646Z2H4NfAVOBomIaWirPrg0s4UslDUIUK5w5mUgZe/F4X8EwjsdL
O7Cbs6BMivk0ioNIO/McaqyddZGzZ28D1WnG1uly3LiHdODoldWZUU4eKXxJc2WupLAsRz/etVYX
oRUTjt6/51sqdej5zmNvPqXTnGoVGeufkRyVTWBVFXL4p4mL97PRZcB8uMyWQSvnA3fix3H8HK8k
SHfZdOBm5iz8ctI2KmbvsEMe69j4qHKtBVss39iHkCpEn1A2qf9r/ipitSeaE0tQwfEsNTs62JE5
O6246YqOHqLZwnTyn1WUJiYNkvQd1tklGHfkxYZK3kW3NbIYLp86eF9vzY5pRwpq5seZxmoJktxW
VlQzuNdeZh4n0GEJJAlSADX4EeoAVTla8+TIu2e1NVtq8KsbXJwPVwmSLoZquJYonkOAJSz3uD74
iwSf8v1eGDMGy0jbQcyJ/FkeFSkVKy3jhNnnTy2E5lM9o12GlSW0Z3jywAczCANK/nRCqBktGcVP
X15vq91z4BGFKxQUDHlUVRn3QErZw/VP6glD7hER/FuJTZQFf6w3fALXU8UpQZsVgWxVOTFNE2+Q
yCUBRhl9RIeCavsG6mWuyqX5i+OOyv8HQ1cl0OuvOnss3B8bZM6ha+xI5IE1jIaKG5F5jQKiu5+T
T2YIekaOlp1zBR9xi5TWSEaab1bXcUtHPVgTpw3nf9I7MZhjOKff2lbZdiuaWHsAH+WsfNmiei13
yaQ3VbyUDnYlSSNBV8/wsCVYsunVgNk8eL/jXDZnp4ha22lVLCt95pysPdKO1Oyc0JYipcaCqyud
sWt04IxOu9VPeAa+pFKFa23Ft24wHofeBEjhuxFNxo/B51E0cYt+if7diD5Y/DVrtb8yd6ABRx9Y
YMvoLVVgTdZOedLyOERTmzVvwZpKL6p+0SIAwD7Df20iZUokb9LdaDnab9VvUOI9Fjb8yNOR+Quh
Vf88i1z0LVNo4cDatqQF+qc3MxAxPIcwkQAqoqhs1NE9ooCUOHCxZxCnMPrwrJbGdDL0TGjG35tE
OGfrxrPRDWHao4n2yh2j08FfjUyb1/TYAFsRnCaGFtIfFGqFqZXCF3HfcE+qMk3i+gVSab6dUOa6
MR3C6ZWCIfGw6VPp/kIjbkH4QwGj9FdqZF4KgzMaTHK6XM/SLsUEbYDATSMAV+Yjkm1iR8hxp1mJ
u3iVO/1QuOAWSzEpHIgFCvuHK7nlKKxktJau+IKVw38zgms6UqKAlf2JVtGMYNZu1kKm5j0sIPaJ
YGIjKY4l1qpOz6OUncT9KPO1IhLvvWLysfFwO+/TzAspgYUWluzcuOhOHBkISuvnODQevXxi6R4U
QVISTdv2510D53ye/CVOD+XeDXs7/BQ1BwvsyI5/aUx0IzY1Xe5o9LV00Qw1qyRuQMOgJLhDof2D
1zLVD/GhCZCJWDcbGlr6d23pJOQNv9JuUZ5BHBIeAh2onIOgv6x+TOCbV7lskf4xMcgI1f+ti1Pa
yAeUYK4B9vRadJsHJ6VIYlAfbY+Ah2Ph0U8YExJSVhkgbVDO0259Jn1FU2VOGNHaLi2NwbwzeFIA
WcABhMo7SIcP3vxjzqox95kv6Jt47brqfUSZHupK3puM7t7+Xl+D3uGPRK4dOUEB8OITlBkJlRJh
MtNiOUeOdcMwbtq6rPCSCBYJyxdJPWoS8SPUtEsMKq+7fhW3qZxH7pQi/Etk0Pt05BzeF+Zj38SE
C/0Tjz6nldRGtKCApTk4XtY59SrZojnrduGVQL15IuGoD74lDTcJiEg5oPc7e2rfHPMr7rQk88qv
EP1UOCYLJ1qujFTpvOcExW9+O7FVeNPvdyt2bx5B2ZJGbUZUrnYLyDYM1PnejEJvOa67H1/jOh4d
fNAG9d/5n06b6Us7GazfMKsEUilv8xETX1UOyTcLZGXQ1q58dvN0sZPHxiJiHi1Rp7t+l//THpHl
dFJGs12cLj8ZqJelazkl3qUdg1fUGgf8Uk9GbdhDUeaLczc1pJVvW8+tIj834DmxlW4TkV62LMBU
bdz9iihITRSQs6eqFTmu4LSB8cDVxYR/3Qp8v0GOr3tFoDrZ8a3KPC6n4Y22bFIlAmDkh75r5t2c
nnW6iCaRkWjujHMBx5tG94UpHdQ5Y4ZhH3vt47fj0IftDsYt7OQwlk8IcXVnF4FZT0CYZt/cez6K
SJU3Vip1kyQ6FCeWyI6qrpFLXyPttCmB4GFjvDrVifdp9IihgMvlw0bbOC0fjZqGSjjjveJ0BR+P
5kO+Ke7qVplp2KbL8BHwgHMp0NwW8YTOjXlbp13uz/8YDt99s8HDLjFFw8mwnhaP7GuC+Yt4lMio
o95RoEs15UTlYQ7bPziOot4TsaxQbYEqBycg+/+nQu11FXNkTCI6hNV3G9ttpJFYTgg5UqgVjWCj
KRWppZYqMSveVJJjeppxYGO4KXihrzrFj5UvAqXScrA+aXbZw+mPqgPh5iy2kFVswiTlg6zUaKE4
VRdzWByrZCNiy3h/UWhp/9mGqJW5kp6r6HY6ulJVYDebd0oKmfZszPdjjuPrn+/Qn9zZPXmEXcFo
a9rDVGFFoFoyPbpLT/5eHp8Sq9nfRprjzWJz4bQt0+7pjDmInvlcIeIZivv74I60vOGIrW3m9LRS
vhDLt5R3xQ/UzAnUH/a0QXyn6PDDlVwDjIOu3rXY+FsZqaozdHakxBfIkxKgZDGgcUV9oOo5Ir3G
EDkiHAFKs+fQLPu1XF5Dqm3my3yOZaRRADaYNVgTx4mklIfbk4+DXkhoU7whbqh4zDTqAk6flp9I
tq6lqhix4AqYEmpdmiS86PzK9gv3rXPvTjCdEVnCMl3+AY40J5BzLcU0ywz52NQx20R8eNVdkApD
0fER7Kt+kyiCVPO+0sb/WZaF6isnLsUsTbEE3UUyhxBEbEXqdsU0l7xJb7zTEm/nwQ/5HfEF4Vke
Ff3aK/0q2HjoyF1s/ZVi+vQvLmYredEMFAHZ2aCC2XK4/kb6svOZP4RbNnJIqioCaUxL8RZpf6oX
CzMeC5IQinJlHPMSMeqLNi/xnXsO0CWQhIul+X99f5CaYMUrt2IJGaoqcZv0Pg3zJFvsfoQKDjnj
YxCEP7gVGZzJfs20PHY2KXCo9m7EcAqsgLbfUh4MDMrb5yho+n5OJHR4MM7ZnyGA0jX9TFiimq1d
TJNpEVRt8xXGGpgmJHpp2rE+xCKwRuQA3vy1Rw0KimxIcLEnNo42LkqiwApgAjVd6gkWI/7a690L
9gJPY7eVYSKqwDyfLfokytqIU3cDWM/YdpL3o9l3EOIpw1O2VJCqxv5vATDWsMs4MYfEWXGXI0H5
24l2KbAws+H3wwyyAH2eU+vh1bkGSugcRnNP+K3YGZZ6jvJwTn8nwJZY2MS5CySXUdhwwcuIB8AD
R+BuncrxtGiNn8GlGTIxDpQ0Xqvu36vMB99C72yDzx/NIdshJSno5GDaWa4Zb2PsscDR2+qf0cSI
Y8knsZfGt4PtQOfyXqEudTkobFwtgWlBGP/2QzCje0Alvwbp2wNkEKEt0n51KS6so2KFbYSSD4wh
1143HGDSz1edltA64SnlM8Ff7U/CRLkXwepbnVu6ntmPl6ey2bUQpnKj1dO4KDTfyJcm+ro2BHQc
zefY+xJYiWRmbphatPrQESJC3wjLAGcpNDY2qgA0zKLpbhHQUN3FVDzi7uvDahB8MUwrRCKv5ilL
YtdFTnJ1HoZqBJykbb0pXsx7iScfziUcsHhPLU94mutrXbWFif3/Kz2sS9rhQzSi4T3FXSZXATJF
ugpah2DpDaTB1hAu3YMIXAhQEKr7JRdRRztbswb6de1cVd5eF8TNjQSv+Q+RmOyoD+09K2xmgAjj
rvucj0XTrWB9bTZS51DbJUHosCYRc16OgsPqRW3Ebm3JtAJ2ZE4wpaCz2pokgnQXEdfJIPPqtfpI
xWFXnIxxj5Ft9+mmHgsuGyV5m7MLkWcChNRyaoO09Rj8RKOHf9obN070RSbDvjNHJ2/FgKCIu8Si
pSdgkrI2jlIILqRQf2jm6QJ53J8L1Kr8gn8ZxCt3q2U4ZycLUy3MpNkCa7wmDvA9zo7oSB2ZO9/u
g6/4++NFNKY3fPQDHNIhy3V3E2up8WK1qLxeuPuw4NOYs80ff3GPRYMeoqkv99AgBDw0b6VXQ7yQ
20fxt08UXxGvecFcmKNbho6efjyDSZxnRp2KCIaKRykhTr5QGO5ND4DELvV6rchrU+LHVYBBHKfd
8vKmiYRP8/ZNuqUenkDXZFMBs5mpQ6vREhidDSaeeZbGDcUdFDIW1M7JFzpiJqV8QNpIEVeT11d+
dvKRqSzYQ4U43jVHhApKiA1aV8A25xrZXm9ZV+5QKlJghfl7zcUfzpIza6GCiKZ5PGTGFC9E4/oD
ROs+ZGTvSmS2gobUZoGW8G4gMHN1iYQibpIhagXIqoofGgIEDQASXKavYHqIyzYVY4pL1B2V1mJb
H40MIwYcr3iKxROlubwzb6dzW/aP8LXdxajV0sDh7xVBr8FcP2Hb8lHi0794sHftkFMHwHOCh6sB
LZTeywJcelgYIfyk+WaKZJYOgrzRPswq1kqJEBH7UJtplYB2q9vYPmtNd5HCDLiY5pznXTc1M2iB
VRr7DYFtysivoIpKFPGRmcoRp8uwnRMxvfmXUjuK1GnGyNheIKulkAW9vvJ9FaZ+ppKs6C30k9QK
xT7ZyeTDhVNrH1WUzNRfZ6nXWsrXhV95rJQwroIsffJLYwrEwaMX4jMw2YLA0ty5xrh5Kjc8EF2c
Mrr/4Duk1GOXQqnrOqbTf9KTqirm2JHS8JA4xuZfS2U5H4wTm9bKG1wYmI3XKyCUq2mjd+nRKCRj
IySwnwe9KX4ZGQLMmWgurq7XIcmBge9CkHgF4MEkVG90CpQctOSVMHPjw0a2F6OUr8QLJ3NPfito
QZFVRfy8xpRHHzo9Qxw5dn549E9OwgIo/Z2q/hscTlUJPAbB+Odr6l1+zR6qgNj8aV7PCrsCC05+
EqaFsz8sSAsb1xPG+NzilWF3rLO951sHNrqUZFkW+ptic/FPk4CyYCUmVwfr781QrJICoPF2XIpa
kfyL2p+lRD4RFdzYSWc0GkRZTteFnGflDYLxw8a+lcEx6I/HV4QWZBpQK/NdChnbFOIFzKJbkfBc
jFmxbJ4aT5E2zIDhn9l83RYp87BcFhwgKHlftO/w4o4rN8eUUM1fGF+xkNJow6Y+Xia0F5zDrXiR
FAlyenYYGsHHaiDQV+ag1ECVicuiF8bo2dIhlkjt9HS0dEX8ZEfqljJG4yipMqsIeF6TPWKUQIUr
eboE6M2AHwpYcNoIvnAq64KvKqfyXF8djssiPqyOQMDB1FtErC7BZPJcP1AHWeNgVcWwdhVWXcWK
ORTojJXz2616jtZ6w4Msxe86msahOpH71BcoGhGCytNJaceSibWI+Vkh2l74sJRdGQQrZ2tEqcGy
kxaPRqTfHZIGI/7rEHPsRYOHdlqS3ngkCNIziUXMoA6W3eDSrfPxsM7r2lzoBcKsV+KHe2LN1D9k
OHlRkz6JoWzcbaCDSheejZoq9KpPshLtf6uxVBqiWAqLQqo+o0d+LJuvDZr8qZ/0dqBoCeJGO5DC
IFSpELuj4yKKG2kwCymZ7KUWpgxZrNpNuPRJBl+JDafUQcmpJAZf8i5RY74/GFJc9v5kPLbGGdGd
qXijO9XlSWyR1EOC4hOdBM4Cn/kzI/fkNSm4flAi5Kn+V3cpi5WUUgbGN5A+oZuZPYWeS0sV7wmp
3h8pWU1eLZm6vM4cQ9jVrUJwpdz9giRJzPsQlH7hpkfhTmw331tKIG2x+TSenHbax6Zz1VQxNBx4
QaTHn8rsRZHa8hnMPUkfjHRteY9B2Fj7k+AicXWOU5wFlBU55kjP+PTR+sdNHTdqf/WMRmMN6ciT
RildXSmK1/pB3NOeg0RDWKZQ4PzehRvZuIyZJxQgVwKRuMwWkCpjGpfaK1J+lZ2RVG6rrh7VIExZ
Zm7Yd/YvW5jQre1lvmoTVTY6IuUIYxn/nh9zZV39qxPuLVLA5VRycDTu0QQuNrRl/acGSq11nmoz
hTNVlVB2njXhUUi+by0ZI99k2zAhYAckE2HgbY6PYzbIRLXglToJYCV6LN7bTldruOgbj1SYzynO
YMBDOCfCgwF+Ox8z0GDb0QLdLKn5Ce6pk5cyzAoRITgj7mCa26nbuZEkCYH5z6CfCW2tZGlHeWFY
nipon8EHQagSeqJ5qWp91mjdIF2FhXBZw9MnEdncF4LdQnZ151G72S3GMwIalVqVkXDg0tGhkdz8
iBsOEftGyEbtwb6dD2awNdD4L8/ca74nwrYBcuISboEjVs2UEi/2MERhVaC/bnemjK9S9h62jZ/T
qgOpxa50d8AmzNa50VtZe8qU7VtT+QQZrPNfJnEjpaFh8/GkYFmQeoKNOie7G6IzIBUa0Zf8+ts6
w4Va8dUyP8PVlhoRNvfAM93ZHS4Np2kTbKKDGjpEUE5BLCCgBDeOmSTlKL35jQ1zmX9zKsmdr7/Z
LfjRWmOVN5mlSLgggkYGcuyJHuBvZjcVpse9m44o8dcFmOr0RBz+TcSJGdL8U50HTBvzzxvDPH3g
c1eFhZMyhvp+BBgvKDIHvu1X0fXpPAEjO6YWZ9LDn9VAtzTZ4hvOKmZFR1OWTB7pMs6T1mfpPSQs
DHZhNHNxe0gOcUBmD4Zdbot2e/4tZHNFZfXq3MOWijkmdQGX8GYgP7oaJrQ7LfBGP5ExIj9ozB2t
3ZVcdRDP+QoDQBdFeqZCkQSNNkY+KdU1Xi8XF8m0NjBYbbaHUtBS69A1TFXsF1lgUjBF8OQLlrzM
AouZLrBY1TfjxhzAREo9HDZvVr5imiFar5C4wwiKZtClk/FpPQBpPCyiUt1/XKgj1pnf291D0feo
JhEEj2YncbBjdhW1SNORXrKV9PK1KbdPNtEalTo4IGx9WSHdvdnhzx3hbcUL8sQEX6JwJbLcGqeJ
vUy8OyXhfqsf5iMkeCVnqe12W1jl25TI+klIlcvRT3gl7BIHEEjzrm6g2/5p7DZP2xROgEGDYCNR
Vo86saXw1ORjvMbz58e2dS/YZgNgLn+pl1c2UK+IPwT9HimsWC0ADY0MWwA/3SPeyaDZw6O8WiFe
My/GTrt62kZm5bCkAIAtMIq6+qUv56mZxQ96TAIQ+Dd1Tjp5h31vJbkfCNw2ic1bmrlr2kz70Fw1
US1i/8MTLKPfopMiv1UKDtJtCFvxsOZH8KbZsNiLbC/C0yBcaeRlLOUlxnsXTKcvJ9lLY36VjUuU
VJRDuiH+j710W1kin8tqfcm255jI4iF8wslbXLYFOv2QFlMONvpBihcyaYJ0/QLrBtQtPSoTH4mN
qM00I+Bg+3gZpJQIymRXwstC1CBhv7Mcqu8CG9kb5ItG7r6EkANrvb1BOcgxaJVYgwMfoYKH8v7E
8tr/C6tisYUOVdHhS3IZiIR+IVz2Ycq2R/niArhgUnxSbBfCw91R4RNrEEYCAmaEmkqC3LQ/mKVv
45LHiO2bmexDQ5wIjRo9Pk7wdY7URIvjKsVVxfByYBVKue42AZNBvxokHu/HrXjcZUbw+/sALd8n
J7Z0OcKkvsO2ROOdnF6GQ/SxIhVhlAl48oXe0BIkDC0l0XcdZSeQWca77U4HoMDOx0STq7t0tTP7
GrJAJ8yjwElnF9q+Pbt8URGkVTfvF93L1tvO5zTqifX80L0w14P/sjWahdIxJsUZt93S5N2EZ9ME
c5VeHtR7g1+EWciryttItpMVc9UtXRF9PDOrZIhOSLeY3BlgGtXdXVWm4A8LeNx7sp3FEW2GbyHL
VfIA/EvxjpkBrhkFOJN2MmKfaAzsSgQTxqyGc7jIa2yuhU/JV9G6vsup3q8XKDJSTh/KG0iq2IjM
bAr5lm312AL9FSw+hQy/tADHYCtKMzCalCGC9/pjwIiE1XLCa0JPlVk08SUyBbFklCVCjG4SnD1d
+H+j6+Zm0u8MdA6oA39Nul3Doc2CG/+mIsaLe/qgAAaJFflwwLbiKZCU+nhgsxfwBuZFLWzibIwh
Va15xIB2J9LRqU8Pd7irbJvOaJZ3Kn+b3NAUdJSoYjz4BUilG4KlrtmEifqcqOK3qyvUv8NDENln
gvVPxABhwCttJrbFLGd5U3cRYuCl+BpAgFYD1S7sHr2vIBS+ARZXjClAu3SDIBCwMk+hZ83zXMwo
dLvHn8bff/Ajh1wJL3tnwS3a6z3KkzjPQ8yeQZtRL5QC/6lhUoVSAQr1m1AMlgUJsSCEopoFP9+8
DCaEyOxRmLToX3rv/vgZ/aWamlMizvothmAyjfNtc3PZB7PuBopx+uzlLAEP3vS6blaTBZYYXWEz
O67CPILKVwxQL+cLHI/gpFdYZy+x450CpbxlZE7DVVeEMq5waQRs7ttoHj6/hgj+C8gOFRPA5En8
Eoi2n9IrsXmBh3ZzxuGgaoJNZgl6aFi7iaW3E0uSfL2xaAiYXzTnPms8gdzlja7fXqYsGSZxxO3A
NcKJGzffZwX2tTSVdmrNsVVJYe0pBw/LFP0YTEw/xJAHy5e39RBKvxoq/UvF5M59SbUCmjSErXTc
Frp4i+IFgI+vjeDwhVJLVkwdEwh+BX4fRQSQItHQnGSDPpDkkByXIm/eTewcAvWxlVbh0m47YC7p
EiaZNg7+/1adGSFecqd5qoCeBCPzbKi2eeW6puHKkNJtyQz5mxkSAujWMTOgBydLh49jHpwz0Bjs
bMOGhuWxDaUaRBq6EmobaNh6noqfh8Zk4Fk0h7rJZcVh+PbmB+BEQzwm+AC9ZL9rWPubT7rAxgi8
bMEqjPeQ7lSstFm1nOr3iyjtw50o1cqLIBOYYttWJLr9RUQ8NDyNB12vIVGljU5chqvOvf+R9kxR
7bozbll2CjQnqTz2tGGHpEvbwB5ET9PLAsrjSZL7EFdklucei2ZAO1zX6i56nv8AkdLavW6xV/Gb
SNT0nHSXKY5gVPah/hTKcCeaA3rg2oKDxA7UUcwSyg7j4+6xbsv4FMk+ZkaM8spaBNopQkap8poT
gwpzH1JFfAhKR8qedygp/S4FkoGbHAZYD4LUkYwdJwdM2+MWc6aQJzeycWxiP+JB0y+ql8tD7RTY
5+Qxl/q2Kpsrkdde8DUsYpYZ6JY9rv67x2G0tFqp85XvsoW+5rYzk1dWGRLLYdLbPm2eYuhgSCHc
oDz9RrTd7dImDCTCJ7hVElWC/k5uNc6E+mBuYhw5P2M4ZGbynb/ubsjLiCjSnAji7NLEQQpw4KIz
dudTn44zh1hAdtnEiJ5dLGOAoaLw+7qdXlfZYyTjv4zSCGU6yzppdvci/kaLeTsl2tNbR/mFDlid
kKhpGjYV0HSwo22YVpL3Tk6/QCS7YF3b4SjNZm62p63Y7tuwEB3ysl3FZE5YrXW4BUy17TqPvBFO
5rVsf2SKsxImxeZFp4K9pmN3LW/Bk1bezMylB7Vd3sD6W2AAFSs28UhqCmggq9tv0hpp+fu6lUWw
xEfJfSX8yxgihB4RGq5HmpjB7MULv+p6ypHJCup3T5llagxaWw93peAsBGmjoGvtZldsOqYbgGXI
VH6CaLAzz3JkL6IEsFdBrtHqtXmU+wjwWo0TCVM4QlD/hLfzmfjNb3sVQ483tWyacvMM0o9iquv5
2T1h+tnGGcqOnLHbMZx2MMuQiJwUNt6t8n/RsvmyvvgBv5GBSslHHXRnnpO24nhbEJWACwXsCXOn
ZvBlXTlYljTaWH8MerMzWUruNc8IP2oGr2BY9qHfVM30dc+i4r5P3ca2hj3RqEmPhRE02ksZ/Y8y
/JmvKX/h5Gn50FO8slSvbKXGa+gNnPPS4A/zeQ9wFbhmqkeQUnWIF5x9AiDqkRA7vCgcRXPzm9kd
VV52RRJ5w7WaNqbW0KyKi1Tla8IXCKNNCDhk46XQ3qYnhuOz5jTayskXv1J+t1Ywau3FoMQO842L
2NaETh2Xno/SUdt3J+xo+0U1lmo4ASl6rxBeTGGrUuIY8+FZ6xiYU1L1V8zjgFSRtzBIHsgt0m7p
JyAULzMNYAbjVocuOb+0sQRStxeV/8IrPM10YTws9hClNDkE5owZsHo4m1tC52MfdVHTqEf6hG54
OkGgxeAEvqt3T7vcvCdKYiz5RrvIojekIWJNwL2MeRIWGvGNdsAY3IW/phWgE+sQ8IG2dKfvWwvj
PHJ520ws1H7LCpXfKV3ubDscdAyfhbkqun5c66nXrmTGb8hsW6EwTi+rndk8UBtjOy1YmbHoIDbW
wXGBzcii0vOaKQu1eUGwG+lcPtgB1GKCF0Ql9meXjxe5fc9A4IiXW8zfuchQ2yfn5c1yRDcLUeqj
9CgOEy5mY1HjdLpand8AzS7B1f74rG1KbTEhxuubYEaOz6oIVql0s8Twy5qjNmHZKOXSPvayu6E4
Wd/JdptDfR1UXY96yw7nEYq5j7sPhbwcvwDu0YbYdm7pnJsFzDqe2ORf92IjfVMW3mTrqRjcc1qX
aG12f8Fzu74CEY8UXaEj6EQP20Jl2LyTmH9nnDOnopb76Dn0+rNkzcYAsbsxjnGD1D11UCuxJhn6
/q6iLpu0kbdZHNL9d/kyYjW8jfsRTih6ShJiKKXGTZM9swSOKLmfnH1RdlxMn2dtprLRFeAamL/x
mdbW/QhmBQ/RViY2ALuy4AuE/A+eRF8VFvOVuqYbJ/tS1aM/aZN01fEXjBMvFHNoX3GX1xGLP+13
7PxGLpjAvdZeORR5/qyfecrJWi0mlJJeFhemQWgrky81jJVTpTypDD+g+keTgLZUQojWhz9VIOh+
1aFapzSjV8d2e2Cozj1XZFepWy/JejVogeh2z40buFuCmotgL3JxbUWwqf93zov+wuu1vEMd+jcG
3qSzQ0+QYkqNjQaq/Jg4Zb0R1Fh5BX1zcIdRY2sty9yQXKKoxuhoW+pzFBAU9yUBS6kP0p7mqkX7
Rlcvw2cFwA3b37JNLp3Bh8XvG2/IbDJVbXV4JTRRWeQouXtStdzCqxBmMlIx9Qu11gp3IuUobXtB
p99r8LeeozQt1ygtpR8LGn4ikZNS5KuIHEIcyc/C/v5AFMsw7G3CY6BvkKH/q1KVPFtBFxn+m9hN
SBHnbVzfiFc7R71odIIcovHwSPdXEWO/eMqDo3nd69Z5frl7v4LwzGqeh5srMb7bThsyDpB2theu
ygfrHSncJRRkJhYHNZsnEmZmRV/IGMaxvB3BuDJFJBI6/9lijX02ERfHaPogTClONTzSCEBTXKFe
EfPllfIWauCvZKuoNeYe4myjZ/HAibWUuapQNitBnPDDjFVgU4EfvkyMtk+VvskdFUhMZu4jefIv
+iqVKNk2E7oPZvzU8uwYhBevzIHoN0OCHA2oua4SSLeUg/uuU27Eqe7zSNv0AtiKouj3Z9pz+VcO
UyUYrUknhILEgayYGs8L3t3wNlo08GV3Zi1t+Lo4QacUWLL+BJlTFFxuyCD5F1ijV3CltF78+s5r
DbyhJI6qAQfL2N26ab2ttV/m77pYg/2o6NuqUXWDywd0R5kcOk1AFOHVl4AZpX4YcNSWT6YFyl2s
4tg9lVU8d6cVo4ZQgOfHHvmGCqcPMWw0YDYAdif4NoB6Ett7DYk0a/L2ZSsUxRBsC5GBpFejwWjz
r3HhM25BOPdKtFWsx9i6wgV9EVX5RVWLCjsnT1XCpppJgL1U3iAqfW4y+IL6QvxfRdoYD9PvuG/M
2Q3gzTmtBz9bCFPq5X098j/OpC2xmsqcMLdiU0dDTIoSB//WsKjftu8RvH8VMNuBeaRAQ99Ei0iv
nGYfb212sS01cgF/inwYv6d2Y/4OmmRBDKYTcYSsCgUM70XsxwXC9SaZZQppwvBxQjfs2XxnGeK+
g7+F/VcJLI+KyaKWkRRxLuVvJ4SsF2urE4Zfu8D4ZESIQ5OcwQvpBsl1w0Xi04e+N8lWxd5tQyfY
HNLCoX+KGo+zpKlz0Jifwq5D0+lC3BoRvHxRLWb4VBLPwuvqo40wjIa/jZZYlS2AF9P+QfB2Jsep
X13ZiBu15OdUjhPZoSVK043ioh4dB7z2nwHxc7JOEpNDSRJslMkSBi+s4AUDYT0Xo0Xs0gnlBEkB
XlWnNgf0sofHc3jrp/pG/jNxk6xfz+wjCc4ukIktrwH2Fqxqc3S+t7q6OsGR4SbuB+L6e1Ea1die
euu1iG7Ph0UE3gdnrWX/x8+vGxVy59zqjMgKncpIiFySCv9xyTEj7pVLjqjMoGrXQ077soIUO8Hy
QGT1zpRndjThSIPPtbP9++O04cDvR9WaWzq44Py+itWUnj0XqgJXo40to9QEAcHz0AMqGrZkkUlK
/mB0H1tgBe+ODPCXMIt2wUg1CPQl0qhlpqy0oawJRGv4q3nhSHcEeg1XB6GOcjDvI0vodX4WVdhF
Jis7X+yK7o+J17c8TylbUc63TJkJrLHau0M3WRb7NfG65T4VR+9kAGcLaIXEhCDXgWpxJ7lahuLh
W3etPrkmbXxo3vefds46wgRkVnP0m5hWH0RVM3vRE/ctT3g8rYiJnq3NViLdWyHGGTqS9hf3bSNC
hakCvlWooRqc6UMICz54kPZWPlW9wgWQSp+kti11pPFsVXfQaqhzYNXb5mZ/zOaxFunFadqPdBKM
Rs1JAwBmvxV/1lPau1FWgmoraJ23kkUYJGOJmz3VxaUlKMbjXzkdk4eR7rO7nzeRLDr/fueAxOQ8
0/jWGvc+nEQmBb/RtiHkPDmMVoetpJZ1X9tROKWeGCanj9EMU2oxWOMZco0SAnGwpzQx/oApKHI4
o4gJBPMUKQawrxABI0vr3Bzjdffhhbbya5iAdI6h7ZGDh19sh2ASQOXMiImYU/PT0j70hYlL8dUr
8kMFaNJyPi1NLTPtzAyh6W3wsl4Qhug3cJc6URtsgUYFt2CO53O1T2HaKsefWWwWr8o8pJlWkoqs
oM0vUT9aBTdSeNl6pgmKP2PHEzXR1ln47Cni/r+f5QO532tFA3cz2FgRoak4BG8h6HGPSmZ6ZBZ1
4XyBMhr/ikqhnN/IY43Oc1Qd8ZxFpDzmI3lnCMlENZRnaO72fpTy/aBOS/dlYhIWfHlZVDN1eYAh
N+Evcp8wRWO/3Uho0WXt+LdTGsP5Ex7JK1U7nbnkZa5ysaSS5a2T5y49O2LLElvMwp82qb5s3zx1
qAdINDaX3mHxY9ANPPcPIlMctjb5cJwP/VrX75ltGR2o5erbljtAqcEA8A62PhMAUidZc9eSUrOd
Q28TqtXueyWXe3jKow7puaHfCJ5F64ThW5j+CcI8958RfVqhWnMvywizSwgyX2KG1ZEt20wAeI3e
oiQcj5CQBv9P4yFBnBj8Oky2JsxEOkMdPXcnbszN2IbpLegqa1P+dvbpivRWydGJLYJ66aEk5kDY
Xpjjvjxp7barYj79YynL8JFE5SU0v5Ec/DKfrLQ4lWQMvcN6CNvTYOic9df0NGOpRJG/zEam8fSu
WlAEilUSBEtl7BcxgbjUnCijLFjWs3mVcHQSI3BvuVo9ooBnNGUPBgHxOfhWqusCcNdFhEUVYsOq
mYkCTnOM8jYx8kDWtBvgCndm0vIwpJebGiP465I4FO/OphENaWbuJ7Hsz+N6cOeJxiQqfiM2ms64
8RmJFCfnxLCV2N4SI6/o92/fR/SmGrUT+fo8ZhQ13m0OgIHXmPnnBL4XN9xVavUNaM02noiJq4mw
r0Gpm+It1PGGaB6mxhwJcZAsdHt6mF2mTWq6RoxN+11lPVUQ050+zvh7X+j1yFKR0LEaXLzrs0LW
yXbl+fyPVetjnPgfd9flFU0aHYMEKDfxuxjRea4PwIoL0h1G1o4D01qSkh9jt261sE+FxgPXkaAz
HcSm/3/jJWtII+qTZLai1z2kkVsJKDtkk1fEZ/c4WNbj/i9LsMQhbcQDaZ9lBgwXtr2zKHsdFkPb
9b9f16ZIYXR5M0PSP1YDg10SWS0qCptKWG4Enj7cSJ+dsDOlvw1Ig+7oBxAuPOxtpPwXSSKBQlND
tOOT3h97Fkxx53lCaq1+N10UdqGj0g5CjCo9OSsJiafwu/pDN1Eu55t/MLeDs6Kwrp+PVUMCFVDh
hH7gZ0ha3h26tFZ2sWxYhHlP+nR8ZRTxemFWC1jO/O6vlpFCvAMGv++zuUp0WwaDHjBHMjVRPdnq
TUj7XI5n41+hZYCJweAS/IB+NQKgsgCr064VRUWBsWVyZD9N4Q6/pJcG9YE2Y+aZqc6+1dBHheZZ
lOy2LkO2uWteJVu5wWE9h/2Oo+Pnr51/1iPeLQ5woWZighlLkEpNECC9vTp+AupKRy6LAvM+bc1E
7VcSrlj5dei6gZX1St4m/uOdhiQJixe044velA0r1RjIsFuqp2sgR7LH2QZjiMkUZuQSwV4YG4YI
CNIOflx6w/lD6cxeHnp6HDaWO+Bodah25ODohbp7f4D5bV1GQtEHO9NAEhcdtuyYLyBARnD2DmQh
4mEvwCSnBPgY7/+KLEOJ95mUOlBhaR4U0Ae3s2uZGJucjfhUx4K/GpO7hmOw9T+Qtjkq1RvDyj/y
I4othPYDq2LDkArrtWDlwnA4M7F3uYaTR7VxKaMe5N0AHNLeS63NRannbJvW3wYAR6kixLwqah0s
PCGaC4fh0c/grhJapN+VmXwqG3s8jHhrNi2pEYECc8z/4jRS3ELZyU5SICD5TTHJc/eL9RTTi5T8
YOQqmCn8KWn6rEDEFgHctIQm6tuGTG24/Ff3v0i5ulAAPDxxVKMohKasUfFuji+Pv5P0qwQu0SX1
tdQfEdU9hxjMYd9tmxom/ZNmpJHYqOtYiqu6VORbS8MIrVZLAswe6X8B0QGpXDRwwjXlgxfgvr8u
IxCme88XKY7YP9CFC3P4vnCnQp+4Qu1+I1BH7BrJTjqVLvepMk02AA03X2tFfVa12BUg3PAhc3sX
It4M3QLRi4uSSN8HpkOSNyf3AikzCHljGWfnHhMC5dQxQQK+zzrwthOakR+4qAHTVmNy+BFXbyUO
ViZ9nXNK2GcMfXyhjLi5Dt/C9dldOjSc1CgRcwFcMoEdB1HjzY970i4P7F901krJIIp/YldhiNp2
9aqs9rLILWGC2DBOG6wnZeVVDgUgIu1JpgPBiWQbwygNwiZuHOYjwjpV4EeJLE6KvBezhoCZXS8n
wMF19W2z72eSf8Awsl7gRhuFuc1d9ZGic1jEqgvV0Q1mlVPKFAtb+yIys7m6Ure+AI7gXNkWx1Y4
Ogxe/+5UiF+VnBWd6Qa7z6bxgLt+THiyRm8H7j7XmMYmNxT2F35BXUY0r2T7R7CAbFmM71oBIQwk
+iESNaxEAQ2libEhv58XFyrFBi057cxGxEdhuOFGrN5T2eTgJZkHle1kcspfT1s538zj1iuxBhI2
C0P5Objl1mnZ58Y6/nwQ4e3y8Q313G9mx4v2LsPGvCffWUA2SkdGaLIkih41jo+MA4DIWDzKxMM6
7fgx0qb+NB0AZOPhzJX1Fi+5+mdaeerBu1XpfUAUnMnjQAAh3VaKUHSo4LuGxQBBFU/jgY1qJnFG
iQwFiLik9NSKr+QGqBYxTjwTK+Ue05ALEhoBVxXBHlDOCFqtrR9xbnfeOL+81OY/35lxDtC4mkN5
ukitgQKvcgaXLms2sCjPeSwLBXFCYJNFCrvsv3O3wz7/BdPw8axmpJUKHGMlf3GIVzJu4U3//j+x
7T2tYc/puK6eI6eUO4cCk5aBal9YbIgJZWgqmtRn6e2gJjtkxmUsksAA3wSJtQDy9wHDwCqN5hl2
wy2X2alnjWGyqmHmRjpMP2yIhIBUbUucKgL03oaG/L18TGWhxCxXOslyVQ1Vn9pHefoEbYSae9bu
QU1jjcxMlpJFtdnDejea44HI6S/3/TdA6vq89554Qk6BWP8bIqqbSCUfExvEICrTXR5nHNjhTmfv
QLd1o2/bFFTIg6GjA5tLndADcMCwqbHmTkommiZ4ynVOrI5OuQ+aVnhCLq00HXY1m4bGk85Y0Li5
oh3f9H8ZHztZxlsovww6jCn3AUWPGPyZBc67d1cQ8JrCFTvQe0PON64ahmG3SYrFlbaznzlQjqqL
N289gyMjlyeoey6Kfz/Bh4FB6l2u2bL58ClQJ1EE0XGNEUUXHKlfbuFzXd6p9DqfRghWFuuO4vB2
U4K0ozjNFyEj7EJAYi+/pwAMcLzYW2INjWewPF7xXC/0RngDAjJm1/JQlav13ufztQw4sWTesCEO
/95Ycc+vaSlxECkjWACrALbA/0id3DE32AySXzo1OBujFJJHjg/F0KsrB7muRf7duPGKPfX9+ClY
+Gf6icUI1nvzYTbMwksmt1H4uZxIdtVENt1gV++T8DIz7JZg3M03ily8W7tPiIGqr3OYcg94ZGKB
t5ZxxbtDFf7nPscyThAPQHf0lLp2wevhkBu/AMx7d25qcmQ2UoLC/IqUBDKQlP7MNAoE8S/5vhkJ
rQPEoGme5wtObC4N73k/gOoH9sOhpn6CsCY9ClSL5GmrmdFceyv1+5c68Yp27E6rZUa/DtwO+IqW
h02ddDilepOIkbMeSjr1IbRj1bES3zQk7N5aTKhTSTWU8Y5i692QOeGnPttJAlO9+Xzdh5r4oicM
e3PaqezvU6mMUJj9jM+IPrLeEVpZ7fUKgvXKuasBbo10I8oLzoJ+VlWxOTsDVR3vu6RYXmIIQfKW
pGcuz+rI5ZZAL2cz9mGVoY1ccZf6Q5n+8ri6lx/ibO1W4p3nf1blP11MWDJpXVt8n3vQ1epsMAvX
PTmCpXpSwtHz6M8XGJpaiALGGPsSI9huDNzF6v8oyW/AinHmGZM7ml/rOmKsxU1Tu67H1+zt1+ou
VCgX6d8Wfi5owFU4kes1zWrk1Z5Yn8luV7SOi+HOPK5LEmIsKcebLJvdVWXERQtSsTtWc6AECvsa
CQqxtmZ1IxLvLcWMe/UWt9hfCwVnRNzijtq1OzcNkWKNwVjpg0iU2vWQEoMgbXNIr2SMI/tKSNeU
eaJFUQpKf1TL9UKgvPHh1tGrewYiDggJEQAGyn7eAxsvTFVybMGcvmF8m+rzMbyZajKfOGDLz09S
hcTH6bsd9Z9wEmpmRtHX4hUzm7sXouRYD6jbhKDeoShMwdNozPCihHWmJUYgilQQgMrFW1Xvb19V
u2eQ42ubILToUDk7uKJVM4oaBu2PYWxJhy7RMG9XCJGUPqtSSKyZJH5FPl1YS0VNvUTFAik6zJcc
kMyFPgBbFaGJ1oKNDK+BvSvH6VNVaRIbcA3Ti8STiXsSl/////3T5KSCyqN7AWG9sZgauYNAFIx4
27rD77TBWAWen1DbLHr7sXKVSERWGNLx5BviRAffNy8pgOh/F7PSo44pyozrNe1tsqe0DhuBPz37
cxuCYgnu2jtCzZ9+GcIukhndWeO/EHFef7/1uYnjzRBBWLN/kPI3vfPOd+0bMCLQJ4Hk1IIKxVr8
0HGUETWTJdcwZYnCH2UPyYCzvLifyEehTurH3bXEmd5E0VphxtK47LTuKX8AyZyqfUxyqa7Of32g
JiXwwQ0pEoeXtFWzfTgkIVTbtiIaKcZuaRnCrOqACmph+yFfzcV7oJhOyQmtQcoYB7Oiy+aGT2WA
/IcD0NNHyxXUcHOU3Ya65arFG+pLBqGBszqV8w9wbH2Yoyr8vw4xNMp6ZBkfMLd+vAB2xkpQP7F5
CwJWs+Ba5UYamihp3bPQhtR+s6nD2xyZEu2hYG6wTRph9Sh2DmqMiFgjfA3OZGppB72rl0UvA0t9
Z2ghOGhviiydjit/wlAJ/Zpr6HZeSx22s1vA5AerpuFenHVPejjxJGuWKNkPtNoLt7TZXCli3GZA
rRzkPSpLNaMoeuavDRjeu1kojSnbWvI9wn+gswkJNsmC5s+QKq76kGI2ruVn1SMYXWOc15VpHtk5
03ShO6W698xT3/ZASICbp0IA9Twnbm6E/w+LY3IQuzBPjVlLNbCHipCeNUvtzhLkpUzcO8tfEJKk
/lP2/+hyKWHRaKz3cT1zBB8rO4CZJjX96VrPVB2kNFDKqtdTjm0l1z9QjUs8R5SAZaq1Kcg/B21E
IK6bFeeLGGfpT4OtxF01QbLXwyedJ85wqCvsLhF/mJhqT47NIyF9w8ZljH7zQdtDu/rEkr/Ai98Q
nxAxk++TotQKBCzoRBOKjLexOlucbnTXLbBovf+TbcZ0U8xxvDsgm11UvhwjeLJAADbQZ7a/5cGi
CWnZ0b+Z5VtNhDDGEYioNv/pNfwgsnwEBxWB9gxn6onAgRegHs0Z/D5Y4w3VXrmWkMV5hOEjFJvm
tjzZMQwfZGS6g7tLy6PW+0Un296u09zGcXo0uv1lX4deFSPb9AibdjLY07SHsEgshEs2iwKt3UNi
KxW3XNhxviAdYWFnsvu/sLOSUpdrcMaWMFtV/KIuYB5dyc116T0jYxC11oJwmdHa7DP1sTeilF7m
tay02I0CW7tOaTsHEnZscOGM3ctnf2SofXU53qLkYuHttStxdzy6RhR+pj8ThrOeNOThte1PfeMD
hlXilgpVeKQU9jq+R7KNE+DwMRLQq6CbH7+/uljuqITHvBKCD5x/mDuecGBjcNCAIAZHCFV03iaD
kIzTj9ugaOAWN4T188Ht7A3Q/f1jDCvLt9cIY6YxzMjqvNb3hD37IieYLWQYbQK63CRad2TPyAVZ
xUxE86Aik9cl3fueVNEFcymrDqmL2Evi4727xKz3cu+xDEtKTJOpZssdPY4rD3/0IO9UFxXZvhhb
7clLfL/QlswAOHg1QPUDjU4QEVqJbnfoOfe6z71QLy3LAE/7Cw59cCjLttoSYxGMpRW25GAFhvzq
4HGCfOPLwjR2Ly3/YRnZxm49MYQ4r8USzYt9kCL4RFrkuqSleRdSSWKbZCtbEflHMLhBnZ11dQiz
Y10974Sn3VQ8oCNeKAgW+DW0g/xi+Hv9/4ZkvFnDm6XodoXWL23K8d23URzkzA+TW3s6iGZvzwX3
Gd09cFBe/SFQuXSyLg4hf0HP4ygbLHvULbJmzPZZF3hnhQ52D5nVyAFeioCpVgCK9S15zbTHGIwy
BeowFOhP/U3AfnZWiXtGVkH0yFZvqHRFTaj9eptzW/Fwa+5Ip6WaQYX9hKQvEyFUHfE9NjYtcXiY
T72zu5m42CQRiCYRmRGeuQ6Jq3b+U5lZr8fMJExQPaUrcLIHT3PBe57d/PVE5d/qlKi0/+Ix9Lmh
C8wr+tWyU7WN78SFhnJ6/9k2ISTphTo9nNbDN6kLQxd7dJGcp13tb4DhE9WwXaV6nKRgkbATNgKt
lye3u4/jT33V9tVvytu4u3Wg1Mn6+r2x6deoOUrsh1K79PmSsUG+bvZ1EUK0wOsEUF/FgTKJnIMw
YCj0hqzpnlaHTso8WabV1DwXUaT9nZyxoPKyPQNIATrY8RKuaYDPqSYuhO0+WyUgTupujKTICp2m
PduBL/lx35fDULFZSNHLF9lBA7XE2PLRZYH3nEavXPMAYOr0P334lkLXz7yQdgcLq9fMAffFj7u4
+52xSaRgGw8/FPOVsuEEYiaC81R2ovxO/dkjR5lS+HRWq5Uh6Z/dNXEKGu47No5KKrzVAja+3JN0
Ou+VBXaJ4RdtnrDmXTi773YtcRc5qsJIsU/fxSjVR3iOvGLtbIIT6wZvJBYpPAPXpgDO6HVLJsdz
hy/sauA/KG4LuQ725xfTXLjrA2ObbOG5iD0FFFJWQd+VS9RHZFbUyxqfqWXzejBySmPwMAji6RoS
cndB6lOY2XHzTQX9F8WF+NgLMS0qToxnZsVhU2KWQz8Ic56RwY4SJPRGtxGwtwG6qP1qU1M0kGR0
40oGQT08SNsWI9UqZkFvE8SqmkNeK26Lc8bj2dDPnn87IrS0vwfeSuXQssi+F8skCT051UxoWOmr
rIiXR6KtXIzpOWE1k20gzfTU0AnaJe7KD9qZzKYSr6sbidd6k8prFfrPwkieC2oho1XBL8ebLheW
ZJcQ+73nd2xsWUKhzVxF/aIGAnh6gjOEXXh5VpB157ZtR3qxjYYWHEPPFbPE3O/Ps2FvCn6SoBra
LXGdyOYDM/7j08GKXIppQ0qJxWc/b3UmEKus9qFqbB1PhF39f7TKXm0vrlYZS2LGbrHwjpgZy3n5
cfRjVGC6MnMVmUyjgMV3bOFmE6rMqJVGu2aaHePtA486GRTxrVi1Bq7+bmwZ3sQfMMdUnfUuVWHm
xY3L9g7KvMVJxPpKQkS1c2wgtBgNk2s5/zHZEYQQhwEPpK18kf7HluwM2hXY2rDfYdM27Qxcx53U
PHayH/BjRDtFig77/LiRrOHrzDi2KB+sK8TISfg9pK0I5c/ifEGyI/N5T32ctbIt6i3DPKNwUXyO
mY4rFOJThuhsljFwK6FZ5S8odGxsw3n4DF+RajpPpcI/p4duCV066zTb/Apsufn3xBGc4MG1mW5M
VtFYuYvX8aX0nPWldVTXyVZliUcqNbIfnh901wLVi5885an/bnYo36VVcTl68tdggK4oeiibOT6A
JmYnSDduri1JhrKI7zCMzXMDbtbxFGoMV2WvAzQh9TYodFQM6tK5kbzmpdGG4gXajOoF2vUqKrdi
aTgPEgnHW2i24u+5wY0PoxuqKhLgWqJhuLpv+Yp0ADWer6umof6IZ1U8NSMviMzll+Iy/OfFv70B
SMDIpqNBy4T/akaQU4pkjmM7G6sJteu/rym56LABlQG/j2EpzubAIUST8ONth3UCFK1ltvrBg7di
5jUraKco2sDTjwn5dNtqqUxwGNw6wqlZPxRMLiqY9ET8zDNTHLKEIKbBykzlI6mYK2z9tYyTE2DB
6WgpC5a8vwBokHgMIwHzH5HPGJv4vNIuaKT2NiYCoDRd3VAVNXayxCtXva/OsNxGIqVsZIvun1lG
0Ag8UnThZMIg34Zlu+IVFa5ssSkkqZs9rGMMwiWQb3tnZrK1VSi5crLyixO98t1eFPO0GPZ3/kCf
C33RBuJaXH6PaYQW0qStix+B1ygmzNc+mc8QkLQFiwDx0tYBmnkv7j5oNa85dqdE1FJwiBKI/vj6
e5pFkWTvN7K4HByRb8uyOtVNPo2IdY7kYb18NxXcHZkOm/qiUNw7t6irI0BgR7PAPvaCi0oOsE0X
5uns3Ylc0rF8oTz95G7qn9GnJuhv1sRDQ5y4FNwjw5hQb0gLbSWO0rTK4ehQTlPWZmpX8TPWRy7w
zcUDTalGD51EuZjU6DxNVIaW9FJ880o8xawNYkVnIMXSm+TYQy2UCglAtdCan+IM1NjxBwfxIO4M
EX1WnqT2KseWFTNMwXCWvqWAc2gkol9aAPvxV6QoR0to0L86Axpefz8Bk6Nrvlxm+giQcR0nIe76
Maa1RFfjruTEstpdatxQbhDNwMFiapnLsG8uN4DqkkHuhmlQ01hhxVXsk8sn65N6h2k2KztW+yOV
rB5fj/faxMrmWtIumCxI6hg68sTgWaNZRKwBSSuHSb/SsYKIYMpOsw4DjA9mmZ1R3mFsFnflL4Ly
sXTCNRD3isTKW+Avg5Yu64LLnQlTekpkFozKOjqLR9yUt/AFMh4OUdwYU7uZNwjqk9c/GC5nvm4b
s+wXLqMCQJqgE0DBv4+KxqzRwEJYSR4zLYkdj7Y0DAAweXg150GM47Znvmxq7cW8Wlw8lKhv/Dlo
asUz20a88lCv8Esj9O7Yk6tx2gQqaErwXl87gi29SPKxKGscHlBvEyifmiQPnUqa1JfXI/9PMBd4
VwT3CzcLuKnX23owY2SodUqrGuoCkGycUmfLx4bcWxbE9tUaa8OGpDdLHoliS9FNq4hbyHgYpf5P
m/o5hJe3zKqy23E0OpHldFC03G2jHkobwHkpBtuSKMXKPjo95prlcCPZHDGvlqX+P5aHoUOpOOcU
6qnjGCA6stxqrP+YvlCXnQfj7SJtuhZgdom5XrjFte7wjPlj+IZQqXbwsiXeHBMfKwjCMAf9s5Cp
C9h3AX5ECoFGESev1QXcz7QZhWmeWpCiiKDE/Hys5e/in07jkC7Ni0TCZjEZahJ4CTeDC3/NQ66j
ZlVBMMvANPfI/26BRjJYBGIcD57eN5odMRNmLGayLjGTU+9EiKhttCfuQXoNei/IpcaWD38ddp/b
9H7CcuEaPim9WYdipFRmxd6RiCFfETXyzLva7/LJzAJukMtbe3x5U2P/T+YMGpMStytTo4ACtPcS
/uhYgTM78orlPKyQwmaJBa3y0K9xzWm5cdSRTLo0G22fk2gPtfS+p8RdvKUshlPrREz5mT1OJmQE
iINfpVhBptON2qIyc9is2GEO5bx/jwY0sFpr1SeXB+ix+nKb4rC7v6QA+4tgoFuHPn0x9g1RtveK
OfZDlZojjDzaiJKs0smXJe7rfwpb0lTW8Ggqv1UIErX3nHdUmQGCpGtq+ppRbwY5RcNLSG/Gha/5
kR6I7v5wovfV2DPC9p+S5uS9SDA8TmhRl/Zoptyddjfcy6NLCxYtGvvx7LzUDt6iBxNqRmKV4icd
SAYNAhDhY8XnfCJvSjLANL3X9bUBQFrcPcy8qqezHVc9uX5clUeiMtsewFha7ApQaZ2ompPUpA+9
iIoQkH8YCyFAotQxhG1ii6bkL7tUbuWB74PoNxDIrjN8F2gKhQjWWDnwMWch1NQBoWRdlcLxGoSE
CxuMKyJMN2VEQW2dudNcPN5zsZrLYTOR6AkMlc/le+IOWsGMRUubbH8+9bqkWtamOP+R3vs5qILt
b/M5s/Q4V+mbYsAHgP2Z51W3UKrc6yVQYfx9Lf0XF0szNtk+UXSvScPbSw9EFOIkEcNUpt6ad6Sg
q6scLtiXqZrviDLCO3r11gGtZGsStxUz0/EetKvhS0kIub86kf1B6nCJXCKjW2vNesvvMCRC4RvT
0R9BNsCbOpNMLg5/teqhMvyYfTQiTlIeQg+4dQwZq1NBiNxi9qTQkpDQxaRSstBGOlYR3DO/wDOX
Gu2h6BnkHicqGvkL7u6pEn4zpVGV+Q/o1XDFQp/IlRz1LyRmpNWp0jYqcgelOXHe7q2CHRtPbi0N
C6D0YKMX0PFRx/VJGauXIjn/a6SMV7CpGeZjiQoHcEHqMDOKcqyfhveBVnT5CJNyJlkqdkHEcBXu
+J/xXJAH9o0IMFRPDG1esjIBMHc8VrhVKQEem7sOYWAx82d8Yuq7b4qed+w9XMJRMLBbFb+rQyDq
OGp0tPF4zXpouz7L5Co7htOR1/IjGv22vsPMjuJAjR+3ZBUKm8DZkoeUZwCHFppuyU133nD7dv9R
ekfApNDSF80c4GsNLPCuHOQSiXzktc30yX4Zk8HVeBoSznTVN/K5WcxKD0gE1LS6Brl6WyizF7ta
Fi7q5pbl7UkFzC67BWSEtRU0zfs+HOiIgupfwOK0RYOFwu90JGq1ZoGQmnsWjlAS43BrYv6KEn/5
4YltavjrUFbGxvZAoYoAlBkSxYzvDueuU+lXgeS6iB6DH6RdJl6TxEKpVNMFWYtmvMiDyFNqwSGy
4TSOiHLg/ENN4zYEn3LwefO8sHh2DYWFV03ZbTmC+/mmuu+c5QGfvfyD5HqDurN2TJXHdrAZqj0t
/H0k+qMf6tcYMPniCo6fslP/Z4UJIKwx0jMjeBO6//IEGAX1vZxBm80fAHXCLp4EX/nGL92o2c89
IO3aB3/E8SWYHRNlB6VKAo4iw9ugGOUOhEPrhRaTvUkm0TgqoEhN3sbl3fCxap311kiX8mfERy13
52InR25fjnWFz+4jPUAkvzxg2oFPh3ewTCiz/Jk2Cc6kyEnlsYUk9j+yx0aZty7u0YtdlnfRr6KB
yoIVnuEsV+Q1bsLKu7LKMTufhGJeBkBvQJAFJxMhHIpUXKaJhhU112R/Ut01avSSHR2n13cZFGr1
Ydirh32NM5vZo06XkSpxz9tz7sotIKAL7NdJp6paXos5L03Dg18DX1q92WJh1TIPhka6TlXlTjBr
mNXU8dyaV/HP/tKJesFm1Dpad2P5pDYke8fEwQIsuqq4tiMlIqGs/hDbpChdfZSRxlLK278VW1BM
UJOFabJUU0iAjCZjnmYMgQ2V714T3kpxs/X+7zB+T/+C6f/Jh5nCxXMpFGWNK08ATNXg5EaFm/DB
H4e8Ru/hCVh+GpynnI3vUZuT8GSsJIPJ0vOue2la6W4Cm/eSFn8dWD/yVYs1PWh4TIg/E6L/R8x4
K37xgOJtUmXv20wmQTsFZKnqVXmE+HS9hgfQDKursRxcTDD6glrqvbuIYIYGGmUy+kLXtAz1WX3i
Fn7mFm9ok2EC6HhOREy3vLIjAAX2zts1HXARBXqlkBGWBUwNb2fBYYL/G1+SDmFn+3qTH0vhRbEq
CcOUCgJA6Tzm6FfjRHc3ospOmAh+k6+lcu9iKfQaMwr+ySHCjRrIzYyhK18AuLrZCzI3Ddyq9oKC
XSbv9jTs77B2JnRFYsqiPDdh5ym+3pzBlmjH9LWZzp+CXTSLUzRZDJ8qIThkzZcl7SNtPdq0UVEV
VNSjFgNzitj9xhYQKI8m3usiIX87E1tXUrZfe1aJtWZVyR8bXcSZBs0axsRcu7B0Qu2695EaoIQn
XO7vMTiXOXAI720Us6Yu+aiVPIZ7JP6as7qXjZpLDXNX6v6xWix6GuByiZU+EwGqoIdodoz9OcIb
fiMsY7l7emr6pm1Y1sIPv2e7OSSUY5WyB6lOPMZf06aRuQrYdc9owtedCP/oiNGEUlVf3rnmtZ7M
a7GyHN5tPLxqHa4Nm7K8cGgY2YNmjy0VBitz/C5QFz5z19nHJwn6dcEpx3ZMh8+8RzMV+zm1t0BT
T1M8KqhGl4PFcW11xUKpkEjtGfShjGgEvCslrAlieOZi5yEZXzYU3KdkirxhVtS1Vhngwi+KM9Cx
etxYsrt9Ig9QqJDweFEKfu77NIKrkM+yXr8h0vCScWv653VW0QwYLkY4SgwTBrTldHS2o2sgcPh6
x6eL0HIaEtsfQGcESDNkjd0BlvR/XD26SaCboGxs0hcrNy82+hxExxEKHLmcRZGrIAlYNjisF2ZY
zLxK4SOUDg3p5GF5VAnKkc/jlLCuETLpHWktJZENvgSIvkIt8FnrmpC0V92KXqJ3pRbGbG6Lj8ZD
FWA9674UQ5xN3Hddw29ayYutbJq78S3SM2rw5JoA3C36nDpws9WNpCWy9ovj7Eu4JjAtZ8e82EYi
TkavbvUQXMAF19K0/+Pv7yRZ9VELx9rWdqOMX7Wqy/1QKSQMSLEqHI8xb0fRvin2WKNt/eFC6zdz
kBp0/+Ls0lUSIH5TpgXMmBT0aUFjh1zQ3bxOKD3+aYMDTgrr2Ey2l3v4oAdXb2VURtjDbFhcGUUy
gpa/IFvRTZ9x0a3K9mjRp78eK7J4NXl3PSCVKeSsK98Q7TKQuHC77dZ/Vunfb1zAR/dnqfRsjakw
uAjiFTVYrtf0PZaqEjP1mGVa3KIQYELB7JU5WcMJs4GZ0ftgMp2Sq6iBAFXiyfozYIyOCDgDXYc5
QY6yw+ljId7ZnOPkqmYwMd2dAPqZAw4viHcYbNmY/1V7bG10hUjjF5kbLOWtU9P29oF68sEO2Zxl
bIwnQFilh3PKnq4WmCg9iKIOYCiZmwdmufrtYzdsk2CWReviolwgeUlQqMxmbIykiONiVkrxNPfH
LRi2+XakWtJhsoBBnyEqWD/jIWmQGuEdyW9fbrS2dT3rGyEd9TirlxHN6Gho4Z9CFmQvah8hg1VR
5eJCW3tq032QLEt2Mcm7A9J8wDZ/ULPGZUyFRqnGstkCgz69pW87us934ijmdIqxW/eZzWqFnCyb
PV7PA2bKqgxQ3G0BkfWbZVa5NQlCcchi4j3+FFDEYUhlvw0qTClKC9irG2PAoxh0xogcUED1FiU9
JGVcgBsMVQHzJt70EgH8ygccnlX6MpbWGZmF5chC3RaYAxeANZHiSAJKTYaH0cF1WwulDVUJaIRH
OKt7g098ujlJIbb/0BJt+SCaC0ypE/jMY28jRzWSPWi5OlWmZNk3DUSZHOiPKQXWb7bjuOkYoT59
O7Ie2GTUmeZYwfNG2mIijxucE/hUJOD4+32gnupOYD6G7e+JqfKrlbb+71CgXWhOjI4BcgPSIAIo
kAxOWZoY75/9PM2rvZx9BbwEr6Zu3YWxxfZ4sdqSzzU66R0zeb07i93LXm80aIaKsnKgMz7o2Pzv
4J0K6VvfZ+Y0OL5O/HQ5QqwE7Sncetsd9pYR0iXH9eb94nnwrhOmokIFxqN9ZCLcBAH+tUWpWWm3
UKhI47FrxZSMrHoCn4PyC4gNp4fEexkGCghuCz77eYU+Y/9LxqLTiUxVpkMcgkFXEIXwfkYvm2Qp
cZTnZG3XL7p03VtumiuM2xiHcr6wCPVQzslHFZQE+TwTy7AN6hnp5rBtYq4Z/TMtRYU1U5PcMjw0
wa0zbbWoRUpwRgBu8LDZiLuAt6J/8SBuzyo9PpdOkbHWdiY0kWcukp4/Butl1K+MDRYZ929ToRdR
5vnEe2K4CZmXKTM7aLcjNfW+A2aGatJlV62pAy2VlmSB2+kThFVaMpMoxtVYbA5c4BIsgoqBQHy9
27x+cWkC+i7OMOh71PmUJPRuQORVwK4t/xcip7dJrQ7bl3mS6W4MfBXc5iN/T6em/NuTOasdgr8h
U4xpRFhlFSPK1oeSE3nOWJdxvMePMHQUZYqFDeWdI87keC+cXOYSar/grh17Bv3qvOwa96bQKDmc
SHni3oqHRbR1SDZrNwVVgCMvBMTjRIWIjJyEKZeOJ+qz7n/3mCXMHgdKx1yw2sjaGyyWUiQfJOVs
dWWzPqOruo+3BNG3WvzZ9AgC+K5TeBpZVMIrbDzq2OgrneM3bG2/8YuXjfUH/fd4T3as/kfqdDpr
CCkBOvVY1Yz0yqQI3CNN0I25tTAxVj680KPBisuqFX32HIdmUUEvWP7cRNdjJ53KZyqcrlaYRCfY
+7JPT/FyURJdGmAaOZoiAjiUvuqB6quYLhXZX3gKhtMgxUXONMSqRnloYQKkgasys2h8n6L8joHX
BmwqO6pZC2TVUnXlwnZX6wIZXjtF3LW8whVYLlChclO6VhFfLaBXDxkeSbPylCyokF/5XyHPkJPT
9N/xpn5ZCd6jcy/OZtj/zXLht8Km21Pjm5mxuUSYsu/EEABXEJmLk6P2HzwOzydGcLwCORe6UYB+
eaVJf05wRCuUJa8uQSAi5twhwYbxp4d/x0KKif72/4RaRg8F69QPJPI44T4X3LE1IaQ1Nvs4SRpr
JQJg4IpcwJtPkuMuhQdbwuWHP95/TImx2vfcxzL9d4q4QS6yiE6wvbNxCAKcmK5s3YpM8KBb6PGo
2fZ2S/aObicZAbd1RBvQhjCCluNNiHCs7qhiVjKE+VUFnii3301QwlvAJbNL5MP7UQ305nSKEKFZ
wY0zUfaWd8WKO2pMTBemEvND1p+HxgSjploYuwALRYe2rKbJ4KoL99/KWiQKLv0YCv1z9ZtX8/H2
8d3SzxeDmLUKwQ1xwyHml3qI3hTJYfyJOKCdP5UdDK6hH26ar/T2dYBBrrMVNxS39TAJDl/HBFTn
fgRzQYIRx2viZt50A/u/qRU4947uxM8rIIYiVGgZhcssUGLigXJumMRdqkr1/E7rZ8sd6DSuZP+e
cgSB4E4ShL4KbGFyEpmWhutvvfys3qRL/6hoF16Z/vDv0WkJX4VeGhJYDf8Fpkl+GQvGwKl+GsHS
o531Fn1cvBoF1yVS11ZAlWokNkiRKjXJmYI3W/BfqCN7AlVxKuiT6Jv+TbBwdcqD9cHpoClOw7tl
/p+5cinwQZdu5i61TLtRVvTNRb19vsLy53GCY+uMyI3X1bt37sgTWliWLzn764t2uPyJKlIxFES/
hjlRVU504aOgLkyfrs2udTpJXutj3oXGRuPIjFpTAph+NwW8uf6/fkpuQfPfLsyuKB2fi5Ifq828
qHSXb7ZUApWv6YcOv/aByQ0cPWqOIuoFsPE5V1FjW37Kal+Qu8Fp6dU+EaEmBZy0v5g+hdgrKNmg
dUglA87feb+1SIgxLmzztBYHzCK5AHCnaNqIFiM0JFnPPFzmrQmpUdUfG2Ypz226vQEdF0hiOiEV
uOeuYFZ+z6xWDp8jutNirGH5PZe1AyuSqBd7wP2xwZ4Hr2sBpmnr5xp/GxvtgNPQPHWn/OdNjqdU
DFgbYXdeHZ54R97vReIArdbvkawN5ULOCTWR6OnnzZT/XaoDV9XYDO97keJ+tdoP0iPIHlQheWYA
HzL9b80DlJUbdhOLrcGIBCEWK9LsZbXVrjPYwFqgzzHtH0blaAj5ar0bXvwCi4rTYwmWgwB5LxNW
uur/L3Scfc29zf0zm2cdr8wHdhGQFe8qQL2t7gVdokZ4UnkJmpHWlM2HMXAnkWF/qKPpKNY2KyYT
R/AB7K4UmxJzpaIni3hH/tHByEcYsAiaGa2QU5eL5BulYK5OU819vteMZl0oYBt/rCicXOsZSA5o
RvEH3q30wubi3PnofkbGBYiMMdtCrEUNQ8iOzi5D0wX4yRwR53CTmhKgaiYBGk6sZIbAIPpX3PDR
RmhY6GbNVLgROIjyB0l7lBzz8NMKCyHUfzYniDudhOGRf4nG+OahG+aJPhX+fEJTQwSwyoB3pwl0
77JmC6jw3Xp/yPj/ZX/pZjwanmrCRVWwSX3r5Jen2Wky5ixVqS3lu/mUYxXYWUlTHv00QX3IA1BU
0C16tGNsbB3h7jzvDjknJUqWkYjZuWA0x0IDe+JtWMWD8AbXjnYp7qm/C5m+uzaD5UqjSUN9JXui
p4VyEjxfS24iDpynVywHIkptg+eiU8DjcFbPIEV5KZcAo5tDhZeXItpYy/T3E6S+vUEEub83vqHy
JUyhGX8o5p5h6mq2NChoG7bsUqOZWvfNB48Je1nLrB9+ToML80fKT22LM+b0V7sDd6gyruWJJ04F
aNYmB7sU5lHlk6doQaYTojXsGuQplkxxMKix/5khbloGPCHYA4LdCXWSEGFDt0TP/RwZEKXFHHM+
3gxDY/w85BjTdC5KO1+ax4kaQUQShLjgFaf/wEZDhfU8xPc+RTtt/Z0fvKsDVZ2t15TpnLprl0LE
ClQUHjJSArAlCeh7gAcmF/rHNUU+F7YAD53vdCeqAf0EWcYF7ph8Wantsi1k6LixTBK21Nws8cGz
vcaOQG17aayBYaXuSHJk5ZqNtKzNC+JFJAyQ/1u8bV17T+aolkJhjTZ6jr9gr2mAQwMI+lOQnPRE
CCC5nkjHIQv7zyFjVI+mAoIeGwqSymzahhGh1Jpf8ZDyLljcxPEcrJCkh0aTUyzplKHXQo26/sI+
5wdqMM5JZnhNH7JqfXQV/s0C1V6dpcKoAvoxMPSZ8Syiqp/E7AtfjqfhGf2zxwOkCqtBndakxKAc
8WoyrDYcCkXKOeKbE0kOaIjqwjcyAxSiIlhPfLvsobOYuN5GBV3wLiV1hiNvjOgZ7iqTYpEv7u6W
YpC+tv67oXtZ1tMRnQ82cQPfaVa0kg0weC6qqq5tpTo8NWI6uJaDfc/zddRWihxfa7MAWg4ODWjh
W+5SlcwAm5CI2kKn9YSm9/mstIYWoGP8w2D868CxzftYbWOIH2hylXci7HA9RviNGUi8PtfyFziR
mkAiAi60WMHV5dF+IxLWs72zqRnP8+g9XxRYonsnNc3k5i/nI3Fo5s6VJxE3HVlIssLd1p+SLMlH
h0r7JeP11d/e7HY+d8eHpgkinlS4tNPptbUKYm6VsIWCMyX0Z1pp7IxmlEXrhBPa2pTwOcIwQfqc
0+ZqbaDFPAm5G2hRPReKCrqSWxnDNLGTST8WpBWCoUxwvo4V5rEauY2RSYAheuP5u5EWAVqvdvQo
wiKNdDg7qSUxGOSSAR24Wc3GCNyQOGGZpW3H5ZppP78e0UxpAzbP5z7A0eQH3842e6m9WPY2gDUN
fjjpEGy4vx/j0YCXy11oWZTkpHR9LgP2S3Wds8Z/Jw1qEYPD1YpXk7P/cbW9ppbKc+Nj+OkPVpxM
H6sZtGJtS4ZW+JqoSV+SAOx/z0mMObaIZ6XRPYPuUfAp42K2i/lIwfTtW2BuMIcsr448P6bI6nEO
OinKQVgeORb8ZVfVSefGKCXLYp9duZYN4JZqDFqHbEYlvJY5ncTVFicPMPeDHJB1USS/fwM0Yk1D
8LOmHdQokwrstAc2v3r7nGSyJ8KtUbloNzmtrd719kP4pIXopfyX04oE2CQcPWop9PnC2+w/dPDz
wWurnKyZ8AjuhIPOnIMkN3gfrGfErX0IMvPSEBbcx1J8y0IhE+hR5peLFWPr/4GiJ9TNO2NtR9uI
pXRsxvDrPBt18mW8KU6fosGImCV6AFwfRa6OrI+ckk7zfam3ZMuUtgjnCCn9sSpzyChEHtlt3ATF
UdKYBN1m5OAlxOadPqIKIwVUgdl9kdbFac+R6SFKV3lUpfMrL8Nqc/QH6QVouhLAV6uw+gX6aIcf
bwuccSDJ0HvAd04Pcw9GqQezExlcjFOEgZy4huT4pLq4aWuZbqXdskpRZWxSep4dfzrzKHrPuPim
fLcCIHbopUdzAnKVlpBc7U635RoikiI2gXePb21vxa3JqVeZ1OCIG64h7rzoTWNmmg5bDmYcJN/U
uFpyfgs8l67246FLitU/+8QedLknf4GOsquSfo3bCP6ZVm15DGjdlIvhaRGoPTD+U0lHbA7ZUmyY
zNi6hDdGfY2T77SKEjQE1RZRYwDGWP88DjU96R6aoVe0GDvc5NTRChCkT0zakzTRNKPmsO4Nfap8
oKz4tQOj98Na9R6kn9i1YZHkYICKuOh+rzELK343BY3XjyzoBxy1JHE2l4pw7vg2jIHvn6Ov8Seq
K2gvlpY/8hevydIiPS4McDMGEHksQtkjeihYqwVq9YuJAot0jx3ZR2foWLG7mCMraMzzSmwSvotm
IhZTIgP7cY0+HDoo6ead2qNRxAPxh0r9wu1xRaUODDK8R6MgNUOU4ZHMEhUT7Fzd7vJZ41xu2mvb
gNT4JeRYHWdCNp5r/MC3NfkEYBpiuCbKSuXi9i/udYYw4n/o7PU49kLbxl7FhU+cVEi6LbGxMOop
5DeWN5IV+10B1ydXwZ1H0jmXy74a7payX4W/Oad3HG358sxXE8kf1vQftIr2BzMLL6KVfs+YHvU5
AqiKheVxuvqDBvYn5c9wc/XRaOIVwz0NU6dk9OZrWhagjIbw0JZw7Nb10sHr2tZA9VdhPIMsuTGt
6WttHvSrrqfbRf3eWU3lOCpNXbyMFnipwp+XDPa8e2tYUi18+rQDV3yAoOTGef7K0iJy+aZOQjIE
p6uTDetYB6RjbrPWikXPH0utlzNCBWp2wLCr2H2ljr4b24snfNT4hFhJPjgvp+52BA1edGl30djG
PE+IB8x1q3gTILH+vL+04PIkbghskmtYTTJoyXaOOPbFAtBKuDQw+kV9YIOhDvS4DQTNWrQFAkzJ
BCTLyuYOTQ4ypK/+/O1wwOgLK5/nSsPIxYQsUgrTO32J2H8qv+pGiM/Ox5W/JuD4RQtIHpWCoCcm
/Sbwm8kGrZQPJETNSU+ljw80v3e7aCNIDDCiG6z3A0A0JpKA0RZ4pjIl7O2mNTxl3lVXLtVOQYMY
1mCeyJ6a4bcXzpRFHVd+3fMNhJtO82iNL74oo7PwtlihdZl6W94MdpSpwqxZgMAIdTPZC8LnmABo
pZLKws7jyHhuSjt9ETwUhSr7qyU7rqGQ8YG9m/BN787hAEtxsDpa93M1fX2qhVn+/lvdsx6JCVeR
7AY2CiMzQqgDB9Xok2TIJtCHZLldY5o5vka9uzhN4LOb/rexTGCRVsOsDVXF6ywAUbm9ETZlMqTI
jDnfaIVB3QHa8P0dzvwGO0gkyNlzrPHxtiCy+u0D2ZNwLGWKTWJqPuL4VUQwa4QYRWVLZZF/xLac
oPSxr6R36glhJ0UN+fMI7KogBckdQGx3fIyNCzE1cgZWs49eMis8yz7LQLVw2zutM4LzMm77ldMa
Thmpi/1lSu0BOGwcAVjm+sYhR/Yzt7OiSECao1Qn01YOGL+AOdvPjs0ZKepz4GypwHv9op7IPJru
ueu1MbC0Vjh6ugigcpUOJPffvOrLqD4MH/3yNRUMvYsRJKftrYKPwmTV7F0+0rniHcbNbNK3kHs6
xCYnM/9xChoycR7cG+4QA1i+f48Jyq3lUI2J5z7nHZpM8DvbLLKwJQeAyvA17I0GP8zK6J1e4GLd
dAELkKH2c3zdKMnrogMoexAxwDN5WQs/avb4ae4mFU3KAwc2egkJXNoLYoeB/iWUdfbDifBRbYE9
aFjdcDnSGA2CiBGuOPTF909ogM/XqtozR6mpZ9kwlkPgxfNq7u+o7jMoMOBPhLlwaUB1fxUG9QZd
as34XwFiTiaul2bjz5JGHu1WGH/wTW+d2hiCaq9m2+AEHpBg0vDlNZGkwltRrf16VuoqLpmy5Dko
SxI13cmrPoPhhg5bo5Oya0789545C6Tay/jsiqP0berUqyVBfnXMvCOTtzAWX0UkrlpE3+d2/O7b
BO+buSV1qL71ZWOZ/8Xt+8xLT3+fL74UvsZAtTmkCUflc+RpQkZHEQfjJbocmCeRwnPMVIPXCvdR
PWLDKOQR95JukjsEudfvLotMjzQ2kip7WJ/9PHDAfSweHf/W4nDWtHKtttBhag0us6xdyp0HqK6X
C31RB7jPTjzdHh8hev5ZcKTXmqGaUJKnF8uQ7btATSv9wYTwx+Aj+KDA2DxbEk2oWz75Ht/7NPKJ
gBJuFUutxCci6bpLAs+ZVgn6vmd41LkZYYPR07i6p0j/zFy/kDl28UwM4v5lMVXn8/VNDiw5u4t7
HdIC5VIHNAB8zWuSLFBlfhLtWI/LmNNudA2lvnIJo9HRbb4QYOuEC9NzaVT7flZw+K56uVtEpeym
YeN5NzgjRol0l/RPNbzLL+DmQ99GE6O5JK+928pIAeJ9roir7e7hIalS2PSGW4yPaNDSN3cbnvWN
pzGD0O9jAM1n2lQk7Y5YMLY4o1+Od5SNB5ZJ/bISl9yC8fCgmBaFFMU6Lywfn/2ZuT+qZb0v3fg1
7DIU3m3hcO7rQ32j2wAyan/0fkZ7srAEiHqlm9shTCeOrh6SxKn4oXcSpbfxiVbioyZSpy8byKDd
DgsvA7HMtCoPrjExcAN3EPztY7qfEwji7276wrKsF1jmZAa4uIfMxoo8j8JeHECafdfmCBf7absv
ZvIZkqs9NE/4EF+JZLNvQaal1/luZuZGOvmZsbyvxIZSPBzt82mHsAbM1K09cosUm2lGxrK+ocGm
yPriAMIsW7AoOBNPet73+89JHa/vth4DXidoD3vX64zwX+F59vN3pNhW9pAW04oz4yhiBcnbDtuo
LcDwjGjzuLp3oR9c48yM/ohWugJFUVRGE6RZdXnbbx/Vrr55qxVNnhy5kMHFR8UU34pfDyJcxakq
5lzNmJCh3Vvwg3R3eKwHjULft0JCr5ytyjxH5qQlYsRFHoHXZJ+keK0KnwLztMDS38rUo6NX/YZu
vu5JLDzLcIMFWVWbjD6HYtiN99mpGNZi1rJQZddL26DT0L6WBPLJd7BSBYjVxEBS4fZf0CrTzsIt
bjy2eiOZ29thpdki3XHpv0u1H63QrTmm9MEv/izleTo6YR7d10VK0l97GxQB6nNsVGT8/9MlvzBm
g9Sbp3Ik2aen4+IpaQZtyIAwO695IA/1osiwchd8tg1iEB7/Zgx5yjPObqFGa7SmG5t+MZsvtOrs
t5hLdZFT+Ur02+pdDzT7HDzhio/R58tg2J3CMaIKjhEhwquKJEW87d4NRP7a2d5ZhFwMxRAYqOnr
7dql0Pf8z3fs2+SyFhTrRJTIq9X0VeOXbopR2cfZm0fU+aQhHt2pl5HpwFHErM4DdmFOI1ajIe5C
xv+2XOLspN6QWcXwqew3F0VvZpaTZv94qdLPEVB0CouC/Ar792co1nPrdEsYQ1tJ6Bb4qQmkXsD6
cctInAuNm1PVDJNlsY5V7/hErya6z9CnscKu4j7j3yvm7fXDRbP197Q5X1nYR10Gh0X7M0GEN9ih
qM9+xPturf2ocpAHS+grW4Vs+nMIFDAhFCza41s21kFkcjqTBfcuCDfjTkQvlVy7J95AGdq4R/CT
Bxq3moJztO1J4crTFPuYe8oTeKtvZMjKzrte2Ubn4Y0SQHo3aHedsHuhp/7UtFRMJMz3fx6tqgs4
cpAVrDQi2dh0SQDsX1dbODl6wKFwZH7Z+yrAyrRjok2ZZo1meuRB2eBqfQveo+zsA+t4lu6DzMpT
0+632gp0EVMjuI/CZfVdeLEYa8bFXNjFnXQxigoelrJgghrC/l+gmeg9jwBVcGWEHevLOh84Zz5c
hbnAToFJB4YEG+Zamo2WsCmiTE89rvVKWtwwb2ZvyJ1prNfO9dA182tJgzx9r9b+VKCOD8bN0S1A
RlEIIZcCsw1Z06Uly6n4Xri/yL7OaoAr0IqJhFW0HXJeKigI4st05n9uXuOruUtWpFHIKNTqVB8g
pI9qdy2SU3rc1tuABTcJeUMQhfOvg9F+ECx7VgXClU9GKAAFlkmlgjcRB8mUgFt+yxS4F3RIPbTg
D9Qj7yI8DYqI9ipnkeWQkmQ7otAfUt+k8AnGp65hP34lw4I0x4rFHmmQw+fd5FVvLDIpDVKOm8wC
dlZJSE0MKnnXvCPS8s7IJYaUUJ7Il3J10drctWEjCvVk6/q+QM/hJ3H9Zj11TGFn7v18lMGmizrM
OHwlYbhwUVe82FZQHTvBz69fpQeQY1Dvc2VsU2g7WZZOlOY3RJKai9wclKdiyypg3ZmwUMB4OSZ3
kfXwuzBkwI0iQIOT9cuWpEmZ28ibJLM8C288xJ5LX8Eb99XgLHtws+XfwRtg8YZOHHlsGAMjJG2F
1U63+YA7ku6P5pjfFzcXMOlADKHp9IyX2igolw/dU1HpBiVG6jaftN6eidQbwbmB9d8zT1XgBO6Q
GIxnQws4vZ0aO23ReQLAveGz5/kIjUNff2/cebvIPRXAvbhfHvDpC/JKd1qydD9xd4C6cXAfDpNW
n1K7Zu0lZPbr6QaLM/rw4z6bssMPV9Khj6ycXppVTr/4c/7kAITYeyI4hOpxms9p2pev2F8BsYe9
4RfrJQgdovgZDZ7bON65hKUjt8bGmvLBkwcPly5o/W7nLhZhfCKBYADqn9azmaQlaXb0OySWiMAJ
2XaMm7WXWNNJK6LMa+4WzmAiYt5xSL5A2EBD0/z9XlgQO9V8OVR8YBQ3LT8M/5FX6Jt+p7IkyQTy
j2kWGeDfsXzTOGzcd6UY9FeGGxVfic19BlI1e/Z6YdTb/YKzAvNgecAidE1LFkOMkQX9oAIVA60/
uoUhh/jo5dONhwfRXml18LiNcU9AA+yPf+xzC+xn4glR04kYTOFbozFYcwEmSqlyunL0qmMHLsbt
R1kVAmPn//XyVft31PJz07fC7AzvTe9rckqBUFa96q2IuYb8Z93+JzF2KqOYU4YcgySskqeze0TV
6uvsMX89QnGf0Gz1FcrPMI5PfSQuC9Gur+ILzH5NzcKuKwpmHuLXsJ7zfexArcjQ1pr5mAZCBHVp
sEQfSfn2d7kjd5fR7WxiPpTmnl5f0UmzKgarvJldykoy8m1EnXvZ+9IH3PqatGkTqqCohlSUswkR
+cZHfGPqzsVKuVsjDxlRWCC6KOW8xJuqbuhPtk5UJ/h5pLaqSyiuR23cwKfxPHao46c0dsqFMK56
8E0SQ8efHZn7VUqOgHncKWazdOvQnl3HC7oh8cGRVf4viiW5WHB27FqzFFVq17U1MgElcNrIyVNM
kvpdY7ytkw7e8nCFzQOR/2XhZo4fAnZAx9ZrFHq66G0Hx+rqo5yP0aaNO6jjpYZGiPvLNYIUEtaW
PJmn7l8NfiAX7IdgiRTXYg4Na33gfXA3KY+EVKi3jbU5U9rVF3AsSkQumu1F9fTUgGw27gZ/Dp5o
aJtaXuLZZTnbH3VNqv3947yU9EXaDVmmN6fg+89egotrv17OdsS5wLDmFSY/x4CyolXZZ3RukZVL
UCSyWXuj/upIT9w+XWRhRh9n/3FlfYokiTghTl6oqQ+CXtlQ8kN1c1fBnPcQ/ZiiYXkmna3O7L3+
noiRNL+CWzBQxAFEQZSOXjEdx3tfvG54XqTtzzF0LO4olZdHh8pBsoi1XmMmCXY5QqxouXyk9neT
5kNifnSHPDEf42i+0OlrqOsWbPH9daF60arB1z3+AGggyBFopYfHw/lI8si48Cc0R6dOV3yqmEMN
LslQB2Y0VdJT4EE0UBfWtA30Ya2mHndGgJDSPKoNGpeVohTxRv/7C+JCIoDgKnS+NT+C26OsymXw
b1HiW8VPJTRumixwlip2yv4Dp1tVYRWRATi1bA4THSPdYyNGGZGrd0ho9QX5ZNQCcldcMD74utCa
6AlIS29O1r6AUxkN9w+23cvo3gBPEuxI6Nxjt9tZk1pS8cfJKlnvyh5f3WkbsQDAvUSapPQyuVxl
pVSIcXwPIDmrCdzfqYzdjwEzFUKIq7xsEWZK+y6BzPJoahjjYQ5Sje/4aEt3+frA58tcJs1hPzNx
mGWjLH0DeW0gz6WbqrPxolCmXWHBiIZbd6FXAdHbmTehIhqYM0s0JzlzCjRhx3wtvpg96/swU5V1
MavHYCh/JWTQlfHkmHPSE2bO+uuCRlucHCRvEmyBALlgo9+LjFASi2cUv1rZ0b9CrUG+KaAuw1I0
E7jWaxN6Z4ykz8TRY1mlZFXiI+RyYLEWK4vbJBPb9SSApBm7Ty+60kQ25So7eQ/NIxJTJWcFrF9v
I6yN0+RIGroW83P+S695ud9git6i42PRxN77gE2cnlyzH6RqZNrRHPimhQtl2kVisG/bl1fNhV1o
0Pvc9slZugCLUnHHnsWiWRzg2lOu9rXHJ2wkb3qR41EEMTzTvyJRB3vFJfpffcwkHw7rYg0+zEnF
APbhGQZ/CWpWTCAnlX4X+TrIcEc4+RgH8DXWUsNeQ2YygTZEtnBayNZkxAo3u1KUnXgTVN1SQhkB
fQoVqjSqXeEuBtBreMe5HGaJtcvsG3QiE+k4sARzsmaXxW59AMJd0w9mSzkEoeIfTeS8OyJ3Ijxf
IzTpV8vFJqXS+xQJsvNI/MKZXM5aalb6VMDqyIvCHB5lUzqRx1/WR8UdTmuTNjN5d/sizto7blC4
z/EGt2itWEoI+S2kNUO4txuT8NW3u8eu2mq7jPnb5gzBhVhB4mduQsa++lhQZXcdilvqZNzvUE7L
KHkxsJId4+3Cd242gNLKoQBXi+2E/mtQhf9GOtnwftfShb9nc3WhSSGlE/1oHGF9VIkXI2UUfsaQ
slIf/mDa0yTUIGKExhNPSTXLwKSk6TzQfStUyw8zWECwBtU+6vbtEMNAoA9uvnIyY/KCE1IPKHeb
ct9RxQ1mXHk6Zus3v32RHxkYCoy3lQXI72biL7S/fpLkGUMAILP+6/YLEyd3sgdYVxsAjRki1iOM
cw1/6FG6Dd7tHOjuXWHGqL2YxQKEIsquZxsAUS7rVkwVYoLz4/yHTEO1Nsc3CQee5n4TtU8kVF78
vaesvxOpfT7h7Qfq7YM8hRiNXtXdrC2o2n/YusxoiYfgQiRP1O8JWEHxf2EwceR1R/p7RP7XRUDZ
nWiVEaBp9xrakUYr8nWnG/YsGkL4XS5hVjR6ICErUjMhCSF8aQbF4WcUBbp65Em+xy/UKoqvnIuc
Ck9GWpu2xn9+0wJKHeUw/9MB9MnQjOaSES9pATLFlp4m/KNw1OTZK8GNbuVBeXBZVwdZ8i/iDo8S
7aWcfBYFjLDYN9+R1Yuj/LxFDiV2F9zBCZNyrnc49WJ5aDp3Arf+ILMzei2gsRAcQcWwcu+b1WhY
q/hKq6QTZuctKeECC56AS7KEIWvst98IV7lIy7hPgsU0LVMuVOKR+2ipXeryvmao3oyBT+MO94Q0
F19IL6b19mMC/1EQv6xKAkZxUaXOvhFh233GqSbgy1yvLOm7INAE2LqAH339Ugyw2+rgNQzPnw8f
zpN0wYMQO8PaTM4FiAeZVyzgujIUFw12ILm5DMwajFCXNfJLUVIlwUidiQ9JosVDXZCtQQJCsGmX
Dvrb7ZwBIvTJw5f30p1opXRe/g6o+I7JC/HmHYMomZqzGBd4G/nfW5wm0jiqcFkVAfZVRpk84SFZ
IJdFnAx9uPzJmgLoqPZn+tpjOWs4A5k/H50qB0D/VztQ7livccrbWTn3m4XrQNHCwGnMOjRfhQq5
vbZckWPw0W97AP2t8c6rDnBA1CF3gXNiWxlfKJD377j6KreYZo6J4g4bRBlsqLBpkqxZ18UCKFf5
cJf6xNKk51hj6LkNBMVTarZRBL4Lo2QRq8IXwjWYD/TFC2mT5WWVcBxWuUBnTxEBK8yQdse2Aad4
tA9tsmUsxp83sTBlw2Dpm+Bpl/61GWNDpj5u14lbJ19gUD5Z6yIAdwo1vw6EJ+jr1LaN+oL3qsTJ
Sz4Ard01Z/+Vhd7xQPbKBxWiRWW6qC+B+krWw8YA6ORhVbRsW6t1qF+aGpTBRl90YWL5C35HBKD1
UbPj7daSAZtIzcxDmLR2bfr3OmZv9MO2gotFaRGXhrRXbsSj31PUufS6MdvaQ7OWN+AduQ+JXIEz
+Lg8SRPcLZ88E+kJnyGS865ypMh9DOiCAZsDNm9TSk2uDsVy6nsYFi27AJGNskrMQTZM+nQHehty
4FupZ1kp8tkQBfPf85heeLtM1D9DZUZpvUNoYBVQ7Bb2+Omt+O3LWhhHwicv+7/PkQE02C32atOA
LnShbo2oYvIRC+TdJj7GzzrxlxEd8/R7H9mYGXb2H2m6Wa58H2W4JVJpGrmeLPMu2p0H6MpUAsR2
5CaR+euSP7w5wEE85AZKN3vE43rgW6IpL13Lk0gZNynQ4n93RwCsZhxGrWD1fSRUfUT51XY9OKxE
lranEWxZKs3OZg+Ek8lz7r8aOQB7+Pe/H9PUxWafyFyl0HKHG4e091Dwzfro2ORdsV474oW6VzXy
bOGOvsShWGhwysreAsWpOx6/AvuF2FNOjzhrX6kIOdTSXT3SmiYuRN7YQymxq+EudDBXIb09GhZf
YG7dj0AMjyD1JUtswv4gtfvqGWLNcRC7/VlvOBA9K0nEp/N9C20hVdwVk8vT+HrZt9m89W1ohm0q
Rq5lx05P/0s9Vml/14GuVZyu+Zg2YSQZJ1gtw5UtLxIAaNJI5Y/RDqpQ5mHNhSC/cEmPjOLQ5kRP
Vv15GNQXVOdp1jL/yh+sBgAYZ79mb2gF53YpRftxK2LCNNdCRu8f4X5FTq4fWei4CX5F3uc8ll1/
cTCWq4kKnLWA4nMNYU8rUeqRoQ7CWXLmod7FASx0SKHeJbMWEsoHMZaVnmZuxxbsiXUuPdJmmD68
Qiapn+DxAgrjTdTumX6mo7AWVzxYYkVD6gLUC0v78UDDNe638grxR6UN9eGNOjRnQbYsP8TwfXKr
NpRGSEYwZpA/+4l66JlIeTn6ASL49C2FJuMWdDs1gyK+pRwtUQj4Ijx/PXHr0c8MMUV17PMHkMhP
Y8YOCOF6JXxUKavLs70CmtVhBDAHGnytjFQhXlJNeZIAVgZmY067fwK0mioqRCS+CH19x1ihvUT+
XDP5UzBqQgPqHnLsAYtJzBN71odVlo/vuU5f21IakvVEx3ePty9sZXEXEWA7HIN+zjH8UHg+HiGO
iThC7VJ9GNUe/lao2nsWcoVe5Qwbb9cjifq6UMwyRJrE+b8G13WPKAovjhDKIL+0h62GLKF9xd1y
1dDT7limCK7KCztgCHESsPwVB6Xtwq8hSH3s3Y6aQ8A+tFj99gZY2hzxvupFUh34Flzz7PyjIAjZ
R043ZMPxBVtCCf9WvhyhXfWNW1wdIPdWLMEIV/Mid3gugwLwe+r0rg3qu3KMuAfmogzzGFd036Gh
K1iIpgPTD1fjN93JTZOfpKCgObLPDCtUDIJKiY+upcu325KZKFsRSnGb0F5S75Q4OQh+wqFOKF1/
CcW4n3frAf5RhfP6NdxVlNzziO/OcYFyQ/ehC8mO1RghK+9S/vGVIhcsB9XiFnXHeTOPqpcplS/m
ORA6zPi9zpRwSoRB0raq8vVkr8kj9EZn7AQhXgz4KgKbu6pLT/jKd6ZzdzhH13KTKWXjztaYaIYO
j4KmFriGgMfnAQS4UnJWlC4S/AA6OIEtWlk3PmhIEQahnrzmPv07Q3tN6gUNc91Dkfv6/SkZRp2u
ib2WemvLVyw3oYCC6Vtu6bOVfrlgrD9OcThIjgqwwtSHLzAFwUK1O/MyYFkIzYup5Y0K4qopR4Fp
7fcfOf5+jE3+OOlOjSGYp/GAeRyBPRQVgNFKW7N3HVrtCDcyTEw/WFeDjvqPRSpDR/2DdzMSOeih
rjhF6Pcm8Fp8hqWxQOcderBB7j4j6mbPFDYTEJ7X//woWMJU+bwdFdAkoPSCQDLLFR6F7YqRoh88
RfDj9IT0JYj1RjfGeCr3/uSpdD7Zk2EGcTt7D2bWC+G8wpzPp/PPqURN1daJ5qasriTZGYDLxMZZ
e5ZdNWszFrWegQ7p7971SLIlGmOIAgsgkYBgxHt9/KSEKQqiXU6LFmIZ+wY6pwJWzmu5gaUNW3os
VRBgfYK8E5c8CjmapzpzKchJIqd+f7kAk7AZDIDjTnCrW4rFBJJulbOOxqiO5LeT91SgR/bLedjW
F2dduAVBuAvs+ViIt3D9VVcYLydeDQ9nQdvlvjXPk8PCZDAVShH6gW3HfVOtEP92nLHUs+4niRDE
b20EfD0ZEJRKJ5EUZr2lcMxLhjBOJP8vw+Ci6xMIbNpfSCbM5TyMykLRIkbmnHFGlT+AgHrBRfyN
GwP0gZmAIwipSL/p9nM9Miogwg6rWOMo40iHlHsOhxr8i2nquFYd9GAoRJJXYXK/DqJVylZPp/9U
AColRT86NB2ESbnq1tbjGGOBo+du2C+7/OqoDrWp6sb6Vo23h5dkw9ri/ky0jxe+AQK0hEMd9FFy
yPfOABOlbyL6yWfdna1x4Sti/CealFrS2IWL5YihXYkMi2ic6yclAkDAAe2nlUc8kzlh8rS9j2Tr
U4VBMaZhURIDEaMQ2Bkot2kZAiQKN5MImGd2q6uiIRkRDFp3qrHBzib/q1MurGzNVhPWr0RAvcb0
SQH+QwmrT6W9i79H5hIJo/TKyOtaQXgNrZURXIlWP2LOIgrfVPPIx5Ri5xd2BGru7BrF89aDe9Yz
dVwbCTDU5FK3zfRC/a6bvF74OL5b/sm6YMDyhnWYEQgP6DfjUaRV5V5BZY06HNEhlAsmFYuB8I1f
S9NIBJ3/v9AQIBEe4EcqoCBO7fAzVOPevFJJyvNlNjDIh1WW2dErXyyQtMoONtwY7xOTMklZ4UsL
XQ5Y3pQs+XS46VdVQS5kBzU267+UFzJLNgfMhzx6huEWjL/vYJ5GNVwnZc6Z/IoTtu8FmgCUbdUs
y0CSdnwPjvwzpjSkeWqoYRG4pagcfO0GW6TB+rNgERwYoGHUe01oLnPQggkaJ4wlUqQvCxpqWWN9
4BrJJxS6jiHaKW+3LjP9PMoQwG/l0QMzxVHRDojuE8Mkcz0z+TgD4NThO9W7KCiLTiuC1cR9fT8t
Yj6VTcZIb+JlLIxqwmyss3DwodXaueABsELXQGcqdFHd+71MikQZNY6xClPjUAQlxYb2eXoUBm4i
XW3gRle45Qktt+ISnulI3N73A9T24dUT8rkdzAEJ+HNDDyetBDdWs3QPiECDbd1v7ZrxC7kmVTd5
BIlOJ52j9yforA4eh3tvAcBuDhnOOrAahHozHKEUUsebZQsagKdvINSRYsQJI4TA6L5V5GSnT8YK
jlT0/FWYDZ2TssQ8DmBT+BVXTG9KzME48jeOdfYNJJgHFDVEXI2oc9IYAHPtmslrJMefVCH3/HYW
nqlwsFdnZsbkiq4VRGIHePhHM2TrxPafMf2MJOW9z17nKN8bTn91iSMddcRGdL8bcUkA0agF3UjF
slf5RumY/+KFThqRNeUJdoD9koRgOOV+omeHJJnx+1TqNoVFADIaw2JOczu2405nmO6TUY/lCq3d
yZHtc/ZTzy7OhhVp3951kRukOx0V5GI/CKwoCLBj4vg8eBtHKYUlzMyyJp0J/Dbb9Yx0U0+KOFnD
6k5OlQkGKPAReOs7XsT+xIGZYYqW44KE+x1kAl70EVfhljwpq4EQ3rWs6YJC+hmS6sjzFnINOQcN
97hI92VdWE6s4ZwX5T/nTAoTNrFm01tcdmAKe4huyz2vqXLk4G8OeYIuxMHVDH74JNxYMp9Vx1h4
ebFN+Q6soSepSvREZhsBPsgh4vmglKIPRWEymEDMLUr35tehCKFDzlMsktp81qejXC8d3LyECpbp
2IEDnW8wE8zRf6QP0fiAKL6J5XJij466gINfpIjm5ABbo2ey4devihWXaz66SDcREy87L2C20+zL
uv3t4CXRZd53wPJe4S5gPn8Bed0GOPkSk60w3KaVSqcubsfbD6BSVLXKrqTOoztkDLjtouNMgiam
IS7GapNakvmpSlXrBpqwNJZG2JA5YwCJcTsISFoQHeqqKXhkp7jCOIv14Jj9UzFUK6XGvZakJp6E
KN6SZ041QkJNZFknvjuiXl7hwtYGdnkA/vSDVQ2k9skUiaM0VxBusqjloNL87sq8TF05uPd/1GX1
855HTAfvrTG02XbVdsxzxUJIptwjiEhOVMq5zQUg5ZYuddhlaPp8NAknt1exnJFzT4avNgo6BTcw
2V6wfnpIh/uKMKVMi2qDXS6QW54RmYG1p4UAOBsmeO3nMQZnAsq5keZm3w82ice5hg4wLrLE+RUn
Diwchmf3jZ7aLiQI+8n0eVpAWWRk0nqIuqE9VrFC70AcXzaYbeflVue2IUB6qgSNPnwwc4srIPRY
XnMVMdKaGDq4XCt7kvU4Cvk24chjpPbOIZ6MnM3xhxSbwUx6n3IsBcSO9lHSLJtA4fzscSHv6Vdq
4xwQTx25lx2kjeOOm26WLfWIvlz9nH0DHH9ZWxwrMhAwmQJWIHRd8CY3uFuP47ijmJaoesXuTFGN
HWAxhUnRprfBXs6ATvn9x+hVNBmkiJZXqOgiECUDoVqhi4mML2Ke+T+GHa8DJ+XVL6Ja6zx4bzpn
8ckkk86spwMfAMHkCLUByiImJoqJY9qIeg0EFX1byRg3QKmxVWZGzK5OFcY64rLt4VkYRt+7oMm6
vuZCGVSrlzH0wrzpVCXQRXVravYAl02GkzBgA9jy3/EqcH/njI3C/1Weg0q0j79wABdjjvo3RbKz
Qqifl6Oq2vs/jqnl9xZkfPY8HGMACkxRRL3/eMb4uqXOIMGqmv0ZFpJxGFbznB+X3/IjevxHGYQ0
6w08VcgdiTq8vY/rS+7zgwDXGDiaPGnMPNpvEA/vaJMeoST4m6Z2P/o3P0vbowtvH+8N5duEKfka
VXPNaQBxba0Bi8Yyme2gFVnU2/BGRND7ZdGpaC8MDEmJpPfPCl+TGLQpJu4H3uBKJVvvauGwRNEp
pN5qxwjv83RctOaxOHbsaPSpf4vdR5b0HDk8eS6VFEWy5IfNMAQeeQw+o6Edo+6lgeeH3L9/tvF9
i4AwBAxSVPrakhJJE5HDCAHs0H5K7DV/+8Z1B0TaT6WEqa8zydTmyzOUGfV5u9BvqCzH0lh9vYYZ
iJJP9TXifIPL/bB2dLGU0f/vUVD8qE+Na4Re7Bo5dYo/hZNYTs8e6a8CN1WCTZJQVpXyaKUvWvBv
uq1/h+Ut/0JZKQKHI4O/+UkWMsiF02fKNpeRS3BSiz2350s/2PTpTJ8kwT+OYywrBkPY1cnLy7fq
GszGWxAQLmBA7iFpl/2Y9MzDdrpBrfWQkzxJrYuHMJa+BQ0FMSNa0U348RRld/5aEmCiaoUeJsY2
iAa0Xfr1/faRPwvxOa+lVxcB/OMFvgxVEWl2+WkFQ1pOGPpcqHe8CwiKxW0msAIrmAoS+MeMxnAF
Mr7ckP+XEMrBGptSo1f1bIBVusgVO7Z8EdZ1cAx4O6BZAqXNVZmQ3KGKwpWwEmClRp691XjKP/30
+iFbf1gRUrOR4lKljKvOpCpRliBujrsGzYToLfRWLhhab7QvVBE2LN6YIAmSo4O1XFc4eiv/73Ss
b7e9Fiu/uil8izmJjXGqodYXuY4RDwMuHwlgx8WK4exsOu1//W2+ZKkqqZu3I1ew3PGlm91Xqwd8
V9HbavB1NGoTCG9KK9cqC1VqAm84zOAt/Nx1Htc7+hOwWvMPPr+z2s9gV2erToAthrxujOs3Wqbr
KbC4W0UXV4UNF/j4fQz4mvem5Zd63+YJzQgxoimFv5e/q82lTOGg78nr5kEipmOgFQagH+8jjkD3
GaGZyoQZxgHE4SqXo/O3lJqUh2BhkfyIDEkgBadwaZxOwYbq45rkDbSsgRWu4Y/a/ZHlGNrob+5W
fkaxUOd2zml0RPcyNyoLpT7/CcTnTeO/OBfh8i73fuNyMoltG2QLg1gcnHYk7itQYcvifVubRQA+
4WH1IYVZeKIFdATk3JeUZqhqW1qx9DMR9BK6SeRlK6h/8VbwjQi8ml/0HPjHVgpSENHmIRqO+mZV
IFmVNqWocQpwaeD/jggsrfC/aEqKiK/jfatG5V7MF+5tRpDkHFbR1cCM8VHaob5Tiuc9I/dmbUoZ
XfdvtqFvudkF73TX7G5W5/b/QAyqtRBJxUq5KXeaS7S2DdHXou2/NfoRqKghOXu+bEQpCl0CwJ2t
6QJMw2PCsJ5OkNUUEeulRfsTvPf+7aFxou9kGZcD9z8C2MVx8sbloxxp/H4n5VkN/o2fRQryB0X2
tKLvwQ8mTd29atJVdwKKw/HNwWdDfXEzrAU/rhjs2LgDTyanAEQeCajLYhrlbCFpVHl7CoKkm/4h
SylFFbw0/NYsh5nejv9bxxcimbR9Xjln+jSBkcAj08q6v3hoUSxe42xnpnU1NxxJIli6Aogjgbh0
m3FNge3dev7IBzdhpBu2QujKIEMCkGhMbLoNWOHdrW1DszBLhlBaSZIPf9SOk7lKL1NqmBCTT4Jq
ukmHv2ytmg4ATf3HlVTZJderQ7cIEr/o4rPVFfYhSyMT8jjj1AcnyHcuE/5Z1oXGETXEpzPR3bJI
TXhXuR7UG/bUhsglV0WbEZg/usi1/YqAFW+lh5DZJ5JQnYt1Sg6z/9Jm9L3XoRKW6IxZiCiOClAX
AVa3wwT9WNXC/vs2a18JBsgSCOh8dLxfxKMwhUrCIEjG+oqtgF/5I/3seR6qDO04lGgAcFEHkcdA
90mBtHzNkRSCx9AKYSPJSa2QfuwkfEs8+PGTwDsUBuoMQeVDs2uw6ewHw6kHOmCOkegiBS79JFBF
H70/vVJg6EhhB+YSMpmQ6vOJehq6X6dVEWnq7jwku+1SR9DTePJRBDBJCgWtZVTM5Q/sRhHxswOg
gUedl9wCIWiuO4bcsNh5Uk9VdAQkjkOEo8v7NHad3RJCRDWErtkgj3zZITO4qrWp0UGQKIcgffIV
Ti2iABBcm3bR4QFwcq+6IXC+dQB9wlEf3JlWn+JaULB0DYnUIumkq1vreEJTlnNCkKdXvMjMRXue
WqITSKUJdmk2Iyfu2/ir3zRPQMxrBbRXTmVFdi6LwAgBUMwh/sP+alnDhffrgHzDAwrLR8QPnZNA
tLbfQ69Ag2797SEsQnwJ4PgCPUqcI++v9wTYTBI7Qwn/RQBq0BjYHy9lxDbkyxd9RBnq282XdNTq
GNg5dKuBaPaPnSM6eBjwf+k+WkIyXNrQgCqSwEr7aqiZrsDo3B690pJ2+uXh4b5e0Vyzn7i8Aphm
S4eIi5K/rl9dquo6Ov60RdIg+KMwirGmrS4GwmSx20P2W5uDlwvy7dVIQt0pOjiPNXrkCiserO6Q
5ljWa3k472bXOIWnxaw5V+8Zk9mKzEdupjs5frqgmI3JMgBGFx3GrRNjI3N1uGaqSIvO1lEUVtIT
h2yiCs/oBL/ukR+wEgD0KqiDRwgxnoWYPVKlPyKP3hXI6VJf8fnmru0liRRCyIni9fQkSObYcUm7
G+owlxhrGr0ndxXbgG0Ox24BAiqjxezw7A8x2jX6qFsDHNMpFgZq6envBfNqRIhy1gFmWJnmbhPR
pYTC2ZNhIkGtr1maUWUvtOcChijKX1B7+ITHMpccNZeak7hqZjUArDJChzJEG9Mwp16ZqZcSvp/W
DHzEnTFjyyyae2zeIH9t9dlp30ZxrarOOk7GHkNHFNqDJ2kI2Q5ANnHyiAW9yGUmLseyufGrBUA9
tgJB+dYFjTelbqNjFV+wkDsFpL4TM12rvTQAEEhWvy8lOS+VZCjEWFx0VmFeGLdoTEXPmUvtNnPt
dYgpgAySc3cwUB0RW9+idb4jniLYW+j8MxwiBpD4ZrchvQTQf54OL1wQnsj9WdleuLMJw7/dd50Q
XcK5rjbfC/+ecbPGaRTUCoJngxWD5jZ9S3HGjIwkJFfOcSc2qEpLAZ1Z9nD1jXlLqTFsBsXPlURW
mLyjgah672o8OMLvxbfodvLTnXWApGRrrMqQchihw4e6oA0pQ+J9mrehrCGYt6BS9on5tDxQzXtT
YMk1Nd/se8t5nrvnHw1eiDeL9nNM5ekj9C+EzvnbzFBiHmvj1Ldw5iezvbIlEIwMA/DVRFQzBmIr
7q7rdEVKC/nm8qo0pDzKj7oFe9F8C7/sHjywuRnJZUV5brv+x1VMwSCvirRFySmlB0CC00aCOHHo
4BCFLJhTJSZWFlr+He9NU20+1GfOwqmY97k/v9+I9BUtlV+Mi2u5R4iK4vo2gL70Bqy7wEQwmgTV
eZykPzkfhpnxWTT66PiWH1HZIp5oRnxi4c73d1uEtDkIkWAAPBLDR+cc1mjLtYqRbYX1aaKhFRwr
mEJBpQ0Fr0vVy0bwhBKEy5vQorxKVkgQbmBV3pla8FaC99hP4j8AQkCCRCQz1yRUystfRHNwL3VO
OmhmXuX0w0bFvT9MAUY69xDQTs+Pdmu5FQXnlY1Z7R/1YkM0YBcOOskGQJSh8oDO0He+MpWRkn11
J2NMFbF2artYQe44yfKK/HGJ4gUy6i7/lpBVwDd8ZTEDtRxWwXQNH9yE6WqGIOZfinj+UwtsbAzd
GHC00aeXfR/zCESD8MFurkIUKTGd/zq+fh5e5fxmqXTjhVZ6SIYUgxKdtm9kZt3stCLeUT0z/mFv
cixWZo1Fpyc0mZwuYkboB5gLd546qQsmr+qzy41DXsKh9tm5B9QbFwPKeXUWfmzxidqUdb8dIyts
WfUXx3rA9ANIgL8V9e9A/z2eBRyIckFVLkfctL4c8kKfG+ohq6QCjCvCu6emzdhzBbH54ncRGZsV
5epEy89yvlXy2nHFIhMiHkSKhXwkeWc7zBHDFhayUZR6VFaGrF26kvCk9eSFEh+H3Ap+BkLaMoJl
dhQyOMKU/OTWyusekQTRrBKFpvARE9gO1oElh6G5UTKF+Gp35BBXi5SFzioOMDipNsotDF0e8fTC
O09HNMMXopt9If3gdjbtJwM2dk4PqOGp0SoHinUboDoyvx0cKaL43efAEe5hSQ3cPZ4HJ5saTcqQ
H3FQWjhWjNzkcMurTTwLIp1GqglMapsHxiwEDYi8HDH/PfEljn/1dUXEtRGJnU8fA4lytYM078Jc
SU2eBjc8ifK0QFYYGv3G+en9eWKCt60+SA0aXZVYk3jaX34InTv166j1YEgn7QpM3ta0FTaSGQmu
1XgKvAJ9xQVm+S85gipZWaAtUAMa7it5VJLDrHBnQLnKxCQ4AnIZsA2o6S7CNncMPjodO8OYhpOg
Z0qcLVIvrEoUMyAg0fuuR8m3dfBk/OYhxkSd5HB8JSuPpCQMG//Uf3pAZARTWWP4hsXXx5RTx8NL
sigfSzJUr/AJNQq9LU2+8CaLvGhPCA2+psMVruWT3fR8scUMtBut5HP/MzuYwWdluEExRHOWKkii
rMPTsCNoStHiqEs8v9C01m28i4S++JsNntM+ow2cX8HXJKQ+YEnspKwz3Aj3ZdNQe6Eh6xmUDCMK
o6OvwYmsQuDnQG/7ebFQr5sIftr7gsdhQDvG5LHg0rieKCOWNbnu6eBfsRzvgIIv4+lePxXTJLtp
mbdWUKpp0iqaMgwlpasjP90EHZueHzzbphMqBH727c1F0n3/X3Nd7gd13bWncSUqMYdFk1rC1q7z
PNAmgjr9Byw+UkWk4d3XHVSC9fhrgXcoEznD2nb7ZCmz9dBELudJjxG/O9sQpJ21dx4gSPO+eUp5
UUxYd1o3vM5jcuKGxSYtG7IO+Kbsi+Q5JrEsX1WPJm/cze/yLGVMg9cGjNGsNEsf15MiLA4FPt1v
bCMW0lfFRvhvn/L3cG9TCvHubhCtEfb6g2YMnGNtBBw3dvxUx7c6+ryQVLQ7xllb+W217d/7pHeS
hf9lpkF4nUSF888X7KsOHjjqHBYc8OXgQWvVMWyjGGHEbLPkK2Zhns2bpsiGTqvr1vn5D+9YpuAN
Fj4JEGNLcLsZv7nnKNSUZU3JwaQNryTvgXwigTd/vsQaf608Bv7z+64YFV7R1m9Diy5HsqK2NAHj
mX3xisi/gB5mMBwPCoLq351BHqK6Z2VM/qyVu8HexmAIemcO1JTtcaa+MhZwqlbImIR5y+cS+7Us
4sg3Krp3yoderN6gIbwGFiH0McVaH5LHpLEIdkKgqhTryHxewN211cEBpVktGhKLKybJkCnl+SnY
oyCJsdrBk0gtJlQoMIpELQROgTNUQfc66fQ4/NawkGKKUs5HauVtCw5Bt68zEGGejIhqIl36vF5X
hWG6yfXMDoi3TWR73emKwIP/qr3EgyM+YFgv+WjpS/ryKhqOHGpFO2czWy8iLUxhY9D7Z/D4gMkA
fIfY7eBDsoeiwAKNy1G3LWkuli6vLd4d3JgJp4m+Ezu+vwNAL9SWF7xqCvvEsCnJW9HscdY/Xrj8
w0LcNhU0yYZqbKFZjeVuBhKgj2Eqgqqi/KxPM3Hlev5jPZ8B98iWivmKlKmh7+9OY6IgK0A6buF5
jTKo0sHuBbb+2Y76SGoxNVMNhV6hkdFwENM5lrVNwx2ZIFDdRupnRYKBuSZSEQXtlgNvks+S2fHM
uXmCE5p9uEDgSoYS0nBJn+viY0hT+66gHT4/gNdd4trVOFlF4yGxnL9d8GDJXgNqURcTzSF7xtEg
K2URkCQMt7IxXdrUECxt2E3nKBfpUnu45qH+8stde4wi32oAzq20KXWy4kMSYVKM4cxJrNp9spLU
zmxu9ibfiaLOj8I/csovI8Wn9CQgUdihjrmtC43z7AM59V84VLopKezwvkjttO0Cj4mhCtKO4VbB
QdhWZJKS8fbFztXg8Uk7c9r9Mgcu2PD9OItGLBrozWmFVzjrquMd9xoyyNwsdIg1hJP96UD3zFPM
4ncCsO54v3SkV+gow2DQoxXVKhXsREje729hyDthnax9dF44ydvbNR9logAEspYC92L5p8gT8ZEF
Y/FgLZNgJnWFeXO8mIlR/xAcWyHLGnwSURJTxl7TzwGvqQUZmmnq2MOOH9oqiGrrO2tEa/apy+18
C7fRQJdK/gkg6FORSC4k1vqad3JDI+hozEPRjqKQnwHUWO/vhoCbf7OGejeRAtmgL6+foKiACBIv
L1gYm7/ECdWZBmFrytxIY9G2PpL1r3dq0yVTg2ckM/5IV4ILuH0UpH07VF5gE0FbZcpY9WF9cNe+
/EnhZhftEE4MFgyr0VtcfOCcVqptzg++fGy2Tr8ZjJIi89F8sH8QFib+rTjP9lBFDD/yaeLI729h
E0Hff3g8bfTp1nD0b2sOU/Z+CvqAew8F1rN7wCanJ52kd639//cYAUs/LZP9RXEFlExqjHmb9kXE
VuwmpxIZzg8no6AF9KTwz7Lp1hLv7nLqvTI3sL6IHA6Qg7aCTy04p9nXj12r34i+cReVcP7VwBjV
02nj5ym6Ou1NJMiILZESniunuoioPTF7FCBw1AaRsT02ah3yD+rKrWxBMY/vWeW/h9eodc+P490i
a5FirNzBSn5fQtobjIxLgEKdzidKPdkKlTb4citw3hQNI++q5ilhf0tBNZtOEaXrr16/Cz/wLzYa
AN7LEwqc5LeK5kpl1dKLA6hoOANaowskf1ki4DOV0xvuPbVFXyQs89uROrAXrO1e9jdhrHWpY5oA
5cuWyJkNRk1bn1aQvHS4IB9lMBhA12Y8sq5NQ6cN+k2w6w2sKDFaHzFhfmSLZggRgb34zEIcqA9E
U2M5Az9hJonOUiODicpI5Ct+SdvcG26Zf6QtArGqSAL8pPJ4cKNX1FI1PcjZhYwacOUb3yoHBISA
5puZPdl2HynpjCqcymJszj9qGeMf1PP0Mf/fHjck8TWLM5KJaeQG2Z4mf8udnwyNVRfNtd4rn6So
a1GclKQZa3Uwq8aPui000THXhvPe8B00CfDq4XKqSw7FpG8bySrPAdoqcxq19irWLtp05e+W93lc
nrfYAdeC34aiJcGKzM8GWjnBd5niOSex3jeihmuJmMTmL+lcNvOW7x8lS6z17HoNsrMQhXDE2v7l
gRExwbpkklWkJk1fi7Na5KDPtvs5IGpPyoOxidgBaYu8UrtTtWN9D+w+WNi3IJvuLHAwhmBmX7wk
EKbwkWGi9UUzTnFAwt35aoKlUwaMq360+TPnPERAbov6strEEQ0P8sqP3ItGXED0NB9LrsACXAUl
C7nYyEQb6T5O/ZHllLjVGzmAdrVAMHfQdQ/i9L0ecaL+yezMHScf8caRGHk1cf8YnKHUh/j4k8fb
lBE3FcleUS+OqsBRHQspRUSunSnEMwYECHb7OTZk30l3bxMTe7KvLp8vf6elNdD7zFlashZLUVH9
UN1AANOXKWEqOur/cRgVQuNIFKlLNUxXmYvnmqQedP++jc3KZWInrG2a3C2EdxiFQxZHWHrxF6rT
VZhzk8Vbps0Xn0a9MKG5MZLLMMcvrgpu1w/h3ni3aDb+zyY/FGzqZCiBjZbliRdTAK4G8Fi/ATsH
MabrCs5YgQ4eVbFOBBoz4O6RzwEMlTVng3rGPxXkmX8VC4b0aDrQ2af0IzD0IA2y0iwP8TP0UA5+
gIF304lBSzZn3E5674Btw3zJG3HA3oWcQFDuUmtX6Px8sRIhyqvpAfMCXm6kV/wU0tHGY0e2c5FS
2gOoRQ5SG7UitUwIZ1EwjOM+hjzy+bfYcyZhVSQ4d56kRoOsukWA6xoWdD3WQ5NrEkGojC04QEp0
NRQ9vlJ+M3EXHtivKlwWlQYQyKrerfG0CRCYOo0Wyjsl6pyoZJbNpreLXZllJpoPhRx4cltpXQu7
S9hXivTNbuH6tzEeQDqBSjD0zeOuud3K0tTHNy68Z0WJB7qNwK1BFA4D7rgbN5Qp/PtXkGVaDrvL
mU9SK4B+o1M7ffiHkw3AJVwrzGBdT5z9KhMJXYvB6e3ucvLP5t0qOOSRR03553N0SeaBLZFVZrrP
boBmcfWO1/zU0Y0EWjAjge9gdZcUgokcqPFoXA6BjPHsDe/WgV7mppnIYIY/hUOLVXXV7iBA1jcb
gDTiItqN1+SnH/U7iROtoblTJR3VSDThE+hNqS3rmOaxWP80AkVT/ju7JC4lc5NfeYFi2aCeviFA
dBxIftW+HX6sQMeg+9SSsUL2NyFXY6/2eDQ6Mv27HwI3GXjFmgt2SOz5Z2Av3sfu0qDmtlzJlvkK
/MBtbYZBUDuqvguGg2itmr19DrRNWp0Gxq5wCDsR9LMmLAwaO00eZx18f/n8kzYwnFWscEwEUL50
2qCHjczajRBxUhYp9cH7Xmgv8m/Vkc3XzIixRcDfwW/APIW5LoeoCa2gMgG/uCEFJLnbzbyIdsSg
60x/W6Aj7C2KojbzGr4co9mTN1lKpqQgmrq1w/vGZdKUFTU8ji8mlGRBj3Dw0hDp6pBXxrhHTztY
Uyd54OxOK8g+G6WIf6GygI9+OiqCqTmBMBuAL1/wsaim7no98fr7vh2g77cDB1wGr/Q/g++CQZz6
XjfuQcGPU1cJ5kWBeNM2sHhBThlESgTw7AumRJ39hsGQcesPNY/IZ2SWSIrUCDsvVLYCRAkPpEV1
hvIV+85QfPPKcFELgpqDTb3f98twHsJb5cAiaDpeY/rPkD6+kNtnl+6NEoMuiBN+vEFRaAAQXLbB
srPwwy08qr3SzUd20nauuwXBwL3XSo8oGUovXm6vswmilFvgJQrG+PM+AfAoym1bFSecgSFHFTuJ
i3IpwhfSE8O8E+5/cYjHUeqx3lpswvHgJAK7ZvTB63IeU8O6V9EQE5oeJk87w3WCGHb/OFkbhHI/
F7bZ+cfKir7nFtPKlPP3GRJv/fMI6MOgNasT/YWpimQ0rAqL9rwCIWPv4i4XhFyx9GorG4RfoUyO
CHT6fRKiLguF9YARG3uzwtqHRdDbfn4aWnd+13pGggZ7X81oxY9GRQeZcKGai7xgT3thb65Akjpx
2BG8xVyeo9V1gYLhHFtB1ZQ9srNzl3S/ljLAXccffQQUd3/ZkEUqCxeuXl4CEKdOcOUofIil/TF/
AeD+MYPdYvixDtYjoKE2VAUZTn2uNh2hTL5ZdeyHrRTUok740h4953nQywS1adUWQlhIyA5N/dgF
uN8zfcIDS8ew+l9Vzmb2S+lkY4EdaGbJr962vmH2HlHsFOpYpMI/9ghlfi4LpUXU99obAsuT7/ed
SHk3e2wpPFzJ2arlJ0BUspIniBTAk3zPhGkIKwkAn7iWNAIaXauw0EKTkVE1tQEPdkHm1RwE6oqJ
+YoqdcAdb1deoG+rt0dm5qCjAKpOx/Q3exOcfKcJYvydYGpv3qfWZJ3pi0epoqXa0sdWN/6GniLp
NrT9yrfKlnC4Bc0hYbfNTtMEzyOoO0o7/KnfjsLRu+VjbJEtZStG3pX/M6NV5UhfYzy65BkVPR8b
/09kvr+u0h3/W/EwZGAj6WkPLDdHwSHjJ+X4rQosQvPXZQkYlQnBnxm1ZUwQzUsF5mCZ++iUoc43
MfaTAtdmJeN9ajhgOe1dq64SBs5UrRu+N0JsfYd1L2TZQ1TaQ8E3FErht4Pgr6IFVP5v0tV8P4ey
dqNg3XLQrxzBbPlifvexhU8CYmU+9Js4XiGU5D0K3wYCuRsu7e07c3iJyhIdxh4O85cbSZBZ9fqn
W1bv6XnfmRIcJbCqaFrgZIQ5EeXCBWw2izXBu4l32pBCZ7S0doBIIEVD2RbciO3mFaa2/KLrr7P9
Cd0tCCf/X7a2ELESUfpZJITwauamFEkZG93KaYS9iFe1NxhKLBr/v6Bd9jRZsbpQAI3rQBu99GL2
f22GsPJYhZVa7v2KHzuBVB0GHHiczfWsZuI8XqVuGKYd6Ssj5Qfk/Rprv45E/35S8fd0/S/GWk0+
JTM184f8VyWlClTKRNoqUZ8YHseAciTLj+rJhi9EMHfEiMN+aDSYrFQOcYkI7a0jzpThNZ2fYUGk
jT6n3ZupoIW3gvzhCxUgWbV6dHZs4fzTZFGocWf3sddWXpEN2PLnbXQFIhr/OeuNPi9Yc9MDMhNF
ftRdD1RhinoePY1t0LghEnLoAzwVaZZjx+3EksDL7TbA8IirFaoeqaC13VL9NAz5JUVkbkBhX3SD
CWKYJGbSKue7FmO2O8kmYiVgYixwc+Gmu2eFcD0gYE5t6KvYQT9TIBbbLWEjp5Baia5QaLhK8aui
/OinCERE3wbo/Rx8gTSvSPWIS5HB5PlMrHAQyFGI37CIbK2gfJbIByrW0tO0ty3T6SxcRVtngMPs
ehP824uvXAiX2b6FOZ3WgXLJ+ckgBiT9ZEzCU6XfT+spnQOXUxw4LoqX5Pjvn1J2Ei1I/T2hoorG
CNRhpTdx4usnMRqcPnZH0ukmE5gkwaExGuAhP0zBwImHJY0k24F7xU7FTWMqOp1O8YrRV9H+6LRX
jaHIe0J3A184yCsZLcuPCx1NdU6JGFfSw2Xqqv0G6fmEYy28NjNNMK/1t+5NfuxIXnbmuWz6MonQ
89k2FU2I2hb8exNv3B7bNz6NE7X4LuS5rz4LvpS5MgFAZwQLMjxQZsJO2MXfsAbp8TiU2VazoogV
AnQ7kJhD4d0UlbZcJ5ehLH+ToRwvw6RXOdV6xOcs+ISVrSKXxz2U60vpbhZo7DasJfjaEPzLURyG
971fkQ9UqiKP/MmWaVpf6vtRAU8CRGYRdn9Cza8gSfPyAptFYelhk3DEOKwYa5OF5okSnDffhzwB
3M6GUNXUzlR1HbZhhUNtRUmVIzwGICNCwtemmS85IJqhcYXglDB7kh2ESUyfjEwXBaOs4if+NEcU
dQ5zEz2K+8DBnE6n2DOGbF6he95Tu8u3RYKlq6JnGsdb2ch2dS2PB5ZrukxnJaU/Aj/zrSjykc+N
TcXWwNzM0XTrjw+oEkkfMK9nPkcG4GQUftFZnczuVt58FnFXyf9MStJF7lZIyGrBia0p0morwKoQ
28SFyToM1nEwgOPdDe36AUYTY9QsSczZtzO8R9M2WGuYNC0uoyWlya7x+J2CCi7DMEVfyjOfmgcl
FtwTl0oVacrmR2mWUbg99PHoX5Y5reYzg8Jj8QHowd8Y2nXKlk2tGkdRBs9npEVsj0gF6A4jzq1U
lvkIm+mrmeItFAk5PBX5UYse5zkgC1jOc/JMEQPSzNbqc8/ykp+zJNOZmINWQairrKBdqFI5sdC5
bGIUvFebK/q/k+oAUWip82netKrXkVmGc31jGG99Ui4OHf939cQb3pcpLF0tI/hYGNnh1Jsfib9T
01P9KcWu2wZh5x2XjEMKh2ngScnvDKQ11jCxENWPFslDW1eZb+6k3PFTBE3IUmqEtJvvQHPyf9WN
8UphrBX8jdvKpx64xnGQPoT80I37dbOn/fHg5BT792xjjUsWQH79aIFEA8swgWgoMpMNvizllrfO
ZQ83+3JxZZ5Y2rBUnpCoXZzxtib/PA05+H0hD2A+vfDvtd/5+dZsX0IRVaftwMJqNWrDbQ72rjAF
7+P45WK4RQE6vSTdF9y8bPizveLtFrC8v/CEHyKW6Bw//E/HvL7rHsBVuWyljw2IZpCAM/wuzHhQ
H3LLecz70WSgQue3ePUeRKYzHrUUeEPVDqCMsLL0R4215E/sNnzyaIcUkLA6hK8ecmr5Faa/OpSa
5fayvpgQGUjB/J1pclci7b2xKr1WiLgcJ/sxPgUvCgiHMWyQ9e50M05l6+Wk5PbPMcay3kRRWwQb
Pz4i1OeytzvKlPYbETlvtcv3Utc81sJ53IYd2YtIZJnbqh4qvxDI7AtvOVF3mdo7lKFCysHNwCvm
6IT+7T6t4pKKp+y4JaZUJewnRS3wko9NMuF6G/OfkKfQk4LXr/gihE1ugR1VkBK/x3qrkuNEv4BO
85VbKqXka7Ta2gf+O1VyXV+Z1/3kY8OYzwtSNifCTP9Xbc7f8/oloxpt3Et9yA2Z5D6b/ROJ9ndb
ch5X1R+/fzRbLT07y+VEPiY89trv2Jp3PQYNeSrU6eiA8pl3KpvrMcek/epqRVkc9An6PXD1SpsH
1p97gpFe4Dgm0ZGjnayDXZSMVOAec4bmjffcUMRxJdbQ+ZQ7CrhPL9nKbp1KrR3O1jHj6zN8hrOR
E/1FHiXVY84s8LgMKNzrmfOFQQCyiiu1tAsbXWzdn5eLHGEGBxdEhD+Ogcs+lOJejLUxZNvPkSFx
BIKYeLPJcdd3ZbZFuFxxQrimEk21FvkQ+VCVLmbRiL4P1s4ZXpDoSHMIF/jzs+x90DX7+vzGVYa/
LuxSiPCh0zkWi7zAWw62+HoeeQVgcuwl4aGvKrbwBbuwzbNzYsfFIMaNKkfeN/46zA6kjraXtl1C
6aS9OfaAqcXIY7j32y5KlWuO5Eyi/sPg7oiA7sqfMJ/8zG48gKBUEKSuFyDWbLzKGwHdvwrlYYJC
JvO6mtQWZjbKZuNts3OINdYObNCM7hm4b9jL2PL/I3hJqF2SGqZy8sWds8xUjft+jE39EFV7+P8o
i3lVxKc2Nj/WX0wNd/+IZi8/zKBJsFWRgLPeEEZps/Gnb7BED0mjUPIZ4X5QSBuwxigYmD4+vEwV
zVkG+XkBuKRX735zteJ9Ny+p40gMiHwhX8+y1aYiCbXmY23DcyMGEnDxlC8er3fDyLkc0A92JOFx
B+aWjTiYFZQwcAREYQPwbMgdxl2HFZZIPhA5j0Ar1sc1yzKeq7j7W97V/UD6VFKOcNriJhR8Bbo1
Ra0I2WdPZvP+uVUU4K8Zmte/xoZtBX95oaDtdvd0URmxiHQzY2D5sv3ChnkyT/ITBnGrHhjEBhAS
QlRLP/xj75sOdC0gBR1KU2xzLO1msYZHvd/kW2fvvQI5AYtLKDAQW1QnpKxIagaToRWIL+w/8xqi
mc8tf235o24HzZn4O+gQrWc6iCzP4dYw4vQKT0cEMlhgdOqdZU/55mmPGB3oAAxmmILHcE29XjTt
YmyMCimfXg/cOtO49AZJBSmYcxvpMzChKNMIvsA8ZgcatVPlzTpejZKyXjWXR4wgUipJfar1tKB2
wJ/r0fC4VBSpCwOxz3/kf8TcotQePrnRI6FdgC8H73NYHHsGlt8fykqnQnUPRklMJAIncy/b896W
L03ENpyEqfwDwua7Kwc7AEuYD1W5eFLXXdn5GZW3woQYowy/GnW7fJw5JFtw/ghYHe42QGRq2xv3
iwthROmK6j1sD9q4yeAqGE6Mce9ll4GfM+joJge9Hdb/il5GGH5rryZjkNNW1NVnyPvA6xNXso4t
Gsm0KOoC91fwJgQaL+wGNQnRxwRuzoOeG/4e4cpP5ZdRBguIZHAILtilNM9wXOmOO+7mGYcKtrI+
BHIHYwVC9VgOgT0xsKTHKUaVyJDh7J1p/D0xdDY0RZzw/2F9LuWcysHv8eckjFtZIT/64imPEuH+
m/aUwf8ow0cs+pUbMhab0438yZC1Z8ZC2057mRU+0x9mE9UVdU6dzNsumrwbA8P6FCV/Six4jYRI
HYuzuvK7ZWWrsVjTgIJDCK9Z0ScyXbfUlfdAnBGDqaD1hRetGQrv1Lq6Qjz/6YG9FUuCi8nJsr11
HBQjTGw04/kIoz3ZAx7ylGJOUtoxjJyTl84SBrr73j6CoY1RxfKQSvhEH2JO3r7zEHAuimWkDfNj
GfUVrNrct05ghmIhcQlnFNI3BaeoMr8j6L2RSWIN33jwPMR1FK3m8vgySUSlHbra0fHCGtBhS4oI
fmcn7NlAL6+v0wzry+lHf/Ws+tFg85k5JdIknQL7R1wc8f58JK4VlM0gWIIckAKeaNVIEBhO1tFL
LW+PgGy3WDyn5orrQU1SCkfIBI+/GJC+5qOmA62r0ZwvFEdxy7aXGp890VQhJ2MW8DKUPSpT4vX+
XWxdY6bDLL74mJVAmX4CQp6WPmYozngp5Hmy1YQLEKx11KcXsvHz8UeHuFxkqBhJhi3OlS2BCd5b
JqQJ/1Ep27o0jD46XRB1j6Ibkzg4DBMYOZKLIuSaMMhn1QaYqzucBcy/q8NqwaIKsK+aJISnK4Rv
EkQYKjtxkZm0552wblC6kanVTd5RM7RiNkQ9RYp5qXtxNUrjPW8XK5i08E7vZrskSugPK3oAkeax
W4roTcg0IwC9SRUIj4uGxgDVMJbeinVlnM27unKpqGwOFn807Zx6ZdCtQrVk2CsQ9DZGJFvtVosO
3RzZg3vhgA/sl9iNGn1L//hW7RMxtiBgIon5/+szNn+FXaGClfIwTnOZr7y+dwVKsgYV2bQxSS+m
ODKPi2tUp40t31sjc9uL+WudkcPA5drrlAAD0mYg95e3YEDArEzMg/Fr4I4xlzQShIggV9+Eq9NA
k7Dxmcd4tGUatNrmXFrtgiQhKuRiqABrB5EV9gLAnxqorxBx8PF7D4tfh2N7FCWa4vefbrUSnjjy
aoMomm9qgE+pz1iHDjrlq7LGR3LiMQXJ8UG3Pubaiz3+Sq0EZsrE5FCs2XiyHoOAwI/ZXtYKgGdM
EuuRnC0CLzaM+PrYDb+akCZNHG1v/B4w4hJjXgk6GHsf6Jq1IbxJWDh1OxYf3TrMq96P8+jsnY4H
tP8IQvBRejXvw6tvdWH0j9NsuRfzvgQKSp6L+IIOEkVLApB/5TM2UFToFwTItbX/vYOnrECmkVge
z1JLhLZB2auWIUPbvzCDR/NHfHhASw29j7ThkmDz5hdBKxXoD/iARJ/csYRXOjp40e9kOOP4rZda
kpTBHREcD3fQko0KCE1L/0vW2WS5WxxVGHWeL4LsxuxT3J3ykPhZk7VnnMV2m+n6gOTBzofnv6t8
SJs+09nRzvHb6ccRwI6vzkAfveylOEdih56ReQmGrA+URcRri0Y8JgQFgO3DTrWB9ykjc0xDvNZn
lr0yNEiTaO+xFNwvRadxmhsw2TvmHYFY4pTzwu1nRjCdWyTIpNlCJXQyDEp+5k48/JH3Z++AD5Vv
ZMrOuTwwWMiG+nE6gvAPMWsZiln1s9K0coEHmo+v6DC+kOC6JAyYuDShUkxNzjV/ePul9B67KsGx
DKFdL7i3pGdKfH9GJa2+CEsG5mGlXsMUeZ4S14yFydfhDYGgCSS0t9kP2AsCSExd5ZBiC7HQfsWy
5QQpYjSGwFChZ5aWAVxs40kzMMG+eLc1Vdo8RXW87AIQs1nTTRKVr0Wj/zBqNeUV+uVAkQ0MmsSH
K9eFUJN59kWrUwk6w8vGKgNcwPc3eGysBNhCTRuWeAe21GSADQiLT1SKoVnup26oRGeWwJZOnRFF
P+GJmX4JYH+h0AnVkia5gxsgG6Oj6anjKbhRLaYFz138lYcZo9NwLohaPGaPqF4rtqZGOcS5N7wK
Smqyr1KW4Rtuln9j14oXDR9oO62NW1ps2hErRUlN5Xfpgc2xM9AWepYXN7goDrlLsroRywB7jOGW
jU0syluD+EVg5B24rTTwQzDO7RKnRafi2JWDp9kbmKI/VEsfLujOEnRaUEffY8wZL93Iq3Cio+2R
vxPxSwG8OwnpdSpbiJZeTzTr3juwy11+sRb6In1VoOXbhwB0z2a48YfWSDtfxW/lr5yTTTadAY4W
2WmEsFJk/It9emEgGmlmJCoKL1CtMqzLKcO1CmVBzNZScrRGk7nT/ChCYiblThc22gseS4j4+CHm
nyOw5PGYG77zmh5lgc/Zwvssq+PQj7V3pnLK72ba5FPiCOG9zpWmUdAwxmmUZI+RLXzo5rWNdCt+
SL16k45PbK0zNmRCOhVZ34MQyOVrGC9VqUZAWMzh8SRdB9ie7Zf4T/7AizafuqwJC7Jtj6JJm1mA
SJt9cGz6IErkEDiKmZNzdiQhLyMziycSW4C2BECHLw9RDYqO74eJF0KkO3ZC8wVSAhRZsjW8kgoY
1iFa2XIakFDNULTBhXcsdI21t5AN3QyOe3jOSEVnI55Qt42t7rQvHI9j9zyGGkuJ4m6Ei7P2IbsQ
MNXLFrraPWt3Zl/HbxB7Vb8fiD7fyfqLftRBoTaPP7/XiJIGXYiRwChqyQ5VE1irLlLjcFpA44qm
H0PTwTSlsRe51DLuprkqY7v6hmU0N79GW6NvObah3XENsKrX0hdlZll9bG2ZohS3pC9spCsgDHMl
/10W8jnNH71VY+z8fdGpwVJOKjZsVOFxIYBPzrNDTcnjebYF1BOec7wYUtKFqXYJeLhPdWEMzFuG
J9DMXl1ZQ9wpv9y2EyRLBTMo5o/RRdgmlsJcIYXRa5TqeMd3Zu1G8Xa0UpymrlnlIEm91/clxEkJ
Nx9oy4gAe0Ul1l+TdeuPYbzLlUVxqHj2ZmcN1+GGhE/uxdB/WRSsHttzKWtLtzGPVZws6dAEnNvc
sV9rsrNJ/KO3A7g58fV0PFdgLHIlllQB1jTS8uzPOkapd2EldThW8z+YOrR1ZbP1uuSHX6iJ1Yq5
kKWz4hxCoLH510HphT1uU7QZmSBKQ4mvVlgeWOS04AyH+Z0zngXMAismdwmMNTPh6huZS9nPKuin
IAimBRO645ApEvKiXTu21TxOAIq7ksdwJiKfclqtxbg1cfsRTXZAhqwJtBwiG1wf6PU07x8jF7dN
Qbg+KLM6FnkEe/68KkA4jFHp50exTUhMt/+5NnntGGo5dlCnY0+LRAEoNlZQYfvBqyh75ZqKA7bC
XUsIsna76fqeiJON1ntyLlL6ULNd+67pqLITJu1Jw8DMQRG0+p/0l1+l5L8VvgBRNvbo/0pDpzfW
bFNpMabjLRygXqBlL++ADmQR/MTIRXXLAVpeIPkQOrqKArrjwOlDGcuHpwKM4f6sO+TdGG3vOsSY
b/n/yecUOWv8IVBhbYsUGIDdxfL15Pq1TDx0njhViXXC7quGE/QGzHd2uIYh5s3mVjVKQ+pr1Zg4
Zolb1aSGDeyuMcVtIE80KkhYf95ux33B82uNxsVLvn4gHGVGh25KcE1kjJQKC+WE8bGa6H8/Mw3k
hRL9XDQ/FAqJ1N17yzg8TqUnZ8BNOIW7XLNEPlcw790/o877RrJMNLvvRY/Q1W3lo7BBcZwoyekf
d3ecv2HEGziMQDlaf3bG3AE0I7EDeVMyV8vmK0ijVySwP9M9RTyb7H3G1X9sIE/lAi0qkKW0ugqm
y2izCkZkDck9yzG7fEVe1useydrJgie6jL/89Nv0Y4HH34cvF9hGYIYyWsM+lV/x3nPgRaenY858
MSM5OEZd1qFLoeP0GtsUfanWl2uGNw2VAO/8p+rQ3Gge7Y7eQcbCRGg6uxiV5FrNIm+vEDZlaTpM
afCqTXgVYGU0kKtcqZTYo/w3AT3w63AVukjC1G+k4SJ9C/ucYcYyl+yqsB98ODTnWiwrGiBeB2O7
G6lns8UEw17LIVD775hD1pZaf8dS/ZAoB7teCpalF2QDwW1750Qj7nB6uRkZcLACPQNRk2wrX98Y
fuIIrAyy9u6yTmiNMfFW+spBs1zKOpqJlS4KJeVWH992zcQkpFIBj7FU07ygXxgC2eKEKdisNO0u
f9/cxpglW/o1hxWVo1l/Otty1lX02p8U0c6JcRqP914LHX/bU+EgHTRAJyAbCK+vXtOqhqIy4x8z
/XuJjgI+daE95GtEJByG3c8R2JtohHDPHtZmKuHdjKEcHOOAsM6psTWkdwsFq6GYpGwfpKdTBH7o
xqTf1gMC4q126Ft1KdizesJYysmh0GDu9VQQFWfsV49odBJiNP7AziPEmqwJe+zlLqdZDpApl028
Bih92ZabksWZGD+Qb7uzgQ+dYRt9zDcxeciQbqpn7b8MwErbs21G5FkqoM9u/kJhSU4UziOsARHk
NfQqI4zhSgUHuoc5x44GuMpm3Vgaes931p6wKP4+8aHmRfrSht4vrRXW+KjUXL14UvoOgzWlm/Zw
U/Mgg8h5Xl2GKfkyVZlghj0w2rUEBBWT3zrmji5ssGmYRFB9iDC8ICb509497AptRH8O2831uJnh
cj+CZG4esen7PXAyekC3Ac/UB1d+PZc2OO3SXp4zAAXtrsLgX2NWHS+cE172cD6y3wREYuECXWnN
pARH3pnEIeuMdaAY9x0oPHDRaHc8W1ECavZ17oLCKSSzeMP3cbRdxN3xU9p44SF1humUtx9Y90mJ
pxN2YP8tryVExbypdGbNRl+qEYolf3bMZdkSvMun1jTLgddLS0/2JzDxjcRqoLIw3B93m7U5RxTX
rTOZNoGLIORXNN/Zr5Aiu9laVa9fKyvdHp5IPHIAgnKcwnkn5BzLnJRUqzDdnqmdMd4KCQKWmmq2
bl1jjvDrIqzEo44zubIgQgcXZa8r8h/klgtlW+v2GiJ8apbPRRSbtUvWzvk55aCH3SgKTcehaDAa
NQYwPqd6C4vXKviOus1u12Nb8SEdYHzWVDNsRAX5uRGCRh7eAm9JylKN3OcdwfMr8LpMQkP3F3am
9jPhfTtZTIjgS/Cd8JGCfh6hMQSymE1+LSf8rKdiPnayxqEt7qAlwGWP+HbJdJKxCOrdBnqm6UR4
VaRGh+QXc9nAkVDAdeuJTTVL6sNlViBqyurrYskuf6ieSVYqRINf4vQCRxNIX8uwS7gmYblMsSbG
hhgZGyYQiMUxnV+bbKVrGPAVEhX44Ge6tEaz34EEXdQRqFGjmqIFsJJJWa+c+fOt16+SU5Z5dN8x
V1JavFGJ/hd8fzdCN7MWb7Xca/G6JQjW53opgFNjGfTqKxyHTA5foQ8bfrQhTI8lP76N/QDeV2FB
tda1Z58uJaTzt9UoyveTV3B578ApGEjCmmioItkvkAZfzAgiFBNpkPMShvv+tEc5iXWOusF5UUlF
oSASQhbr8r+1F5UTJ5tmdeYVXEz5F1lkdq7g8pwTmRZFPuLv6wv0qlxlM/V7oy1knVVc4QZibxTr
YyYSTBEarlrGhxD3nn5RtY76EdpwFu0iYfdhWfEY3i+XTGueKBKMyROQOEjHLRw0N21iwYoN9Dg1
Qn1b9x2dvlmcH3FYOeidJ5KxgIo+e4TLQGp2pei7fNMKQoWXuUWGo27Gr/6ZYop+uIXyCNBeypgv
fHxqjaWym7vsydAMea2ZNY8SUMk4tTLDrvino6P5ycLHTDFmLE6nFxcrVzpq+eb4pcAsz88heOom
BddM9OQZg+jRrvB7t8X5sUjEHxVrGAxDkSYwwh5YLuzt09vP0q1cBXGZK8sJC/kgKpwTh4LpKBdV
72qi0+ZzIKrILhAXc9DBRhRlK5i72tY8cTMIoYu9VYuJ1E7kYXKnISXjNM/roy151eaEItBAxYww
nCbN+VUUcjt/93VqDbSuhAdLujYsGc6tiqiWED3d4GOwYPpyobLBqDlwh6FqFRLiWgDH43Oo6Whb
2Nnwp1y+LjOaPZ5nUgBNXB740zEfxSngIYfmTF4+yuICpCKwSuBa0W2CUTEON4xiAqlcGdSvExcK
LysvcF2gq71TW0i+vR+Q5R0aTU3m9JVTwLfgoyh7OxEaCjDfRDZ0BOrR7oamKEA27ubnPq44hg4s
bHv1fPiGAQcfH10sN9CVXPM1UTR32RlsECIfXd5VKYa+9DADU5QulT/k2sj4UyMOivgD//YWXLOl
gR1cB1Q7B0Uk5hPBwzpnMOiM/JpabW6fcJVQV+QZ9ST0Ra3Eq1sfwogE+nxoouAx4e2aX/yX0ews
og/6zsMCKT9iyTNop9gBeXBngU4LfiLPxhVzX8o5ZAVy/OIN4p8vp0e8aU5b82XP2MYsE0O2xbOb
7+guatjES9MSs3VrvsAplfrGhgs8PToVI3gy7fH6OlaAV1t3Pail9EEv39DJwhbXOpqqJFOZGnrV
DFxVmZPJvd95EoQCKfUc1fuw4CUBEhwtxr93Zy+W8z4zu+AHM5tAFFywEgWKnAl5fGwK+Pccum9i
NkS0IBdLDNsC/8S6DEdeZYpLt7QvknYdcXLyZUaBcprVrxUYxZ8Tg67AU0Xf3Dc7GjRqPgV70uxK
WPaUjavOg7CSozpgFQhhCLNf9shJwtsJGWf+qo/0cddekMmHuc5cq9pMjO1/RvSuaEiuONgf7Vvb
LpCqFGKmFOa8NPCReBlIaMDICs9qXE4ej1nsAgCzg0JiIgsM2a31aM0JaUZ6CmgKexIugbP+GOYz
EfT9dG6IwRCFoMgMScSvSX19/PbGg+KEuVZBHxpxI0tfP9kMJ87mySDYiVP/H6YT970xARfKGW0s
w+eUZhhpA4wXPJ2HeKvvxMYqYYyEKlCls0yLmc/5XCW2dmb8Y190u0zSeien7POPb49G6s65QzQM
mx9tG6eFhv+12YD7JRKbH7rLwjvwNLxEKSC5rwnY0SOeeEgywDfM+rXx28pNl/SMk6mx6MLSiHfW
ZDPvvfPIZRuTXuNEjeeqrlaCO6dadDYrDl1ixgfbfBKFv6GPU3/3ofFu+PWeUJxNU0iIYMRJN+QU
+5t/3bpl8CVsUInJEgj6/vuThjI+zsueACQkBkvFWzn9QSjTzJ+VAXt5HRfzPxwlBOUynfjnAf7P
TvYniCjyxWvDuXEgAreA4vuegcicSTDWfwRDqevSCBXdNeCTuEDWt2KYOQhdt9VTgN5dlgs8wg7C
+pI2BqiMj1Mxt2uVx+ctMf1bbnLymNs9oOWJxBER67mYe4Zf/ri0v/aflblxXPitSaA9mu+w0TS5
5iquUExrzzcL/leUIH3GhYlgwMom6dRgG2V7/7XxT+8nXmhaeOscS2jeTAhFdr8qArG74Ue90b/J
0Zt+R6UCNwozVFncdvkhBRsqxX+WVa1fy6F3IG52znF2YIlPlaF9JIYsYCm+Y22yRrZhvZSl35u6
WBjwt63j4ESc6tcGM0RG5QpWoAIA6YceRLuuNLxhPxJx0pSdGvu68oaluQRzl3hXDi3g0xU4Gfhw
NgNnB/cvU0ebehGji3AhygkRzNujO37MYU+6fGL3qKiDOpRxU6aU3yrGzJdB+5aUmtIdlt3KDTGx
Tb+6fQs1kqPVVS45sA/mKCnBRI3UHx+/Qg7pFLjWMXvbhPAMC4EKPPul3Txvc7f5rVVX2kE7xDh1
qtJP7IvopD4EUHV+9JvHZt4LiBNC3fvAz1+aAp+hZtGdPC+8GiXzWJUjb4bHuo+YBXRKf/Jq7HQH
cs9USftnZVtIZjAZbX7Y+4SHaZA4JZ1MlANjYST1jEObCBNETQw31fTfs9+/fADH+KMng4czjpa8
QoRIlL/MkSrfbgtbulyDec1yHLnpdNsm1fpiFvYOoo/BBZIvdTe+GXnawoqBks0dCd/+DSM4qHUU
VS+aP9ghCCcfPg4+zQHKRFSYRGw5xgb8bGNErib2q144HMJkTXHu/1sX80WbfFSQtjIgeh0/7iBr
EQm4D5+/3hKedYHrBEN3kkiIVgQnG3oGKWUNP3OQ7Ua3wJH+e8rFE9t80eboJUVHot0qdiIm+jWw
+00Pz3vTJUsYJKjBpv4cPYGK3iwzU3bM1dPlTA+iPHuo0l2jiuVEIsHoXbyMKH1p+kBu+awlLvHn
hwh9r+QcGgrChvby10nsdfPE8gmE7nvAunueDPmNvaqoI6TqvYsktaVPrT1YQ7san3MSWZOXoWcp
5nJxv8nJlyDvKpc628K4Kj6mmx1h7bVafYJ6DzNIdhJNrrz24ZMdMQW4JMsh247+1Q/wk6ceBCtN
cJGo/SmEilNge5Pnpwu6ISo4HT/X97G7JJd8y/vvJgcY+NP9hjiodu1U/HDVUJdrLBVcAh0kzLVO
1V8xbkK7QTu+6MF5GaYAq8Yiju/X9lkxigWhqqhe4PCqIRhPxhMG1P6iNIreIGb4F4r9GmZj/hyc
MEKrzdQvUwiu2ZiG38t0gXryCCsJVPvo/FLtTVaVMCUvXGrciHTtA2kY/4zW0vcoH8HZJyaOoxGs
2XfljZLbsRi3CM6m9vuWw9qpUGWQ9hbLCNUsaniAS1r/uUnfOrXX8Tn7zGqiWelpM3v9nsAaWzcd
8vMhsQekHTPy6D0yRsGytJ9Ao1yI5Zhy3zg1PnBbGq/iHWFQ5MHyk5UkHTolI8QqGwbYFq2ZgeTM
e8gnmBpzhe7SIa9VE5LosZHMZIhSFPukEHhsyivqhUjAALDoCvFpHdyO3ixnnezxv7DmwD7wKce/
ytozbbRJAuudEXAew5cemj4Ua42kZTY/6mamHsDB1BO5bInrNRnV/qDu5mW1QwwkpI3dBDGqlP9J
SjQUHwNHk1dlsxaxNGqdmSOyqbh3yWsNp/zrrrG5tlE082KV/ZQ6UI8HuIlCq1btS17idgvMtXaT
/4QFKsMxUA5cU75diMj5iViNSTuML6B1BBm+/bEzD1t5FBbTyDXDsGNodVWz/3C7sj8GMEMtffFz
57WMAYLUrwM/tTooIpTvBIL/Y7PZ1nVpnusQznmqQBCOoPObjE4TXQPfkiSXZskEOb8kAxx8SVPq
VF/CeWWCPcaimCb5YNFd5JxgdBD7R6s9yyKy1HpJy8bHMAaTshrEIyKx4tXLizYfnC+MWhoElIkk
hOiTdeq+L0LOM4TRpjgdJsouNP8ovbX3I6x2yhp2tU2Bl52DLs/HctPw5LU+8OOb4eJ5TUHTM6WP
HS7btaRj02WmHWEfJfWQXZg4xlFnNPS5VcLns9k0WCzs+BM8xulcyifbrgC/Rpj96pngH3EjsKkD
rwyCELsx31H74LDq6ok6QVZB0KQPV2of4ZED5E8BNtlrrt6g28iW8h0KsIW37HlQ/fQeFmensZh8
YK+QvMBd+vw5/uYwsKFPqXviNfAHZINYXoUj0vpVFE2HUN89G+pARL8mTZAoTbrgWuCERZdPxZkh
MC84UFT5OhtN7b1tpSZBlB/yE2DO/Ej1Lc0RA5S04eYx6uU17iNfqlgC55+dKgmVhBwp9cO/FKgK
fhAcGRXnuCWp7O031IjcDxVeY6lvAAsvJ8xTg8Tu7LQ58Ys82Wau84+ZsgGONEKQSPmx6PtGpMgq
DcPdwxsdHE74RmLOLUQNkNKArV6oENjUOp3U/LeTN9ZnB3VxKrVwahdZvxRcqq5ml71gbyguwVss
7l8Ayg8fH/pylrq/wbdHj/Ju6m7Ml2OeqAL0OGskylnoJsd9WXzlD2oUGq+od400AEoIL/Cp8dwS
zzw+a1QnwLvRA/JZ8/sMh3inWfZEPG7L03/+mT8cFYt162TPGpbJ2wWtSOtzeUk9WlgsIlmHrTOd
JuLU+RIxKaDN/obynVlPxKa2UaIUo28lwQ/hHt6Zu5esrkcKpNFbZvkFRXM78ov4SCFgPOhjzdoe
AjBw7NdnZ6Wd/k+b4ixcNsFABiitjnGFc4lZ1wiw6YvjmRQmSob8spNlHcp4QO2VtOEJAOB2IzVf
hWWHJtNoBqsjfWm7qPxiP9BfQcq3dLKyzhSpzxSPkTIdX7la73ZhqFv41+wHYWzk/83zw92n5Dhy
yehD92jBOv46bfFcWlUVBfmVkzliVRMFZ7ucBkVz7WnFIIvKP6niDzeLYituM+Z4gp1Tj4FUP8sV
wzsq7Knv6BcNQ36VfWUDD9NRIZlxRDC7WvOK+So9X6NCZB9LRO0N/bCf7CmwIw+G2JWxveVS+ekE
HElNIjkcRZ195VDFSPyu0DCDOx5gtmd3syoXHSw97Io3D38AjhWAU3xPHmF7OGY/5Nnd2cHeT3F/
axBeEUqcxYrmrQWeFyi76Xtu/sjDm199Mlfb7AbxuhpQkyTH8AXWa8MyLb1xkiYISZeTcDAj2+QS
HbrCUPFyBgTHsMUhx2AcUWSCjI9ITLy29ndZcatQz54OSBYcRtbUeY846dtqdGgwnCx9vy+4A8qS
O+b2+aUb4r7x+f6UxjDsb4sg/NjE3trriGvM8CRBupPyLi3nIftm/h751g7l7K60kdXWql3lqUZS
tbWiy0IG/tSMDaaMzgUmgImvfDQJrf5OvorivvFA+N4+eRWyz7kRMErxEvb8cbT+myB5UgNF6MFo
FU2FT4nVOvT5anShr19osd5UgcyTem64QrvrpPmhp2ZmwDZX14pibrOqlZPYE2FsitofchWv/2K/
JQVc0Fw8UReKYMrPF3g+oE2WIYjEdi4B6SF1FE8Q/oV6M3JcQ341BmgSx07bRqtLUWhejBSsc2GA
oBUdhJANWoYt6T0VtT9rW5ibdmv9sDQuJ/XmJgbZ9+qGoU3CCrNt9V4GA1ZnaCVH+X+I1KcXCyO+
aJroZZLUuQoVNCwtEktsezECgl/fVNU/Vb0fMAHDL0BYTI1dhTy/6ceB9FInGe9MUl44BRNqQPKY
BdHNn2TjHKtil0Vs3GX/T6cQ0tAjF499+GtRIBKfedMORXBNBkU0NX9ODHLp00dMcTv2AaiD7+0I
iUO7gc7ayUSOzEjcfE8ev1qdBquPs9WZHIe/WcZKhlYIktotMODtE7xvVRTBZNlgATOe+3nqVGoP
V0WxsfHeKLmyJmj7ReljUT9209PFslss/n0AdCMJH26P4yEinnNM4UzjC03M5kb3614lgZr+NAde
61cl0oKjZvg/kxxr99HPvPEFiBPcovvzrsbsgWKr+Kiis999Ftjc3fG4VB4/CWzAt93cmnSS24uz
hZHWDrWJpvPul0Sl7EyjX7rH0tno5ot+hATPl+/Z5gZBFNBmzwsB0YuhWUD/cQzX/cF0OsDXqPDJ
aGyO/2z4kEpFFS56PE4C56J+mnxlFwfpF9iBiPrzmpndLqRUfM0QxecaDNYKf20RoLpI1bTLd07O
w3q2G1GIrrg875L9KehQa3uw9KiPorRkhmjbvmXcBsVXhnhKKumoZHd1srASppRnfqXu6lGg+ffe
4/Ulcf5KRl6w3UwA3F0d5V0mbu77P48knx3K+AvjcLnHQjrl6JI1LPTABB8tPvo7nBKHNwkioXwk
9cKAxWWfDTGTI5YQ7n9/63rhzl/3rSCN2Px0Lg4U4VlH1tbZGO789MUeSOlDN4o/1KBhKZQVDl92
wLWpDtepDIbTz4TZ2jD8OJtjvKQ+TxQz6ypRzB7KL3H8CC3m2N215BjyUbQfqqseZOBrYKYZA1G2
g+rE6pB77jBMNw0RJakrqD7/TgvC79zpmJFKb5IBPKPq6kjwWL0t3XiyGGXkBTi/nUu9P383cMEP
TVQ6VOCL7OIvv1jxF4gC40cz0HOsDgL8Fr5SROMt9c6xlX/+eJoRoEdIUlHU/t1zomSj/oydtIvo
G1tu+SKbcbdJ5DSvxtVQ/whnNjDlhRrDNzIUspHb4SVcMzN0sBgylMdb0R9xxKYVapIXJNDyNTw/
EN60emq4aZjFiNO8crGPCJ3IyprB/xnrkKL6AlJ1vOUc8pmDWCPThkhsWuL572i5hgrSI12g3w6r
QOUSdIGDzQetC1vla+6OM/nWohwBbPenfsn5tYpGV2/HM44xQvv8JHIh9KAZ+H1cgJM+TN6+Vioe
Xxk/EQ8Q2QxMdVIOw/7nlq6Bwz0PDKqCAVkBi18Mw5tOachD7MLQ/6tSbjBcSXR4sgyjbXav65kS
O4dTn5dEhZ+ehehwHuofsezdseeqVH2f106fuHdyPQO+QbdjUV+fS4tSpIoAFPeiSuqVdrnYtoPq
4bU9iSa2LC8yeW3gE1OzuEQwgSnupxBOJsxn1WG3IlWnOw4GkZvxWK7oAER4kiUAXnKqy5D+ZzRz
FanadVN+QsQU3aiTap5w+azM5u/HukY4xVr4AGbZsqlIvkF/gtzAcNydTUfrwj//yvqs+uqfwcrq
r/qKbk1rq6XZ1V+yfa4KsoQEZenMcYpEiH5ZWqcw9fEJlEsDaggy1YFn3TqL1CqQJUjKxxPI0Yyw
yow/Z/J1KvvaaB6nUaUuPP87y74vrh2Ju2gjVeuMch7zaJp7UMtPcF7ktpIr9SX879qtP59/RB6k
kTTzWZ+Ber4ByAY03C0+w4dy5enIsXFQOMcX4Zh7TMadEqXlwXpvKEgV3goWARSomWav0I4XFZ1D
wbLWPHc1BbTgDPUc2J7eOb/mGIUwIAor3qVyeCP09ONvuFPOFATxJ1gY0pmPsT9dtj9hu8ZunkR7
RsO61KMhpHxEQjknopXGU0DyEzF0I44OFwyHpul4FgjA5app4JnV9AJAF2ce7AoH+rdPDbMVxuy/
5GjRPebPvo3YpOdJzInvt2JGiP5l6nEJWPlcemMszL11xUAIiUcFNdzICK6kz60xfIRs4JWWSks5
ALliVb7nPtGoZ8/xT+uJxfffI2OaUwHkOvHmbd3R5B89uH1qlA4ZBb0rl42LKyuYd6QsI7iYhzL3
SaPFwCBLDSjkXVXkysZaXmN43Rw1zcPdinXbPIQmfqWzMEqGk6Ia0Xdnr50Q278wkf6fsnoSjKbO
j/UWqaDPjMG/U3fIz6zU+U2tvoK47+5b+FYN7fV7dX1PAqli9N2pCI+MoqORMBu+Fe01jwGcuNu8
fgP9S5klIWRbKqkeHZyUj/VnHhJCFQkJb6VCwuDatY1UJcur7WgR65J3CJmm9ibj6YskM112R6mN
pbAJpraNsGbhHMDOpop8kWKfwSnjaIvBlV49skHizTP4vCGifNVcw3o8upXp7fUBg8fGViWSzthk
CAP3vWejxH1a6Uiou1tuIyRVDj2IczyTp9ebGyvQ6Lb8rcHCuFSnXzc+sabSjVYTAHfrw2z0sNZh
TTav8oHmle+1jrqS3gErHAZ8/5vQ+sH+j+YjtlBZjwjOS7qiNWtO79BjlLjzZk2z7YFpaBi9NXUY
7kXRC+svUFzLZiPtBkJHoNtgPRhQ/CepEU7I7MN+2KG9LBUAOuu+LXiwyrYWZUu6KSxjNJi26sqk
KQfl1J3js19DSJ1BGwAAAJXY+7TNzUB4SIwghzu9HOQgLmsUT+yefgpkv+45wd/8Vw70X/zLIcvT
SlHYakoiOW/DLyrs+2hRFunf7bznbpPuFureC6Eh3kDpAGvwBaxWdwiF1EkQM2Y5c4238fNqRMMR
zxLhK5aSfU/CPn4NJ3L/LjHe1W/E9ZFG02c3fO5w8UUH78eAOStjnE2DpsRIOiBkLlY5uLrnh8+5
UCJbYxfTDJJZQRxRgbb/i6HO35RKoFPj3V0TJOQ/g+QlF0inStukCM2B6uW7SdhkqRsT7R77S/1F
wpy76FpxKicCkU6b7x0W9Oc0jaYJVdyyivtxI4JgpPKS391m5SXHt8esnu5vAe0f88SyUq6v9Vdo
+zFy4FincKTkT1g4DxVW6WbQN1dGwK5ghuOi5jJcjeoV4cOXuhbR6GbEqT8eABoK+f+TW3lEnM9e
u27gmfVeW2vUS49EIGZzw8Bf6QNt5vkzFK7Tl+L+1XCPBcIRPKVHJQLEFP8hXuYKayZjElGsjyXq
gBNVdW+A1SgOQI0zGKs2uKhbfYBWCPjHZvbtIq/D8KVW7kaJzP2QtclZqHoDuynbSMLRnsNI3wCM
2GzPPEINP+9mf1Za9ry406LoNc4Fv+jSAlwm+n5rCzIsQEAB4KXG7CdySFzY4Ad0T0kWdnx8e6ff
kFH8mr/Fmeoz59wsmRFz5N1MEPi0lOJXL/ukbqIq38pzRkTIPgAK2qfDloFw7BtZYi4p/XttT5XM
++u1a5ExTLLV1X/Vjd/ZB+59D3HSns/7tRlm+1OWOUpbAzv6LBKSWN94Oecdg0vzRiiJuQNh23ac
S36Ri3VUhgtJ1hnDMLWU96PZY5cOFyp/4DxWnNqIAEfje2TEIQBtOdNcDt5llUEAH4jlpsDjNy9r
8mgIOgtPIF7fQXgBPLmTb/bU2oopRS4a/8s7GWq5FCrJzLY691lr4LpN5VZRnio++wGJWREDMYCX
ssgFb2P6nz85TCWBmlee74IZJyXMsoSYYsrPogqRL+XGFlVQilkpaX3TYD6Nn1WYA3KH5QmZ9XZn
bHWbfKxs3WgH8WapovKQnS85rbsrCLSgJofwwAIy770nHMUJy5MUPNLQY6zra4ETLEq6y61agO40
GigfbavEe84DBQcqFa4Zvgml++wor25swbKdk2KMi4E6CBxNU6mYVOVi1Es/JKEol7v4fadAXxZx
5DI5OR5zs0qrFx9Pm1Lbp9u0y6dFmHBSEEwWf/cNFUCaHaip8GmzO2PAwXPHTL9KYszjkHojvlyP
lIxaNVRnYlFAZwO7u5liEh+AcneTFKWeE6ikKge2QItEpEFCcZP8XhaCWyinVKAUtDZD5PP0d7nQ
e7bjKqQRbHJ5yqqm1PF3HaMrbnD62tUOurp1c9d+tt+tybBKDw02DATvnFBQG4ZCpcWR9UKpPmMw
/wnG4KLX99XL1TKcnhF41PQc8Qa0UYiRVyuo4cGMJ/xzKOsYOvxKRZMkJvo7JZHrQ9T6CH3qeqff
vEJ5z+kLPbX4d1UsxfwVeP343XO6NoE1ld6tJe7++AbgJe7OK2evQFhefYx8ot0OyF0j1/F+ddm4
B0FheR21OSWDA4ykIiGrLUo9ldnTEUAiTXfx7V/I6s0WtM8/QdXmL8DSt04ogvRfXtwM4+JuRDz/
nGVbHEXmSzugurdW8p7qRhI97Q/b5bq1syeEyZTVd5kF3JHIsEBwVxrpYiapRrRGMtmlw/EYF01c
ZQmZI9VVy6gq1nQJDvH5El0w6cc3obglfTND5CD8UTaIZxs/r8Ce6TnCJ3fk0ycIXP5/kHH0CAIT
T98bTI+t1S3IsR6UZAC6OaqEawp44BfggZNm7sK9JCZImgd1feM13bFTIAg/0UlccAY/BwTQgACn
bn4UjP1o5JVBrF5p8nE2laPdAMDvXHPYsNabnzOrZzMGHawrMECamBPZ5Oq2JehhNamBDdig7FCU
W/qz40cgjhE6/2io+CRfGbfYjXrs02szcV/ONC5WmJO/bmtZQJisvI1xas3OuSwPgVqj7qhUbeF3
ac5unBRgKN34KxlJiFgD5GsKLibqGzlSK1ZUvcY99Mu57f1wWoPbyu+yoPELUiA64NrouGaAlMHw
rJ3POLDFMCg5mvum+lXtIKZAQN82PVii61VWb4wUvXQpzfeGg9kYfDNeybPD8aGIqlKcXafMA1ix
IhH0saVaLFUmxqhUg1jUlAiMrID4nL6ogyAHln2GWjywz399iDV9w6rCQASDRSrNX4kXV5iKoLy+
pX16dag+9Bx+lFnpbn630pDEHUD0NFZURsnZulozvDlHjKmB8Gn4V25pwCZ14OOA0w0oIO7RzkLn
WxIAtc9z988fNfXIiaVYoAOkzLNpdv+Cv4GTFepJtON3jZXO/c12aCptSCi7uxx9iH4VMFNNd/Jf
yZTj2xE3p+RHjKr2u/UMNVitEju1YdhEh7p35hzstGfWkL24ZIZB9ZoOpe/METXtnos8p/cNq3TE
TGuZQVfjg3FbMugugsXgfJIKGuCD8CyIhkEduFimzHY5ZsPtNZyQ4N+oYZjNSt1lCO7Pqv2/Gt22
tag8Gu4O4pypcULYuhe3thoeqYoI4l4ZM5sdJ8XsabRG4MCqm58R4rQYsGR8HbrDBrp+Qrqy+j3Y
sBoW5IYHMPHkU+jk3C56kP+T94VCgnp1VrK/qp8V22GBhJhp//IleJ+ZWAs6sPJ3c8OTVZyDhSBz
BefJh2FUaYUbEsr3/ziXjO/wXts2RxtKB70aob9fj3S9CiL65UdWSymD4Ta0Z1Jx9G9EjGmIsU4P
MkTdIdroO/RfAd/h8byZsXAWUAZBPyuhA731Cxi+X1thtBOE0pnHVRRR+02cFaZhGX1UsrZRZBYy
erC7VK/qjLgMt7cJqFW45/9a+KbJ4ELf/8Zp7ECP6yxr/W9dfzVq1dX2+nnEzoQg2cKmv+HJMRDJ
LmgDd2wEiai1y609kTx2zaX0Y5YKz6v4ubABqTFupjd1NX2dvDN4FLz65ffnzbS+2byrapCvFCF1
88ygazAqhrDS8Mf1BC6xvZhg5vRITFO5s9J4X9T2Y7EUVT19JTN3MliqKTPJ2fEFztsTPtv7Lp+Q
LVECcmmkZsg5S7zDChL7eT+cFXStqioBCmSM9OwnSjRFA8zQCQi14P0cZaViBRFyV4VyqGXKmovW
BiQ1IObCdlSf6I5j6iHbKL+/4QeE1l7cAlWSQOpWU4pKGw13Eo0Bz/w8TRdOUQDHSMq1Pwlfng5q
0sKnr85oIdSm8kTYA8SG6J9kHVAxmWd3M0JX4ev2egj4YDvUibrPEYbkUgnws+CKtQ8SK/zD/sEF
FQ5LKn98ljms+EaHGfzSeQ+rMYbEUfcgdmDfTGG2rCMNTtZaXOb7RyL20fRnh7RyaXlBpF6HeYly
wiAQ22YC14csmMLuJLyV6dGUrpSUl0Nhc2vCUTC5zfXgA/pt6LysxQXeA/WQRhtmsjPKZhqp7KpY
oc3933hCdM54bxAMJExVpPgQDX1d3au7/ddXOFHvnLYlQT5aGiCetdaL3TLsQJTBNwODuSF82/jY
7ClQeRdgeLK/ymr66+H3YFrq2tkP65AVanewrA66pNVxOOr5Ds0EXZcU1r/JIvzwPcOg0v0MGZLB
NmJt+YDdDL7Y0Q+9EC85RpH1jvYB5fNP2rsXPyAfIZrSqzZSdMdBidfncGXvVzuuxTvFkN9HvEU5
TomTrgnw6OsVSi0GAoCFFUFb5W8b8BiaJYhnW2luHqcSHnios7StiMEHYULXRqJOqARUmCtTnRgH
hc/UyWQC6kxaXshQkNOgiOL80Ij6NXy60cDkeOJNxBAEqQ5Wtn8GAUQIE81u0gj81R0O4St9xKjT
vu7zESv1ovrd9/vAGw0rH/m5Zal6HLYH6oRn7BgWxeJTjhuLfdOAe32BDGoiAS4N/ZFcLU7Z/zWw
lZT+pBqnfbfScAZN90duIW76mGlYYnnIcskprLxSXQkK9foLaggud15wlFlwvS+GFdfHavbg88+X
MMXjWJxE/P9a8O2F5hpyBClTYI5jy5HQEkMkeT0dU8s2cJgbACErlnVXZAO6XAWcBgp3x4ZR52J0
Fs2jxvb2xvMzH/pz+8DvYIHObezGRB6FEHzqL1A92wxACq5UiD8xp0Dh8fg7g5hrRhHd4Hs48KWD
lba7U+v7D2hPvyONBakgXxrhZfm1Cglsz+ts41auxS5JWy++bTbjbG0f8797BOE6gU+4UaRncx3c
fK5gIM4nIcXwLmWLiGbBJsUx6cZ6IoioUgJCdRM1qZRYbbfNizKohhVNKsYi6djWBwrxkD1QMuUd
kfNTOQ+dQrDxxHCgp7xl2nM/BQpqdwNefb196QRJCT6tkMzIY/3pbyOhEHGdgbdhF1VQ8ow5mBgY
Xupl8ad8MT+/+ts+NkSr15sHuBkahVp0yFdqkwcdE+OlgCmSdhn/cnrAUq5Fddmz++QG0ec9fhcq
Zt2QYrrF9g5DI+cED4UtZL9JHUsZxS+g4u+JxrH7c8Kr879zOjQ0w8H8H91QfhwOHKihLDddLSSk
soh07QqNToJFi+uwZu4BPcBm2DV3XknCsKemrJ1YJq7cPYJmeB0t1ItVrsiPrptj/wsdgU/Iejfv
lIr3E6JbyUjCAROsaxOHrCnaD1HwFiqJhfyHTRyyGITtfadpuWfWIe6XHlmS+JKrAMk5k6q7dLKX
/kDSDhqtqG9tdMkTpt7Y1SYFizoxVK7OOFUkrLACW/qwuRZk/Cv+JJFxRx8bwJ36UuJ0DsmwJoLC
Z7jvXEADQHE0Hn+6oeZS7MhSC3g48bv37EU9H7ULYGGkxTv/XiqhND16gNQfV/5FbYa2zVu3KXnr
hXsq9k39x141DEKKhie9CaVrIRDsP50MMcTVP5vc5P2FIJKhn8B+6IQJYT5micDTQ3Ol84ljJE7Q
vAszwjKUIJlhfssGuJrINUCVagWq6bjNXgp24uX37ZHMSEwOnM9J/V1LDBm8HkSFPcMA9MOPdhSs
WtyOk/SdPUJvD8SS5i8cFXyQteMeW18Om3X4BWlhVs6JypgYLI1P4c9jbm6G9EIX1y2CqJ9TWn61
yo0ny9USqeVOUpL48ROydF14lpzXxIfp+YEc/clvmAEzwH//yoArd0mMdFjyqkhL+zYF1avewMOR
y3LwPcOgWni+Wb8/AvUKBi1mLADhSYEtW9odLSEfPcG9l58EedMo2kDv+WfJbaR75+HDMVehKGyn
5y9cbsncpF3at4BV0UbZN8FXYtlQE8Ei9mAnrV5inU+3UU9pieQBcT4LObzydShrZGRxCrs4orYw
FTOD349Z2M1Tao4mfnoQnxlHS5anpU83ET8Cc1heVllaO/aK4XzF/gHSyQHiDJX/kvCSiecRJ9r/
V4/zeIcQSy1Y2vtsc4HPjvYjqUI9OfQyxI/bLmzG/k03oLa/Gh+2qcRYxswLeWtQtl7xwty2FJcA
NRDoY8z/qWcbSqPIY5mFdiN41aD1369sWBtjiu8Bf0NeT0ykx7kIvaayviLUBn6xfOljqLsL5mLJ
pyrHXimUWxKFGBnJJX3A3vSdOpPY4LwJEf6PVTeYxtgv5EbqTxt1pAbU86fjh25fU5MqviUWOdU3
xGp9zjHZpkriM/2gq3sgO94LlTcFSQKP2i/4/jucCt0XHibe5UbFsGuGEbagWD73hA421rF8KHph
lGxY7ooZ25mWma4gFScukTO8405lFv81QUME6cisZAECKzjkspKKpOPOwyPsxr6OIj6EYHHT+qN9
GHVyfC5z2Qv3KDdXEYs+yRyY0gCDExnh78dl/1wv3VNVF6hi36+xUS9IFuDVk2O7pTHdd2J4IHUO
cjdHt6ahNeJyMDN01Vq0uWVVrkSpTcakuXbWHzqVypCwfGbI/IODPJx/WlH6PFqJ4dayabDoa3iB
mNgY0J0yt6tmXypECItycR+s0P3kj3m0nrAA6od+V0Lc5cPfsD6ANLc2RgSLpRB2YzAeDv+8Gnmf
umFnRMJOrOtkAQfx6Av4TQRRn2ftLdFZ5T9XyDdD5mSYMvfjPPLW5TW09pBu1PhcJcDK495WntiY
Lum7N4cCz1HSIqR1j8qit2/gBp+jsvQhS8M0SqrRx4Nwk4Z1jFJqcIh0qapHQcom5+B4zgsZ31qT
/I5jiGBACPoQGgfyoD4uiu3JAiwhXzsD+948pNGRNJtz3EEyBm2Ds3cutaT5eqslQbpn3nmvx20Y
lMXzf647+O/1Yl2Goc7c9rQkap4dtu+H6vd3kuiNf2d2CEBnbml2I1n8EXKntCxpJ+kr+PncsAUJ
Q1wzbDMLhQz1A4TViPMyXvFAD+auN2Vqvmhm3ZgeezJ3tileULTs8zEeI4y4faQPzGq4GU2faQTc
pw8ZgX3pwHbtz8oJ9C/IHY4LOY/dHwyHciT7itst+W2k7My9SI7UKoOoHtxE7mSFP45jq65rSJwv
/6j0mZ3JlgqtKagmzwIhP/vv+vQqRbwsSROEoewaZ/axy5okapopfK4EE+DqGD7AteVKiOZxKI0h
OoWjBrA1LuYePQov5B6P7OjRH5PGib8iLNNBPb+bJpl337FVCkK3LcHv8Zgthlbs+kZjV+bEHhCy
4BvARKCDQI6tUaiZKuDGzmAUpIBFcF874rzUBsCv0c1UxIEV7SaCIbQ78jt8G6ux9s5KTPXkTLO2
0FfruFyBT1lDwuOqo2NUgiODWDJtOwiCfqcJ/S0UpPWd+zshukc1W1JPQ+rDqONusHR9neN63n8y
FyJU2cQ0JK7ztRGRRyZGHxnPCXa0LgqwPvb7pKKElaPT4kzc60wCKEj3hHy0DE5GLe0VB9tV+48g
OVDZRKRB5hBF2cKarH3GOb2g+Z03gEWOHbxPsyBZKUVlrK1KxoDXIPjvXnOQ4hKGp3L9b38g8uUA
1fTFLXvMxuuewiL8vs8azIsiO+JuoTtCbOGvjIJGyweRSi2P8dTKsVAIh3HMnC0PQWH9boTdLgW0
iFmzZmU4a7vSAK5eaoCUzzBN38hnHjaJH/Uu7AB44si1e8M5HnCZrj8FMsklEtxklKhAkny+H5Az
gIjbMtsnV8t4ecPGz63fVUPIskFaKOiLNuG8SO+lXmIHU+AYF4PXjG0J+h8tSembgwKPq4iMdBSP
hGA3RMZh9ftErD67K4tMwADsLAy2AhQ1tnZW6LmG8tGJNYuvB0tp3SdQruwE0nxRODeJO//2J6p5
DA7AwYyF6cUcY3HCdBBRuMHB84BFNTKIJusoK1eJFWfOvr8TRQUDrOyhSBj10qb53CqmHEodwEeZ
w0VJ8vsH0D8DUxkWRgTj6UlK6va507/EkIwRgrhOBIW24gW0C/U6biIPmp5HLDMgJo3ClIzgOAuk
rsMuQl4N3AUv1xhQVke8VasqnDpYDnPW4AoRxpkDiyn6nkemQ3/k67M5oEVMMGIK2zYpzYWbxtv/
+ayxk9V2IqVLwjHo90Lm+ZADkq+XRnD8/nnJn162YxJTa6pm3weox/9cYPiifI25TTfM+EO5p9S9
iTYMLuaSPYwnz4EtVcYX49knh1j2C01X71udRG+yFAMrtZbfFVGHSTgPMMbTcP9UHkTD+dp2fVvy
PcydL/XFC+9uvl3G0Peovb+l788LgZWjc7tNpo09+CyUDwOORR75wpR1znI4/F64QAVl+X1kV9Jy
NQa7SqzOq0U7HMFja0dCGIUmhQct0iIPPLrCl4eWrGPtAS38TsWsWKXQLrGU198Q2kdovuSXUEDQ
LPWgT0JidsGtTPjbvNgn/UHfLTApgD9Spiyy2tkoJdlUXEEnUxBZbUd7EWlT0Rsy/DfOBDBpNR3n
r3an8rljNFZS4yAnzpiDVGGP0Gt9mrmW4m0NHGTYC1ihTE1eLZvCHVAIwJ74kr1ef9Y+PmwQcP+l
4DViP670jWrhkdAffsFyJ7+8UeU3Gzc11rh/0PkNjRtd4BGSlSNo+/oNTSzyibyBC3grX8eoc1mH
2+efnkFgVDwtvfoEtR2raCAX45SgTVk4VEDS/pABaW07byAlifnhT/C4eMnm6/hZgEyowhvlvnNu
UpfQmMKx2kf1RwKLrR3cLI3MSvOlVbxjrEzsonok9LAV+6iRutX60ECb/aONm/Wld39EjeQT/rur
nby6X8QWIcuApBLXu9Zl6cFogL07FoFWBtVWxZG6ixmGPBsMFI2TSkZfk+5feNUsnwDGUUSsMTxU
aMx/6MOIo8JnOjj1EG9Mkh4+zQ4BcMQVqtnf+0q72cJUXryLekU2c1uNKYllj2xzurCggxrfem0u
jqP21UlAryz4cHuX48l9OFyqhQeCIUZewCnbBiyvtSsnJFM7ijzRazi0NvBL0kVGVU951je+6Utf
XJwQFNyPX+91PUy1SVg0S2fJWNnDhsZNaPcAA32FiXeY4srxuqz4n8XKnDfY6iXqGmSDqWYvbdG2
zo3Lu34xV7FovI3xMYmUna5glBJkJoMmSREN/xcv0SEhR9N2qp4Z1Tyt5hqr+6dIc7/03qcKxcv5
/8li7J7s0qnHM9LnWrHUzI/LvOs86F5Qa/TwCdecynuKfO9Kg8gsNhFvuLBwBiu+d/bO2cHkAuUV
cTVIvQQji7cAGrdSCuVo2qNaMXHNEPC7LGodbALlDAf2CMJrhDWUvlD0e9VPpQj4MdOly6IOJbtm
TL849xlzlLyHuavyNdQHpgO+eHRh2YsQAmYI9kwt4GbeAe0/LfKPTKwEKO+mcPNX+3ookK5/ncZQ
gS9bwTICuXcguWhX0JGO8lhoDGbepBmGZ7bfLhstB9L5783glEowRXuX6Gvjt1kZUBHriv+5Z1bh
yawPJZXqj89miy7btzg8PjT4Uml/FdLfzbCsQh/0kXsdg21AwzElj3kA7/ysXL/2qr9D7mO7TPNn
OsJP5ORxkt8tuhb5cXH4qbJ0oNCj0grrIYuPA2YU8QDr+vbLzIzdf6dSQVRffiD7N2GKtbGB7Kf6
PDd1sg+V9TU039kl1SnE0z2PB2qleksBiUKVDidiaNHOA5wOLU7m8OrCKOm7adR1zreO3Ty9PTC8
sR2ANll9Y5hu0JRxDQ+sr5iPkTnopWSO36dK3tlp94SyuEV1sCvTCcB08qP2lHRr5tCfypq1LzkM
VKz+HmGkj/CDFe95HV3nFBbDnh2OweIiacCllALHx7tzC2sn8rCJqVsaMFXMKEiyD7hHZRgDzUD2
wRw81vqykyWmH+lue6sn3DsAQzLX+ri/26Q19+pKmU2qOMdv29CfTmxZYCkrpAM5WvDaYg4luGCd
ULkAY+FloTjD/mP3BH6d4UP7mJNLXv/fbpMdzbYPeR7J0M9pbvjkQndxbBHw745umzxuo3X7IE3z
Et3tUKKx084bKFHzbD/3UUhUPr3n81hEl4yc7fc5xUwKjsr+bmqnFCEuhTsn+e7l+RgU23XJ8BFY
ZZFbpgWCRP/myhX9b1ZuOTIFiEiR4e/2V81HTzRJRkX61VXP6Gd3o96gImv4oB7yljmphI8XuufP
0P+PWy1EUkAWKtGTFsaAbN/PfJKQP0sIyB+uiGz93W4+Yd705/M7zxuikf+oIjLkhfc7zoKJVeeh
x0QdXTKMpV04R2iald+BNf4dZL614IccCUCJ2dFNMBB1YGF500OkEXnScfYpwGh60e/rh8ttYeIY
rQorkvbDpF1GTZje7FDQ2QW2aUMeJuWJIwBo/xtuSiU3pXXc8EzPJWXCwGozFDytcsF5NYH+7bsT
ERSYbyiMiaEyXzZ7MKhMAuEBtSjnwhVKLBxVY9Ly5EIj9eFNhIeu0jNRh+H+NtGhkZCe2gycntZi
TexEYyCZavnYJKaTEDWeoC5+223+aEI1llk5rLh7V+jDEVB7UTHOt/5yjbjUtJ1uOgMC/JVImRe2
mzGoHHCyiJ1NQkY3LssLxDrScBP+G8auRheWBb0W6gGR8NUApp8T6eU3Tm5R8fOxGdDV/fsQaSMe
dn7jm1N02tOL9sj3+RnEulMh5k0qmFII2KE4xVHZPsKKDY+H9jaeS2jw+HGlC0oe4lFrYnY84vjX
O7pHyaq1VOWrwtYqL34ekHZS2PLB7/X1FcAhHvTz82GfnqwcUsVd22TEBuReZA5Eb4ETW9wpm0BY
0oFtE9K+DxD90xrn9ehOEr9V2EI2Dsk4YTwta2iIcI0hneWMbPItMoNyQSDF1uZCLk5+QRsSzzoh
eWNF8sDRVAIKXiKZJvhESD92mMOur4RpSZMEOMie99xJmeILu9DPyYWIl1q3PULQ522WaYsO1uH6
mH0OTHgjCaO3JnGT2jtjDZpOV2aIXpHOf+N/tYRJEaPcIxkv5r6x5v0vIp2iQSBC5gIcT9cIQVu9
YoU4xfPsOtucmv8MaWgUjY4AxqEAwqeBXfpKmxn3M9MXh2u5PJZiePTvoRjOcIj5MB28isTyb0l1
uK6Oz+FhfjdQl2nE7RRwZADI5bqAmVFlU86OrKFV4Oz2KjnyD7sYPiCb4GHrgGbdvlFyf4QA2RN7
sB7czPHpixQYgSNhMCGd0I8sUeivDyI3fJi3FaX8yR2qhX9dehHrTbiPromoMyOxzBV/b8UFactw
ZLBga8mXmX64wT4MOTnIcmJdOEBXtll+O68ZQXLNZWkN/ehlU9NiVMUjPHQTviwdNVrSca6uLY1R
A26zQqlAXL56kkVFraunX2S0apelLhCRjM/vYL1ucTc34kg3Svu7xYv2/+EPnl3RwrWvCPiu1yvy
UM9cNOkXHk3YkXx8qefKIvMKd2Fn5X6sCWODNXB6+8TJIOPY/W6Ce2sbY0zlC4UfwXCo9DxvQd9L
O4wSsaxf1AXEswxZja+yous2KgGO6eFmIIufpv0FMHRc/9aos2udvCUTzwUajlx/OKBmgnApdWQ5
Aa6Fk0A48CEdiLGe8mj0rlnZ2DTCNdE9b9cg0ogelXlIUvJVD8LycfgSbifLhPGz3oruvMENxqPe
1oXxETEK4P9wP9nFJ8fhD6kXUNjYMCgVSo3LOV4vofp0nj8un3r7USZX8bodh4bGSvr/6g+UP07t
+bt7Aw5E2uBXQhQG7LyAggqUz7azvRcqSOoIT5hvIJl6k5GDx7otEyYaWBgg+BeZ9ClfQQAJ30eR
fz48sEoMi6McPXsi+CaHfMLOtRRLEY0drWcnMmX6fFYj4SUore52uB12kPT4RMoz3eDQye0C9+/c
Vc5tL5ZU68qU6g7qe3163PMAK7YkRtjrLcIleHXl95zFq/WWLa9lcAEV9v/GvfOUDNLFctGQnn0q
VMwv7MbTLgNhjgBNr2zUPG0kNGRgy7LOmYWg8BAL8+AzTTNwoX/mk1Vun/op1TnJAJ+Lb5ASwyVy
T5GkC7Et4n6h4UbhiDbMvT8uEEehvfrHrykFJjtjv/1H8cifqR+FV/W1lUisUiEnouq9jr/8vXts
MbB/Oqju4lT+Zuk9uuWWGKk1R54W6AJfjjjD6mselSn2Y6E5df0+9jsNn30OZMBo5tCJ24nNwSl0
FimkdbGBAC0ndSPt0Xz7vr1Gsnu0pCb+CxRDScxO3K7dTYo1O6TIzpWN4CaGm2CxSVC2CTu5zbJX
GLIZEBZOkokKqfZVs5h86Nq9O0yFtLNx73+0nNSJMtj5/AOxDkcDU2sWpgbGwtlvvrwTfbTPBTDg
VxbNdEeRs/tkOp9Gw6bAkuZnS+QJG3pzkkLsF9FVpPDGYOi6Qjur01yGRow9qw0v8TsF/LFBJXvU
p8v4kZ04urID8AtVCM2M+ot+mfPPK6PvjBUTq/lM01SD3GRglaAERn6jX3fUI+bA1+jycA8ehr+k
gvsouQgcXIlUYqjpLEtQ81oOaL2CA3DbKw0Vf/iWs+wMUb4q78W0Xhp4ZnQoOONezlZWx0NYGJhr
2/bmJxrNtc6QdBQzWJ9Q/osFekswvjteysSCe7UCCg/dm4wwlXILusFTF3cwctnmeREDEEaoMay9
CwAE7bma6JLYWIISpQnsW2jwjPli7+8PPrxcRR4Mat5nOLq31HI994PKsx8MYUNj/Dy/4UfYEzI0
ropcpxbvioHopZxFqCQYOtlF67xM4+QQtn3mjmtAyw80fjovSxD0mnooPnuuILhIl6J8solFc/3f
oaVcwNYsfOnKvltPkakbKm7awIRKEfzv677YhGT+ScHdffxDeYV5rv9DPx612EX3WkLYjzmivr16
iOyItOxIB304INfFk3SEJcQvMPwuuZjIqcQSEjm0ahXOQpaWi3CN5lKYRuVlFhoGIR2D9cTQfQh4
r5+JSO6NLnRufrREW0MFFzXAoMQ14dez0LFNqNeR+nMegELrSbSXj5c+bKmihz5AjpBhOPZqhW4V
FAHesNrwOKzHpKzUwQaEOoxEt48CqnUXbJUjRE3El7NX360UZvpqvtp+A/OqlvOvk6FfeOTnpiRx
TcHM+JTO16bZZDL+dVeD028VB6pWk9l3029TCjET38n6riEggZYJPWC6PB3WSdzDh0XkVipHaccu
4gUoBm7tb7YaC9b4NFtNbSgZs0kUWcBXrGC026CMj1TbG/pSmHIEop48bPVDH2US1Y/I1MHxeszy
efFOkL4HBty4qqC3hGKYhWnyUDcYg3rVy6JA2uaYUh523R5r7xWcEbbh45qXkXbkmHoH5e4FFbUw
2oOV3Bd0bIru4Y/bkkkBpsQTSKTh5Z+SBsu5K1RXYAUvS8W8jJyjMXqa2pD0CTzYUyjlBGxcu2tO
q/wHVRh0M+Z1RVQsVrgGYcYmfiId/7rFo/fWJlDR8wLQGE/uknfUNA/j9kJgLauzzZAfemPVkrFF
H6g0fSmDrYkg+oRabKSyvhlYRr5E7ooSPw2N8gGJzt381t7AkKfuYeao6vsC1Vk1WPQAPEico4A1
PwbmMYlvvEmVXHiSE2iPvqZUsWkmavqc6Qkre5/T8AFcRw5ofCTLeVeLP37Mrxc5+kuJD5sbNVJE
TdVxs3dnS4mXvorJ7T7Zyk9/ffGr3OUrpqM8fVr0rjPwsFLu0gxYtXvY/0JjYTi/QLo6u4C0KHiO
BMlhgGE/vF7KFKPVzA5YvwC81kTvd2QRGxcg5+J0RIkX8vR2Xl2beXSL2EfqIEXc6CbU+yaS4eb/
fKaqeSDm/VLlU04b4rSWoeznNlX2SIbYn0BsgLwTaxAkAIt7ncQGBCT5IkHD5RK6owVl+lYkGMuc
ALi5Hu4VS/N7Rq6QZGiHDCmQ9OCdXeO+O3QH9c67lqJX4qmJKOA1QpTS6HvsbmNJPHG1awhtW4pf
qL31eyEjefJBU6JvOldQe4KZNMq9uyQXx9AVyWsZVmAXRCrnhw12FGd+otbWRdd/TQ/2UyI90g2D
xgMwKJpDBwOXHEkwQbpO41WXqOIaCtf1cDvzEP+0Nl0zn9sMmT5TCAVO7d4wCEneuXYwkDjC7N8d
sqvXo3mKoDmnPaCLpesr/tdQ5QyQLAjhEMOHR/J2NRchAH1ceqbhFt3/IOTfM69cx97PCJABYNRt
uDKj67smTvH0QfdFxdt3r+Ia99yBWk4lR9k+GB33Q2DP/nuJUJVdZkT//cTVdv7goaCQpxI8OQ4j
VH+ls6Rv3bCh7p330A8vhs3bt7oqYSX+m9nkk0hRnqN3wEzuKrKY/JNZ84UaEzrkYv7ycJzWZBzr
O4VgSsCH4dJK8SkPQsk06+eJSvidU3wyh74APmhG9NwUd69AOuk92kA4iOSUUipUFhx8VTEsTNFa
acLXLVx7pSE0Eg7ayrtikrmrxX+HGXQXtPRgQHQMmYK5X573k2KW3Az0O34o87vtqoT6disYr36v
07+NOj6jsMaR379zbU6rcw/M3/0cBS+gbbl4ic5F9QNFMKlhPLFJdoT36bZuh+67VPoEYazTJoWl
CO7j+dITKN7/sQ9fcKKENx6FROpgRnj1CN6xKqbWhxQNe1kzULiKwTR/WCTgnZ75onriDIaPwvtb
O0i8xtXvWKDKGbo+G1+iSkGiu3N9wjFG7IO4O5WuE57wqRisLDkzJhQXPGanMMUtQE+hSlPw68T1
kAUEvwGG0F8RuA1FuHeGV+7MFY+UkHBs3WoqvaZIGf6fa/+sPgXixC8lYNJyL01GfCI6QcAa2ra9
QacQ8anUEvovKSn6ZZbKL9NuB1EMhRdY4i51C/bcWy70rKxRru3Km0OKNG9gb8KrOdONBzJMTX2Y
gJI682jWxJXOYfWYWFM4HAUiCUzMKwhsCuhdgTTQn0xW8GSzpXgGrUAJ0AuG5Ike6Pp/sKZx6xRJ
+3kZXCeEGAZ2g8qHkVoaUtp7Az8r4QbinFfPfiYAtqo0ecxM22IuExbjJqjhdfBirUoa1m6eKRPo
0kWm8M4ojf9C9BtLuA5EaS3XPVFL2fHK6SIXDkoltAWkTlnaUctqOd6Qz7hPHinTmr3fXRXinp4x
bxqNt6usOVs6/54tpKH3XiHKTSB8vyh7+oG32/U6QBhSKL7S1p7UF0hzJXCLFpnyJw4yrVpJwH2V
4zp9becISwDd0j83s8reEXv0ixw2tg6qwYMYQEvNuFfV6dN3pcpZIJVY8KSX2++juNtK0JH9uUOi
REclwi+q0PWhBmO4HBCwfi35j6URfmo6NasM3kwbDEAfkbJRMj/U1TF9nwbe2Gkcn8TttK4jhLpe
TErKhh6CXBzCwgOC2gcXVtZwmZYQX+p4uomA1/y3tzbKde4ukKL8nDKylvWF4hFMNW1DFaQ1BJPS
N/M4j1lpyWda/gxRxfb0MgEiltDI7c0MVex/m4oWH958LRUrvT2C9JvuD90fQZWr5s/cX+gkYLFd
ZmIYUVUoWMVKVA0H0Avz/hpnhxAliGTFV1Kc12+0JITvDrAYgWtLcuqRdnF4EsEF+iINgH8KU6DF
ib6sXr0vmJ9cNwQY7Oi/yFoabNFikpV8kOx9Lv/wNc2W0oWYOU8JCvKHzFQfgZMsxYqEWUOkaN1j
YVqewJcKJvy7f9PtKInF7fD9H3UpZ8Uzd3Tw9JhtR9Itb1iExxR4rUZ2LqTxtGLL2tbzO6nE6UKC
GgwMRvzafMw0DSHdkFg4LxJeJNGwCMNYwVHp6nfNl+dNlFO+yU1dtxnd+mOwTv6edKJXj3lZ4iY+
3xMgoNolMjStVseRD2XvfGROpF9XK5njQEDio+fwrry7WU6BRhqQDVMqinwhujhFgbX+4H73/2eM
NgWDQwS+2pGyTAYs6mU3HBxjr5B1Hhe+y3xmXMcnPGUSQx3ddeCOsz6pA4jv2vjPMS34VBJ2m23R
Xizn/36dA5tR1pT+wHB9mJm08+ixEkDfabela78SUGmjEVIKlvUxuVxg36AHx4bFEt3cRoTKb9T/
r0XkFtWjs26s/uaxrVGVg6PuJTdf9+zeDJAO14NBj+/qO711auOLc1qJk40eZu+aDK4JlTI5fin+
cnQwWqEvUrOFFaixjj5flTjC1nOhmy6wnhF+kjc4rZNjGIjDMVs+IoT1PN5BGxDynreeU+yu4/03
sVh15C60kqHQRo2EMb4/hn/QYOXPnB0vRfT+Ra8/Bo1FmwygeML7TTlH+Q0KO0Re6k6nsdKRFrJP
nb+PIMyqKFysbOH+/ojAfomHizImg/HNd2+jf4F+T8jyky3uH8TkPBgSSGB5JIiPIJGeECTG+UsG
+aBSJsJwx4SaosoTdRS9TC9BqGBFWECaHrOIQ9VW1EWz1vcnO/izbKb2E0b+fqw7UmoJB7/DQu3c
ZfFCRr1x6TpXwESGVnGGj5e5OHQFVzZvkvHOuqDfD9xsN+EcWqSZzrA0XillZtI4uB61Bjwud0sC
gRQUIu+8ZeMKDqwCokFnahXeTbMYWKtsdWvdCTtFLO4HDdM0QSkPqC3lUJwN68HX5iAo4A6ua7BB
0j46fsz0zPWm+5QPUPekJeV8cHUbnzpOAm5Kduwx8L/mYTUsQ0Gep2Bb4SMsFawpvSBnP8DSkM+v
D8/6ElXaFFotlvGvz8lOjETu1dmPtq6xCzx6nSTCmd0+2QW0Ea3gGidsTF9LrFmG7omkaCQ2+b8p
+rcCYcPvvnx6gBFk+15hNH6yI4OUpROQbH9c/px9lEl/ZTp5XkmmlGsTcvZG7rL56zGPdHEzfifm
xWDt5ulJ8WIdh+mnZfrEc31tv+bTXLBwnf9nViVy6hiRub2Aruqh79PBxgGxYolIV8oF1l2G+/te
2mj+WXRHJgGDIY3QD4LcXy9kNCw2oXDtsMAMZVtFLAexfIiEX5jXWXC4O96+iZRVluj4QW+6aN1m
EOvZgjVlLIQwEBlampNOaih8+PixIswkYcXphVy0BWkEbqzrvOgx5JC87brWWzTN91lgG1ZVBoOk
70uElWhO7/TJF84W/LJ4EXfxJP60dpmOkGw14lkaV/pjFJ50haOZWUTKswzOWfsqgmc0bgF/WgtP
bRyAXaxaMBCVTgZR2s7MEg4oONtvP3SY2qjFAKVRLDTIOMUs9HMMCSsOUERMhTahy0+zkpJ9k8Yg
Cp4GSquQ6qFwl3vHTa5DDLXOQooZcKDWRoifeRDndo7PVuSGfDwvKkJnuBvglXmlyKZmsz9nNDYb
p9VdvQLKkpEdQG4/1Vi/hZhEvV+fNmciq7euzihzKRf1ZDZbqFbU7mG9ij6Hsh8rYy2sKJ8WpbFO
cRW5vXB+q5XkSaCMbKbyzO3hOG/k5hTVGd2jRlRdpsgba8lMEuu4fWXA0cep6BB87cAHwt+pK6rj
WL/CAEO9pmT575ZkC9P/56MORxqDQmAhai6pZ03xJDsRCc+/7cEja5nWs8sYbDZeEcqVv7aTJbft
Qis7AUghEAPXj7OSsZHMmGyiTNdjE+2+vyfOuqRuWA9UV8fKaSORUjcNCIT2KCeU5n3xoJ6nFPjF
4ev5nDet+oLvx9zzetPou3UK2OsDvKdE47vRNeO3gRWCDFIcKA4EUL6+I/q/J/wD7U5EPKGiAVP1
5Fis76LUnIv0b374G0YiJGdDJQ1bFKjT1WU1SGEB/IKRVNJhPIbxCGuzdksVO0zZFnKeRwtusoQQ
KKqmGhDfs3D0dO0jxsYtKMIftavgQsxCM14gKJsaHGOG7tlP/G0Y5u8nFwYveNMAxWXwGO8EdnhW
1zawupu5KUXUC9JBQGBVeSdlh+/Zxzt9th+DTGKRgOFDWnVzXTN6YOhWQxsBXdTRuj8NiBjOeAhO
7fGozls4aMix8ATNkVeJssNBmMPRBRPT4hJ+xC2VjejAsr2B+JBJIagf23wI8YQeXmrV+XEbnjX7
EkMQP2EXbXgtOAndyyoWBIlSIn+pE0EALzKxoQQa1UzkN9Ij0nUCHoToc5B7kWejOw3Eu1EznAuo
j/wfnsuU4xeDTep6P7Vw6GdvHIlVoZEzOmCGED25qvPE0SJE97SzDg/AhonZLYJM5EuuilulglwM
Px/AnDNm100uUZ99zBJr+t59Pet30hkcGW0z9Qu+EUl422rgqenRv/tkHCMkLjgi7frEC0VXHJP0
TdqiT1j7VJajB67lmE1OMN6lHXCZT8vBFdzh+tUW++w/wpvzQyl8ST1ypB6faS4ZjUUYWzO0s80n
sEaP3zKbaOTw8Rfgza48AgIu8eJcRF4QwIWnYEuwFSewDUjt1N8eh3lESTNBJftK9Rrt1gPyoQXq
NrX1L+vw7WRdGzRz/b97l2g2vsZXWcqN3DDMBXnIVgcFsHZ2FSzk0XzDyWYA3Kcb0g7GtNXArD1B
svtkH+Rw42d+WJ+b0miARxKqGZcnh4Yj5G2Hyn/WBDQBCMjbNQGZK5K1+sy3dlP8akinZ9oWlZ9W
jBu5969CACtu8QgAbyADkmyiPyI4WL+yN2i9KTCkGHdfNbWIOIXqF1vnlVQ0EXjk/ptIXQBv5vAu
+AHywqLvZDqOPRxVUVaraNmLJG3tCih+EWwhExdJXbUhNfSSDyvChLYx8kXXee7fg/zjIkrWoD8R
WFQWWERdg246xC9WVZAQG2Ag6U9oTbaaDgKWiWh10j6iQqbekSg8Fh7X6X1MGo5cZf5wLFpg6ili
IWL0pqD4wsY7IdJ6eLJyzfDWX2N7e+KpbpYYmV+M6mPhUR8YbZa6MXKVUjlFmfdcJjZYX1a6P16F
88Sx55fohr0D2ubEHtbX085rEahxpttcYsI14ZVV2/JHWk2LbeMUGBAov047zeVWMzkuAeiHPqyj
eg1+JdjKbmsDIQu5ZAmRBEIEGYVY/OBgvYFGNMiJ+tZKZFQaHqkUOBh0QY0b2fxUdfs3uvzdmThk
/Y1iKGFgNP2sH/cfMvAGPWgnE2tIWS4NprkrP1ttlLdSFNQ+SkNHbb/B1Vz+v9iFQpsNlC0x1K2W
JcmcwIMkN36C1TuxM/iIzClEQ0VV1WyWPcoUNBBwGwBQ5Z4pWxK5qY6JgBGghaWpM/Yhqu9RYvI6
oXBWfS4s8L70PtQXhpt+i6o9HxIlpe5axxmu9nrIlOkqFuPPZNsbpFtfhRvOwkHVzjkwNvBLF8lS
ieUkzfCVfEhqLdEHx4nCfOmII76/YVMDE1zNRvwKwRy/WoR6d1edH3m5BbbhVCun2ta0oX+zf1cG
pbsSnZpioGEGNsifwa4sY/lMQnoakBJi0v+3Sw69HCNkBYWk/sDYiLVNd9lupq+uvvCQLEdVIqNn
kqyUGclgCUJA5YoRa9k6t2T1Gq422VQeKC9GTMQODmbN8+P7Wsx4HIunmqR8EL0Peh08Lnt9BqbW
lzpJuYuCBMPq1Pv7xiFaFNnXDrxYqBKlywKHFEp5pJgrjoniIF9hPhdN/Z/uyDnmroBoBLWa9UHl
M/HOA6TRcHwNNv1rscrxjsiwy6ERR9POqpsZwV8UvUdUKq7u6pReOyPCVELLJ4NKb2nUSa87QcZa
eZpvzAsX8pjwyFH9QfnlG4X9mQw4OxKTCDcqbzdtGqOEpfxnDgNufOvjlQvI+tuN0b5t35v/j97j
HYh6X3imiX/GyANZxhW8SGfBNggysgXlGmJP7WkprAhFHxpk0dRBXDWE1xZMODMD/h+J1toqQ4LS
xrDAG4cYQXGRs5RFwoRAZl/+8zRr1NxXDj0GC9XGm97fxlAQmu59im9n8iR0Z7qYtGXqNZBmw45G
JpFZM2Oz1WyZQUfReRcdGkOdaT0lBBOUhE7+9hGXJr3iKtOjxXBl2X0X4OnoB/HUJRwsNToJ4l3D
XCqZTWHGx90oxqgyI2ej8ZyS+q62W0tp95YXX3fI4p9Luz/7o8Hj5cZpMAiF/F3GBphT8XaNq3US
2HVHV11wJPI35fJHYQGLJ06TAsCQUJQDVgkWkVyNVcwIgd1hGaTP/as7xU3YB4zLP/cNLdhWJJS6
VnmYbLo3u7T1CVvQT+nSzatqAH6VQikrRjK8QEZkoO/sp63FoN7h+hmPEoNtVSRWQi8XQ8BI3TUB
JuI3NZ960oO5aC1TiBgUgDDDYCoD6fiC4VmbgecKR4jOFKYh6y90Q8k+DasIl7/BJ46pwfp1lwuR
o21WMYNQzla+3xhP8qO/3vGkBnfP73Uyk5BrtQ5LznW29GK4+gzn1EnFgi3CmWcSN1AiIZjyjqyo
9MqvRdTFoM8vp3WNWnRJjtCx1zO6ucrTXY6OCCFa3iMcwC9a007V+Ud4op2BSL1dHDLwXmxq+3Mg
MU0/ocq1SPM8930v+IuYTPFrP+ZEgid7wdZwDyUr6Y1QKoCQ8NWme3+DphmDQws2acMNverOzaLX
xJMMakNx0paGRTG7wNi4h+KCIZcqXd+vur7lFHzVErAJgeM4DjF/55oEnsYebVBW+n+EMj3lFoz/
rX676sC6/fI25N8b2kbueUAJDmZA0CnPRs22/JM+0oBKCTaazxcIoKuUUfrJP+X7t5U51JIWDFfg
hxROJbe76Sc2K3v4UJK0dAQyZvHks4xEXSKHjyPrg8qDjihsb0E/Oa9r0auVywOvTyIF62/F7em2
wo0u3sOIICMkhQxUBdW4EaMHYW1rpOKO4dMFF7exBZ7M4sz9IKD4gu5IxSPE1aPKvtxH0jCV3RWD
dUNf8KGQSN7HWpdQIndFSM81a9b32jnrVjYZQU8s6xl8efR+K8OGYxVhsbhBob6yEX4bg89yxFAW
sdIoMrsZsG4s/4xjgrHmc6FDUJ22jAxUegnkjiwnN6thC5jc/mCfAeQH9GoTwUp7Tf2F9B0ILjOS
Yg18QBlHZhodYiuRGzMfLrNege2NVzzCkM+gG2yplpbAIgGterFBEZdD6dno/CcG5kPEDMfLCNpb
vzKi+58D7HvVRiJOnO8VY/wGSLxGxgkdBTxyFETnLHNfrOGWlG393QOonvsjpW6JKdEicrvs+1b1
YYQHji4wJjS7YSgqR87WbC/8wlG0Cjs464k2oRAl0P/uoXTRDoQQjQteo5mDcuMmNgFLnK4nJRxS
XlTIkt3mmRVR/mpI7k+Bb5NqwonxJ0nNrywIbm3cOn503eJVDBTYFa18SrxwgB8bfAZ4S3cMEsTF
jlWVS4E1tl1DwA2dD4mbg0MFR4cFMbjljo3NnvnkWMxs7blMRtKrKBZXe1InDAjRfqB/Aaq0gSi5
uDvtmThcPcRZbUSJjNcw6IzwIJYbn/h52NYuPQlFkMitkoBDGqVNcpyT5gynqILK6eH9cfAcnahu
9qv9U8sQ3P6q+J1odzwEkqfv3HkCyy3BoDI/w3L1y7kEEIJgg497A8vDnDjCkBb6qDPM1GIy20EG
e8GVrPPgBPkdvXNUprQFyGMRRzj+HaZT9h4qGGDyWuKvjwSqADuxrreZHMy6rzGYm8Qdr06ouCyq
pVYYakONA1FzqoS9+IkIn5uFwRKy3leFFUL6BKh84temlK8NnCD7RxT26XGe4KjtQ4qLbYRDVbGo
UGb146/rd1z1qjApuM/XwEEvpu7LTGSWS32Mz/ssshbDinMwan5NsEtWUDs2CohHGAtpNqTo7qV/
iVgjH/Z7JpYTROG05Y/8IkRrAzIk5vXmiWueGfG1vwYnkHoKyYezIitgprT3zCKMOFACgHBzwjB8
b32DFC+DT54P6+k00plMUkdSpGKRhNRlxPgX4fs+PoxnYnrWsxB0LE+lyraEtjUtgUq2O3bAGS4t
0n6lFV6Aux3FuHYyQTYZZLvJlB7em/sgLpXedSJLMeqzrEDiOgJA4zi8sR/rIQV3Ti9anfTGIvIj
efcpl2JR/il1nPSSOlIIWKyrHoQualSMgKJCahK9UU/lpjGPAuKaTtHyxSXWrQYIi8G+B3h2Wtvv
128v5TjDGgA+BVvQ87rLipJnVoVi0gu091uvfmSrRpio6eECWtsvMBcbRtbiUskvUkHMbid5hkAD
Sxdno3ytly1WLzyNgShqBmbEWgiC/wpkvd0wkp1M47isTMFtBfV37bUVEngXfW4xzQR/wV2k7dxW
J4A7rlAQSjn7evjHarCyJ+SKvM+onRCFzcy1SD9e1ebLFEyiCYMCfyjVd7fkIYXAbaAfKyrxdXvv
OtFZeKMuEXKAt1rsS0JPoVIIdtRLVzDaw42ntm8P4jzDTviAKalGAwaNsjbh95/X6et+Gn+fu82y
CqJNm7liozcf8QXUe/aWkICcBrK43dE64FtJOaCfE39zAIy3SW9FPOa0alM6Sd2xH0ge0MBSsbwz
PjmvYL+ursqshzfExCxRZlz4FvGBbNxfWDq2+AyFpXLKd+llyPSnanamVurYYb4RsJ3U8Gv1Xfkd
ylMkYe0jbeLuKKLYDVHxijv3Ed8J+R4n2Gs8nI9uCA7DDNsDxTrX9WkhnbHdrKpRVs2OtJAKgDSn
cfWIMAAnx8l4qryUSi6y6L/+Gs8V8Cp2MbgdBVwrTN8WuYxOLvlkBo7d4sXQZWA0IfVod9kj0AVw
fO/wWNMcRlQNKmMFY6Q1MUBCWbslWqXoTLut8o4Y7VuhidvkfEn26PafNW9FWO96BqcTrqFPstb/
Qh0gdKD54vB9IDdQq4WynPl9h0Qi3BG53Ngkmv3Q3tzSOp0RaeS3NHdJbxCGldX4IlI3DyXh04o8
0pZsXHoyQP+0BnCb39Te8RiwO26vqQhd8q+oHLlzdvEdZUJw7VVdaDNCMj5/2qDe/mtMHHN0FGC9
0Po71ILfraAZQarBLxKleJxjpkihXr6zyxALdThRuKxQA1GdgXRlAVKsqWrFJDTaN39nwJj+lQvp
KHQrCg/f9FqdVHux+dML2teeibjeNVZDS+ogimNCcsUNBUNYPN4yEs2umszvxx8DUmei0fCm7vNO
jWl5xdpL5DP8MkBkEenOfH9QYLJpgNCCaiwBrVqEodiN3zaCUHj/0tX355vFpgojPGaXRloaWbH1
yqmM0s8h9zHN0iGZGnd1hdxkCpkSnai+uxO8kZ/7cg521vsOpM8LGGd9YKHQ/Am7KC+jKYTz5t6+
QhGS9TBG0MTpavn2qLO9JmuCmKT2O3OcwCE89PZeU9/o2n/KLkDeX3i+H6kRk1KH3LhTJTjJYFs8
3CUHI0gH1nahP/QuxrnoJparUcRBVFDvuYcBhPoIhUX1s2rpW3mStZ7ENsPU6QBBJj3IRV4NM2hY
SIz/v4JUV+GJ+ZSYQIG8rQyppVXoGP6bVuiypBHH8VxbIP/BtwbzPUYTdvfjQ9dtVP1nhG400PDg
Vr9udd98Ebo2X8iibtEJKdu2mwRHFoIdzbFPhOBFwvce/wmVlmLz9xtAgNIaSYqpFEZgF1p7eHRx
9JyqP3R9JSemUdvzlYMuEyDa0hbme6BFxjF8FEajIP5xdbjCxdT2YiNVmmrOHJJ/+lbLWwOe7sZB
xds4s4hWRMI9uLAr4Y+OFmlOeu6KiwTbCjuhnH6Odhvr2dhuRGELuTIYva+Ds1Z9syRiA1UeISFt
L2JZs0bpa3QfMpzPB0oIo/D92BNFmM+e3JZV9gPvMkq7NKyZjG2KC/umgUwcYwgsxKTRH5tFBGLT
wu+UQL4byWZ24RM/0z7q6WsEp4nD6Juj1aPYHCogo/ClLiQdfDZw2DsrPr07SKgPK53KGXVQ3Qz1
8YQKey7ToCWocwWaeacXDfGGOAqkpnJqrdlhzVb7BUUunp60BEciVFJNX2V52WU51tVp4k1pJ0r6
XCb9S0+y7reretBn2y0WNqro8V4dFItdAGa1DZ6Ka4KiUu4GLapuGzV52+iPfpK22KOCBrpQ8sHK
bHNotQ4x9TzpGBvxR1XmnC1ZCXorQparrhKxgGq1A1f3t+Sawv0UDnLGzzOHl0YZY0LLqdEwhvlG
rDjc7ZOOykU0Jsect91CTqAOmbRDJN0dfGBYYT171H4R4vQR2KYRt0gWxRIoNdbaBsksehyJdr7S
unVQxB2cG7L4UC3wwQ43W0ZxvBgDFD1IclDdT6ABkrGMN9z87rW8ax1SndMpjuxA91wkFi4cV0tH
jwC9SeTPB9JxXT9ObZ1tY9fzwZxNKVenPJPzdUYNPsKYKxsvHG/VTezu5LLU2tM2LgcEjBKmwn3D
LjHEqM5VLS+Ytq0RHAlvsu9wAzHob+6zxx18auKHOfyv3Kh07+dmE6g3kg56XZome4/8V4mypNpv
/HMARCPLMr2ceurbp0s5m71y1s+54Aus5r9CqmiTXefBpJWRAwikDC3BrDb3GqsNdgv9G6g7YLAb
PsvW0FinTxsCbzqrBRVbaVarlHwZ3QaymZ/16F3zj7V7i3JziydvjDca3HZnR9zzALVGt1QFofN1
4itPDIthdqoQlcfl4PdWccraAPS76pkvkTOMQASUG7/MPzdCGE3A9dZNZEySXOYA8ffAGQe2OfMM
YmlXPjzJSj/0VztBJqGTVtS9JHxSoBsmhmr/qcYuiXu1MA201aoFuCcgdJYc+obyAq4lQ60KHKLP
TAG0v9y0NWA4ByPCOCPnxuLcuc5QSxTaix7fnZ8HfdLgPsZsKojnQeA1323QMtIbSlBymQnhCq8+
nWUMwzosjpfnnVBt5yRxUglYzwwUEZvh3s54oBUYGKW5ACG+1XHexUem8xQjR1qrHXhoZyZ7WgTN
oYue+3uTQ2OrVoGn4HLu7JuSbWGxWydw7XVp6KfGv3AuJyaJPP0tD/q2LDIdzopSTSQsBZpEA8rN
CR2ShoBobudiRym1iWSxbQg6S0XvImjQW3AG3+E0UGn1yUGPJ8BoLU9JJmz8e/iZ27rVWfMLs73w
bXOjtWiyYahxymfO4rcWp2TkKg5/2lRpylXbiS2O4pHmIPPgzuR2h+BQCwo+tD4hJ3ypN47/wF+B
okLuntpRyjeCiznYHueslv0xqyzZtAKdLxLP5Uzsh1oR1mdlzELPMawD5C592K54eG2y1Y7qOGSE
n6SbANAeWXsUp1K145iYu3POuUh4fSQzhpN5mrTpPTq1vBlwAuVPMkzeRPW9h/6JCo90lKylpERo
VZShUJ542W8R1LH+4A2Q1GS2ly3fu7HY7ljpijCMdm2HTxuRVcPejjnWaOhHN1z55KirQYPPqqOW
Q0VEXPgOfEXuxd+FnvdW2RUMU526mgmkfcPtz5YLdbe9dS0vMdAXJIMJmoAF+pQ8ZjpzCkGugnt8
qwLpHXaD8ahEVZ55g6nA43EBC1lJja7qiZPQPokgEp5k8ygrwtC6JIbpav5ZuhXyW3YUJuy/hKm3
pTJIWy0zpT0NlWFCJljka6eFghUxZHzsj1rE3eWFHoiGr83QEYM4Z+dWfJ/LxeCl7UJENO6oCy+S
HxosYTYpfmyVnwoZUfzqwCSFdxGHWIY1/L+5phF6N18+sliBVJ+m0rYFWNVANVE+VZG5m2TCLAWb
PbQRxgnMj08yF6qhJnwaH1FqIe46iea6DK90C8ZZafAYoEUsPpwm+Wj4a8xhqj9LmigKXAWR3xyd
y9BunyyBhZwYICh+ehG6qdlI811CRE+njsxk+G12oauv1Qf6aLSnpSGUn4CFIXONbPaWvoVopfma
nYAd8f0rm1/sFvpUGacuEhh4Cvr3mtwkCnYu28zwVSnT0DcVScNbw26EoMCuI74JpKbfe4SMKZnG
FnnTi0MAaekBoRyGaRJ99qtbleEUJMn4WRBZYu7o41COAKcu8nyor2ta5M8cdI3VnZKxjbnuwFzH
za4YT32TLBi5ntfdzE26Q9HuCeKYDMSlDX1j9FKga4WrFE2RUKWNtcvM0q8+rSfMlbB/sZCH8yUL
Mhod2KYpBhUGaN2jrEb9Re6bnZvNjzg8KY5ZDLRPGEkXIlR8nf+On8Ww1Zom1GfMYaNvVfe68Hjn
ToWxwGS75yu259LQuQbHQ6lubtyRrlBYRzB3xAHmPgBHckvUtN16mCua2xmx8ebo8QdGw055SvcP
07xGxvd8KB6BXW0JMo00IgoSxW5iGexp37VsCKCwTYWv0BemPZi1/gtilXBT80+gW2N2FgkXnyNQ
I/W2qhdVQh9M3K2SzAssu+409wLnOIbAv0+ioMurhGvuS+gzmP4UI0Zi8Bzt1v5NtMum02TaQWgi
boVmdGr1NqWpixFL/lLpCzQ3xSHKeNnU26eDor8ug9dexGF2oxWW72x6miB6GoM8gbT72BuPT0Qy
RjiJ9mexe0zp2RpAD9fFnEhvYgb5qSzCpI7yTQYG/hSoJtzAwELK0q84t/BvzvADC8RmrAHiAqfW
s3HpQyuQApri2IV6cL5ux57PTT5lnzVsOBdAk3BLtPYZVz03Ynz6td54QrQAvYF25sGgqQ0Ts7Ni
lrZYwCA5lhnrcFSd82jLIS1DAwsQhH8/7RnWEPMyFQ/NIn2af43u2YEV91PGiVaINrxWGWVeFDIC
vx8ReuFmCeIb47KJB46LaKoZ+K9zt6gAf4FLFIC/ODvkDIJUzXBQUJ1g2OXRzfVuRBZLtcKwV1BD
TZIr+HnJaID64fxZi1GnDycvFkSa6KMAMvnumSSpObFPD8A8IWV36ZKPgeX75XT0kInPJ/TMSFlk
cfzq5uH6bgdA1ugeW1XCMUln5A9pnZkAnCqjr3FnOnZFjfVQiWy8qoGzlS0hz004gNqjqdKh7xQK
SxonlvAcJGG/uNohFq5Xpvm3XnDPw+20U3WkWz4PVqgXq6oR4TmYuRO4ZMbi7vlxFXoIA4y/f3AU
skBzXvGDMP7N6BSBzf6vBwEnKb0bJEmT0OMDXdZUV24t8pmbpHxbBGYihYNn3GI+pz2QWMceZ/KV
XVMmlXYQjUetAjT0pkUQB55dyz61XY7UPgn9iWjZ6OtrPguWdS/gTMxipQFrH6WwQ2DtU8kZ83Om
IYCM9GNc6dX5+/g/EAkvCjjgchj8Uvn6eJW6j+Ed/dhUafZ1tL25KejSpBoDg9/aKnJGe/rkn4L/
ij/n9oWo3Z2IkkIquZrKJsSivVvnkfmMCkSfbf+JuGWZR9Hfh+e7T6trSSpecCQ8HquXJpfzZ06J
bVII/G641YdabL+cQDs+C0O6BqLE+aeTVWrYPfG3itC7AA0Lx7kPh8OkA4ViHddY542kb6ZsjKMl
raUAEJEn6htMITd6CSCPdDSoFRkbadxLINOBhb+wUpebCMjNAGgP3rY7sJP5PTYM8TBDQnYqVro5
/bv4UV05DW6J2SqbQf12z6xV5xVVvYhQb3EEz+EmB3GyNZ7vs3aMUUe5apDy2ZKR/KlokZBCgVPs
qAVOtyCrUtdpvzXYOtObdNRvst/xTZdGbMniAL03OObAfbLbiLEmCeSqBCgLkFmJZlIoCCYYh8bO
o8xf8TBCOPTXrr9hqtlnCfQyjLlxGuiwrSU2xJhJruJdJB3ZY+AB1k0uMbZCmRU1/+3vep9FgVjF
jduOssB1aSb1MIRZkqYHBgts4PHLbaqhezdccGvbN2EA6GZO20DxQH7S/01Qo/FBMaSKFBTDDzh/
a2gwpdbYgVShJhxpss2/Cfzha4a6AggtxDBLldJgBWLQjOZpDOXuOoo7YlPjEDjli41p82voOeVO
SmGa86ZwPLmSiXtOM9Owh/QYG69o2oIbhZS36jxAuA7TYzbWwRsnx2YzpjBZc+kNtfAbXo0vdeqo
KFvqZ/ywKqlqvsbvs68zvcqxyRL3N1EaYGzf64NJs0nZA509Q8P8M4MtFulr5T2fwkQqSFOVGSAg
jMae8XDWhWIasFMLcfJ4DvVOjZfze4+ppOlKWuzZxBfSeC09R3+X6+OLSySIxe9JrehAZHEkpGHZ
ruAQdoc78RXrHE2ODif0Ltx85DCHwz8UlKXIZWbeenLxcwsYrs5MtCnHlQk54/kKnZOzTYDiq91p
hjsnGyHnweaKbyoAA5ErUG1s4xPswOFgDlZMmKVT8XnQ0eXlS1N86mAOrSvu5Ib5YmU4PJ/aFTfd
C/Pn1V9jT12539kzap07RV7IOw2BOZXylJIeRgYBTTakUOwXroMpOZdCtWDN+92dnhtt4cJpVapK
fhKOxWBZS35XG9TLPkzO5mIVJwyaCnl512Xskfgaec/SGAMSj/ujCo4C+HshjIv8wOsQrHAXZqpt
sFf5v10YKNAizAMvmmWj3jNDKXi7Lv8d9R6Yi8Gq3qeZSuvLTM+22JGdDJADIkOoBo17dchvIgCY
FG5MqCQWB8fXem0lPWXzirZfYLmY1TsyaDke6MPDuN3GXYyNddoG2hCTsh19byA1L2yMystNL/+z
Y3Mh0MrMauI95G0h7lFz/HJ6wUvgER7/6kpFrGtzjfLFXB/aYcCfd87igKFUtysYFvi2BD1j14GD
wB0UhF8yuM4pMux1vM6fxYXSE8BBqbO8Q8Uj4J1sSqxKjcR4/twfV9SCS5fd8Vzsp/PzvSQAlzYW
tu/BqFPZrOsNyl7gGtiJT3ZWRi/XFatAo+EqxbHIf6QpOAYM70RjCSWIVcdMl2EV78sWiYmhtJJc
ubKvDgxyEW34/0TtKlv2qekCtPJqInBofHP1+xN4hbpXR2BTq2Ox9GkFUHU+4tKsqw6nEc992S1e
OtDzGwNh8gZuSqTSZ+plbnlRDd6cFSC58ssf6b54Qhi8Ac2KYCtNiFdIHX/wbF/8bMw6ThqZwFqK
tHOnBMQxwkJaMYjUCY9DMgwHjktA9zlMYfcVW61dCNGzigs3C24yoRYMeerXssSSdzirx5CfGY1b
tr9sJsXoCR24NpwoUrMjx1N/I4K+ZsYxYNUOBzwPUwXPWtciQYOxKfQb9pMzU4j6RamBd/2ZPlbi
23ukaMCDENAcACmL+pr+GUHs6lfBzixk4Dr3Iwg/HNgH0jQr8OttRiVpf2WtRwSojbZTZJQMX8lL
08PrHZsKmaqJhixa+asNvM4gpBNx1HfSDCGquU7tex1+KHGQZxI3BWBMJogzHTRlpJmMLespbTbF
XdqJuIP+3/R3NgvJb0/7NxzwZfPXtdKuogsa4xcwYDuYNjYKiE2LuUhTCyOBUWgvdvQl01uNts67
9K91MbCe4t3xg6CqaXSeUBVA+V38U+Yt2/nPVpjovtjv5eb8TX3fx1igd4IJ5vC6SNEP8EWeS400
mVb+5YzTfBWqJWYqK3QxtyEuxWz2cPmr+W/bpW0DCAxiCtlS2uL79B5UjTnsYSu5xql0hGqfOvRJ
E/kAhIX6gaBoe3jg/Oiayp7HnQMDcyM1Myvm80mMtk4IkSmvf04QG/kkcCCfVt/A6hCkh6jbegZm
pk71xIlpAHoTeZ+FsdHi0P20MPTFxatyALfPsFLtEnGI8PNJU3lynGWLV0sxvNCwSj2YEg10MohD
HnagcE5V8WXH5gUYTWn8FzLLM/6LwS3x2Nn2p/JUPrmErxAi6l8PAaHl5sav01P+8mzVYM93LOmt
Lrv4U6BScMIjxpYYBDfo4p0WnCiDgcfo+zXUGATjeOjAwd5QCA1dbVpKZ/n7QPUTlbxt0NWntbHn
C9OVuKe1kiF7PI97bJjnkiZXOyQf8nIldz8viqpOb8GeOjuH3CbMSHOKjKIIJuhbDjYdRVHUTjtQ
iWX4cnsD1cXKGLR0AAANfNnGwQh9eWbzYGVVGXBKKo+Dl9nuPEt9Fot+ykBCB+DPsv+0Z9jamROh
TKBVN7CHRJ6R+OLoVzgl2ERe3H/D03gDwSywjervS6C1YLTvm6Ytek2pL0hMHbZCzhMu5TFMHu+J
UakleimCEYqgqOoflH/VqVWzsFs7WZ0JYtfgDdXd0ED4RPj3Fn32TGJxzVJxUNtCFk8kVU7WEnLY
sH2x0oyYdgNOyFf73O0TeKo0PPumqIt4BE2mZqidMYXdCvuAbwQQbOpiEF4X/yMoilWL7mZmz/xY
WNCG+OFtaTkoC0FRm/B7DoRL41IfXfRCCsy87vsonxtKHE9nshelx6QGskY4cPG/MWPwNQfNzd2r
koRMFfjb8HjuyrQxrd7Zz6zG4jzAOAbITmed2PftLsbdDO2h8OuLLh/lQrKs6hyMx3HK0k2GAKiA
B5/9Gu0JXS1g5y6pCPkZ99mQpy4YwYFtXFN/kp3E0q/DxHRyxi8uIDd41yAo+eM9IQma0WlrbgnO
H/QjFMb3PwqAOyjPWMppQVrJn54rqZA0flTcw3pfsCs3mBgPs/Ut75Zf1999PbpbSbsa37/ux8I4
MoPFOI72Pg76VzZMu+qeivvanIHZA1G36mg+o5ghIMPJLMjQ0x96ZijVwFRTASlQyB3n25TyGKM7
tMXmQyWSG0cMKfuoBXN6tr/z2IscLGEJsGyT1csVenTj32LAviaIk1GnDPOzQSgK60t3khc6CVHe
SVwVeAd2aHcbsO9NZ0uUNld1fUevirhdgwvG3vXw1XLIwOwspt+GM1XkHocDWs8th7PfB1lfZsce
Idi3mbkNJaDqm1q6jAOPlO47YWk/Mi2uAe3F0/jbbysbqBKLZoFH2nWGG9ZQcUyOoKeJ+UEX/Dko
IvFDT2NwJMHgagvyszCdT5Ns7vvwIaUhanwS//RAilbXJVzZT6W9TXLZH8LIHJnmls6Hj5bsebHb
ENlDR+LdvwfekP96SlEw5ED3zGtTQelr+X9oGoDMiOmh6DqiDXveoZVopGa/A5ZTZLG3L+bF4IPM
4ZFOIXmA7ZJJuNi7NTIT7u7YeqVz4z5oWTJZWOIeJqv3dFP9wtvqTG+g0lzK+WkQkspC4ENwjCiC
/gydzV4FV7hOob7LffcJsJ5iWF+85AJfrZl3qmV5C3p4v6zNn/3l5HqRn8DMDuGQOxiJIPyL9QRQ
9qccU2Yb3ZxwwGz+ejS0dxQbS19qK+txhVF0n/axqvtqBHB8gjJJdb7fb8uVb39kcO3q4iwGMHdu
N3AyJP2sf8dETv2HGRMiWhIoYeD7e1Sv8smGeemHTM0zLO1lq/lxD1bnBIQRHrRYL85PuqJPYxOg
KFJl5uJhBjv68E0i4ax2+1Gx0KyIYnc3hsTQoqumZHzOz5vE0opT5VA/Nn7ou6YaZVYsa8BEepPG
5csJRH1PPhfFP1euadNvx9V2XcDIReMjZXXCturz8o7BBhlT+WSQ392GDr3D7DnXhfrHrLPT0MlF
lK+Ctn2LXAAjRfQOr4aLtJTjnD6V0D6fdJGt8cClqPDlxnw4Q3UNqUIACRuo5sMcmWWqAZ4y1Vx0
dX+eI0IaJTm22wS/XAyMkiJQkKc310rUbAoyf9TDV6zfjYNPmwimPkZCPUB332EvymxIG7fviaEY
C3cvyvonmk2VNplDbS5+bB+OeYmwBhHXCnFVyFHItwdaV0XVN9bs7JT4/csk5qhrtHXFv22VAdvD
HNwbe9edvk3YpC6w4FypTuGtHBbZ45yZbHqwUV3zM0E4R9QpLBUtOZiMny+/G4mOupWyWiYpmJPC
v3KgYMgHGqY0buVhasy9yKV8gXCiIgDlFI/w7kL7+koCEs8Aqs1VcNLgDedFE94fUvQaA1IYN09F
mlLBt6p2lTSZKYvzLjENPCzZ2gfYkAGuoRt1+f4MiLBBDKciI3mUb9ZWn6wkYxcdw4PVgPQKdERy
G1/EZMau9MHKMVDOi9bwqR+AUQlOHXfmCQ5oGVi7aQXKvYavwQCyWtYlh2XTJ4HcrfnzR7y0YtmB
XIwm+lYWftTG3Q3MlIQljxlWHy0v9PtrHAXAsCYiyNFgDTtRsMBvcANZbW3mpw6gVh625BulVjGW
Fqy3Wy0aZe2FtxApZsHB0ymLIEoZex8mEoeFJILKWtvMZxR+WIdh3YkjVMHMPzbqdtR1pNcdp/uu
f9KpgHe7jxDzC2py8oG1Eyp5YJC9/X7x8lwOkSFzJhklDltdF+GRLUqauONo6EN+B+6TeusaHd1t
8Lul1JxLgAbTwm0VG0d4u+Icl9zHkrgbYH9w48y7wz07q/CUEy13kqosKRNbFzI3THttFFjowBT2
2EZWLjdXxkuS/7xDCDSi+m9tDv3FNdLnym6qxkocUEVNjUoHlqWOjdDOBlnWRK8q4815buYYDWWJ
YHwMfpLcpYNLb4ye04JXz3fPexiYDRnlnz24ez/Sixgn4mGzZkyBo2Fg3TtJzEnH7cw0/X5k7ria
P6waN9pPgYlwpcn8dLTFsnIlLctH1kFx7CzlJ4J0Djc251uY8Vw7CxHvc0RM00e8MTK70Y2a+lQg
ZPJVkoly0AlaRVGTlyRhchpJ+kRiEIWenoEM/VUrBqfjshysqgmZUdhkD5cXryaqf2gJdUMr7ebO
08+NTyr9ijtHuczWWxDBTnjs7goxn9NdKkBGFMMqBSvd46PuP9wTZZjqYlta6nsHjBPyBME8TAw7
wtpiJOxmCHd8T4ncv8fVHvbA/jRAH3O+KqbrBb0Hnn2K6alIHvfv9dr0G1sZVlBQohjdn5Xy0XEg
ZAd+ibnu9XXpwGHjCAl4qkJ3afBE2I/9cxShigMk9PpH3LD/PPbffHY3nnTd33/o30x6v32vLiID
N9hZKCB3lL1i6hE2h5YAJ6oqlsrzZ6LURBn4b2MeeOOG8ty7RR2GjSiWIKVwG2pmGfmuzJnGblde
ZM9SxDFlh/Rk/aTQvR4Za5G9vpeoYojKb/CMu7DEmFn9/M04j4K2URSaMAyVdQICUP3Jc6qZSTx1
NapZI4UnYoGJV/PtMNOGmSX+Tp+CUkUw44jM//RScYhywmnksim5lL9IqMYtIJSF2G2aG5+nQgRj
QcR1Dildd8HanrfjCImlI/VnSgYPRt8BzLp2qIh9jwlKwguIINAmYrgA/QDMCC9Et0l+O1LIWgQx
uSg7dl2K3gBhOBHFlKbQo/9GyAV1iR4XeA5H8KcoNEYTfN2izpQUVr5VaudZyXs/WPXgeup0v2hK
zPHio/4qZt1Mu6WYlijt2sbpI3nc9aUZMHvbq0o10JqY3r/xRC/Ivgwpm2FgK0Wp2nbVSJvWnPLk
jv14C3FUO0oDPo5JGu5Kvpk5h3WnsOe20Igd5Pfwqt6YENBOqiYbDW3gvbN69ARaqR9jpTp1hGSF
3eM3WDgJFUVnea6KxuuIzsXm8xWA4ykKL5h8H5kGSGhauQlqfP2GuWZY9DYX8jwenbCRUKr6Xnr3
a3e2pB6mhBFqkLiEEaadCI6WAK3ZiUcb+QVAtuCqPKOfZMC3NEs0vKiacb0r2PgZXAsiQK/1+rAE
x25Oj1kNVqpPmA7h+lkGrNFHbjiSqo3QlGpqPOdvUaorSWYkVYuRokFCoYkl1W7sXmK/EXju67EI
UA9euy0wCNTzTCXckN3p3ddua+oUVJ6t7dhlYks0ykufoktAEJi/ZtcecFSzdVnifuGhybhbZiD1
1pdFZJEhhK4CN/xtOUmYMSf9CudHTG8CzHpBq88BoaIPuIZHm1W36UaR/OqEvrbSyNpCGQ6DzQ8A
gSRG5sNWDZfPxALBR1kdxO+eTVQfAwgRdIEj7mc+ltNQW54zfWmUVzXBiZsMzDmtFhDBvqgP5jyI
M0pgeSVmEUPbxImCYlAan0ten8Y2VGww95RKeyHaK7fS/PUnFZQ9GJiBDT8UbHk9Bf6DGdhyMUbK
KpMhY8URz34QdLidly4pCrtD2V4dO9TxKgThymz6xBWTHkcVtvKKm+ioZsvdfTHrpEibEz19MiMF
689WuNnXY3KUvwQOERgI3fmO9irYcuiQXmOFlM3Kl1IAL+IP0khemAbNXazcdGWPrgj3WTAvgaQv
RoadA0GI8GVQMCo50e6+LF2eZui9Pp0dP9XeIGp8vCyxWIBB3tiJ/cWD2WwWvy+ephUAwe0KYtGo
dM6LgzVRcIYcMgCoss4ktTKRXXBsbB4iwi8cjSoK/+P0xKvNhuP2r0w5KzGuFiwIr12X8eYOKKBi
0nLHEmrrFbP6xJwIqjSHntn3/AHQ8VsgGr8Vsq2/JyPrb6TbRtQYFOmOKl9p4X1bm8BdFkweyRS0
LCP3xiH0l6b5hoT0mpHClBg5BsN//h20rWigoxNxHX9RRASiVLkKoNN1yl4BvC26OKt/FgBdSnO3
GA6TigE8oVMxT3Sel+EXe03fbR2xusy6Ged3csmfV5O6OPvFRH7OpnvblQzcYCAGZ4gxE+hAexin
JjXcb571pfjL6Uk5ZVhK+3kmOhXlj3KWPr0I/cpl/l2t9xDqaJjtOCDQ0Uyz5vkt9KS2uLg/YuHK
Gfx+c+NdKu1MUCun3funMrP9pLhmnDsCs2Vl6D2NmUx4UlB1VXLPV5EzTmJvQ90nV9SBN9jwnm3E
ECc6XQUhKeZoy8/G7boKTrMSPVFzTvHnEj+ZSeHDNkRQZG3bWWGM1qpewGlhMgxysp8K+GCfUTsC
X3zh4/bRzLrKZu1uWtSwnxyiCjjbvRSzqIhZpPu0QjvqVs9aHuOMs3/Pj+7MMeQuIr2az2jUYENP
selFWI3pxeeYYlmdqSTa37yXBwbjt9ONFcn65QJq0rz+6zfrZ4naoMhfFSDBPUHPrM1CwhYhE8Oe
HBsEgQGIAIsHvSjZzTUnqO9FF7lg0vbvE6uvfUflZMARzRl69ejDIAWDXK5M+kx9NHeDt55tnnHj
yqu4/7TqUnQAvm1DNO1H3WFO85WNkZTR8x/LzgmJz0dwh8XVSUNLijvlGsjAt9D186+8mmKwkdrz
ALhdoxKwR4qLvaZyiF8hugOdaYlVt/IucPXNUTrBG7tR+Ud8JJDQ3ApFpQrB8ewOFGtrOrIWUuku
zkPjncaV6x1uVv4OqVzRN8/04cLZa0ELFpr+eOSCP2K8PekDvBYFOfphBereDtE7jTAtxz+DvHrC
aVd5WozflY34lq/kc6eN0D6hnc4AjWqKS34UQUf4Ceda/AkuBV0xxNVQjDNI8kM7CTZ7x+akxIE+
FCqP3SoOrDHMnYRclM1p12lwpocz3kGM9l3e0CQviJU9p2axaUpFKYSTpptzxuVUAApLzAVJwuNE
CCpPx5A8g30fWTs2gGMYvgsDOV2+7tfdzUJ/FZqqTIOOS+gqwTEiYqq+9mnY4T4DdRYGMlkXYmEe
AeItxdFPIc/HAQ5EVdObEtPpiGPH/M8oHAa7lICp6SEbgN42qL2cr6sfaVG0CY0/sQEC02T7jiTs
WREW9w77ss7oTP2DxHawInhFqqJCPUJL/CKR0Y43GJOnrop6NNxcuVierG1YDSdXZGVSc6P1BhAt
UKTRxTqO6i0uVpnbn36Uy/ya0cPTmHXe0plnIacHn3ZL9ZueTeRbvIbDPPjYe7XBVxdZtMrs9CHr
BCIo1oIAygtOTXOTIS/kQU1SYmYD4zJc4yYAFMR6Tmat7xf1UfZpNvu1FpFtvYrUo1lOSY8NYIQJ
2d6B63pb6evOlgTgL/6zg4nWsrDjdqjtcZxpN30C6iIe0KtcrmWDjz6iJw5FehqCe7t339ChjZ+H
FvfQuQNE+dEx2tbp4Qdxd/iVFNemNRpFzv61W780KqWvnxAcqHggaujyegHVooTc+1+hfKSnoGvQ
ieR96lHIZ8eM4mI+AtjqI4TPat3Gk61n7/hEuYW8aFRnGEQSgqglaKkPlkV0LOCW76nx7qiJxed8
HsvHnH2jzPGj8tdtqmmvSRkOHO3nvpwn5sVEZEtO7hUB9kgCEHhDMnjvbhJelb9i+cx++pQjK9dT
NUuyXf8Sn2GfjISxVFcNej1uf6OjLPK+7NENBK2BMt9oiFNDeIvhayQLdcTTku2AUJHnqCwSRAC7
Cdc0ea5WYqDPMfMXy7CQuzkf+Umxv6m0HzfExpw0rRl8W3+zgffqdo8ZRqHcA6J9z2KErpouyKt3
+spHd2/AhT1E59HB8hcIyeIwJ8Na1o91MvA5T8PANP0z+HWNIEfo0v+zxbFivM2/s2D7rLWiVXd6
8wEQUTOQIoyJJKZoH1yU6eoVBqhV6ZA5qXr7CDZGGhUjNzaOo0G2bpXbyk7jU4e8oFoCHcpTqy4q
ob2tgNyKJzvr8R73yYcFd5/BRNH7A80FYtPCePGehTD07heHO9Eu9Zlz4tw5JGrsWkFsbtj2+s5U
ux1QH2qAjhxr357wySj0qsQgA6q63wEgY6Gz4uvC4R5+fkHM4c+gQs1GkJQyBhN9k5tw1jX41a6L
z61MxH23dK1bNq0MprvX3wOfMgdzFq9GimwkT/BcsItQjQ3ZlpZW7HZd1+d2S1jU6Bgr7Ce1aSQQ
zjC9l6N1AHlMKhaAN3C7zC2rgy4IP9EZvcsLxfvi9gNLw7gjNYkx0bw1wVTvXkLIAva698Y0RJmX
6fIWr9BSCEqdYchMWU9/Pqi9iD3XRhWexj1QqSaBF/WCS8kYhVSoMNXlHNmpEqf7eW7j7ydJfblv
C/CpI7WEzJ+fkWsohJX1vAvuaAPpQI/Y1E+yp83Ci44gU1iABE0eIPIDWL5bYtMYMoSMzIG4dZGC
KscrvRedQ5/cBvR/SQWyRFf6Odc3CXGXFOM0hf2G5pDn17idN/DeX0+9cP0vjwGjGaq7VrBhKTb0
D0Z1CJKaCmpiNA1Xlnns2MqClAoTZWKVl9TXTvCb0KSnOTELo8Tu3zLnmIjqDUzbCPjD0MlDdsLB
KLrmANrATnaLPEPDmPpoyyUzj0YO2rrhCixTrDi2VjYRPenq1vrh6KzlQcNA2HmZ7jyu3uqFJXyQ
tHDDiY2rIXwdVguuA5K2eAdEvSK4RPMEXTPZTzBy9NVz7qdBA25kgNXCyWnrSOfLIagaRg19wawS
/l84e0GpGyb0sz7NbZebc76Ho15q7OyBNzBD4ab0jlC6PKBvx905ZTyZYNYVGrbI7xzaEXJfJYtB
ane1+nZDQgeVlV38bLLydLNNO3JJYE+A2vTeognwZ/jYVZUC3DsTa7i5FEmFezIPFgJAZX6nI/LD
DMD47PYjfiSUZqbQ1rK/huOqNfoQ5OIJBK7+z3zV1EswMbhm3bg8guSdhfB3G2UqTu883eJyXdMf
QpHN6ZSCJp2woTXGckyeNKEYGsGUCkvzLbjeljHT2iLmC6vXmGZto4+9Bgkjkqk5mbKCLVMTZ7rG
gv0oEMyKv1Ul4WSRR1drAAJkOkRROmVLM5mpC6TEjGPyiu1GHqDmcSxVIetNdKPDT0fALGuCbXhc
o6u+nYNuucmHJB6dGLgr8gkf+6WVNiJ65izko0U6bRThSffpo3cr9gN/TpypYUD3+yjzSHywZl2m
SmIFEY5MCw5pRvpdo+ikn0XdGMQPlf7xjXhCX7nP8uX/ueQXyhmhVzWeQmu+JXlFRANk6Wf9uqtQ
vQcxx73D2UokU0U8OtxqGKKpkZcpUx6Rqr8rkbuVPlB8C7edXz5zH32O9WYqiYlZqHQllLsWGxNi
w8UeKsodm/MkJvihXZOt2wTxrdnb9kvlK81S6uWIs8ydwIjOomd8j1Skk/U9fFJIBsaBIKs0VwrR
hn41o8TSwIx4gr8ml9W1Z9OHzHKUJdp0bn7GvydsBZpck68sm1QWMmN6pysh5YwPUM790K8mBcA0
vnl7PdM/sjTbfmcjTsfh/l0dBFBoiV6yR/3dBSAJ+7bgKRbZUxligPH5PdL2zrDgIgiQsrPwIsnF
8ENf7SN9l8DJvkWhYG5FPq2PJL63OaV3/Wms3RZvOTxApuaK3fPWPNQVV4s5zi3inD3mnNpbhr09
CN7r34WKvplaWvdS7I32EeC63Bk2+L9x2ykuF3sxOupbd2rvVzzZiFYwT2EK2Iy0yOk7LVqblEwn
tQ4DHgGvawEADywNVLXth1CnivPP32glniksiHU9IHCdhlQx+DncD8oFCjoT1TTp7EtNq0YzCQIQ
tpjXmJ7hYWSe1dk5z5MkdVZ4DzQhiIdouZ0Un3hQuCop/rdPAp4006qbbxDZSsGb06EA/NSovlxP
+rZt0TRqFXkuDJT+88MaVoJLGlt/TB2sZbe40RX0Jvgbgu4QKal2O2guhOhDQz/f6axl3rGFDJG8
jz0BfAFXunTqS0/5Mnki3Mu1rqx/zr6woT0IA9kXcTFSMh/Ntmb/+KlgmIqRgVvGOF7oiPNsmaeQ
lKgsSadZcXrrX9rnqi/r7kDhSbGZjx0XqEtgAhOd5iJ2Py7C5LJ9zJk8tw/K8bAdZFkzQVxKOTwu
4YHfskFRqM4oIavAL6ieABvCNJ6g/+vP4Y9Vo9Deoc77UeA9RGynOLimr3iBTDs7lc+8ibnJDO0o
N6JUP/1PsPnzjwmaJigqMaK2rfcpyIzDKTXeW5IBsxcYEFfhR5eQrkvtPTMqXGVfzA8PSY0Stn9a
o/E2110Ac6HNaZzyriePZSHzreTr3hMzRFh4DHKdMxxzV4UVdjDwEIphAN8oH7Jj1IS4Msvwjkrk
sdGdooRcu8z4saOM2Q8AxiWeZPNmThuN+Ey57suT7DTcnwwyRK2l1osChy+75tkC/Scrdczlj3Jv
NcU1qt5Zpsw1Q/HY1JpCYeaWXfg0NDwNZI9bKhwZhWF5/dUMkm/hvjPmZ4het864hSt/JMtMvT+M
4xbXRicxezN9f7BZXWhouHSEquQUK9Ggrb2sBP5/MufVrf54WIOIk7iN602LY60VzB0MiPe7kR8B
4MNQ7u+l7XIc7FbRtkuqPKLGMrywk+QaHUM/fTQArSnZDGdhYxKLxaYWVspH6zZxWzHdCnRdavOg
vojVVtucKijroTayIsUFEYBzz0xcB/IIhPPlrC4J2mwhZsu2rj3FWIOnWnCr3bz9vjeJ5kg8xYLL
r/VIcyG22KaeZs705fAkhWpqeL/s8hHeIBC2cnOm2joFsOwyvS189XZP7CgsnXw/hwsQYbxLVVZq
lyZNqk+qTY+0wd3r2xcQ4nQzUXxlTgU1wpFhTnGB+IyiWkb6MD6KLD3PFPCFr86LiKmFKZ9gqzP7
ol/HkYj8w3ct1unNxzcSoXoBGqblS+rCYJmvvPd94JXCl+7i9Enty5TrvHxOeHGDps2Q8AXxG62E
zF8OiorVTS4vfqGnFaGvScMdUhdLFwce+hf3W6j00R8zHh+ILLbcuqQi2AhXUQ5TAfqgRv4ESaFQ
jfOGexZlt09vmaQzMz/1fION3ljW3yoW1gPcwmrQFUvwGx7gxeswtNAV5vr6sIxk1jSCFwzfJG4r
WWJUGG//AQzsSfBc4fsQd7Zd/A+zHIy/ewPYhGUNWU9taV3Ssc4zNbXMgiDNZGy72eKOvEK8u4z3
A8taho9GybkDvJroUk7ePmQR9+nDju779VT0EI0Q+/m3oF4K7ruZdy5iL6zAtsnspkLjYf1oWDNd
rtpcDUUPmKiZoT69o46qxL8Jav2vQ+nxJUM9RKe/3qgQ/BbGKV158ZvB2m9G8g6hTsLnQrM953yN
tyjK6KA0xzjnIToYvMpTsbNJMdQlDEnp9ZIdPxO2XGhxwEwPVbT6sdCk8aAowkGy+vR7cwRv44rJ
PkiCJI0rh+SD7HsheKWwtrnnjBBIT62en438m2Q4zfxiJNCqtgIEHWF2qk9M52onNmzhFvqaSwec
7zvcKPQRwfrXv5xcjBzxmQsJeYC+W4GQFyYrEIFfocnFHKuCynmjyIS4YllZH+NXl1SXDBh3nKbb
14wZNXMYFk1wDNnf7KLjPuEqGvUVvCe4NnPtOZ3xZ5+OT+rX398KzO3cWq7eal9mCz9PbMl3FqLz
yM+bk93i3WDqHOU2Kq1L1R86HRVIBfOx2ju6ps09wHxEkEDkNKmnH+NwrBfZ63HLkmr1Lf/g+aw/
/3JJXbxh/0Do/0e8GEc0fkEydoJFiPL2kdA1TyL3p5VGrlBrJKRZa/8xk+F8FOSPC66ZLe1cDSCN
IdiNb/tzM0OcB1Tz8UTWiFwIDAMWs19mMsjGJjOgKp0yzkYTdgpB42YVYCPGiyfftXAhKUwzJCRv
7UIfWSc5uD0exIs3MaJdAb8r8DKVEZuUGDRLGovAvVFD7kgQ5JSHyeKx7zaI9SpV+hyw7+8ei71n
0wrdLYlWVCnm0kGwE8x3HLuncKsmvpQRNUQr/Jq+NO7p3yviU0rKC4X+slODtklcQyEmwj371NeU
SWIy0t2Y/5bj0HMXt9U8Z1UBpF1LyxIHvFMxq0cPHV2M9khn6CRWxuKXFzhRYxcUSIbG742YhbOR
PEMiLLHX21J2bgFq18r5z3SYl7k/75S2tUmvX1R62uux8Y1bNQLTCvgDJDBpJWyzGc6mdn+kI47I
bHZ6kpHnC3ud6zctJQZl+an26hQvqm+0BG9NKNAbr8spADLjGLyKE1byxr369qIB4DbNX011biOK
Gp0MIPLcHmNeatqA37QSyi5DxDMk4h13wVTpLC4g6oAVpspd2ZWQg+BF+6FTQBGfK8C87bPYANpm
ZGpsjmzM1GiYLs/CjnsmqrJXiR4Rr0zTYB/EJ+HAOG9cjpMgPNf4M/Ta5mfQc7vK9/jrDav7KZmh
J+IQUNtBl+jmO+QgUFUuMg8JQhZqBTAVWfTxAJeH5dWIFfZL2CEl6fA5+kc0X+RPjQP2JB1h8oeE
4kt+AAKfUlNqZwP8CbhAmYTpfThTUCX4LofptKj+Bx5nkQ9HDEnOxFLbPYfB2R0Y+kLcbVTj9ZZP
wA38gsjXQdYyS1VPHb0pD97mf6Wjs3j2lS5Rk20a0/bnRHAlVAKS81HS2y358bmCeRHr1CKiwmXK
7scqYgvEP+Yfe0t0P7lxlDWpXPHSEPmmHoyaFDgW/XieEByX+218g/d5ipSkKwcM0A76RqpaL20m
RfgMkzOI2iSLoOGA5+AY341n/pQRLB2fH09BEcYJqCQRIshmdEkdV1BC6nrzht6qpVF3gTM3jeE+
Qw8QL0Vck/4EafjH9qeQpg5460kvx6BFoqR/NS/mC2kLE74oo+yD12iopePdDxaoASLpCRBFfTA0
1nh1qVnHrLufTWL2xdsguT+7TE22np+dRDipcMTqXkuLl1qhDPa8923jW5g1erfgLabcGU3xSGJZ
XMgcwnMt5CwgHnAP9NHUeeG8Kr63j0MmTdW5PKZr/Tas09sfXT8C9onje/htw+zqShJWJsbdCmNq
PTt2kN9w0cWJq0HMNqyoS+PAV0rg5IjaSU+xxhASbJtlLggOncML2Xj/2Vhr0+Zk8qSBqgdO7sen
j6SaPcgEMg0PSNXKf4byjZWBKwAUZmyqQL5L3QU3sl9B+Y0vkWnq0R4su3x6stPdALoLWhq9ssEa
r7DF3H7IU9e8LckfQwMqe8Pgb9ctB5He2RHY35vySt5G1e3wT9QEEZqKhGFalARYL0jTJB6NJuUc
/yX4MJ4jUhV1tNu+5ZpB1Zg+G9a8v8d9uC3A+5044rKqBtxOWEThmcGkQfNVKkgunw8WTJwW8R4W
1S+e72gjrEl/PVwlW/MrwhZ5FDueGsjBXx3rtnTOifvQBw1M5M7gSATCqWcyMB2utA3/CafmpUmI
MObjKTj+s/6qeLzZ/TxkhcKRhOUAY3SRoIMM0AcZpFL+HWYbEWw3WmWphRME12IczbSik51mECM2
jAafDbpjEyDFEZvuWbemNqVaRIbUe0NnKNaQS2aZ6xh4fMx88sSHYYE7C4AI1Cb8mI6sV8PYUmpQ
gyZv2ZlM0z89pTeg31cVENnU0jWfxSmVAQrL7FcHFhuUXAASRCwgN0QC6ux/mTJ17umEcy1EGNbI
XVMUmC8W44uT0e/Jl7YKZcpo4uDPLq28ikzoUOzF9eNSwL8immpWISnE+TMmuIG3u886162i7d5a
dC/usaB5Ezy2ztT/MPxySQYRwGyHRFwdlL12iUa3+qDAy6ekKh8RVv2fPlXgjj1Ydcq9m5EiGAY6
BHZwk+ywrwVDJ7pHxwgU/VUvzrYY6s8YTSBeVKDlpiXaHTp0qlnkNGa7MJRbev/3isA3CKxp2Usk
apq9Lt2s0NU0rlOFvu8j5f0aOhFD1wB1B9df/cEeW81GV8i9nIm7X99G4o1bJfhaXemjGFkzh5+9
ipiprG0evcEWgdy0gx9Msj5XXv5meepf448HF9o2qdJ9aocGPSje8+9bEa7uq/wT5Tq1yz+QCSFY
kBeuAMMt0DlsNp+5+WqPfzZH7ZMVQbUy6EC8SlO0WKWXijcRKOO5+QA9oz4LmDNBQPyEnS8IaidU
Iypi+iOqRNg68RP9ispaA4+O2dlVuSgcLsed+3y6HAXB2UiUZkaDtxPjQ4VFh+5ijCkeSfPpW6DO
qZ5YX49A/wztsipiQO+1Z738Z5J5hFeepzswcSjJZvDKdCpLBxhjEEQnXEobBRl7YU+WVj0mvOMu
e2w0wbqQPlIgeY/aynKjYSA4bdU6Fdt7z0Sb7M1zCkeQe32TunXBWN5H5MBnT7AXzAXV1fpX5kI7
3vGN5+sG4PwWMsFvmWCtMesS2kl/e6GJZyOVGXkfhdQA++tMrbhxiwkpKrELR5MrKiJwbLbuTnU7
1BpFFCNsG3CN/eqICMIZm/IYC27WP5LmPDhCmAJ6Tm2e1aujOBmg3EVUfTa+D74GFjbFpCbqPkLM
+9FfmbfLSb5qIQMXRLLH7HlHg5wFDj0rRj8nC8f8dGBfxy+fQMNPWG71irLDCDAkWmTlzSo0AtN6
P3gPwLV+Ma0CTuQIcSyc7sQrrg0qSaqcYJT99O2HXVXzpPxShf03rDxW0mMkGk/TontZq4Y2a6WP
EjKxNi+X8PaO4XYO2rs69R7CKMsJLVydIqrqXnpnzbeDqFeTeZYx0lFOp16N5g9yUW2+x8U33yGe
AmK3okwylXC20LQTDHlBHHDubHApo8J4QQ/x7+bpM3mxtx9DHQztPVtKkH23PNUPeBTa5a/VtLFc
QMKY5JeRULAJ9jhFtbT/dywqxbZEsP85iNMOrILTCNvpKdg/3pVH0pL9BHzNtOwoc0UEycXKFhCr
CXrNxvixMRbu+mD4cwd/VH2naIqhZnxyoB5qPeHwD2K9+ccoBnupOSn+DgU5DwtnBcwOo3FugTi3
h/nwksP5juvDnaly48fQhOJZr8YY8FIC1e/xH4C5kNdxaNfwktLr1SVYWRQziZVVhAqYU6hfpihX
Z9Pl7TUIyxMyqraLYxkBUlDtUdH8bgeuftyfH8ZrL1rbfzv3sS5jt2xUbva1ly4vJH165N/rQ8Cb
ek6nzKyqjOrGVEbz1ac35Sv7VJMc45hqTSnC1c+Eq8xsq1zCnqroZ0HqxaiS/6YINuU8RwuTffhZ
15IWGb0k1VMs1najKHJCNpUIS1DJ8/kl2CLSnHlBUXmOCUwL0R2fN1frlV7qz6SM9FWXfkoEhU9/
Z5ueaxI5zcmqDdDIG1Qh6FGrKmXAvgHM9/z14WukJoc/SHyLx0/dVf+FOuAvYbTrg5iGKFzoYHZf
eMHmFe2XSCmkWxRhDIivQxcUiaAJrs47V4K5fQJZj9+OPZ4QOzCRaid8kzmwhq/JgUxjQd8LhIyr
3JBzTIWRCB2TE788WLzR0m8m0ye30FoPy56fHO/p2/F8WZ8XMVJvs6n/iLrFiWpYsKDBPSoM1MK3
dGEQa4Q1camNDyjzxLE7/NEXNCjWx9kh6IAUHuE3H88UDhMgfoY9wpKQc8a+g9/eFPw+Hrd2Vz6e
2glmcLCSXOhn9JOiPhCHsUHMSDDn09rMKZ/3FK8h717G3/oQ5278yhb5qHO124l0N0G4BDapffSd
Uq9Nyt9Mda/VcxvD5ys56lc30soJM4wHLtVNcSRXcd5y7Mi1sxj9tKwJTZOGFzx/3ColNx21+oWC
/QX/LRCslvEAiI7EjAneZcTaiCcIGIEQDge1GEIH11+tZDQxESnTj/fIg6Jt0tpcglj4HjTl1sUz
n63PVNHwbZk/4UlmjXbHfFNuUUQE3emWXgwutoMAWHVGgS3+aNrk7qRg1pU0jduFRy0Wxh2LoyDt
1QmSlZnhojEBL1SFnZLo8PrK1Det7GYgqEiE/sXI47EtvDLMDCeBT7DbM3p0QZNk+DZYW9TPToWt
W5KCjfYHPQmyVwviyZkedXll16r7PHtFhJaBnXwHiBx9jXlHQyRZxa/bHB8YnzGhy4CPOjM1Wr1Q
GzBu6F3fRxysxpqKgZNDYfwhKjLFj9r8poVXccQifVQxJPuHY3XZMhyE4Yam3IKnK1X1r9cw0ry2
hA2j4OxkkofLfhkEP44y1p199AKFqAyh0YiymEuH4RYOCEBgB77YCZ0wg53vXCNvl3QuAEMSX6oA
CdGVx7YtxBf4U6KQyxmsoJoz3YbKwPaukRLXyRi3w1nZt9WA+nAbFf+rcPLZSA5W3/eeJx1iFoaU
c1x6kha3NBx8TlJ9LD9rm8KlASRHYlfrE1i0zq4Xx4gfIYAzFIo0ZY5PkCzGGzUVYquKLYllfgqb
c2ShupxOm9p8ddmTdbAjKPdPaAu4kesTvHbFjBCApHdQlzEtRwS0B6LqDIbXC5ivJhL2+1eAnNTp
FhYmzIiOPvUos+/hKSKRfAg6amQkL/9CfHbtFYg25shlyNSP97cNmBGnCNr4HWAuEtKoZxvZDjnK
3V2V11Zu7BBF2mal0AS2P6aJ3zxg7J4zdjTYJqhsQWSZ/ukmENzWrOdCiujjCdnUBTkB4gRHS9SX
RAOTTgcefFM2U+rAjogrP/b7TRfnF/c8bbYHZhCPp75gVBscGZpQPkUzOQMrWCyZFYNXhuVrwwIQ
JrvWgk40gKd0bor6NnYR4mOPgdAHPRV3BrcEeULe19+yqotBdSUQamErnMJmkW3Tk5bIhIEcjBl8
Cv3Hcy6dYg0PswbgBFNnYk67pqEXjZOuufg8fuCbqo4Y8N4RxsjxqMUfSZlBCMQPDVFZtXHXjpgZ
ZQ1gZMqH8prHywoqc6wuOT3tWz1QVDnD2U75Yxt/S7CxXDKRIMRGxtjga+E/yA4LQGim49z0fgr4
4odhtLjdP1mjz6pNzfJWiySnvDnc9YNV4frxK4+pjAg3lshzKbQjWU0DX3p8N5TlkvvI2EkiVU/D
Y9D+IckuT0ZIeCm9EIzY1hp52Q4mgoMzCbaiC0YGtUjOK2d17TIszIj1V07wdAa7z0djYo8j6aYy
AB0zDWIXZaCuBjBKbZleltLCS4WfNyjH0zbuONFNGnYHw1++s6HEP2ZyBzN4V1d1tFecU+clJw/k
mAMCabBBS+nyCgQ5BmS+t8vTZr9nKHjLNTJExvVLrSqnuN8fx7HUgmdm/2Upu62xBK1VBSJkBDJ0
54ii6cQivpUOOaL/lqBdZKOvSoa1DHZ1qFwK65dECude8AhE/dMHELFfR3ZQDA437pNO0GDzd5kb
07t4iaxHgNEwnTAFzoBFO7mGEQIosM5vGcr3L/bTC2V7ZoOw0B3jGW3mP0eAa6CPHMxPZYxUhj24
CaAvsGQAm5h2h9k7xDVkPstTQm9TG/K8mzCsWT5zjguoyHrqmJZycUnxXhttal192ADSGKZm5edx
b8w+GQf2ke7vCF5b0hPgUcBzXrEirX/avkiU7tvqplSo6V1VH2Qgc2jUZU0G9dPltVlQtkPZwu9v
DTCe1Pk7WlV5Wwk7Noo/TkqxHkEjUdGkgFlFtD6V1afaSsZF39v9av+gvZvPMOSkBKrqU5iQhCRC
LL3pHoJVAhB5N7EJ/GXxbICPXLujWPNfQjvqckDRfFGfqX1GMHivlAeeM7rXd3E6E5tvNWxqRoZW
FhkzIW7Qj6/PPjQbbkZmDyHOB2TYtHog/TWjjGxQuwdS+x7ddO1neyZ/z9svzmJBKCw/Nxw0TiFw
0bz9ecYq9xPgTSqUxZnyTZJt01F3GckVHPIZlfqfCFoanCv4RTZeDcEgRxX35Rpz08lPI5Ndzc1F
ygYESz4Av1Tmc83WS5gBbCEiLYqVZ7WxYsKop5RS2mDrof+nj/wfxJc7sesszehApnI+gyqi475L
CRFnDO5i3uyDw0jP4zZaXZWZbU5ZN4T93THtBU4N3U7B55pGQ25ETx715dU900uBiYGjqqXLy3Rs
Wa9YdASDs2bdF5YvCmM0zFHP2mF3QsTwaBvDHkTgU2OCiyLKYGBJ/5g5UcgI8hsAwiqByaiXxHyq
esPmtnsE5Glzz/eLsmvCLTizF0d2u5pl3hHT4jLzl9dEiO8nlrUCbUM6nvE7MX6i0eEH91kObvwg
LJ9QVD1Nv0BHWHIJouZn1QZyE73wJxBQknluaTX3pJQQcI7Zf+ruubysAINGh5vYMgAOI5E3vLbP
PN/Oxo1WwTRhBtrBd1+lLQl0ZNhHinr2MRQmx5P9mZPBbbPfFvrEqNOfAuZZkiMwSlk6tH+sPuS6
YOl8eBTqpH/AqNbDDjK4MotmYMy1nQG1pOpL1a+fH6RpRyxR15CD4jbQ6dTz4t+mI7L68NUMtzrb
wL2BIuvmFRaK962lgEKotjtbxMXMUI0vj0hQyNJkUiYLUA+IDHEYaRwXZA00yhD1F0vc4sNs+EIn
MQsovCjw9a5zrV62uXuhl3ZV8jqyRzSBo3Lr4J+RnWbW6he7NzBD/gf2+7eBhoT8IVhm/82Fqxbj
gVYpMdSEOK7kOMS53/nLiwy9yLhixBVAMCcd5UcU+9cUzQ1iR/xgwEe0mFsLtMI7Gx9g//y3phsZ
UFaauxf4FI2nN3KjA2JxLc5fJpCpO0lLUNXVIEKVW7Z07k7qie3ocKz9b+P8vh9hGB9xcL8idRQS
sxhElrDtHxeoEp4dA+/f7le79BMc3JwUqvAkHvOw33u1o4c9xhB01cYPftyZAEK8yN7Iimj9raT+
GTJguPUFAyil9vHXTtU/pMBAQ10DZvXKZF/uPhtbqF2W9QvMrAcyBHYjSfmrEMqJp6juBXZGxYAx
zdsaCmhSRN0mwh+XEwPL+/Sad/JjKNSDu+Rg54D7YPnjrVRi9VVqY8+LrnTLwi2gA6AqWgV89z+g
EhpVKGOs+OsHfbMHnkQS7DWHw4bwsW8W8pSDgFyLKwVZe5Ii2fvbptVH7oqK6CFG/bYoLypwI6TG
q6+B/tahFM0r2ZzGdghTJE6eOONr/UmlCSVgpfzIaAXIRA6dcnwS/TqVNtxkzbELE87lbtoGfvh6
7AMSc8gG9Z3ZEasT78dZTMgWiujgkfDaVilDtKDDSJaq+9fnNTATsZAxypPyWsrQEVHPZbZFnn8M
yfF8imRupAb8n8IWE2+qzIGswqAzI0zos/IPzfTvni/63IL8zBMLTBpUlwHMTZ1iDn9iHECkExsu
Mu+c1AbmlOjywhR48pYUn3/ii+OGZ3w66Y7OSm/pbfIbX4Euy/VhIJ/8TZLKtqF2ioSUNzcTt4lF
WSwJrsdbd0B9+WCNp6OANVbRyyFP+iq0zZvLk8NzalS9aMqpcSjVmttKguHRMK7jTc9FnFYYMJO1
outE2Lp0BK8gtNgpdRj09yt4aN1gV6aRshkm5cA3V/tOrBoQInEorBhKR7Kjt6HsjiVLtRHryPKj
AghJllsWh0uu+NfXIK9GHFqB9k5rJjfFzDnheVGj8mfxUNdHi7+XQGUAlMM/McurEWMF8lY0EKSv
GCuWrwddQRgL9eBGfQZ8CXjnhF0zPk7L8Tpbu2IeB4fuDOGI49Wk0FWQ4pKhx12J+Luc2bceePWL
eNt0DAIpL/+p/muFO8V03P1+J4b2Pd3q+gyiSXu4qvPGNfHgmoo5xAUFpQf3bv28DeIFJmrRe2sJ
zmkSIh45UHOE+cO8eec/AuVTUSKAcIj6LhBqSVH9ShmWZlONYvpTptKILEyf4xWOT1c0QwvemFDf
S0F4L4dvo12KjwE1aCF+RXg2WiVkhz8Dwdsrxz3hxCaRHOdhdcH+4AWxTwW1mBotvedQeyoPh7Bj
kmO6F+Dd+X6ASxX85oDJkjzzkgKo0mu4SuzI5QL73SVmmixQkjsfcF4fuZXd6v1rncGYRPNkfS4N
aUIgbO7jav4cRcCRrY3Zfq47qtwKW03xLtToR9N5gc5eCspnLYajKrQXxO2Ufh+eMBDjF61j1gt0
54sQ/7AjQ4RgtjmVyZ7Df617zkmm6U/iEtkHdD5RRDvhzw1zqPRb2nV7E6eCn01fhnidozOK2Rt5
tMN50z19TeEsKm2p5JI+xC8TtXx2voHPt6Xv08mns+9k5XM9aZ3kcQ6ztZbZkBSJjz9INjVn8gtb
/dqH3hfpTiLip/tE7H0hEkO1zCW48w4s80YzInVYFN/aOO8gQoor7kqFykILbq0l9VSlmrvWvsct
0A/0SzZNXSU3nvj09QnRvjT7VwuIw2Upx9JZrgamW5AXyJiKLvnBQMtJxOtCR5ZTfejmXj+XWY/s
WEMi0zhU0XoaUJAWST5PJA+HHlPT6jPMToOY4AI4pXaiNo5I03+ILdhB/GGuho5olG3WASUqHsn5
PxFqt6mtoZndK7t1SUsPro5Zc6ywkeMYHtz4HGc7H1FEBFYqrZk2tidOrbN+N/q2xzBC/E//OiXt
Xzo15Rr/abVvttytcNdUBKRAk1CQj9X/19MDUrz8oQ7Pejd0XEL8LpAjmevQgEJOmGME9Ogkazkw
4O8sfC5ZzdxOAfr/nyrDDuACkKKs5E+HUNRrg2F1fIQNI6qJiTREQiIYpOCPToKRX1XjyoCfKcsX
PZDX7PkEgfbr7YslEziAX2wbb48gBPphaneZrNjbZgt21DToNmoTVuv/+F3+WyJu+MEJMaX1QXDE
YsW3pvPqnoOdCN+gGr+SjuKW76Q8LZJBKXiJqv79kbXv5YmVKA/3j2mOkHEQ1W1xGctOPbSxJyb0
JKUs31kHveSaFz4ZKMGCru36u7DUduCpqAOvC5L5RfRtBaUzaBRuO/sWsyy03SfLbMgWjpQe/lf+
7sdbsKIgmoWaMwIhKoopHYE4dKNGgKtKkGW5ZISp33z3A6OiDnYTm71bfdClMC6pm04yB2qzxaOr
RDcBUKoThtf3lQARoidikaX+pC/A7J22cXS64ZrFnNFmyq321GrnyoBBFSEtG/dEHZyJoCPccPPD
/QO/2r7F8hZT8XX2yvR0f1MvU3XJ3vcjNEPOBzXglM+GvI1g8E/kudZFLtSdFw5MPgk84uLmjppF
oYgeUiteIQgyEJiutR4SphbKZ0LaWvZCFEKkPA03N8oHt4rMlTJHg2sqENIVAokkaUEJocqaTE7z
NhWtBYeD4brA+UHIxvdYlG3gICjbLpPAUyiqFGxXYcwD8L7Lo5U0wEf6Ol1ZryGc+X/RBDmc0Gtd
MiTUWwVSO363gl0DkN4kMValmA8Wz+C5sCMwM9SZ46yYygLw7d7xzw2DtRmR7rTBZ56pdZax5hfw
ey2v1xt3Lc2Gh8jG50USOJWR/UZCba90r2XwWtjiEhpgmt14ipi5qurqeyGUKMqemxH5lHRWLXmw
7A6QKJ2ep4MsqFNNBQYD7MRZW7RcY1CvgUNiwWEcz0nxuJnwS8TttwSZ4JqtZcgJHdW5ccIgZhuZ
waWJuGJ2TjZtoTAB823gm77zgWDO4Yjeox6OekWaobnUqIxvBBMcOzfCVQ/yqJk9cZTaaKZ9FBPQ
vmfjUrotoDgVsdFciCxrRqJ4RJNU4WoqYUaz7mL13KwBIaVfPJuvFLNDQV6Z36jEgXUQhS/t1gap
UCujczgWqGiDRcvjKj8qI9Gz48gQBex++hGLoGe+AUA9f1bC67m8xhY4+CglE0jhhebtOvzHehog
KmOjwpP5bk3qnEqhJowO1wOtKt9BEuJGL8rGaNObfrAp+2YJwkk5Fh/Vstbr7JKyTZs2wkO134Yn
Urw78ilb390vnKbEX8Vxobf5pZZ4RUTFkoo/Baua7iCFnpBVVNO+DDqTBb5S0BU+a0Fz5irX1sDJ
wrjATh/ZpLUpTwJf9XWOU9KIKpEEwUsy1GUPijUy27fpvqZSzk2MtQ07+lEz86JDpr7AoqPV/LPn
0J4Mxaen7bVOFITT9FkTSMsDg1MPEzbIWyXrcDE1vQSlULTyWmyPTTA13QQ1a7wy8d/qyl8mhFXr
cW+fjZU+B6II0h5HiX2e6sOY8Z8HU9WwN/oAGLSyKUSm3m3tphJMK4bxouNVaZj5rLBB/tE2RDcf
Lzcxj+NU5bcNmGFm5B/J+XZ30sUIqhlMPrXWG2okthGyzTIxHH0nNGdhVLW0kFoIisx/j+78/746
Y8+maBs9SmyzpB6XmD7mar8jNSGO8/7fE/7iVY25FyUJG8SKjlFFw0qU1kblQ/POeNJJLxCPmCDa
wCKU0B1u5ruFqnSMhJ706hxs9SKFKVqY0YBSw/gbvSNVKXL5PSvOjJfxtGN754W2q1c2FvgzcKpi
9HBr+RP98v3crIjwdC5/Ui2BsH6bfDCG+m1bPQ3Sv67PXOCRVnZPAUXcBF+yIbBZ//ZHvBgZDocz
QgauZ9URuks8jwY4YKFeKBReIXcLDsoF/pN14bTp1Ezhi6U8hsvyKwrSGYDHsiCt6T78Fly+ugLn
ejs+Ju+M7m+YfekWfPsI5NtDuYpD32nxNpeJsszogMImMES+OPYjKuRl+CX+lylg1ssJjKwgt3ef
UN4x6+rZjyKi2NktY/yQapygZSQHKEeIa73DdGjAWCN92rebq/fjHQ6KEc6aoc8IXluFVKJppd0t
fboDgf8mBrvVppfUWN4oxP4HZpWkOJJila+hZrdlFJyQii+s1BaYLZwn0DKWBGWQNohW/fuVWDUt
6LbNr8MeM9D9ZB5LMf3/r8ktJUZtUYPNZMtOwK1aDm7zWu3X88iXz/fUDRaJ7vD3ugGvKckMk4jD
fxTZdsTdARcKMQTpNgJ8V7ktmk6+5cR1ut6LnqX3T7rxEXJa6dCpyCS0882rTNLSKYcoFE0Y/2MY
wftXU62JeLMMOrhO/xpdydQLtJ+8zni/lpiyp7DvEDpRXzfyeNE/TTL/WpEIVi6k3MfyaKJv0ful
NbyHAIrH4EH3+xgnBJM0+eBfrwGkDPvwUVKCp+1tgjANEUXtLZLAVkDjX1MW6Zwr7fYSuKrJ0xeA
3nfwqpkpBaHXt2H3vNDcrkOKS6jiPZwqeO/quiJzmwgkV2pFvyBcbgyTuLFKgSKO/VuO6WLJbobZ
V83aWy3IjzyTkjZCp3Wl0SAwyVhe1lieYcwaUo03sSM0tj/yuziSa++w4XtsQiwofRboDJei9AK5
W/R+jAqbVaEgaYD+DqFWPzXdc0dkYqqw7usAEUgE5DxagLaLc+h0/WQuiK76sy3dvftxRzezzjDJ
1HR2ppG9FDRzwA6ta+50JjP0IB4+cfvPkpITUBBISQy4CyIIFtSq/Q06o72BKz3tsjNCuAucSOMr
IhvF56EdVIlepGe11/za86LGpP4AC/Xy1WbLkXG90t3gMHIZZc4XMik5nSo9LY+zdqtGQST77HeS
KzzpiFG8hdgT4Lpw3gCrNI8pZp+VlGgs5r5tT66OVaxjeVUhnZKOnHrG+nL1aVaqD2b8oYV9sAdY
U8ZgD2We+2ZO/p5lvd1yjtIv9VV/toTHK+DOIZuzfMZvvHqk+BvX5j3oOK8/UVrBUAcRkXQZjum0
he/gJ5Ugsm1Ypbvc0K6uycHIJ4pdEKSEDhzAI7AsetKRBCFbb/UfXFE8cxQ5XwcmhsrNZf2nwlG5
WXtBsFIford+xcVTShV1ke1KvNBXtWsmC5gIXkbK25zI5KXwgqJThDgIeN/h0yEqSuGk9eQ0uq9h
aRVeI8W87Ku+nD7nJAiWm16/MbfnQX28fXnLoY9KEi60x29RIbK1X3CZeeDz1UGf82dG1GlJ0NXQ
K/rX1WISt0eS6W4EalYeKunMOdjLETBkDOXeCHG9EcYC98yTihynGz//bjIUM53o2oqa/Z5VajVU
M2/OB6iii4uFZ80ef06k0f95Z98ZxsF9x6KH6Sid/zHeEj94WOKU1taIl669HNJXY+gQ9t9LMcjH
BFJJzOOz0Rxd452v3nFqbdGIQxOUYlA+QwNePCTCv0NGZ8Q0EBiRTc5nTA2iQagH8ugAa4pV9IM2
nQlP/v9OO2rCHjEiR8bv582BDU90HkFRdiijX/KmKori5TRV83FG3zCB0hEtPxY2cnN7+aIoowT4
9uwad0lYjPqk5RqtVFdACAOqcJtD6odez2LlZczJdCeU2/XDbv2U00xQFHcYhQQWiLvBYZER89E3
XrYiIZZDRLBTxUSzlPH3ISzOtlGyKTJtnI7ZP9b0AkGlbeNYg4PI1WknzeHIX9bdzDXCeLXQkmXr
93SplXUJHL0I6LI+lkreOTcNF2h3BbeIiPmcExT+1X6hjL8Mk1BoHLza92LRjMkA8q+CmZwiaQ+A
mpoYXyV/pXwpf87gFgbV6ekgk+PZG1kmDwvtRMJe6zaeNCsqmbNZK3vawTTBroCDsZsdVCZErhGx
/aBq0bGpXoslMi3MFikEgIibvaMXHXTBw3cbkTEj05PmFcbmxmhIYgwI5+0rzepQJc6eJTteAT48
0Oo9HF5r4oYk71pgBXDH26nV/8bu/u2jCZGNizIvHTHzCD0T6XFtHmbTkS6EhIQChrw88FaDiQ+O
4dRQJ6OUce/3qUDcHzc82+KSrXSMMpwqdpij4i4Bkz3lN0+kF7G1P1NO832POWoNcEQJB8031KmZ
m84AKaZIqMlqILK/K+sijhXk7Jj4cWUuQkyhVfeT8ZOL5jpTbtsdQvjlrEoofuipp6Ly2Vk/XFhJ
oREzd5HoQxm6E/+vy+G8UJNlJTefnjdOe5nLdQ/d1A9I/lKo//u+HIRZtYSlIA8YSIy+dQLFxiDc
4v5usD0oAr68n6acENxixld5gp3KbhrlaWoVc7tKMoBpqAcGU4nv/boWtD7uKSlTxUvIczEFSdoe
dphzOnS/Anodrb/pGG580lEDE+yfEcElNDe7CgrUHyh9ogm1N1mDdJ5uPQlwFr+JEo//Kf9pyajX
9vXqWQ4Hl4ppVerIZhFKi8q3qi8lKhnV9pY81f7oJjLpy2sELCTrjdhvA4Naj1OGmF3vdAJ63m8W
wTuoIjycIOhqZNlhnBZYuGzDMXVKlBZ9R+D5ZtyDa1TGfwtHwU1bAthynGaUIOy6+EP9rRI17LLV
85iFNdGZ5LEYNlOhXbBm9B65rBMXdyHdmGodUogs9RfA63muAURl/6l44MXTCv0fX6G3pjjmr01l
a5QZNS/9qNl+gpiX23HTupqRK/z7wIer8TH8SSGrxNpoTSnrzDhLC4t8tei7bH67cpXKyCaaJ8y5
ZM3LdzJuSDR049cSbrU/jqkxikl3xNJEnuFBWV6quBYkCoGgKjVK5dQ4rlfoQMp19uFSGz/YPf/i
v40WMNdpIxLoMp1TfFN+kWTKdv3RDfwA4Dq7aqynqTEE0Yaa2D4HwM/1KKeDj/QO/pyFCExehOQQ
hXgXdsAKjn7St9LR0uGafkOB/Plkl0N+vyERQLkG8WeQc7zSIoyOGkOP44Zw8NC750urmsYxvMUD
1buby1CZNJESGNoixMU0LG3zePOalpqquKWOmzT72jcsCSSt5met134Wmv09agyO5p6lY7nET11q
0c6TXEUmrqavyoEInbEQn8pYsTQcVsktIxp/FOfqzLS+eUYE4MoRODtHY8yrY6QFy1MgyFbYevMB
CcPDoRby6GY7JW2ynJkcKmsU2ajREqQscsiaW5RWTpUH/xuLdVXclT/tLQxLnHEUXNb7XQxOzELd
5O83etODjufv6rkLOklCeSdCjdF2iRFS4bIIVWPJ3f7l6PL27mDz8gjeblpd9Vpjr32GxsUHZxwu
L0nriBcM9qAJs596Gv1sSKFZDus/4VQedJkjmjEqD4zDFSbmmaC1N4bSyD1tUai/Hk7S/zzVgWwR
3uVktP3fZe8STgf3X9ni6kQiaQnME0A8/9gLek6TDoIC1WQBZCgLDyVCpEB6FBNq7vbSj9VE0Fq3
X59s5Sn1/n362vqew1fPTnxkKCsozVuAWdevThEkUOc0hl0mBP6mrfR5D9SaAKG/HFeVlzDys3rb
3liWVATHa89ozwrQ6i+4vUyhpBzdb2W0qNlITpwmotgrW9jyN25sNfhao51gTm4Hz0XHeu77blCU
d4f2tZQhQtPEv/F2WKA7bP2Mfu2kf7nfUvYwFcKu0WARepVWsCCbYjOYuQ0Fij/Sl0HDO8zR0Usg
RGHc2InECOLu6hE6iXBmie7q1l81jChC8E+U0T43CDvg1ZdO4DcognCum1fYpdy24HDX2N0JnUQw
vuNhn38Rl0EXA6H+ESlLL98pyV6VjrdlfmBUNSEVreK3cazRISRqCttGFPFrMdNep6dGc3c8BL/P
g5A1h/koMByYiKnY4/SY5vvkK32PoLyiT55v0/FjhzBFIdSr+82ooE+5iEAkGU/t6fQ8xRtO/Hy0
GsZARGHBrehU92WU7jauz72BM/v3X3/Afyh3qoFBbDFXpPWUVppmdckKocynrQL4zpLB/H6EB6FX
Kls/xol1KtM7HrmsO2xXNhUr8aO/gXbi6ZLxjgF4oVBq05ds1OxsVUU6fApZ8BKli+me+SXkgJJy
Z+MVFLI3ZnYgHbXBKzkYp9+H4qMnLQcfY/al3yk7KQQEETgsuN/TO50yc+IBNLQ1RYbB7wQlC9eK
4bRlzwCBV20hSxKOWl0VK0JlEnCUTAaNb9XNQe3NQiH9rEQMkFTDT+v8AzUcSkKRaxZTidl+3BOk
cASF2218YzfFzXwfYQkEJNWFF0xJmlB/giNrF6XkbUFf1dx0EIZbAiZlzZ3Mjs28nfXDbi6/jhGa
Y3DmtHJ//U0VYWNOavRxWwj2I9M7Bxw9aMl6c5yy9GzAqJqa5IDdhpd0wxCa2h1qPjHhUo7J60D1
v9sA9+gFdSucLGdmILLNc4VSRoMj5xzspmJI/nQmimTq7Tu2DBahW9IA7+NACRpDwFIWyRUnDzks
kIlCKM6suuDkFauwbqSCtI77a8jw2+ae4aqkv+1vzYNNsb+fcJ2b1l/rZxksJtBGVGIwTbGdFtGm
LLPBCqjU0SBENKRPzpJwCdh2hpQZfRD8pb2SBf3ichmu2/GrFAgzc2AeyeHNX0+94tv208fenchl
h2RfcaMKIIpXVj1OAvQfikkPOw/rGAwVHrE1ERDEaeDv6+vK/A9LH3bFqEgbd28XJILpgBzIu8U5
Uy9scdG8ckSwhgCQ5SJOVWicbdljFK+bGKZv8pBVFQVL6TOvZzTgwY6dMTKgia+cLUW1vwcrYYCo
UnVwOUaq3f7QYo7BicyGqX3EClXM/sjgqKO6GJ4jXvFNhZWZZfNBAL69wqZ0IyuHsp/yhZQv0p0v
2LtO7yIM2dyF55wDnUujKNulHZKAyORFEpUgwuSyisGVtI8Y6N4EzRMizuzUsJE5V87xq0BGPlwZ
BTOHqCe6wIlV6M3+mNvoOhyDVsenrlVqyKn+vtHDTAVArpEUJLIppgdaAXvEuqiEXus2GgvFt8rf
FOqT84CzB4oA9wzPKbeFeZaS9+/s0rwIIvWKBdsxbCQGR19YPYNdROzVvXhwbiBjTLE/AeMfUxdT
G+XJ0iNBqIgqclkQI4lUFsOPRBSF+Qv/ZQOeExEXZBvK4ln387AaJ3Xe00EZW12u1qtajfTtjzPA
0dDf1Q2HSxN4kYPJHJyXEB9gk8JuEhSvjgd6zn2v8P+9PkSstVEw0w0QTluVFjDkUu8ObnLHYNLL
IfeDEyOY/G0vRp52vWsQk2frYz5+PbTAw5+ZNLSHqyRppSGYAhQsQqotgyMRuU2fcJBoKyRk905j
ZGjkdJdzjOWxJEPeve+HZc16R7c58t3hJLPe++nJmboijuvmh+GWOGsSVjP3B9mFg8zuPJYv4HH4
ULRtT1MVJS1MM8yXy5bFpD5UxSZ/McND5kAiOb0OjlKyyRQNSAeBM/C6MDf0k2/9DsdF4Y6vG6IA
8k2hvmaD04Th2M0wokj9IP/Hf68f5MIb1ZdQ0nq3ZGEedpDRWEdYXBGg+nBIu9jr+xCaSj7Smpur
vrwiPBBY11PxO0pUdTBSkthsI6Pkbm7v3FhgslbXOvb1HgAHkSjfPLGvqQBhIvqeV7GRWcLkOHDj
oglemhSAApbVeM0ex3d7trBOMi3iPqk7ZF/Dt48aTLP1XnG5uxeYu5K/sXb6vofZSjiqLpYKPi7o
2F5INDDScsjNGM+tBkr8hoAbDwOtaWhEzcJlqOx3VWVzdkqoeidq2CgGmHcNqFYSOJRbuhxP0hPA
p+8SALzO+a4EgelFwK7XTb1K9Xq18Vr/jBXA0V8bZfXRzu7w/xnAQ0TaYXF/95O6oEYOdT4Sjojj
3X+NnxRQk/FPZCiEvklrwrbfURpUQKFKUW+H1ArcWG/Dd34S2QQn4X4WGUKfyuqCBkDQzkO4tLCR
jfWdyqV4DcIf3xFSLM0eGLe6RUUcLXpWAT0cxQCSYm7Ew9MZPIph/4kdRo83xXpixEr1gyn9+QQB
AnsjuIqKQZMs0XNK+W1Kuibd0zSvqhK22FiJM1j3Q8rAYGcyQf4KGOyQp6G52GnVjmLXXSMt/lO8
f5JVfeQt5Bwp4rqjak5TFvoIeZcGMfdBy8JQrH1TPD/DBQMSMQ0TulCoWVb3NmbUJjw86qB3i/j7
WNZQ7UjFWtNm2YlLOzNToGINf49ttGOM8KDxMPsuLPSaWXzfufw9CqFHQMTuY0laOEhuYw2NC3/l
XsJWEDMXFXldmE1wERJDAVycGwf+JxEmKfOWyx+ildyNE0DUp0pezZ7I1T2FOjLTjRYDTmahKlvK
uS7aMjEOCFjGLDOu2XHQojvqx8w/RfPM/4lhyF8yOcQ2gKVHSi81Fl6nKnygBuI8aoRSu4siz70q
9eB7zvMmo45J34BuIO4K3DhzPHnI6j6NUHh6cpBodieJ9ngCFtAu8FyI1IbzWP8ymTohyXaJPI/0
DaxJzYwCz8d8r9rQ0aBnBCXyjlgJbzfd+ust5kYFkdvssOCSvtaCwochuawvCl2kPD0SH2FHv9J2
X10WNIh/AvEAXXqPhFXFixzRQkTESi66uvRk/SuMP/dD+GpuD48dEORw/2f/eMLPJKWSNnap4pqO
nJ1jV4WMqWkVaIhSlMINp08eSlpUDXUbxr3hZMOW0CLSRHeJLfY41UyJDADKDJDXObcOuEha0iSL
aew/5ONxfJqnpspQ1t5+9AlsL1NuTcr50b0w+Gw2cguF0KIwacRWGj/2OzWN+rkiztLv+sBw2x4F
s9aHpxxsmCEJ2vPqMqCJVgvTaIrw/fL6TunpSmRlt3YcOrbJZ4bKyEtkf27A9SMDMqMAofVxB1b3
ibrC420KytCU+EHaQ86d+MLFInbncnJgW6TeLCImigzVTH0jjFwwRlyKFP0zF0Cw08quj4tva4jF
oDMKjy/kunNJKsVIuMKhF5IS7vQhsweCXy98Hu4gJJ6zwkZ94YE0I/oNq9fHOvw9SIEjWILiJwM+
37fdkE2VVspXgdtOXgNjMYiyCHHobnSWjzI1Fpdlo510KxF6epqwdG0lPJJT1T4luylkhUIJ8auZ
3rFChZiFmGC0EziiGU498jj6rndakZDvqOI6E0AgK6nTn1Nnm9C9rA1RBK9xy7N5U9eEMqsz8Z9I
lH4C8ikpGRhQtuuxjWiyXxQU8LLMGzroOhkCbY059gfNmGozzJv+gmJXgaE4/QWrLpzPw5OskptG
i0CkrfFoasuk/mfxbciHmBwz7G5f+dEh6CkY+HrIS+LraCyBAy8NjRqEBckQ5IImeBu3fYP+pdgh
THFD6ezy/kVJgh9KMLYrkCS4jkcFZll7/2qCo0ITXo5+Dr12mqhkvhv2YM9nlL0W43Rua8bPGR5X
El43ZGkuPIVdJAuIYaC0UjMMhN7jMcXWb8EuQpLV+3WmUIyrB8iSvYBl/3UynPBPf+gydnh7wJI/
7e1eaojWzGmVOKfS0t+YjuOjK/ptxmINkp4zJlQ328aAZQPvD2Etk3XJOK8s3DttXB7mm4bCIvUT
KoYqgL4klVZMIXiw60xUg49WWbepSvQsqrJa55Nu5j1ijdI6cRV50HBMR9lb9AcGyHy9Jv+bdy/x
7vzEtn7OvGPIIkyFX0cP9mGbOoqY8wpsgKYBvZFVausJxoM74iYgJD3EyBiZvU6WPVU5RzFZJi2N
+7M5+do2hrnF44B3OKHcOg1Y3/tEBp8iGTcCWL8vq39rWv/seaVa1w/XO1pzR03WIBp/pI8R+q0w
1R4yMb2r1rNln7+cb7GCSJ9T0G+Nrs7NkIHBsGUvk5M7yUWsyG4I+sg7mwppc6XUPB67pEIBIdqi
yTKJMTj+TFDqHoynqq8+9IyWttQKXHZmgBZevvjIfuXDIO/jk+4T04Am2W+UNWR7kS8zCLew472F
DqxRO0AQy7yQ/aB6e7U4r/WPOfAKw8XnidLskbVDrlrbJFuEDbgyh7vRB/XqEkBwan8EDMaz8bFv
L32F+mz3+Wzau9IJniaVkw0WXN9JeDDkgAEdU5ikR6eKQJiRx0Qh8lGwwYlpplRstqqEoo/RGSu/
JuQPiDVZ7YlaK3sHRKdc+m1N0ViAHxZxpl/2W+VQlquZhhTBrH6SPEbiVT+wQ5OQjIRhJsqlbwR/
2+htmty5of4CA1apXDBFXn+TzblzuhDsdAve2EzXovemiK/ffMD/lZQbqslAzPBaGVl0I1rSzuZE
19r9BR2ZXX7erIV3MWo64y3tKKGieha2ANaZ2KFHnKdKk2R4APUyAKKY1/N69oIqE291JLR11T4e
FeRVHfO9eu5W7GG3zi0uRKqA1OOKU/mxcdD3bkn7/hnIXq5UJrDBkLcNEMI0lyDqMEpabKnSn/do
Fi+Wq9jKGjmE1w/PtIGMRo8H1PnWK6TrRe9iASyQKj9Kt92MxQYgSEKlmRO8Oy48LQFfp81psVew
C0dVREPYwi+f85EZB/g2wGLposgsjgk5E+vMSUczfYxByzZbQBer0zQsBXBzZKmntkFm74AvUz6L
QfRCG67dr9UP5U7BrR33X0J1Yvw1vNpp3Tn7q/qCHAjf1XrV+eiK45DeONkz3mROnkExmdFBm0L4
dzcoCBO8uXLXBks0Uyf1iO6M7z6BY7NWFH4f/WANPSSDW7MQJRYtNp0hXCYZUmyeCFd9I4saxBPM
n71E3NJYcxoXOOfyvMkPUBHyrzZWhN4aT3tmmi8Dmws9s09wYqqtxdxaW2E0v4mnVIHKrA2bgg43
ob0azdxJ0x3EtAwjXMvBOH154WpXBkIYqmoGHlXkQHzgJRuwiBDjY7ouLz9CO/cJq6QQHGIOrAFY
t7VNdZsJTiQp39ELWIlpF7Dm6qtZD8gHy4KnRAGZHpHGkA6jzzZrfUW00t10vDyNSJDSsjTOjlPH
mYI/6Y8KLhII5Zbxr4Q6q9ZWEsZYd0peXLMSgUtHtBFZQ74CWGohdLyGgH72oxQucrw9/qgnt8j1
F4WLhjbHPSGxVIibFQa7q0VVWDfe9Ge+mBxECrNPjfM1CofW/C6ytOiMB/ANGz2+BM5qtuvidSQi
RVv5Rcm6mROoQDnybvaUa8wfjSmwe8kimVku+AB47hAYpaplNcG7qO5P8PJ3kWwtcCxGNImTeXdH
2AY03L39dBnp6tbry9aMAlSl7YoF9VuqvEjlNBf4HzkdasHoLMlopq+1w4PpbQBK7lDgFRTe3C9h
Cr06aDV0M/ChDPaBkCJoC9KClC3XDPKsu8k3pNCVqWro0wX3LVhVp9o12oN2zZWgHfH+2rHSpXQ4
k3QdXFyskOX/n3A+xEnlAZ4+l6aOi05/74w/UiZfZb/PnqjK+BFFtPXXtwj9XX02BxdEsxutC37U
QBPxsnc4GiPs9buWHnolkVqC1TFDvEiC4VD4cqGZgmQjOLBIil93BqII0KYTcOwsbGxPcaKl0yxM
Q+XVdaKMAaR4HJB2l8FpLiNYlJ6rzjuozsoiggFx+sPXR88Clmf0gnm5xzxFdm1LfOEMu83tD9Bm
cJv8GpC1tNpf/YCD6n0ppScmc4BsPScYDPNhSZmx7QwlgwdT3s3O4pMBFFk4zrridQ3/VfDPIsNk
20mh7sHUSz1flX0nKlHcSgnieLROEJGayUNYeZGN6pDjucrj7GEymoOTL/B3SNhOb344kkz1Htvy
s9zFJn+3/Fo1G37s4Us3nCGbumMuBVciolDXjaRhkxF9yssE77yHHNqCONQA9zl6osQh600GuTs9
CoNBQwWHIBfgmwtFMJcuTomYKKLcM3M0SV7mfWwWuYOj401ns+GkGWupHoTqS0lu02t5Ui831Ccd
Z7eXuYB1Ppv3AQduq/wYukjWMiRlC4jytGgEhwHz5kdJWneiGnbQxvJBTp3hL+ISuSRRzdqqJE55
/VWq3WGViGIwuDr+LoZfFC/hxCWTSDblTDT+gzMM7Fq7JkBNHiDpQSzDhAeCLGU/+QrJ5bh9o6Gs
ypHwCEHx/3omz7VfEC15zcg4SkfH/3CAMKKJiZt4c1prM4MlRwPsFGiTWpr2cGCM7b6CXKFE2V00
vOefJsmx8dyaAby7oA/7xlbuXbFaNX9gUtI4I+5jUZrVXAQCGeUFGIk/W9pEE5rP4HjSoEwFDI5D
nuG4wGSu7mSr4PVYZT95yQxbXc8D6YU6V0ZNdSE2DSYehDOutPdXOahZzXFqlhBU4+gdYDQ8x1DG
r1wS31MmVyALQs3heaLp12C2U/xMyp5Ilwuq0vkjYnmMiJpfeTo77bqTRfb2lEjzN1zZ2do1sLZ2
GPaTw9Pg2HLKJkpLnWwsxK4+ec3KOtcvd2Ut530zSjLqwSyr3IIEIAFC2JdjMG4RK5SSYRlekEl9
6vFQrAmlQCOLtDsdeBsw7JVG/d7wOl40+YvxKNILQnlwh74Is9lSE8ewlA68ag2/i2x0wE/vwB18
X5qOeH6UFofZCBt7ZiUqdelJ6kpAqfAowoytCoM9UUzZ67zTzbstseEBiL7ZjdFwZ7SNyE/1i8mm
d3A9/OTxLS1OEFzw6W0pQ5Rr47i266PmaUox7uvzKxQgxa6cnq2l1u9rdxjTgYQAlAbQs94TWZfJ
xnZGbwPuiYvgGkiZ9gbo2nav8QXdyw+EgAaNicW9C7JTfhG5iL2xz4Lt8qeFphVAGWTxnkEH1lfB
DN6jJwBsoo5KuKQ+FqBZBb6ZTlBYOtemrtoSXbhpcY5jlyk2OYZHbEm4AbtlOS62CsOFJT/Vikp4
Em4teYA+TYgeKtEOZyCNLIQJMkzPUDh1e8dZkS5wjexAC17xFl2haBR47AIlDwpnbrf88GQ75eZz
wosfB+9Cxk8rwsUxmQUpsNkOh7+ugoHqZ26DxOfZ2EYE9IU02gtIUaozhKoQCZwtpKqgvEHQ7o3U
7Z/nrdTUmniEd359HkR6bHYlrF8QLQEd7LmlidtCrCi2FZgF1dXizkRCL1y+3jBPtVrGaJ2CO+Ge
meXrrn1W3OERcVPZDNkusBKGcKkM07eDuHH2aAllEohscBD1VB5ERVgjWQt0QedWa9hK4LkJFTkV
iFhKej8fHw9k/rc9BTOn8liQrb/H9O8rGSWO2aE5FNjnC3oRj7QvaBzTALYTbHfTTXlhfngmi3x+
KbziYNP9eZIkgXVQbxTDCHq1SyIIzOYA4ENYfGC0xu1jOhApNiZaGF4iFr/NiJFpg1lvGnkGL8Bs
JPgaxibKLaRMBQoQQmjjfu8sWirJ9iZTjPupJ3AZ7noBv8Ss19IqCbOK8S6lmMfSKSCeEvuqfWWs
0KHMkFjOFugMbW3iv7dAPlxiXHzGu/4A60rhyEQGHK6k7+4X2d7Q3dPkQvn5tImPKk+3nW7guXhi
ljY7WhAEs7QYTJiW3bOrWxmveNUi3SL+r1WrdvCy4BeESyYBv2e4nWqyg7XNNVQovfqd78bXgngP
KI7fm0cyuSMxId09UvEy1iKdHgkCXzI+2Y8Q0qjJAvkb0FwQKeHf7BDLtC5D6JxnkzbNlGYzFWwh
4SPMV4BZZu0eJe6ENziXHAQndjFVnGwbczuIf++3Agai6nf+6sklyBjoi4Q8RoC99XL95IJHRS6q
nIWE/COXRLsdlaAsa+ISq6LgJE+YeFoY9+JlYCatz/D6QFL8aSFCUiWCpjtrIiIvEdwqAIXeVK2y
/4+h2K3Ljq+5BsxWxYp54OPCvfFdIF6X1OQlwoLiZyqpdz41gFNoG8iUDVB9YY/FyRoS74Z27AJR
QZgpEDrN5jpOE2CdINzQ9m3RLTwCfXCU2pcLa8ARMW8KdyNm5IHlYotI1shjNM7leybemiY2Il/3
8YKDpd70FP7AuyKUYO+NbBmaCNUVwbx1y70kOQLcsg7q85V2yJ/MbzI+rqET/DDOLjFWSF1rmb6W
hgUTJACUOJwCNjq14vnPxdjO/qdZ/DJdlRS4Phea9LOefbHRP0TSFF/IrpqYcODMtZgGEadbO32O
7D0XeIHr+0SXESG3HBwKlSLYilNLr6lhKpRPIbfxOKFb4/1rdfoErKPVOwY9KhphDXOr3q7yceqw
br+UJu0YGFi2F4E2fPs/j9Ly3OohChtxfeJMUiwt8aWwu0k1vQRDXr2KN9JBg3HebZA9R5J5njHR
IGHM9fMBj+pSgLvY+x4S0doondds2c6eyrQhHVVbqT0+9lhrpaF+dPTfVK8zLRI1XbuXSt2qnj/a
oJ7wWh7aMrWPf03jLMsrNk3OQS65yUEIsSdr2TfK0JnG+m0HjxYltPE3qM33mI0ry7HS7zUCc1kS
YeSkikD6uh1daWOg1nrzVyXCwODyEbYlv8ZPIz1zmNZ2dQLpzrQzTY/fy35LFn1um7kNEPMwhNSy
8AurjWJDITxi/JAT/juV8hotfca6fhcfhwQXPcU9vVr0XqDm6JTE7aNq0pwhIb8aBEarBgXUMgVE
gDew4Dzkl17kru8ssW79pdA4BLHmlRCHbXn2b40ECSvpyOlbLpiiuMVsK+yZJucuyEGwL/c5tE3s
7kL87A8KhSzZCDTahA3V4rFPf7g7NcMxnxLZILGTydGVivq8GJHYNCsSAfd8uQ3IYuxwTK2iltIM
no5+l4bc6AJ5NpN5FbYmQIXUkc5wVv9uju53YBGBudpL7KwgwKCev11pqVsj1lwzoLipUUD69oi4
Dv9qtSQUPNg588pe0JmPtBdgufGOuaHrJPKHPlZM71qUdBTZjpHI2KC5eZd+P9gb40zH+3lIWfhr
OW/sGe33lRdXdpgEuRkg21Y4x237Fk5+ckD3Lx2J1DM1oLbz6wBeLiOO01j8p7LVtv6W9j6JSv1r
8iGnvjRFRc3HSYbESdbb/EeSToAT09EYU5XF6JWuBI7abNh6aEe7A8jx29UBfHQTUAXgjYagDu4r
JUPez9wu2fQe534qPhBXbEE/5fKRVKpxG/neFQ/KCJD9R7Ay56xPPa6s5wm023xf7dzqjCdxYco1
1XXBf0jp7Rh1Cuz3WxD1oA819CeuI9MRG5J+bOznrAjPEttswUYyDA7xfqPNhiDDEd15Hb7I5WK/
HAFiUf6eeKQLkjVdacioWw2sOt1BPXZh2ZsFgRE+23N2/aHBrWHDHvrSh7HWzfL+urTMRspClOLT
4YvMGCn0aNXgVNyz8D8WPMjdbv9i6GkpxKmtXrPeEBVyNMkwmXSDxNTeBOqxOf2VIG4K/txBECpr
YxfeTNUqY8vA5fWnqKM4ktK1ZD8X5B8GmOE0XpZBEFntCvx+kv+9MsEwHXVnD+9gsHhPWYsuuTiv
FrlIr7e2BM8WbzNKD7LyVM3+yOj8sFczVphhFRVADxEasVqOI5Gjlt9cOXGxAjmfouXEDIv4jxV8
nuU094CPKvrcYFIx5OrqRzxnn5QsZEZghNTsULbnNxdihiPE5c9wzj5Q5BaIyeU16r/dIRwTDdjB
vAg6EK1rRGDGzGkXPbhlZcMByIQ0ZLkdWZSMeS5yGoQ8aWBoR7ht7LBrI8cogSWxo3RKi4cut3g7
h2SDmrOpvM7F9WPpFiWc/J2cMzQ8KI0+GFqZIVH1vlboDUY1vIvQ7Ww7DMTI1+915JtjTozSKFCP
we6GY/cRmZa9GrVbPPB/OZG0+42NrFAmSaYnZW3gf4poDW5YDJZIq0i6xTnCvIbjKQty8jkEQeye
7o71eMsDcCZIFysxJQiT7ShjFN40Axv3v7SQjjQQUWrEkcQeaHwVW/3nF7eL+evTYaiA61r3XAPO
XrwUuAnKnlSI56JN2QaXH6nidmbH9p8SDRBS61q60F/ucmTk8+QcO9Z/j6iAnqvoBJmtou3ldDbX
vtOWUz5wD+HzeTNwyoXCjwnrFIL1XxKzKeiKrLtoFXQKBqGjqHXxpqAB/Ikp6zohJOUAiedaAQTC
WWPQxOewJI2jyY0kr2Ix9d3S/bAAMpXo7+DG4+nXba5T2undym6CcpVBg+R8xXx+LMk/9255vfJZ
s0UVKsSb31lgOEfBWNR5+W1bccnFJ9XuhO560jX/JyKkI7rVxo9KVN4sOHC5050+U0BpVQwrvhxv
DYrFLzy4wTsoQPWZJJvXS06HUbQra/8WGDZSF/eajW+GffBt+q2wwOojPRSb23UJ0U1eS+ZXLh8a
zy20PF7m6zBy9xKMuw5FDzOXxWHMOifJ+suwnwNydUSJXetjwtOkZyTY7qsro1gW/mKm7oGskAAQ
xmslDjSCl28JEIAQO6kwXBeD6JQj+ZHcf2KadUVUv6WfQ3gR0f1GsSpWwCOJhfWcCibtWNcjtsi0
qO0Qf9PyEPioWE4s/JITDomYfU5NZxw/697bgWmNI70o0xKcJFrZO2Hi/t4Qa97F5YxbH3RXy2jX
iyDpmNfPPAIoQVmyBsFlzF1Mtn6Gl+AgTRh6qO8H/7BIbSwhGCxuWTghk67QDKgwGGZAC+FV1uUo
Vx+7uitW9cmFYPTU680ehBVgDd1Y/ngq94LBCz9n038oyyysYoGeeQnERQWHszON+Y6Q9RLmpEYJ
dB/qWkgQW6JjSH+dWzR9nJMZJCwGVKwvtDjEt1t595RrvRejd/40TPQKOo2M3HiQA9l2SCo+Cwsj
Rd78Whk0YIAXtBPYwC3NERcqc9yPjJfZjW0CmS4LjmATAc1gvt8gRCURD00UBJ6/b4V+IV9ow/Nm
7tqQAR5i1yq9qF6nIMPUV/S8E0EqZ4h+UeyWcthj+uRpBN5b+jcWtD8jGzCnmbVgNZQCjmIIGww8
7iW56tPz1kM6JgbZL9ZPYYU+m/ZQh/oSAXUxR7oIfXouu1sp3vyWxm+MNMMWiZ46yBR9YlabAlIk
gdR7ttxyz43Q8RhWyS3s1t10/EZoOKkOSQmL148UMJe0jh7humq7/L5/4kz/BoY7/hAFbrNskreL
ri8qRsNoesjn5of+ZJiZNAsi/uVr+IviJLgV8nBqvBx1G7aXXduYFc8vDlceJ5n2SRoRypLpuqTR
b5I19pnasmDQm/m2x/Zvzem5WwvFt0vzp6gNUN6ltcuoY1ql1BtfqjmJZkgpSPw9p/1QFJlX7NVF
pS7Q9lY6fvnMK6RFNsMFz+jgCDV6U1NAjEGnB2decXUMlfH+FaGo8vWPxI1gajOWMKNeNlIkR0Qy
cBhwiNb5i5Rw/O/0c9Rs72faWMCQ7lvnlgD13t2n2ElPRczeDAgYALP+Iu6/62ZsQoM/GvAREiWx
znHyfj0d2LWoep6Pkc3CYIkxZzvYT+3p9bWuZ+z7roGLTdvOcFiiWitwd3tj58pqNxWDY+q6TVc/
wiH3NjT+bo2JwwbkoDAIBzg9iDe97j4jaxMd0Y3i5hwf+hFWVhnU8BZb33vyQUlx9a2HxhG3dCz0
1Y78ZLqeVEGlyV/NSatx/DfgQPIq4NEJDzYUHmGwf3VUC3awbf8wEeYF68A4nDGK/xm6cYLUAq6x
UxGDHJOBhCBb15sB2x6cSlb3xOJmVQdt2nEDbPtfidUSm+Gb9lBz4GO5TlkI9DuBzbWEjxyvEarQ
T+5I4xmRgJcx3Xw3E7x82POUNY9yWi7zjy2bZhi6tnbC9E+evF2Zt1qzOVDLQf3GaU3mlAatIFfo
uBvO6D+qvcZvDDnittmofvO2Jjgu1dM2Qw/8moY7cLbSvxWnAI+ZmJLytur0mFPYAj+Y6P3HFelf
2wKaf4FS7JG3Hfr8v0WabFdObxxzAtBLyzYFnYARNKDG/+k4aqH6S/wF1DpuiNW0A0XQdF0+J1J8
tDiFiAIiE3K079qq8snNyO/NMeEX/ly+37KAn1yGdTo30UJeI6dCLu5eY+PjE2MMEpqY1xTN1Kod
3iIU1Yetu4U0crSSQQuOWFwxUxL50c22cQB9DjoMGi1ELhOUO0Z8Dv7Y9CfBrVHQka0hOE2l42t/
ZOQA3Zomjw9AoYUmbZxyX4pJNydnN4fz488O6WS5fs4y8+NMi1p7xGYvb7g0GpQV5W8InddYMJxv
tfRRWvwGjBiur7KrX/EstQIRB3mj2yi+y9PbHV0/8K3/kIC4HHOwyQqi0OdIWivxoLKoqK26jaia
od8xQoBy1P0PC0uLQLKtqmffLg+r0MR177H4JQ+FnaYj1caYTrn4ppUTcZYVntKrcozyozrz5Jlt
LrHZ6THHZy88bMv/KUVyH18Yrfvw6MC+zQoSxtPZtw1dUvJmhQ2JOQzJPmiRC95Jz0usfCtWhSWi
KCxSkRM961PqIjQJXb/Wk84KxrVUjchFJHRF/UGsXf8cM1LVRE9W8HUbL4URzWzcHgwZ+EhT1HlL
3x7B/qifNsUtiZd0pnQqwR47cNTqwefB8ROVxej+cJCfoAvCHMiQ7lVGTEwR+84wO4NCSaOKuhgt
yX59xS6bUO7nTKHqfvO3WzkKmHXwOgmFvpzTxSvAw+gEWDN2jhQETJ8TDQMlDUkV/NzBlPcXOnMj
LaYy39W4B+Gye0nHCDsDsgqcwWB2IT33cRRu1xdMILJ1LI3BABgJum3K+ddb8mEbXQVSQf/YnBHk
U3Q2pZeKSDxOWCBsnnXjAcATl78hOkN8aJNkq69lvgdSrY0fJaW5x19bUyo69r6Wl/71niZJT62C
SovS0T4wQfz9mYjG6r4p7+b0xdDygYeGjegO/EEHd+0saF8VeOqUxMAXvxiftTK9BiRUR3V7FmdX
tGxWeDdquv6NQR0LBXI/JTFghu447INuh9u0lm6SBJvpW9FyBbkVVuqNl9wEnTwoSbkqnoZ4iPH9
NHtOnDcCQm4zVI2E7Ks5TyeWFzIPjsEQaFHeT6h/xQ2Fq7mdfF3gPfqbixpkxr1bKT4MleJ8x8zb
+W2e2TJM8Ccu6NkK0b0Gq+eGSJ7WQc2FKNNFB8HwpWXEGzgz2bUxkXP9MfDIFmYRvNTye5D69VsY
p/HCbS5W6CbSMmpJNevGwtJqRVG9LICcC0Fm2u3bjo26tuoEOZl3pTyrhBxl8qHkTXjWjMg/x5OY
/L0ptQ30QwwTaaZYrBQT3YmYqzQ+fR8iYOsQ3AxjEcMmxg4V+khW6s27ffqvoxWyg91xAs2UGI+S
awLuTZbXRiDeflSCycGY+m9/zO99iF6hW5j6jWewtCShGe9WH081cQeAVkqArWaGGX8hsO4p0iaY
SuJz4uZq/mqurRlgNRsx1KXYM2a23vLiluryOdtKToHskEjkR07dacJGnudfpKTljCSC2+Pl0Zb7
gAATzTRZXQvN/DFuN5vAqSBlCofZJmmFNkz+LFM45bh/NwMAUIhQEBcjvJPHa7KKi1NKCw74W3me
ZzbkzqvClvppLRbN9A9+8ptB081bCVgfQBrrYUsyuvWfIXaV/pe/HemIqMr7/5wwhIiyQgbYXpoz
vKD8QMdH/b7Xp9E7ato1C6LZyuFQBFBdBriVI1r4GMzWkxLJnYVqfDe7G2HtueXRPgiShdeVmZvz
qk3jMp+u89qjBXmUME3qWwwoaJ8dbZVq3prANMQRnZcqmzhAM6FhGwlBGwK0GYrwfx2rcXU7RNl3
McQ9yOTdvBdEixN5lwSdTcREvkUDLLX6XW8bYtkdINZLA/AkaYZA8s6+UkX3hQR55RXLZKcLl/xG
AW3CTFIH+PqE6nTehgeQm3D69JNZbEztUDaL7ER00HmEL0j0tu9qYvGwzcIDQgzIzhegWB4w6LnL
H9K1TuozkH1InYV4sagaNX1uwYADoStrxZftl66By/cswiVP69nvE91EJu7IeA6hDcmlIYGYrSzy
SQVL+xGgzwEKxQJzAy+sSJsHPdsvWxRNnT5i7LdTcmhZH4+jQt98fa5cPGPEjx3TYsQh2iVf/JJW
3fqDyxjpnFRzcveh//3+aJQB/fJwiFReBpm2lqpqoeNyJfPO3LlMru8aWz4qNceg7mto+xpzLewA
9W1Mpz7HzqM4KuvqjJ4spqGz8rdLZodTrTWB/qX3UrNnQ2k6BxotuEbjwf1jXt5nkEHSSX9YnfbX
SreRDRW6bi1aR7McEgu0eKuaXDMU7wI7yCuzmhxJ56v3GVpK/43yKVxmEHOLIQjGZrhPy/blmCmQ
p8KJdmSVR739ywReD4HdXHqQq9qLuolNql806X+xb5bSshwYbUYALywSFWYqPMo45g/7MeOaDPaT
pf4YwOhCjhGuZ5TUMfuCMboASoISvEz8uc8dL+vns9bg5XeV4dYaMc5hvO3rpHxboxM7F7tQHb2j
IbX4L1MDVCTWSnMAS7ysXTEE4+0qYHurwyIl8bFtld7zDJT9SWlpEMvxSf8LXFwKK7B38vHDSi34
z3JzcXZjSM4nE72GykZnzmeTbgOiwWjs6RHRTmW2GRtUCMWCYh3JVe25pD6yxf0y+9PooM0pYWwG
GEZXCWn4bzhGNLILCC59JxgxTQrDjRU7F5ZDRFcocE38MaVJYV12VikJ3ZXN8rQNSCON1Qgmm7Lk
u70ZuiDM7F8ax6pq8pgRuawKPJawfxWFUBACzkSwKLJ6z/WGQM854iQbWTmYV3Rmo6nRDUPFh8ZQ
+He3w5wxHcPif05Xji65tKr4gvN4s3FPztk8Z7LkKxjyLAO0F3S9SFSCJgnGX9KDwQz9qoru5K+9
LQQdYX0vAcpkr6dtu0Njo+ST1j67Oq5s6Zg/w4A3qaR33AVzGQh2eyAIq8hcQXyV0ubxDsz/wThV
BT+Pr78s80w5DDPhzjVqRwA5FqZBSAfxrvPyCTwkeLLs4hRS91qqgE4SlgkGwkvlBJaMDiop8n16
oAmdi9f6lPL+CbWJYJnEmBrM78j7C4z+Wf4MuCVz7JKDW0ovI300IzgKnm/k7sU2gLawvvZ+QciD
uuR3jfWW9hvk7jCi0SUHj9i4w+73ThVmd1CerAS3r5WorF+nBtdL6GiI/NdSEiAybqIwkcaPv561
+PLHkheHC/NmZ8eUn40U1gCZ3okgwbLlTBfVQDOFR8wKDP0607ZLm/yz1H72+ssorBwbW9SyziEv
KE3DxW1OlWAvsYgIAlUd7GBnvQFaICkpHU6bLWT+G3evkpfUeoEYwbHYcIHxnn6l2/vnlsT8a4JG
lT0SGDWCLiauuzrLbb41+MDXwNzkHIL/urKGrGzpBzR5EZUSbWwaZFwOUBKcepbpRulbl8zSvu6i
U3mnFl15ylqRwgECeB3twrJq3GVAZCPT7/1IWePNwwBSEEGPTWczFc1+zrFpbxOlgc7ZVWCCW+2l
9xYPRXlZeeskQISwekhHzrL92If4YWSTlw0LXTMIAlih8IzRESqRh1hWAZ+mjxBnkI1sMcln0kg3
zsh1FcsgSxt1u4gXeQkPs+n5sAotDHqgJ4/+3CA9udtHnCK9jIRf5vH6maUk03KHakP1AdCZqaCH
7AGgC996nFuAcQH1a5iOO7k8/kJJox5lQ+dPwcpv6uJR6RbfWeZ54MAQNQUshA+cAg250eNC72rE
LLobA6mDdqTCjqqA/iXeoy1NdByDg3U3JoNaOaX/ueN1HrDCcQJ9539SQAQ/zu1+Tt562za24qD0
0SDGpjmEw/uTg+zUsaXFP56te9dy7LHlx/HYWe2eUiQYI5DgXbiHhk1MYRFL+krx4AdyNKnHkL2a
ucQ5F5tkci2NL3OS6zhfEe3ahv4759qcSkYvYi1Kl5E1jPjmPRn6lZFpIjfJKdOS1xKLoJVxJnuB
ri0TPSRo8swVPkMRv2ODbvX8zWaMERc18IvbSBL4PXrDobk76fCsxKzQDgcmQ/MGV0Oq22YHzDif
x22F1P4VyVafkMrDiTBD9DnobQCnVfBcZjpv3BRFc1PskWKNiOj0UrIEy/5VR28Zg/VoE8QnAsEC
Y5iuXQBUKdaYESV1Wvu45TQKet6B+GOX5HXafQgrqwfsMrra9UmpZ1F38DgOItLDFoyFff1dzud3
kJhVLPSz0XjFaNEVfe6bKwjN9vmxhlJUgT+V8z5MxcSBe/lvJLS2I3hJ63BbZl91nCcgf0ilcJTG
VWP7tvjjEr1qns7W8T/BTjd1W9qqpURmawYHLBR4p7QMU803/CLGtW/1IcK0UVlJD6swAy7eDxoQ
OkEDdC5+ZhabEhY0uHhl6q5ymr6uHqzGsuTLzYo32gaGpQ3DWM/WdbFWQopZAcDGHT7e4080oLI3
5WelDjYwe8pjGbMX6ewWE7wwtLra5WpapjTklBnsw0axpLtFjNDxUDoR5kpzrs6uAmnAdfP+FWLK
MKEQem0LwwZdivYOX+tVk9GkU+y/jkRanYplKIY1PhmWl9UcMfd3y5XBcDJw41gEXUiicOtYMCQz
gkQTKXoXGjQYtZELQI8KejPYkukWSVPOY7L/4eVgPAwbCmorsiBhSJHX4+WKIjUoauiE30BgrMuA
4qmz9uvuaBIvBSJr80Z3mYOkrNYAdCu00UZqsZ/hlq0qq84KGt+WuzeRubIRn6QSjj2NgtZTDcn4
u2fhdnou7MuF9ZhBz10V0ZO85LeW3BymW2wiHhDyipecaweCwlI05KQhSv8Ti2sj5ARrDcr0+V/D
NeQ2cBIR2VMiXgLCOcKo5CA45TSkggBgxZ641uJAt0Vh336ct6xyAq2VTTlkY+mMHQCGGhIXZNU6
cP301qsMqPS9wn2BMmGOtIAf1vtvXfJtZGKpbop9cYVAtHAAByyPIGHGJeMVL6wsRmyknk+ArhV0
23FYrc4ONx9wdABe6Nh6yuVgFdGdkwOXTgUsnnMDDSrgqSr1NkvS+MzdZsx/XxLKIShz5Dz1qopL
iEtSbA5PTPfRiZ8cQt80M8722wL3xSDLhU91foUMYH9bhi7TmW2bdgI5+TCalromiqxTNBPxsCOB
lQu1BJJxAnKfHO37G2bgg96VFe3npLBBXFrNhC4zcMTzLeRoUBYTiGaCyRneZMGNosG6Uv+dzZDI
rQHmk80kD20O39Y9/AuqOYX0jvdhWOVsYAqnyCOC6dqpUZy5miSNGmQNEZIlwD6uvlPr8ai1WjB3
macQffrbhhe+rCA78aHk4OL25F6p+U1yzEVj6lwQDtwJaenT05rVlqJ/aHDXhF3rgWBsCo1rksY6
+yaC+muojze0vhvuIwt6JiB1W/GAvBtDSMbaX3S9IYAB1q46lNBnSj1H7f3LdHmj/roxQLAhGk6B
pp/Jnl/DWFeKCOM1xPmEnJI/zjBWLngzKr9JaG+wWNDtRgmeWsk4Cz9XFGsecDz6bmUsBkXV8f+o
wm33z1Ya2hfhmnDEPKeNJw58yXEEBPiu0MPqfwhnNW2DuDOn2KxrnAUBcDpOhGyOPcia/Eyx/1YO
eIT7QXDg3gMPAIc5TXex1y6KOAedU7rv+KjOL3QWUNkPLSBkAqnfcebXgrYDUEzbdMOc1ByUz5oF
ga7DirQdDywM2uEOhc7KQg8bs6AmILAZTqK+o2vCVobWe3jfF+0oP0ivNzdzTI2g2uNn6kSsNyBz
9WWQEZUPTaWEOpHNe+ihqBMh14gI3R8u+WrHVZAH/Rxlbjn1WCCkLvqUshfFht1/ygH8KrT3e0+G
u6vlld4cRVmO3rgWaYZ/KQVl4RqvJ0WVfYJWq350NJG0/BA8u9JrS2JE+hUnlXYNrQeEP9q2uhOD
5rXuYDAfcyV98/ZfKMMkGug0RXSiuVSv9qXy8S9i/LPIBWfudd1z98P6PCUR90hD9hk6o2HWFwFu
fA65M+JmqBDKa/2YrDE0+L8GhDdXWh18APL9SAVxo6yD98ZlJnQZ82ebxuo4NcfhICX2LVGGyWB4
mlSdiO8PeBvcUdKPYcXlh6lnz1ZhPW2KY7EN7vTYSknHfWvqhVRCSESepxvQ3C3C/fnYDOQATut0
TWbRkVC4F3JC4l+muJnXlFFZdvyIJjKjjTmV0Jmp1v+qEHivbUNaVzGGWv/6huW0KoueVA8zJZYE
l35t/s8xUddjUq0FaxI/dslkooHcYRKutuUcsoJ5c/5v4VXIOtvIjgnuTlCWqibrn2VlpCqZh1v+
v2cWsJH9GvDbCbG4UQevydur5Fy49RQvFAK7ixETWYYADNlrNO6TFzq+OFAkb9L2LDfp/dc+0px1
+XNDJfrJSqW0Ff+iDFFwXt3HuXlQuxlRBKkqYFgLUH0Z+VpybRWc8LrzNtumGg34pWH/RK0u/l0E
qbW+YK1WI8KhSwWH3Dq2avwFieAAtMKgKFQyMHdfT0fAjYtTOQn/Q7yp2YQz1L8/8SmIs7ALPdDh
2rtpPrIint936kzWHGMmi8dye+NS7ilmQAkokAapd8CalBugRIryU6xHm+IkOeWGyJ5tijTcSaJ3
qJgJ+ERzsHF65YdF/9DLQQBtKuXahWuOmJXJl80k3iX7k6T0kr4n930Uwneu1fL1+OAHZoxHXkwb
/VDPmNyOMFbfuGUAqirSIEieoPWBgmg1TJoV44eYRudLuFh3cw23wGol6esMgx3Kgb8S9aSQ95wc
T2MRphOVn+22g0XqHmST+c9ns3qeVdEl4b4/SxG7dCunRMkj/p7fM5ZfnfWNF0Eh5Yn7kVOeey59
svxXgnsrnSoDeCEAoSfz8mrJzN1kMAUaQh6lD5B34Ym9lMpmpqKHBFOJiD2/EX8IXN8E+0JdTaRV
R5UvL4uAFfSLdJvU0wIrdFi6lHK4prIy4MuOOYvkxba1+wj1zv9k0eZoO3KlyqcN90/F+qhqJRqs
xe56w4tJxQHNUx1LCPM5c++jPoY1VycvanLclvEHfsC14NJkdWkJ8Iy+teJgMlgQJaX2LS+x2SCZ
enljFcFn9bU6rAG2vu7EaKUmNPwJwqNbHXEMPVsR/2cqXvt0v0Jbi1ZPX0rrEfUpQkY/LJWsRLlD
QLe8+oTTqOWirCr1b/Qy/XKbGCQInZ1QqCE0pW4OF3vtnNmvmDDzZJCRmVBsI8A+2qdN9N7Z2m+Y
6Jqf1QXVfHVjqFiSoi76Tyf82R+k9ZhZj4VVBQMsODe5llGGPtpuuZq0mJOnlIzV411imRL/xPrn
fYmkAOl8iX3FO18UxrfxWK5TWZqoqm7kZ+k9DmCJNB+ttZee0gf7b+xfRUCffMUxGdv2DTeKkiDt
wJoar1qUsylr9NLpMoD3ptSK+WKjM4y7bDht4zPrRGNKp/zK7QNAF1p4ROBfZ2Ok6xWYUPruPIen
Q7CWZHrE5q4TnQod64sfYyvBud32EeWgz63yO4uzvbyYtUyMYwphMvwsoaDwisah/MaEVUQZIlES
aboLk74j4uFwt0OqwYG7pC8U6G3Vv1/qYYp7GRCq5vKDyK7cRftI0V3wW7kYB96yXX/IWTWc9aT9
byy6BO6qxnjbua5nONQV/GcXVhgvBAOHwAk/RT1AYyqhlWVwrfPPEk04XVFTtdEukXMfWqf1BkZq
i84DyJs4piuFP+6xtTZeQaPn2c34kzEQOMDuNu4t8P/ngDIMVeBfmj4rtFqyE+TgMAGXscadVtb2
QP336A4q/CwS8spq6VhuaIQwGMU/a4TZhVVBvPIFK+aw1b+kp//hui4wmEPlmPSepcManWU9HRTH
iIOUYasKgS6V/NPQJNi05fkoJ99eTWbhlk3rJO8heH/yiU5N9Ei9tgL6gz9J3AB+2eJK3ju65r8k
YT7e3LnXTlBDbTIKTS3KfG0ksBON3B0mhY8Ofc20aczFfSj83JEuXvieVMwQuJ973HigwD5KsDbW
5oX+4eK6S09/hn9USDSrE6TzyKn5GwJLtjrTw4jPW+kOvP3+xgGiglnCE9lz1BdUzIKAmrwQUDW9
WqwdyLit2GLSChWQovHCUdYnGyO0Fp3QPRsOmwDZx+4OONBrYNMDbwuzoAgOYJAqnJkujYVX3eCU
h2hHpfFUIIz6FQuGmcE6yZuyK1JQtg9pEMt7EG097ste9HnoV51CZWCu7JQwZv/5d6KLUFqGxSoD
k6VA6Rc/nuJ4oyTUqXsMmie9AKI3EYBdC/FOCIxTEnaZORixh1rffr1+RiJVp4LYjk8FIG91muLh
wwgOoo5p346Dk6SmlFJ7Tz9G4el8cTzPMxFdC+4TjplHlJvPP4R/1eWboC4aZ1w07VOhELvsJ+QW
OudU44VfPcxUGvezny/46SID0/+JwdJ33Cyqs3Hz5YS7lY+9RLZa4Kp2uvJ5pDam9JWMPT6Hv0qQ
SGCJdtAfOCg6n/WA9+tX1Ki9gcw3MFLzdhSlZv/2MdcNQt6CGpykpXN+C06iFU6Zpr4lFR29cOuX
D8HqiJ7ABZVWlYfn5uZQwvFFb9bX4uXJvJyLsCPP/wetXjIFmXKzUZuOnteFaWRMZjD0nD26tmXs
XxYeLQdiNCmwFPcwRnFpXgbDIEPelMhl5vy8YwAHpjvIjLXgQhq/Cwu7A8InhBb0+hfx/NFYzXnK
AWM2KYndnvaNmP6LA3NNI8QmkKQJ9h5qg0kbvYm0fEZZIcUmPNqrz5c2SjGT5t7jHDzJOxM0fS64
ever2WYDPPhHbKdKFGDlze6sq6rXfJJgA45Xc2WrXNL0zM2mtz7rJnSoDGgOdPZjlHLM7VThoxa2
YhqyXrpuJaaJlAQ9wdoTLcwtTby4n2dldnDOZ8lyjcwKC2mbUUYqZEY1Z1RvYx2+KAWOn6gVyJgn
CaLZf5KgzUN4pTds/59fs0tTpcebULtpSGTxnRkY8BcimV9Atszc4UC9285GCOWpUKnev7nn3cvw
o01BCiQnAnaBOVmsALWN1Qob+ebnljYprIawMg2Yo/FGWHkPACKyMBivY4X7QFSkp1O8PJmtmzTQ
VD1IcD8FU/PJ4aiM6YFP2Cv5RK4wSBHUbWkIUeBZVBDKWyEHnLeF10yrtq55J5i/61niIExA+Ftm
QD4fKvUv1d/1QgeXSdoKdoAjqWY3rZq07y2rvXTpVHMKn02axCXDvIt+3KpDMIRDS5Nh+vZv9X7t
C9HnMhbMLfFRN8byK2OAzF9OeTvh6KdpHFe5BHqptaKTVFQxjCjelLXFe+yQm8Emm2WLFjVoNgnO
AVqrj4ombiBo6+t1yo/wKNjSCBHLeDA5ZpyeciepVVM80PPrF+2aRgqzhEsnsgyW1BTiQ2jDz/dV
h1G4uFaUhECGWzWSqMCnBC/wl7b55oI/77lfbhyV3V22fHj+qpoN90Qy+6O0n/6ohR5TSCPPDJ2n
VWDM8ssN8Gkjir4l+upoW4x9Whl9EH41p/N2d615Owi5UdNj+nzoImFo76Lw1+yKD6iiRxECD5Ys
6w1qD7T4T7QbXBjsjYDANo42PFT8R3kl6sfXynjxFYowiUSQ429c7fMAnOEOt4c9dqYf/5AqNVFi
iJLEwQ1jG8D5ApXNi3Z5U2pm+nby0Ey+Sa1ePuKbskL2nAxYWFDZDR647fu00Ta5XUV9U89eVEwP
hYa+/FN98adeepj7QEyW7ORJuXUv3C5x/JpAfo3w67NE6G04KRupKkL3+5txtUSmSpgkmKYD7MDX
90cuc6guSNi+VGtw5D5ADnCfOHmIZ0+o4jGPZxQXoKgdxG/70BwZTxTjj7bViiWnftmZYM6rY8FB
XxIC4IP1VsCCwx5WRGymZgMXEXOuJFfjT4DUwXIE+xtXvqTna8+ElJM+uldvvyhGUaAdMOE9ela3
8IhpJuvaV0O02h3oOQv/4RR/PmXgJKiMoBDTg0Hg7bnhtIETPdsxsY0rJjcR0pqgEB5q2xqY6PO5
Qky9y4jkViW07YXEIAeluXuGDobyxQSGUkcSFGc9DHrssMJ2twTSEibbvicEVS5GZDDcswXNzKcY
GnEC4hgZblTFMTJfPVk5i4S8C0IzKuepMhR7bw62Vi0PE3leFI3l01i4j3As7QpAa3vu2VHC/YbH
XKxNiXvRNoQyZEZi0cC/x35Cg8i2wE/VHdg0CrRKNRQ1kW0Bs7VDms+iLZZs7Nsuc11O/4fuDmBs
zQ9mYjMcwZ9yxu8N+2jktsG/vKtMbnA0CL7PFIih8wioQbmgelnxdtf7PrMoHPREl8POCC8fSc2O
4Y0vENUOMzKAakcDQCa7McWUt5Xblphd/lhXkO4EbezAFS1PDHkdHmSFMBI89qXAej19/ktJM7my
gDhMG3RLK/DwF9PIqRfR0ZYQotQL/wOxDuYRRT4YmwjGOwpUyWRsRLX7l3saaHIkDc76KYNO3eSS
i3p1qMgK7UxGrRXb3a4VSWEEJ+GuMV/9/X7AsOme9yFdP/UKbi4WvrVJZqmIuSlcqhGkVlqnntoE
51jTW+HDr0gmrBIXedXfeqsp0hEhP+k4uSl56LPGweqhwpXWjPmqBFKmK8IBacaiurTV5CMuir+f
lt/Jny3SdI+N2AfchfL91cxZVNGWubanto7NdXULAYIbCRZvoOHa96jfMDLZa/ZwxX0SmeuoyQD6
27nt+y8HBPITQpOWnQP1meVEZc46OfcWKHkLK+y7V1at0uhdvPgv+JH4R4dVCSw/qCuHWynr3Gy/
dBc/XWIm4Z6mkFadTt8BMN2XJiWRfgWfTBO4tIEG/KdfV8O6ObspAXO/qLbKAyRZd7tU+HNI8StK
9eBlyIPcEBoVzvhVPuvUuVGnaEw8EdtpfnmhkeMT9XHgm2fxplDwhgruB/48FvCyffPHRgKM6/Fv
39H1hxNqqBpjlWFMtmzvkkmGwmKSskSYCElQxbRqo8TswFnntlg3AKqUb8ZyXN5e4XLNGU5fMPkI
JqPxZcDj42EF9kauUmLEeYh2/qvbVYM4cmBBp6Ra9dYdby7qVV/eYXHlMZWOUYORvfjSD6l5nh/p
zbrzwzMlV1yhp1WhEcecO7qg1HIXCxu9fYxrLbBb1/cnwsRnkOAUdHWLgOBXMpXw6Pt4rdEeMzcz
t8UiKjBOfHGlyR0drfe1V6g+wBw1EtdRr/g6dnACVM7DfyU6QNR2ZAAjDtR6M5FPGbh4ktYZDfZv
vtfRnBpqYJsallB/bSeLUQZXJZKVSE7ovYPTFhGS+P2jX/c+kO8bcqocLA/OZHx3nYh28QJmv034
BoiZPR1IFICSNQaKNsNFFLWoUfsZlqsW9uwwSLQ0uNQpywJD4v9q6KfGBNgYQJutkLuey9pfI2CT
QyGbrC0HUdOYVfUNWlfgS1G5H0te/dduc8bhVGahZk+2TCf16P9nrlK6aO86LYtDxRDOhk6u9sF7
HE1cNCZBCU9qSkhljEt+NzM0z7hh+BV76tZZvhwkxXWvWit5yzSnV/CkRF55Ab92JQL2i7ktkSE3
1b++nsMNHxs8ofmA1/gAUPguYz1TygffCae0DjEHd7L2G16Vvk/VOVDvFCjb8dYybHWC88C/wtkK
YSfNGLwWn7Jt8R5oSJuMIQm9ki8jTGDY3nQuUdhkGIa5cY1yw+Naes1qREwg7QpoLuUzuTI44B/o
n5pwYRemA8cbXbD/Fju4Li0ixFnIKkYpizKM52XhdQ9g7GWFg5ahRd4oSrHODcWXK4c3KQx6rsA2
lrMA1nuNgfQFNwHn1awq48iaGilk0fYPqXV5gMqAWRIyi2etwrQOHdXjKrdR4Urm4QSGBfwMf12Q
cTDvHxJh1aX6hrsJsCPbodkZL43oFOGsmW7SYzlsei2M8PdT7dwvf0Rpl7IqQEwpXjz1ql15PPl4
F9JVN05e5N8p06bsoBa8SJKHS8BwXFZmwhS50Gs0dDBir/Dlbjx6i7PKIfYA4HwDbfCiZik4qTcv
EPlPtgbSMqJJ1xJczFsUG9B6K1ZkjoQfbpOMyghPTWmZPSBWnV6fvn2vzf962DaXELz3HeJOFq3W
XdFzztACyXyveJE3VK65pgBk77zHQ46BZJaVXvtw2nVxITQfSqh7pfR9AuN6wCKe77WGjTAzohoE
6W5SoOs/nkpqiCxQ5sTezlxRrrOzIjkGYyfB1h0ujFfcP42tkYix94O1p4X06b9LV661ZKFIX9EA
8q9TdxRn+pMMPm4ITlDvvIDcXk5K4mv36kjysgepRNpNmgs+hX46NuVo6h/TL03e8MWF203bHGsK
6L1tunKck12bqGIO9WxMqnCNTCjXTg0VM3dj43aI/JnahthtOHlyJN/lGWGN2FKjy2XhcNIHqEVx
J37XkVBJppBB6fVG+lGaX5xfXlqehQMC3u5jigSbc5X/dzQd9PAOEsvT+QMOqJ4WM4kNI0RWN6Da
3cbh7UnzPC9/QR/nDobmVSoiGQ0a3GZh2wc9V56wYz+1VbbfW/yzZ8coZ0uZVYmzBtSkx0lT90wV
UVXTIsSuw/bTVul5AWcbuEZE3cTMmN3Pz7Cf6gxBsyBfZmQiqLjAK+eWQGrUWVLjtDn+l61VEcTY
V8wT0dazEWbnzsQLQH6SVXwiSwM8kJKk6GvpbXwhlSrJXJPuP7KOVSPrrJqq3iulJU3aUtPL/Dmv
MFcc693D4VYs7SPSJwWt/ceNEpUs0u4kWa9op3o72og1OzbhS3gUKvpoqfK4F/WXdR2HCpup1EM3
NkfgAItp856ZvIc+OEIWi3eKijPQJD0jAXKY9Gdy6N6jlD1Q2il5oLHidSbApP62v1zzxNHJb6Ag
R6fbIQq+QGEbpt3DQn8+xzgki4UtnsUmKALhd7UDX05DFvkk7+axqUeES4mnFeTz1xp/LPkBNJhD
WEVbOIm1dp/cWlIRm+xiUYbZ+QHJhr4RuQziBtq01boH63+X4X5umHohQKp/HJkAw/+e55uopWyg
6vAbur4QG4P4BpeajdneN8kxcZJk+h4Nllni5qj6T+p+dd7acZaqWaRkIwrJarPZdjwYHch8hO1y
1RkN4ug5hijxVlb1l4wXtByV46crXJrWUoQ+r1CCM1qUuBUio0Kv5BLSOL7FuP6U8wEFfI4dneUr
oKfcJ5gPOkfo5XLLBLQgTE4NJrXKjQ0OHuJk8ZjciCrGOD8r+VqBzYfTmswzrqY21AqEPhvRf497
GpWXATgv5GeT1w/KEycMJ7WTAPchdRIIsWYWIZzBZwLfYpJFDblW9lu2PAYQ9lJi4YQ8s+4A3sgv
0vCOws7sVPQ4uOAdiqciuSuwUaaxWKMf1GruAGRCpvcFB2cS7EhpUwaLGe9TrqiQxBwsosTucMRZ
0muBLlVHiaMCLULDkZp+UwfKdJShrpjgpA+Lb6vl1gaI3gmA/Wozp/6aaNcZKKN3wwzq5O5IFUk7
qyx/Ne9nuvhza4AUIuYd2yPzSf4IeT4oHbkL6O3gORQNhntklYp8uLPIRIDRx+CFOD9IVkBD+tMc
rVXH0x7q5UOg6q+vfiM83T3rP4J93jcGtOyXnMrbTHj4YN37H5jmMl9fOXpPYFK4VwU4QtBQTz3l
II89QjVfgdukdi6nMT9cr+X78ggbUGbqW5wptj3/HPa6XH3Rz49jxohVyL9yLC6zppzPRQ5ohBCI
SnxTDt/zMxysqOi5f6gI9xpNqySB8VK/Y/QOwTkQvaI3ruua6WWBaQ1dICNT4vi311f27Klm798y
4GvG0fgtZ5zO+y7KLUk2ZZjdaI0aLBURTuy1TMq1wG1aoQe8Agg+IVaSoQmBcwd1H8drh08sdWtN
xSQ/AwX2QLcAqhoEO+iHNqVRuFT5MrdrAZPeWhHba0dsIqlMaKXiw1aQionxc/c5RI5s15c2yzUa
G+fjofQbdom8mlBvpAEtZnpQy2P7YA0zAhOCVteo2IBwP/EOlClOW4qBJvxLLmXzJCxa/z6nXtrc
mIEvioSFbQ0S2AWX47J4BQYwNMDEfbuxEhC1Fgxf5Looiu45olg0ArBSkVwQ0z+cLxeShgbOLdP6
9xeSCxkitWBuKVxoWZaVBUP3WKiE6sGmglrGuhJx2RY2fLV/nNBaEyB5G7asqtDqlnBWD4KnDIP7
f9XiR9NL/0B6cFE0IPz0LT5LdQO49ANyMTTBJrcrppQCl+Cu9i4LECctuyx5ci6jM0B0OpjfNZl7
N4XIivcJzIKThVj7OcoYCDtmfjKJ6VU+KE3OyL/EvE0L3fRrVf3t0lTrs0RZwi7hLw4wEtp++1j1
nm5coCRaYhvgz4+GKX8cPYhNrVMoKHIbmVtyKT7NM7wZc9SxRTgVWrmL8JoS6g/ZQ7idd0JQcIE6
17tk1GZiQOmy/mm3gwjLe85PaXbubZuieuhfqBp174Sr5cLRmZy2vHkJUDvLeMaTykzyb+v2ITec
4Sr8H4Dr2wB5XET5lhzyXAXLR0muPWV9oxLgP9liqkamyzEBl3H5CHSwCaPxt4itx68wKGjNiMP6
+6h2r+tAC+vmfs08fab/hD+9J0R16z3tyiHyPdOmStpd19wSigNoZVWySyYfWdJwsEXiFxQkpc/I
m13U1CDiB88lZiPNtdXFRepwGrJRSsLc+dAgi7cc4uk/oq/dy33GivvypsGKX1vi8OmhzlZ44afB
U90vqe0xIJrsIeeCSRiYPA3Mupod/HEa09zK9o78zCUGf+2bGEfB9k+WQ3qzSa4jjjc5PT/XSu8T
G9DIOJKC9JA+Dp0ljTetagXAK4K2pcpnexDPTPUmXvmFrFwruT1w4qAjxpAO+hQGwsS3s5ktZc96
QFaGPkc9nHrCV37MscuuY2TvnldtBOHFxfc10Yy/dK/8gmVpkMEI2gJYnQXB0Z4lY0mYMP83TxDY
/svhQOnh/0RJF6O7VRAYR8EocZd918o0aLFz8lOE83WzxB30rrDudI2ibxDF5xvBp/kmrKmJe1Pm
TL5I02xTq1hC+jRiVybmZBrNFKmlkwEFc8sUuEv/D/B17GHMXc2CK0YpRwyBTh/tW43ZSESevorb
8UvU+UVD4VPo/fk/1VHJe2miStRSjGsWhIEUPh7j3NBoQ4uXtpBG2hL8p52+xyV+SvkubprZMdtJ
vL1f3FwmGlL4dN5asqymPs1yJckjHzYdRHiv8DHoB3pbH6CRF8RIbF+KvPmTcTe522ehI9IukcSX
NMSNcjIbWiGS97aqlgGWO9VcYA/Eja/EfBHsmKWyTdaX/XboXXFfH5GaKdDIhnKFk7LYdw3/P0xA
UEjIvHHpBE0qM1+bWYejkoCGaVI2woUiC+lHtoGuZ0i4fmO2WivoAQeefXYvF+ZgL+K7chjayPM2
8UvxIYREMKDnjkcoy/Qi038cSgsTO4l1KwWLPsgdneZ0byPbd+h9A81F5YKFqg2+F5PYfKfOw1aS
BI5ljXyQYTuFPtwRR4x43QIweEX9+lW4iHZ19AuZyo12xyoHSY05EJvgnvSwesLZaoFLdzTrXpTQ
nlERgkNmE+NWG9RdszRdJyo5RY6kWDUmGZX1aT534IFBrSK6COFLiTWC+XfpRv6sWR6YdaXxfYCA
HHhY83uImu9t0DRQHc11u6krdPi6FLP0AeKRZ20PKlnHApuZq402GEtwPnq9sTB6lMgiTL7vmP3k
MTm8kLQO8kOiLIQADSCB/ekSnPUKAbIyl2f7Sz9ZA2IkC7nl6T/kNprjhXU5yrPJ++O2JGQj1VAW
BE1pjQL4T0AZShM2amq5dXwj3WnTYt6yMVPa6C4EP8r4EEVafrgYKsfLsyT6fs5fdiBZGqtDZ1lj
LoLZMWxt/lLP5oMa2e+PAVWGbhsE/DLbPXQxn5t1X145gF7v4vPoRP6oMsI9k5xczEcie6wCIBjB
D1SwcPyrEExUPQFOGiGRoMUOXhWkW5wZzWmvw0K27hKQhS7aSKTZ0ouY6kh7R9dcl5sQNRKzoqnX
x+BYlSk97mryIrZQYlRkXKoaf6ZwgI83YE/mSvhmpuT6Rq6AxM7JrsTDGdbQNV09YUAp7jMS+rKq
uVHAAs5YK0DKU6SzIxIBG4hCXNt5+BE5msYqB8mhidQwFR5X8jXdViotubLSVbLKxee3qg4fAOAa
5T00V6UlhAAANQZawVIpW99p0t8Bagk2DvnzsxYCDnYgbhIc4pfeRLq5YasPAZhR84FBAX+WkZAi
jm6cY2r2SL943bc3TMOBmQmEtl0vbB0/69+yq9zllNtRK/PtSsqpXE5VDdFYh03VqN4tTk9Q22jT
o5VCJdWymKFO+CygP3URWp2AV6lvbqFmmpz079b/C284e7QGsj6b3ISrRQRi+1PFoO+lYqSoB8/h
LNj7PgoxiXoJjWItUrmXxuvefTy2mCn1FVqI1qdpbFSd9bzVabOsJp4fqi/+vBxonnN/fLQgE332
22FV1eU1xc2BK/x4tke26gp/UHfrJjg4MIW8Tj8c4vo4p+JvRW7gWfcPILe7UlnYySNu5cJw6jFb
zJrCIXYwPoxaUxj4Xca+BEHROF/fq4KrzdZFDqiBxLxy1ZXKoWebE4unw0SIwMh6AHsREs8UeEnA
FruaKsozzxtTajyzxdGDI8rOE5LQiEiH4mht/D/WCZKyC8S0nVqmc/UlfpsQu7zYO0nizsQBfjwD
KBHSE6AdLJbkexokLgPPZN80kbH3nYNl0Nd4tWvPWbXQAfzGLTahFxXQXqGmK2HiriUevHeYzn5N
Kk2wmVk3Ct9fFZOCQAxcaDp1287iqRZ4zylUCtCsIi5nVtG5yt7Qt+l5m/GLrzK/VtSoU/vby/Dy
ai7oVLBnysDDGKg8vp/deMF5quRaDFtmazf/rGLQUEodefCn4ImDheTLP+xOyPfCiyAyuXaFr1qR
bmFEkRV6IPoTyalVhsphLwOJPnI7U5PXchiX/Ix68FfqCCQlvTByVszbU2FtAU4HiP6N0EaG9rHw
or+c+fs7PTWnjmkcESHh8gX/P4b6mHUqTe7X7pbKfjEgjrGoPT14glfyApJh54U+5ZfbAzgc0LW7
ABa15gzTO3dv4ra9ecNEAXYnuscCcpaDvt+9UbVucN99PQhDOCOV72qLq/YdJqMnp7+u3CwFa8N9
uDfV9QGMTXoZ9aIRrc6qP5g9py0F1J1moMbXnlCLrVBL+H9llxCf82ej58IpY63u5Ge40Tk4PGxp
K92iA6DAlnx1w1ziRMXsatL8cBgKoXrNfN8bUPLscRS7EkU0/9nbD2FNm3kY4j385yjOBrsvlQ9c
JDNWbqEPbqu9RrYTxpOe5Dveg0iirs4v9Nk/rw2LYtTKV74YOb6wEP2REmiqAO95mpto7DPq3G27
hvGm/M5cGhlftuoSwjJXnxnM3Qk0X8SRoD9mhkblcATPnz8Sjfj0G4IWnGDmizyAjMltVIKgqEI/
4VMckbJeuOSDxiuRjZREjmmwGJ6X21Uplu5WLfwQIPyuLs4uLHQxOSiZf2ahNfrBTJJhZ/uMUhE7
pUrIOVlDsMTjt1OEJ1S2mdWPNmNnKs1+15MvbdS+eZb4tEyrhFO6uLbUdS1nYkrbDixwQMt/eB2r
QZHBt49bM9EV7ryUM6SN/8s9FGscvEV9nCU72jBIYZp4I3nkiztmAU8RTE27vU8Xms+YQJpIBMXv
aFahB59rdcJmuqS6EzTy4nGOOVzn1m75wxmLtxuBueH1XE6H3Ka9oHlDj8NUjxMJBaoGqOi1DDdy
sD7mMR0fDQmdvRDB6Onc1zk5Qmubl11l/ndWQlkSIwSto3YNmiqFTPhHn8GduJ+/bcx257qVkL+K
C2ZFSWTqGntAO3Nn9svcKa51T6/zhqCH2vynR4dwsnhioT8klq8Yys2gyv9mMxXmEFaDjU+TR4Vq
uOjDo/Lfan/6bAqjw/2WND4Cg5mpvWM9YsfTyXh9t90QfcL2HDPYZvCKfAJWYNmfHGlHJOlbHOmf
NtlB2BeHvfYgGvxw5Mm12R1Navr/ImeEBV4fWWNJ/9plCuwi6Nsen5HjmvikQnYFhuJSnrchHOdD
IGWGGMzasS5jhQ7KyZwiOtUSjkWsNnEgmfsG5da3ubPmDPpMLPGh/CERcwQ/xQa1gHm9P3hlcZCb
j1d8GM/K0x+kVnYg4huAGQJNUgpFmg6kV7BQTUvKTStOwmOEp0pqsYcOjKSM6IOBxXYbFaopdUzg
bRgB2aQCZy5j6FJg9Bkh1zZGjPAEAKG+V5d5BzsH0Fqrzte7XyCzTPQUeWd0Z7yrnjUPP4nZv02D
bOXvwH4ArtiB6vrXDb7zIgGHgESIXr1S8AIP8l2Mw1BxdzlpgVvcy8WrY8bHxtKPjxXjDKosxD+V
Z9skBC1ix/an0GKBA5YXR4zSFWG7dpaA+oul6ciNWbzF7MlyJOt2fx9IlB3UGXaSKeNkKpj0qD5W
20D/rwVjbF4KCiAu3Uf5Yphu/AufY689LTe5PQQcKC+xxOSKmL1N8jSTVBWHB4pE9brlNiMc1dX4
RJRzjDQR13l7NIj/iNpRvV4U7410kTxV9clP4SvW8HfjR4Xy/gGmoqbHX+aFYFGLSTXvYFv0IcZy
V/zBXh+MDUnUZzP4dSccljOT1u/TjEMyvzVmxqVcpdeO351rammNLTDDmHenszpD7AE14BBkP0Xk
xDFUF7Zq4IULuNwIUvY3tYvBaGaVit3p/9u3jQUG1P2Y6MJ7d/6yEQ47P3wN+rD+EJlqxnMiBtn/
4+cYYehbCJ1ANo5RjZ3NzX+cIAccTv5nCLfXxC5APmD10JxR3u0i7JR9P3TQwWxeluVt+DNbRQ9E
Vwss0kDD+Rl7dQJ23bROHgNIvDjCDDO/Om6g3uDst1rQNREnLgU0Z2tTEQuVxhzLu1K/uvLTjtie
s2/7uXFderiKkshXRnyx9ITAhEU7pNNkkEAX3U2J2MBrkDmOXf7hWwkHXX8oC2Fo6qnb18KBiCyx
WbAPRESin0hLKBp21H+SLjuhSKMAHzQbQk69CZydKXPO6exXSNQ937j8coFPdalXKRN/N4Zyk2ZZ
sOJkNayxbMerWKQyQ8vLRI6x8gfGXR+4ZQ0EhEkKSy9PizqSBT0OI6IrC4CzWDuv1ecsT5f95MdB
ssRB2BNj2whn39/en4ha3Zrpu0hlBazJ3AhGSokbpbg9+vm+0W2BIsQu1PbmGoKg/+ow3qNHtnkM
jLVFMJ1NhZ0xbq/6qn6U/lPfmOz2xxAhCP2QqWYGyY8ag3Jg5xN2yKMNuwGhdkGPME0AP4kXY/94
FOyOH405iFCJwMSDRiLyHIK76Ldq3JSjOiiZkXxBZkz6zPfz6uL6xKoT1i+X2rNvXreTIg4tp7QU
K3IQKoMJnQCpBJ5+Kb1yclUFfxD1CXvaoyOSCfgbBAsRoATqOQQmQPRJbDZAoIdSavJVcI+xLHrr
Vm9ESy4+F4yFiZ5nA8blMmJ2/Jg0uqGBLzf5lza1b0HCSogdphMrf/oERM/+GpIMEDY3fjK5+Zmh
Cj8V+LKv3LZ5YJEDe8w0BcDlNAHhuxEhJVIQNrds/qgKYewthZaFIriAVSWMg22OTREjjWsWEuuX
vaOAXLxHQb89V5m0/Loe6+69aHBnEQVcIxH6f2NCcS0jwadrFCcJPUY1Xfm3aO5pkXOROqU8uNlk
/WwYfgwj4VjC0Tx/VV06z3eslhN7NeVfkQ5SHIl7H4/5zZB8KxR00noYC+l0q8Osa2dDqW6m5xtS
ASGIYLF8nzjcsnfQN6JYZozRY4ZRAGffjk1Oe1AlBalJ0slKDUu9uGBCQvFMXAY66odMBOA16Fay
O/8x5cIPkYchEzVQBch/2nNaShQ2bD98uBgOpBukZ0j402k7513KbnUbNmFG8I5IvtMCOLTbwCjR
yEvwrYtKK/RB4wD8W+CeNOV3K0lqNcMqsSeca1Pj966la+dy6+6baTHUOYVgINunxPhV/j/NvQ9T
RmJudJEpcAzcaLNOJ4EGcpYIU0h6dSjBkTPWe0Omj02/kG9rgvI1E0d7gj9RTiER7sioMO3TeJRa
u5gJFaNxmjCwo5JT1Jt70ca2q3pt9Mhy9TbcbmY/x4AjrkQSN4zVfRmYjLdbhLcJLHF8hQCoGtIT
kxyvQEucwI1PGaMabvrcyxEbscOLvSpA4zJ+9kA6C0w5w7yOuq/GVSfg6jhC2A9GAFoctcYFD9sw
NQwvTt9LPr5MOQaa36UjmX8ioVH8M07KiwNcdISdaG8LEsirfWW/JhRhN7dhCJ4b+EA6IhvUkP+W
IND4HiTBQ/8R0OW0EApH9Rk2AtZxm5F4XEM7zovhijdoFEfWltKXo5lNwDaIRM66NDAs+btg30wF
8CemCnVnPnSkUWMEgbdIW4pArhwv6Q5Cgs6V2O8HPsvkwftKXHdBOMoKH7ycwUN6GBp6UBmiLwQ0
hcf09pYdZzswxeWxIkO3RdeSzB3msbjzXRV0ID7480nG7leasSgcU15hoINiMo0VgYFfytXsVrIg
Kad2yyXKTCLV05SvHOQpCODBW1QfOsw/nIMjgwcUNueD+UgBCbphCt7JyT1/nBGI+WhSmmkZgvY7
6seVZB9OcuqmCEzAKbRJqGR+4qDnAQmZ0ceN+Sj4ZPghgjcQpMi7sV7VLTOq8LuqORz/PAXuLqmV
5pYcc8xra52LAx2BL2dxY6aM3a6WHhTp3lqj/iDuGn6CfcBaRH2YoQv5/5h36wiQpMZK0tNiI7NX
HM2fGeqAiNTJGp2npj1f88TyB3GvhG2SJE+0ZX3AiqDv2dAC5Hobq554W9B7YGn+aVHdtF30zRUu
SjTPqnQftI9BiTqeLbgfU79U1F3wUCHFb4cKk3UsTkdMRzj2LrktSNyUkkphTxD2SLvxWnwv9h6+
wldPByCQ+OEAgbYDIhlITzviuN6c2BTGxfgD4rM8DkkSvTbMKTEENDGEUqKGWpU3WpcisTCG+dsN
H6+sPMZ7MXM2wL6wenuFNp0WBDzdwqHcKGVWBM1lBzhBaKXevLATWjwD8opay5Mn2uOueMU/xpaM
x+5NYyeUFUfA0TMck9iz2Kaw+PXrWYVqf/PTtFiT9V1BzhkW5q+3lCDoAcE2UwI0BjPPcQsjTGPG
lNQSn7YPULDK2zanyXo9OvCJrIXaYFNde+S7IpbDBqZGMgSuWxU6P20NcPYO3/g7BnILi0pqse6g
wD3i4f3TUVUw/BfG9PW/+qUUfxbzPiLGH5zlvL21b+UJtsfRaStCH0ac1Kz2U9zBB1rPH/nsMSvG
yu4x2/THSZNAJT+UeYcW6tlPmtNiH/fq5GMElq+NeRQm16ihLKBu7bJwHYb7B7Lw1R/WQT7a9P4A
b5MOPRb1nNID3ZgQt1PgGb1hCzXlneZ0Q3RERjmBjx3ZB+tv6Y8vWD51eD3lJr/KJTuPIl5J9cXq
ATy3gQ8inyce4LIrqao8OKF92PBGRIt3H4vZV6xgbs6x3SZ6UjD3/MJ2IVCkzgWai3GpaEysOqBd
vkcLtL8yrMJZWk4QxJBB/kizQIKeDzekDPgEggb8I0hWPYuumg6fyMia/ZvaIh1uZF33ZQ+zX0Ul
XcSI8593s2LBA4iPLfjRvBOpUTT5AGb8XwS4tVAIDx5Q7ql1y9n5FGzhakMTFx9V5pDO9UOQBrjq
2bFfnjHa0Jz4gL8Jq6Oq8O642Xv2MwYIA3WfAJCFLZExpY1AnwjeltXZA+gM9U/yA0PQT2jj/rTr
J5MTQdml//siu00WSmiJdk+52Wi7U978KUI6YITKygM+AU35KAnEc/HpFyUgmmxGgtXFvX2sTp+g
VmqXTeAipLw+9NDuMElC7kYbUPbhrQPj2gQSqwbYj7ERoQfPg0rERP0PwwFrhAXKVOUQnl6+5+rv
igo1UJli0HvRXlFG2ZqgaxUitY/ZDM5RcrarGt7ipNahvT/6IAwk8Apk6tqpciG4qP7icTvZTeYh
5pWcBeja26stJaKKZSoKSemr1zsbNu4F4MpzLIcLesj9rTYj+QCFZT+sg4HHRcAl04mNDpVD5XD1
QAp17ZAYXVDHIngbfsa8H685JP/F8TrJpDEQKf9F/xSDC0Gnvke3BhkV2+R6LzpgX8yYHCmaHsLY
SqRyTjgNInUZt2JCKCzv/+zB6k6A2KWQ6nDpiv0s+R3MiC7zO6tfoi4HEkTG639FPrXrll6iD59d
VpohAYv0+KLbagUVF+8HjR6PN5GZMDDUXitK73k0SBe5oLM+7rn/DXyHLaSfL8SD8v9a540v8JKM
WVw1DkjK/81r85G0dB7JLOdjoXXg//UEk4sGt7jcKm9wTzenI4BVFNsK8fDq4XJ3KJ7P0aYT/H2g
wXJJaxckw7xe5eb6MuNqZuB+Ra81GHEUqhRhsAmadX+kJ2uabuoygWLlqwo5TSXurJAuJGsaj2cg
iZEVmTPdrJL6y0f6DksSmJdIqjeTnXjJXwCcZispvnEPHc3tJ2hrD/J19xhyIxR8VcscpE5Hk0LJ
e+daYu/qnwdLq96qHfYGH9Wum8RZorAG6oetD0kC9pGf+6Xjw+CWjaDDe8ykyvbXvnHzS5v7ADDN
oqX32GFy+Bm47k5WC5Zc/epu+W1S/y/wib4QFdpKpKLI2epsnR8pqaGc+DMVzWkPgrdxdSBKhG6+
TH7LI7TiRrkzgBt+vmdRVls5LfL0ot915ZfiB3g17uYt8rARV6mq44T3nJHhVOROoRqjUzI4dwyG
c2hTTRgQXKrUnm5pTFefS4OP05sie09XP9N5hYp06o9cKancCYBAzMWv+JCcJZpo4GgdgPWggsdG
xZJATNqbQIMTO0TPcDOAyTAmdej+jgsq50CAio73oKL9WPw2/MrMrRbCDP/0VMqJttAHzY6qOIuk
BtyZ0JZV2ppH4wbcLcRagLG56MStyGfGdm40L0J+g2um19h59sS+Bm89WwX5HyspRqBU8xr9yMUb
kVUTGGHaODorO0PtBHzbasGSUa4KLtYZ6OA/svBDwamsx93V5LzzZ5FOAtF0w8w1OY9Vr2SJyXej
qYTyEPgzOVYiFGD3FvHH2jJu3BTRzsSmDbieYK8AtAfzanlUZSky/9DuaGIPXr3/w4/SWzxWNl6u
awzmrJ0oSo3MTn+Wsps2o877pqwhTcWHxXgBcNvhZuWpRbEEkpgSnRKRf6kn2KVHmn8ZscI3xpHr
iXx1BzDqJPu6YZslU9UdmOxeiMwaJ71r+pYeJfp4gwtJ0MYXoNSm4naME/sT0Xp16cttE0noSaXG
BczJXw2Ke3O0w3Xj/ZRM5FMp9LO2vb6sh5sdU9eWWTK8I3gvMExI2ycMX66KuTtbeL709gmk0Xiy
tGoeWs2FSph3g0U/zCFg2obSF9OWeZPQPu6ug9sCnndX1CtJJ+Idoim6iZTqupBvGFYcUep3VEoZ
sMfd8lMYMvJXtu3ksc1pA2rOysr++nrbWlVWukvqxPwXLL1xtPB7dNLNI1ZCKtZpd9lmxpVZVJPb
CYmT7dxgQRy5t21yuAAtOz6dhdh6P4l0+wGy6OktDXfZbqXrMzDdT5q1kh6gmqEIiwBue3RD33+s
up/8e/KbLIcr5IT2Pdm8KL8kXKYWCWyAp7W2cB743PbDc23rly4Cigi1X/lBknusz5dDzSxmWbPa
L2iRbUKLnsjJYo02MASi/7uReAwmWrkX+Eq8rmj5xjYl7XIMkl08J/+J3tU6PUWLOYsggwrjxQ8r
SaNpApSzgQ0OsMYp+Gsgi5wL/j84t+gfH5nE8Ukx8c9cSCXmTpXMXivIzvKPKds4Pf7iCQeaMEeL
9zgxN34heRQ4Ic6JoZN4bbgakcCBIA60eDAIhHFflW1/nyRi7jUt9MSncHiFFJtRIwuDUMPYnxxW
ExDsd/PmsxTGVBxcPCh1B08YoABuZ/SpM8iShMnByo7ysVOEjwbTRcy8Dtbv9U7BV+9Bc1NcrgNH
aWBhRnXxcEHVhA4GX5EQ4Jbmo1h5MwAjNVO3sbSPydsg+5+7iVT2qxVfsjVcP1ZHZGJQjd/P8T4k
j2wBYlHxQimZeWgVFL/9soTew7PEYplo86ICwjf+KAQ1gZeYC/8D4uJucZZiKOf+/QloLhT62d7+
ilzfkHPmNJAL41juVpzsY2TBpwagAd+XZu3agrhO/pKsotJzep8Xr3TJLQwKPp7NDDObcJdoT9o5
/2DE6TSFDWwDgOBi4IL3MBdhQjScR2JuwfWQci/KQgh8ZkEOSFAuS3J9ndKnNpfFVyTs0QBEAPn0
48WEc6Pih/C70pzuNttlqaxV+J3UrjRY8lLloWirZ4nRKSbX+XPo9g3kxOt++fHOc57zzoWYSLMg
K9KGjoHN8o/Rx7xApBlVFZh6mm5SLQ7fdqP61YHqOOgBMMnh8VwPpk9bq/P2poiGs70if9HG8oPX
l7jeOVm/okVbvJroS4U7nZlJJmLAZXY9bWY11YY+L0IpQYpDerCtGnGipnYiVXGDeo6vsI3cRh5+
/F78o8YaG1repi+N4TK4lJgQtShLAG/UThI1iF0UKGROK5LGJ+5gjbnDjS6SHYRAqAFOZ10ubcAS
o0ks/wmU3QtSiXSyiPd3/c+3g9GoMyAXFWE2UKjoMTRbXbeSMhx/5v+gkB82bRoaAZD4kk+vn+Tr
ByZbSZ979jUI04nvQBcPcby/mPczFSoNCRWEcfEGSijojUlOi3YtrXT7ooMz0KpKv1+QvgPywRHZ
37ca/iGGgNVXeSJ86gmSu3DR9v6Fw77/1VCfi7fJLpGJp0Fu1FirwnM/r6yn4B9VHRPS/qc7L4aK
aDT8H5RSkNvHZQm+cQzQdfqTYmP3u0CWSQcStvmoQK04SwcGd+SRszt1Un2gyoFiTCa5wMzBkUu0
qATcB64hpERYsM4XfKylBoE+7jPm5Zf7l5Yw717muyveIb2l3lWx9lJuXyUG67AV40sQrb4L7kax
nLhi39B0EwiJx4Lh6kYTJRqa1MOa3fuK22bOULeBEq/3z1Td494bn9tQG+8+Yn131VZ9lISUEG+q
kLtR0ZiJq5lHzbiUJshqDsaRop8+nvZLovhxC252NB4tkyCY8U+J7bewY8dAimnoDgigHm+EBX/O
kBw/DmK5jzHuLQPo0aJlVu8nn7l18yrdDP+xAdO61t+Rim1zG5zipSl3K+hhRSqaLuqVm508FvC5
1idQ2nmtVJsj20sDnBnFaxwbh32NQbgLFytyY0XhhHskCAS0n/NasetClmgPeXeIqTRjdzNuXv06
3sCzdqiApjvSVwipoIhyl+Ayz8trZMW1O2BHc2caFVk1SunYn0eGZDxlIqMM5KRX9HsRhof3V8kp
6es6JVeHQG+tOaNb6RV5HkTJmOROgChzLCvf7d1ZhBBQF0Y+0ozJu31Q453aGHfaLrRH9UD3T2WB
jxv+WZk5b0oYvPNZej3skyCMPZgOVdRBHV5FTKp48BiVkZQpVuNP2r72dbVubOTz9dQtVxytoZY1
ihOkiKG3TEvZE+ulsPw1x/p3zuzf0EUwM1W5YyEoToqfOIXhaeAErdbrF6tlv/GzvmqQAbrrj2fg
TH7p4krEDSW6KjC+wRwGmubbeJfDGsR4nG86jTPV11Cf3HDl9QSBJIXvNsVCnXI0L2NzS6JHQ7r6
m9HMOd4AOxmCxV9mIRnIG7PWkaI1G+yIcIrb9F1uDpWcenX0YgG6K66oZTxoeisc0LTf7VAvUjns
ueCTwKQOlCeA9fu+35oat4/8NNYHiWCWfcYrqoPJc49rILxD5R5o57kUVS+GdCCP8B9kFWzBDyAt
oR6EToGci3NQImp7LyItn3x2TQu7Bns1G0glKUTqnAbVrDI8bvpmDFJaHwq6yFfBGCEXfvygO2gc
zeCKM/YpEzp/Alz8FVzAP547fGtFW9ru8Ibgxv5708Bzrp694jY5055YR5fkJrcIwkEqnyAW4cCD
s/7B76TVelCEftemoEHQrL9DOpZgGruaP4PBU9rt9GI3g1rIZjPu67VeDJ+pgupjJFs8yVas7P/x
1TdfyhR8fUpXfIbWsxuOvx36WTujMM5sdXZivONxQYrYXZZlW4rzUXxlGZ8CX4QyONm8E0NG0o8b
auhgcGM6B7eijyOr9IxOuajRSZJu1Jv9Js8/FhK7VT6YC649ehMY3ZZbSeviCHjuCBD7K+qh7Gjh
4t+OovFrasFv+drNGdJlolDSdIGHMuXqO+vASEntIcJx15pKgue6SxCFzJCI0QTfbo7ywmOCLq+x
DSEjJciJNyMnsMH4dNb96VgeReD2mrNcqI6+UOfkvwMcuSykOjUn7oyd0xafNr4+Mdqx5kXep29W
P4FyNwtyakTShqCMfZ9zdetfxLaIeNWZ55DBQU47T48awV6WQLOUhpq75WKWN9oUpkXW1xTI/aeK
gMf0G8WjKqmCiuJftetPcgD0mZuYHpNKr3cLF09bY/ufgGHUfRz5qTuF4M9aIJ2nI3EjLvXdi8Qg
Z7OvsUu7jA4lagXEAlSkM8cGqU7Or98QIhL6VaFLlkmmad+iGTAuyv2WIPABRZwVbATH0FGM74uV
Mhtqryd9eJ10V7QeZ6Ccz2wlFpALCwEqWQrdX9l0e/amz2toDnG55A6/nSEr1p9fSKvL1AfP06eT
JFHjSmAseV3GBiiPrQi2iIyX8qHJE/Werh9tEyAlP/XQm2TsjVkSOHyH+Kq6KcA7nX/kMXlp/ujk
emkvWtAsN+zBH9Yp+ZelC40F7SUuCYnIfhTOfsUdEQyE312rrGDu04Am5wwuUVTEG3Y9YIn6y2h9
A39vfqn9BjU/Iwbz4Ch34Fyvy35nTYJg67uoPXLYtcbgntFrVh4Ble8HdtKmcOKKiQpvb2qaBxCj
DaR9emyetqDHOgUhr4cvT6N6ZSl2nLdaMHBs2LgVrkMdJKk8jdjLCKRv7HgzMtdFb/csvPst0x0v
cN+XzZqNEH7OuS/vZYLjU6HASi2i0O4DyeKoLjpg3i2/0qr4785wMHf4i9dQC1ceHVBXHVRk5P1L
pbkIuXaeiUrcxanBA7diuKw7WGW1vAKtaMeRSUhPxVtHfwGVMFtM5GsM++eRoijpyepzm6L8RLjS
/ttbhFaYxZ/eiBB5+mPtjDUGcdyOdPr5ZFJhEeSdzn6N4fIU47WPUzx4sXi60OZAJoShHjcLT/to
uzwgUzrV6wXojiAGAL2nG5N7INpS43kImYK4XizVfkgvvX6bfbk+VTUT4kg3zUYkbWbPjzd4cLjF
dAp0WVnUVgmMV7RrOsorcM+P4phG184zG34XCw0akMAm4Y/oTqsrJJq40xtnBLxd72IdvK4XJnbn
m5bteW+EFeuCaF2q3oLvg6GMhArd6DjlhB72g+wuSKi6XP7TEcESUNyRNm7quQi6ZojMFoC0ebdJ
p+41v8vUfinOhyqd9FUgr7Rb/TN/zTkIMAjBQECEs46Kbtg2pRRvwU4uG4KPxlRIWhpjsDXj3b/L
YZhxP46qaVsmH/u/PQauSiClu4m43K2VLTUECBw/j4cAHTDZBVJoGBXuNmNmEduUisUBb6GAg5L0
IiYaCfhnGyqjUq0UeqwnqMWKPEpgb/89pIX+QmBJtROmzeAcIWgc+pXDk4Wdlt1OfuncqhEDguh7
d61NBFbhTcgGk3biMl8/KTAlh8KdY6FYElgXVNoskR2UNwIrsv/oD0jOkx4Pu75HmGxb+ktWf7E2
6H9dQkN0GFX3IEbHNGKFQ50Wy7mf1DJAeRHwKF2qIvckIeoSllt0K47MiVYhKPqkEIrm8Zq8XUEp
xSdsIhC+6hcmnFI5DitGDPA93oAyzq4JUHQtc7hlUgkNzkEsI1rzvSIS6ijpD+x5fhZWK1hGHy4D
+MFjewI45EYjUcELz+UA18/2B8joF9EqsmbTIvH49IBAcaNc61fiYgXQTxRWED/WkVLBzmIXmnfu
n3+/3AJpvsDV5W3zZTx1wiB0qA/5IJ9R/lY0IIXPPT+InQGaGS0uIfSdBH0Tdo9js7wE8yO9sVq0
Td/Chdb77C51FDXQduIQN3hl8Aio/yTKQrdyye2uymbIXtpPz3pa5jdU2ysxB1+JcGlHe+pHBd2+
IHm93kkG/U1K6ripvvjF5wrwQwPYNyGIHoGviqpT9f+oit7mlD37fRPKim2O4gnHCxMtmDtGSHY8
asyJsU4UYJoSmIgD3nnsZrRYmugfHlb09g09SbOPu8O8B9sncb/usUc5P2b/l5Ug6eYcpt5w8bLq
iVFOljX6gRML0IpwvhPXH0e8cTlfWSCJAJHmvwlQ47bJE0KmZZuDi7ig+MhSzub5krmxj7FLhITP
mGx47TTQLWoNOK3CLVoQ7W/V4zhVLf6NA0vjUp3kZhSnDrsE2nVcD83IA9NJJ8dxHn4DrPp8kgih
eqPFp2ml8xK/YnnfPh/bbQHh4WqSKpUt+cG1uSs+x0ChUJGAg4mvluAGotDgaYp/wS9dMcUeGJsN
3nOQC3SbOcoOO4qlsNOi7V+y8gpijosK17fsdaWyaTE0PYX9XLLnxil2h+aWSxa5TPp3rum6J/aT
uTlLCZysfbeyDIFm+QVruHue8az60tQ+Dd/VD9W8Lxk81eXfRQ+gFze8O6FTw/n/MCCSapgjZDLg
JHvWLhXIgTQOw5ETTOWTxJtBfQprX0WTwy9FmF2PiG/YZ/q/4sSn0bPacUgGwTbJQMDdVuBeeYv5
97ZgSF/UNO7DHUJKLgc2Csrs3H7VbCAup/xrnSszf5ZWZ6Gu6wxn4jTPwSiG9l5SvvUod6XS8gpE
xvS1kfecrPJFXDXVnkzx7ql/pd9jYDT86VVCpRyiDx36w5cC+G6CmK8+VSs8C3SQYJMtBhtyyX9x
BJh0srSzeYNYvv/xR4R964b2fuDyiYICEYN5HkcXHPNh9SErRpBotnMWthWi1ZsstrH+oxL+Wph/
U95COCa1shvL3eUgUP5VF55u3fdRo/25TWrOrOmtaHsB/G0CLk1y1ofWh55B/x4vrHvnW4xlfU1C
qUJBDop2fo+OYbseS8+1l4NO9Xr77HneT1z5/iXhyEYbAh6RpNNfVxzvu2BMVerYDeiEOF0NmgvL
7MaZNppqrmIhOtAcBPBjwjPj145u//dRY5gCXBa1qyEgsGhrFZmQ1A2ITToisJTn3uQr+9ZjONWi
Hh95ySsk3hMXOK83pNRnOcWZBSRfIrCc4UAsjcM7liTQ+ijNQVDLzY91gs2GzRUbt2Qx3J+w6zGE
ULELYxeW0avBzlULtRyO0KYEh2E5W/dShleC/8YOwoPqo9+eNn/gFaz3h7dti/id+ow1j6Y+dJXp
zStIKZrUJbxBZw64JqQWLC4sLU97MrQ2PmmBAsWyC6dp+iMS52RZYcepMkoLO8aYnvLTrjxFP0+L
/bxoxmZwjI7HQyLyb8CFcdFed/puZx6sjDboFVxSqAR3sLyUpnmLjmICyhy8xCizwUHaqTucRfBE
SXPjy+SkB2ZuJAOUAm4PhcTTmP2Rmk6iwIy/2agS9qPLidZ9He+e0TSJAwesd4l6pCtkLL0ts6T1
ljQg509VLlimXIsl0mfax8ejAmFGhdimndDuz1a8B+rmRSKuV9qJr9tG8lZ1zCobal2Zr13qgdPl
dbvrdiSqFYTWNq6WK0Wshei+uq2lcT3J7s7Pkla18k/A/gD5lumbFNKawPIm8l3T09vGdNiTQIT2
6Igrap1iKogb+0s3XkzJsb/JYL0/SrEsREAHj8qL9AXAlFLgYKQWl8un9VwcU/XP7kF6N6jLFMSX
UiTGi6TZQQcQI4B9yQM6q21fUKH8mxt9UIEEXjRbRHRmjIJ6R53QO/DmyJwFfHT4y6nlIKN8LDYt
dEvvjR77qL2ZbJQh/9SjsuFiKQhDgfymYm1IaY7c7C9CyTl40iUJDeuaU23UKrTaXBJ0fn+15J+p
DezT0OjRwqbrLYIGWH7QaKATo3OvVMREs0nkfo0giDyIjbPKvov8xyuWK1BYvDhujviloV+iD+/E
xYZHSanItlgbwZIIsK3yvKCCtu0UcE776lXjYXO19c2OMLkNTT7oPXuGajbDfHB3/Sju+C8BM4Sp
EYVyDL1XkEzup/5INhzc/fjJdC2AbS43L7MM2srz4qc0plQLn8PQ9BVjKsdg+kdwnrOfxAESAVJ4
iaTP5oKSiXvtnHePRKMqjWPkbUepMLgsvrWyFBQi2/gdXVk9YIdQCveysgaoUMl5Vqm+LAm47n38
eAV3y3vHjB0LIWPMR03D5IXgWAeZnOR3b9EnTjiuYzxUVg0OIPmib+FLUU3ZEbnUp4aS+DA9IYtu
RJTjI/mslT1PPBPev/plvaDsbQteyCqJLo6T6VlzoyVU0UWxx6ahKVfiLIMscZS/O82qcWfm/vCV
gM4ciohABMA4vrTNa3+whmVMRNWwxBk+ZAaAzRuJkdAGPLTMpPcRPauuffQSSDu9B337hKi2RgrU
EDey4nEnDm+vNFvsNDq8FVgxRVREu91flejYqNldmlxpssFKxOYjqUcSgxsN3X/OqLvTpBRMSMz6
ldljDg968PAy4Qwl63P9OCzodqbD3gz9AWFde6jQ+r2DMWlHvFxYdz8JofKMrDXzFHHq1AL0YD4p
f3npT7Spl6xid0BFV63CGUsKSS2+XVfWbEykDsyfyBxTGmmpLtMrlEkaW11GkJ8Oed4FzhOUkGFZ
eOwrRX6hLdpm9cDozJjKOjfY2+umRIflhTFSL5ZwQp0XtN07IGmQfHor8qt3LdWQtjbOFXSNtzfz
xthyHQ3S9NAh2QzxNHc3gLdLKlJ/FglDM9uVs/0CIPfepAK0ELl6rCxF/uxbg8rIiNaHvCHLGejB
ZMHJvd4AvYIUSalPB0qCGzu4zPO7cgcnGUFUNYdcHjiyAMpescCMS4CPT8bdIpPlk4ttQnKormF8
U1xelKkE6aP2426jAUQx5xtu7lXBJRYnEJgMxJIbRHJr3VlghVScPw/2wqLp2hjDJ9R+5WeHF1ho
t3L66OVl4O0ccDqoIEIAgXj70PftjwKiKMgc6nvjzNgoweZetjEGL2w8hi2GN7SNzE+qZoOiFbIF
I5tnYQKpHtYvk0sQZIMq92YQBkD3WP8Jq4jBiB4RU15Lfi4AbPE8J/Xtcz6mYfBfzXBHZ2A9de+y
XKtVh3+FliJaQlVIRdEzJWEg/1kVAUW5zmkseAj7f/1PWchewcm5l2bUeCyFQk+dDoVod0kpQ2I1
IKOt5ii8IjtMry10iXGYrbK3obCWiRx589rVNnL2wtWlYZxl/3cD90Qzaf+JReixpkQ6c93QpJgW
pbsCUdHzMDzS4bUIHphI1BQydQpUwLOyp02n6RhiMzDO9PI8T4UhB7EpHE4Ze2cdP+dI7hqwLptP
t3FdGq0R1AYShz31i55tOxCiY12c01U1AAKe1KzlHHs+nbFvXLk7V02VGJw6lZNQVEtbpefXmmas
o0XFxzC5yzYEcw5BpFCgwv+B9HjBPmF6mUc1gSjGa90s8DwIEkdgmYtIiZuvQmXlirq68nvY4UIv
/EmubZPTFDjQXO0rxcdiNY7SXJYltBDq/Bh3QlQDRbAKNlGTa+XEU0lVgkblSIsUUrlYy6kOSO/P
NhLtnpnJUtDYKrkJpqvUgOOEDdKPIwcLe9AJMwvmaxsdJiOB+kNlh89HSmaQ5NZUYZo8+IEwssnA
h49FoXKDT8WeqvKFvlvekWQr/rImVo5dUpETYZU15eJ/Xwo8qZAW6azkcxycCna6cf1mYx7mep11
WeUHBo2AbRSQrPStzu5IpkW4ib4QdO5cUFxVtoLKbwbSW4t41uBJ0PbOSvBsSz55OawmY5HqhOFF
3Dxtdvr05xo9Y6VClBcWWtyuMK49zrFDFXykeR4ZzZA0QSzgxj020D3ozu2kL+aF1nW/HvGVa3uw
DSC54Eqd/uY5AZwQMtpklEXtbb5kH7a79hhJzLeRKNzN95Wn0SWnxwcViABrQHpHtUQXbs+FGMGg
8PwTiB2B1w27+NlD9V5tNieLc3/N+NQC5ItscpuGAbx+SK60vs0TgMbyzyb9EyY2jqMNf6TB9Xk7
UpgBSsRmSH9BoQRTX6hooffHRGbo1WbhvSxLKFcwanFButYQQya+OmR062w1S2O0ytPji1QYmfrB
HeOnn5ZDuQlH4LxEdQLBf1o6w88Eq3Pbq+0KvWWfsKL1HtH3Soq4JPDrSjTWIWqnkpmHCmjVhgPu
j5oYObfRjrmAJyNnEgbR2LUVj0Pgnyd95vRF+JrdmR6vMJ6ukVPBHBS6pLHHPakGXgdYJRiCElgM
algU2+Zxce+hpKfbpk9G8N1l9NFFktYi+2A0EEyife1LWliJt1a0sAjuFBhHgmZbif7PXQwwip18
TqLDO1SZQUyItAZt/gCjBAp7IpN2vXNeAYCuphE2bCHaS7Nh/IbHvd8oJUJ5TGOS76eVYWGFKFyK
9c+ItnKbA2zFih7hDjqY0kt8jTunn7TVnLFNtsOTi0zY/OMrD8LtBznnSoJzqAA85B1LMVEu9Ufh
JlIRsXpDsqmWwCDh0jhvdU5lLOfG3u+wWtYw0jmHpZnw5TA1ADUXh4+m8eVczx53a8aYsuwFft2l
U9lCoJakAUaugj3tx3BomxRglP8JUIH41ykZhJEtRUSeMxvfUIQeRSEspwPAU4sNkuiPpd/vgUrS
5ZifsG5xd47TmYzPCMbRzXOUT5+FnPw/8dno3I/Xna7ZaknfAjZi3hdfH3jKHXQdAv3Rb3jyEzIi
fV9phUyGB1w8iZHsRckOxBhbNx4LZ2r2Pf1/IJdtW7VFuIkEL3ssD1O5xHJ5CiRU17rvn5cvEcSM
kOmAIH2MuU2d43ulNnfEjMJAUQURjMG41CihN8DyMArp61Ewj1QEh1QJdTGnH3nKp2EwpIle++/0
ehaz34DwGj7RFgEd3TbOPjRjW7OSbB61+fdrXPc5ZSe0RFzIpVlghrVndGRgWDMKN9UGGnTIHd2v
ZLrUd82tlOZHcYh8bXK7+Q00nMK+NaEIv3clBdJV4rs7KZsC0uMJokVxi7wDIdTGhrR0W/Lbh4Se
V11jduzcQ+nLwhQoGvQ3ldbKM01ozB6adWArt3aWxSV2fqQ6DfvyUvj+0sFxiLBJVsVhegOVjemm
q0tnCEV9zLQFT08xallFsrqAUkv74C3GotP9HkFvzYoIOH4cUDlxFcm8vbnXsxtjFRAfAiFguwib
3vR7+ZyU91BiCF/IZOcR8pPFuXJHFjYuWjlZHHYK4GCubottIp5d+uJ+OOl6soKGEcXJ2I8cVZWp
xSWfx6CwjZ8Faq75WAOJC8Yg5IeVnaWimEgqK+Fi4VPLtRAZAuaHSo9xQe/cIcCM2dfwh4Gt4bIp
IGTPcEH+Tc4/brgzFzjuFx3CWVdcn5aONIDOCkFSpBWOQVfdaaRv92Q1WgIIfGg1VCNG1gNX7QTN
kDwTb4XB5zLQDXG9uZgxzbdg8xA6X08Zm0hVIPzbEPTFnvPBhoCwrvzup8rBOFmA0plz14hdjBVH
53Wgic6FLd0MbRoo44kkBug8ztfYOX/irC1+tkbx8A0MevSVGxjzVX9NS40HDquMeuRhLkW09ura
5KcbcYAjXEjyfZCYDqplQ2sE7brVte4z0HkMqJqAEn/OhUf0plF/Oxi+UBU9E7paWAjk4HAyLgbu
r2Db44sAqXyvpympUwwo/BWDTTaj8eHowmT/wwF8XJtdGlp4gRFlt7fv9f02xZcNk7y5tDmmJROw
BX2rsd8iePJn/Bxv1kcC0Exmot6uuT6fgiqrfuNnqn9JGnZjI3yVSD8Qwtqd3MdZPJtPIKdKsx1P
nujxBeRdp60tLqEr0yqpaUnCDQNhvM/Mn0punQhEQ/kNG3tqw51wOkRYIOInoVtsBrnc0GEFL/Mu
Zrm+RLsvRdlcDsoj+A1zJkaHL9Tnm01MHVRn1hvD0vh8SW0tBDZ3/qMAIut67o44Jwz5gLNLIpm9
1KJn2y4AatTYhhm0Vrf/pF8Y+pzEbvmbzCJXDq+pRguT6z8NeuK+vtIhpk0dfVb8kw+8l86Eak6F
79M8r85RDHdGxA+U454D4EPwoZyYA5ue+gkgrx/YYbBe99wTQzdyJoSbNEUquKbCWlEWdBOGHvze
m1VAVHzAn6j8/8GCC9c0M4z2EFEhYyS1jG4dd5Nyz3N3ZITPGTFyFsT3+LfkVmbnk7UqVzWs/nmD
c8pZWmf25dapfN/MlSR1LPIPmB98bkOBQV6vOfDqTJ9w5gxiIbChxjjgtdJOaXtTgOejMwh9HeA3
rfoaXKvLskZnU4Rhl9cVcVRfeiDa5i8jhY0Q+I+RDLyi7ZsK4wrzAiC1EKGJYSkRjZlrbUcz1t1K
Klokw2zuX1G/YApvPwSgCT6iNIiU5RrMwuk+CNBNnuB0hlti7C8YmPseqa7hPSXaarwtDsElqVm4
wQ8+ihjjnCxgvCjkSdZgf0txNUpNSaCh9Sqtdax0JD5zIXIkJ5mJRQy+koHtNJZ2IVykLxA72rbm
LBUHUrCTig3kUoiztcLQTkVSJQA5iE1Dn4TNC4f5VmM2pYK9lbAEjOo3g5O6mupzSQGretIdQPFz
omSreOXGIqoTM1JohxmnSSemBjLGu9I6eOxi6mzdvi68zQccncbRrI8EPZBa5iz6DZ0HIictzk/p
xXdVq4nOqMf9j3k/k8rjpjAbUMgm+U8Rt1EnxZoxKYGhB17xNo03B4DE2T6JfSUEYqwZsd3rpQJn
bJ0Rkf80iFhtEGaEbHM1DHRaUJWOB3iEppqYNi3xbYKi91JTsjbQhAV75M2UcU6FZAENFjQ6B/Jm
t/Fnhr4J0IJv5EHz/zOgFXEgHTZEAKiK7jqokMSAwJMJNCylhAuX9G0ktivZwR3H2R5yJq1ErHe2
NHWoOh1OosJ1nAIvvP4Ayln6AYTBsfvLAuA0xgWhbm6CjpQdsByQJDOVtnHmDxKzryBA2dR20aWw
mbNIhKxfh08cXE5aHO18Hx0V3lXreLNy5gVV04XYyvkDmTU3YyL9jUTClv1zIr7Le2qRfVD5fFg+
yL01Ojb2aIWiauxO654scULb2Zv7djwkfWsnAiuCg8j+FXu+J7CXi9ThALQtEovBBhurct/Yf6Tm
DF/o0C3lHyCYzUQiW8qIgL5A6irXmKHzD/s7iNG+yFyg9ix0HRW821RT6A1WgFMcahm4X6tzYkNQ
/UvwfxgaCHaUF/ow5zvwB3/Guv5mZ9bBgkZ1Yo8tmR4wZUNzr1heJu+ifvBRUemTnPlZzaTBnoQ7
eTiPf7GpkfV6W+Dsmino/WUaNp9hKjgcT+Uv3VCQOFvEzAYjtbdEoe4CMgPkohgLB+1oVj/vfVAN
lRLbaGxK+B4krC11XsGr1Fi3yabitFleFSk7uq8SeAkmT2OTWPj7DY3sr4lo8DK0npWKH8eR6S/z
HFPZ7Z2x8IqvHoG5iSr68mM0lu/o4wJFj3h3Xy2elWlSQnvUgmIr49z0TUROJ48NyTOHq+tAlwMv
TzjA8mg6TukQKq+6NUrP74lJoW/0agEcd2MXOebQRkJ5nFYYj1BrfSxTWJtMwtluXI6bFLfiXay9
Kv/zBk3cn6xtQEOKu6T/TtioY4ngrUNlYW/sqZmzCd8xh1AirMcr9JXehPF+RX5Fhn47I5blegLR
7xy6ZTvU7kIKjtnoMlB+v1s2lNeDBck9GSTjudrT3kJcgzhoTp6fmwKe+OgIIs4w2IhBtbiFTgAT
qZxDRlwnMC7b+rwfhr2FEjbACDEYdlUlr4mebvPFAaZMpJPHgdUzzxny7Pq/GWHkk3kK4+EKIU7i
F6B0D/oKHtOw/35a/Bh68RBBvnJ3cRv0mTq9lHVNNrczMazbMrVUqKBwtowmLEyBj6ntK1FLrU0I
nwvCWhw42NyrkFqOr9sG2s6fdY0becRvvJZ/DQASb6VieL9FLG2DgGcOLryYjWneSSlhZes+/C60
GNBGvlbQNGdCKl7I/i4A5jnTNm3Y7OVVD/VmLuLnSArQ5uyCzvo3piW+xgZlJ06cxUuUdiCf3y3r
swldsh3mFvtnj3ZdYhg7zuUtj/f2l/dQ5sykwJSoU2d83JJy1RVQUYATVyCOqvkbmCNBh0CRxHCb
d7HTVKC7Co/0/ZAcNkB7Vv1Zk8hGP2c3T/ri/F/WnWFnylbVB9sxa/DXdzFGgU89dn3unOUCOs9V
J6XNaIpj/xvJfki7pcoOLnkif6aFRTpmeCjlq3Z0PYC4NVkBqACUMFN2NrAM+oZAfbku0sQ3VQ38
PZWazn0y8o/yc+bDWjtJUONsPOspREtSECRFGbTPGQRQumygpSyBP0eQaZMoq2W+kP7hM7gvn7vS
9QnOLroK0h/JVrhLLbNjndoa2jLpjB4oX7GulEkta0YY+XQPzD6jTeP2Qeokk++iUHB7qvQesDQ2
7SFcWu+RbV+uBMgC/Y4niMGw2rnyt2xgLeV1Jrn3qrUnzkNUgcPpEjLy5y3p6O+7GvOelLIJUBjJ
VNI6ZfIIjsqmLwb2P3gxQsTIFtvOJNdPWry80DixToZx/ifod4Q9LNtZpJUf0Az4u1xVqYki9IMt
0DsvBewZFheVNGas0TbrSK56c/e7UiIVyNdpkzwqFfBFRIEYVDXDsWPPGmNsB/oNyvQSzRltOjR3
mf/ub+M9uj4d4TpI+HhT9MUImQZaxt+FvNr8gHg5ZzeUgtFBLmbQ3/G45rrSa9QVRbJwTeRbAeiq
8OH9gMPfZWUN031JHS2nKVHYLg80eli6DXnJB9TRU9advybPfrOVLxj4eWyQEuHb1BxEjC6Rm0YH
u2LEcWc8JqJOVcPrEU5DKEdijuktaAnP+Nh7UEH36uMBSz4rV6FX9zZ0B8uy4u6blvLppXbv3v+h
CHTPMIfKBhKVz8P5GUFv8Mfmpqv4BartgM6yOIsDtcSa+sTU7kfHcDRIR2pZgoGOxY4peQFrWr/a
Om9ED9FCTfhwEFem76upyQrzvXRI+sKPsOwHMUtJZW08KQo2ka5buIpfzXasAU6F/MFxdq3AAsLc
ffPjCi27E6wETN0jGC3nUUz4B1NCS8FdxSptckQJeny9eaKw7Ewa1v6dn+LcUanKfr2pekrmCADr
xJMLdbpfYGRLsmwF9G/gm7oMfaYYPNoxxTfgMzlOy2u71rAk77yPChh0LJXFdJq0/lseQvFV+N7O
fK8CoYHZ9vcSItBpgtiqnITU6qHj6ZIxBTC9FZkqSOyKn4NJZBfbYUf3Hr3zTRVIjat1zEEDhpxW
8LP1tvqqSOc9SQnNIJqzoSe20EZ+yOTirYjCYftKRITPUuNJE7KskwNU0Liwvb5X9U1MSv8Dp36k
qGfSZJJ0K+FtBkonvhWaXv4xZVcFWkR30gve6/cUoglHrllP8726q0aKBAJh2cFL+qmgXHmmn7hC
f01O29RpgkWuTUQEifxRrfmfKnbu8qWbNitAxiu0zYrwOB5SlJ/u1idbuYTFy3FC2iPozTYsSlbX
E1D9iiY/Ee/yMIWeeQlfEY5Ry37CrV8wF+z07HJy4YRyw7eXtoXc0ozo5OkVb2/2QmfwBT8uk6AB
t4JLySNz4fmjAfIOxB5/pwPZj7//Sf58pj5AWTi2/wm0U1f7c+p/nt2b4n2rRGFpgJ1blVG0AHBb
4fo+KM2xdDnKsPCs+t3Abod+GYkBs3axk1c5wDnRXJDeC6M2rCa1WHUoITg3/TdHnJwbb18aIxMe
oF6xXBuTBjUPKvaacuwUGa5Ruj3q+/X/Mm7j14WiQXnIkJgOzhETg3L9hUuLN9nFJZjnKSC57Lty
13w8t+9PgF+huy8BQmDbh1b68LdTrwijYpRPw4S84eTAw8o4hF5k373rIWZJ63Fmd3IhxJ4aEoio
5Vz52UpOPgV8sknWWC+UpSwzzGPXLWFkFNU6cEm/XmSRKLfWArVpVdChBN7u2ij+42is8wGiwQBO
+y3TVq9Y0eZ5bkvgbCxL56Z5Iz1GJbAxLjFQnHrS5p/7ySBV91sK4Ia0q4xoW2BpIiNRB568NXfo
xAP0i9/1hY0J1Oo8Vwo0HZKaOnddvAd0U+6ep//Pt2T/25iw8nymXxGoJBD1m0164/a5Ggp/CsYT
NutLLt2GGPTk8oSdC/fw8zGjuLmnD5BqX69Xw1yEZ/0ENvF+QMeix1kFg6ZbgU36hzFauXs13pQI
hvXFMrtcJJJ0DZhu4PJVS+RNrRDL7wdz+nwlkwBMb8YpdcxfND+yLw76lU82U1qn2m7VYwaeS4C+
vB0mTM+XJBfGlbiZyZIlR1YA0/QJilaSYts5DT2a1R3QL3PKjWwfiZXDrWePIPZUmIsH2UwojrtI
78aDnpAXXBCTpVQdtl0gP0TCN6qga+ArlDRUi0NEcJ0TnFWNKkDjzHlvAMzO7wkJia0B5E6b1iu8
xswFHYELD18razF/GuO+znYn91lilVztXeAjs4rjeMmOtDUEb1jon6VuHsiEBCeW666NvIXbsI0H
lN2BTqbJ7Ba+fMdGJqpm08fxFPSg+e24XIaZ520Da/aNGL7qGfNr7p3GeiEjLZ7m6uI+bsgJooBJ
U2NX8eI9u6w39+8s+XKkOf2gvCG+7l96YtZRRlYWzsxW3t283z+E96jn6cj7M2cuyX1u8WeFm57J
4UxW3pJwgLkgPvn+plj8yUQOryJd4CIBD5pdOXauqvees5F+tuOS5PAOcWWeUmuY+O1GI2v0WwMX
fb/BR4VtmNqveHh1euGNE4FnK2rmv11Y4BX5y+Ny/mzybovdD/YxpqWST6wKWxNT3OE9kUtwAMf5
idanhuRdOj2UziCt2/OWcCknK9HdmOGUntVWi/01uu0oaka1DZ9RvHwvtzh/cIAcaX00/HsNzTJI
DB4/m9STp20JtkXpiARXSUGYsT6To9HjFcqoMWnrfiDi0I2kzlr501JQygJAtF4PKWlpTotWz+iX
rhDFxAfbiUfnw9J1+jSSdvsW5KIHdrlHUp1+4e6a+uCB/FfskRKuuVWFqHoxdU0X05WV7EIN/hQf
0bu2JLKYHwL6q7ViP9xW7cWjepRAIfW6x1b4d5dfC8foJdeYj5uAWcMnhCJwdtfPbEpCaXzi0dzQ
prQ9EVH/g2WV3+Ntnu3VkOcXzba2Q/EmlLj4Yik2ZvuEsWxmVHZ0he9OzEquysb8vqTUuI3+7OQ/
y4m6PBENomnRvO7dwmS0NJmeMZamZYLcXStxmCmAOBxVQDMyG9SLyrxxXNkAX3PLOBPGLC0P3aAW
c9e+UQcOVdUGeG5BXroCf/mzRZ7ZbV6Rd2/GDQvqRBJRuZvsRI38FGb81L+Mzt+3jMGZTyDWDRom
vsM0TX1wDS5aBdVD6r+GUAZ5/Bgd3OO2JTHGRRASqiS3NyrtnpqMCzdVJYHNmcFqWQxDrGameW44
St/h6tOOCR2VIq/TQCywhVRHU2yiWoKLlgh8WZA8FXzEjyqqkFLx/E5xoJ60hWiW8SvQgNsubW1u
HukMzdPWkG4wIt3g1pfglym8F8LbDSLccbn//LuSVYYGBRrqiiwImotWX2VaXp37XNsNir1jad28
eOaO4b0pXVgEHB86XIdm8ZjHZ4299FqT9HBF6NHhNKXboHarfRmGut8eLzfkme0RA/kyQudADnbF
kUZ9h0XVAnIWV2nMCc9qlcQxM3VX7/9BEnPVV7Cf/7/9/BE7mumRBZrm8XN0h5rrsWpgNgrOqpiL
xO7oU2mCqyn3bWVR/fX5uNZQPkTUWkG/VqBlXQSgOiBdEFa+Q5yI+JwnAhtlKUDSlEbtrInSHhic
6Y5jC8bCz8WK2zsW9vISFIXQ6D8FgfsdrZ5PoRoHK+rTaT0XpXJzHMki4PvAeWp0X8fPoJA68Q9N
iofxmvhOJ0zD2G3TAJtq409zOi/72o8neuI96Cl1DuqrZGRg6zVpGKnTV1BOq/r3gPgsB9xdtk0u
kkr8EdaVqTtarZHgHKZF10MKeL+t9v6nBMNx73+PR43yAN9Zx7kfZB89lesmeJuNv+KK9sI4lh5w
r0bYc79l8l6anCHdBwLIqToonaC0i2nil3w54DwgHXx64cqtdn/BJgJrhuMLARrxhVObTo0//xhI
KRB4/f3MUiieccRpVcu6cvDbWoZk5sfRGvszlfyiMn4dPmXUNhs9ZHAZIrRCs3Pc8WYb4wl5aA7T
g23UyKIAzH7v2QddIpD29d813gjOlh3cWU8clF6RaJP+6ew1yK8nkqvBRiahhL490tVIWCSjimdV
U9EfMpUgHyEfNU2jbp7Lbo01oVyAcv1zUjncfBwnbBWZMg5VM/rMkbqMl5tdlIWy7DdrhxBIyWNG
JPpe18THM8cJPIJs68S9hd8iSZYLaZtb9GhkS0yZbu2i3RRwHpTY4rclwT1N9zvND0BYOhwVqhGg
TeGWtPmEWU8I8cmIYyYJktSf0vQWH+a6hyBL1MrH1gVSVxnjn/G0pypY+AJFAMpF796qeJzg0+hq
w0oHJGEHIPFyuoileDneikdb2Ev1Frma/Q/bORL/TrAxN2XSGNUnL5LML1A1KvFYbQh1XVx9pD87
mY4nUp7Qe888TWNZVYhhSxFhDyS2VvoZRm7j/klRb4f6iet4yHbi2/cogeDMfXicOhOJbi9CBv5Q
lV4eDAo7g0oIiKln0d8D7PX/pWnviVi2wbTm6dOhPfMAeFGL291NtGrT2MEbLYBvgklEXDSBa6ZL
lwoRaEmJqDtKlGBdhla+/+ru5HWWiSj4OE4BNxvmvgE6zdN2RHEwbr7Ed4XIfwbmEw3lomGxLS0s
IC39JoyzRPeB0an0SOgu86lAFfMz6q4o27WaVDLrCdptdaMJLCxpJHtLYNzbC3qY3bVaozfHI/3J
LTrBzyeQL3HBy6SSzVF4qFJrfZPFDkzFhyLlq9T8xAPKRykSey+avawaKsq3XdpEgrzslJ87te9i
qm2XFOErPSFBKmNpjAe3rURHrMKkbHpKuQVtMlwexeATRQzmZRBOaIBel/M7qrubpmqKhWuviz6K
5tF6R0rrDNPadLdfbID2ZJGHVPkCOGwwmMbDeb4AwvEzz+sbp5Au+1jUpC/+u/tVQm54Bmv/AbD7
nGL7q3rrxMi0Lt19Hw9Oj3R3Ov1ivhk4mHaFfhAzB6f+uSkkXWltRbFbeDHz9wv++Tr4nmYHcLcd
iYCbf4A+mHnp7twyauay5uiAMCnWLLqxEI8CrYOVkO4CcRI01poEdmOcK77GH0blnU57cWnwwpI8
YHGnmLy8dkJCttZE0gnRg/dN7THEHurybNh6RjubQF5ofq6J3o6DZMYrdYJaKtcfmQMa65fs91Io
jFT+Jw7KQMbBSPvjjCipMk3kVW+83aPI3HGsz0G8Bq+ZgJ3ToJurMdNb+QdbC2Yz9AVfjfK53//P
hqUFx50zsP5ue+TA4SCchk91yS1u3UTfQV+DwALBuloedaXLzN3Nq5Xjo8QwLGVY7iK3m04epVVF
0m4OPJUngGoTXMN0z9+wKqj5Pqd63K4CsrUOGQUr4MAjx8sLl9LuR20K/0tcdfPzA3yqjD++bMA+
CLcjK6cBnjMZTv9upCr+MkueQuojqRtnuYFCheCcsNeMeHwRh8lzOuEg67kZk6/o4jZdCj+xaIgY
y6U3ELHbQhGlLtgNg34FJs3uEtILdHl7EO//Q93uJPGgEGzQvyk8ckSxuHO0rdd8yOaGiw36wYYr
NEnY/sHTNQjMm3aE4TTOWkduROQ1IfwZDPaxXogL8MWyqptZUq0zJ+2SSDf94XgrlhdPTXm4E315
A9GYWIXXzIikcWbXlvwu9p43GSByW1UQQ9rZvO9VcR3qFcww6LIxOdYhcAtA3CqhltlaVzVNTP8E
bun2F3zFnwN0NfrB8qgIpPCm7ahJLZCSO/oMrIPJze7E0ZPmLtPixAd6eiIvxxHsnIUyEmtdHPKe
g2rbD5R/Bapu/b+5k+KqI5pvXZuizbeGm9knTaaEpTxCQIvsP9EWTnN/aXtsEIpRwCN2teEKBKkl
WcmTM6ff9oljeMs3HLVU7ACeKuLB8zzwf6jiEWkuyzKrv/Gw46xfLsqcHnsxb7qVus/1Lo2sdVbA
KJIQa5lWgiojFNwMit/wSd4VD1UZ5Tl2xrE4Bk7bDtSPNF7cKfGpNDUKgcF7WPxpBvNHQeKj7My8
ggJzvSTgy2/j4wOlXUhuE6DHdgt9q3Hl6/VI5JT7ZkEjgsoUyH8tSDBFXvnUnSavyWDhq1XrZ+lV
Rc9CTwkJNDo5rKOlB2hmG4vL3H65ClyWhMwEJsr52eQVeb18EcjsS44cGqDgd5eanBTm1cgOAhqE
3mmLJ3it5MhI80pjfIEYZeKnSzcFwb+t59FXayA6eydlYiAlkR88Ms7Gyudsy0GkhfiF3o+NDjUW
VhfLQokpFhil2sqGYeqDk04aND9qi05ki6GRYAg0Tvhrv4SkoI33h/cqxNJazl3uRaC/3FgPbWVC
TQ+1Wfz2Zm0n+BEs6JbCbFp7LGGr9q4HJwn5PfjagXACFWpJnmZ5ZNxINMFSch/PuWht3LEh7Whz
AUpXBz3m4+Exc5szMjP9grIRNWMTeErUI2VLKUQ6OCOSR6XtIFNQ/dunJRjztDmo0b6y903rQiUR
wCSR5sHh/aznWhr8bF+37SFJi1Z2+fU6Gwq//HN8Yu20PNcAY6oc0YGo6XNozCoSAPEdm+qgqvgZ
sGfTiblTEKL+AxC0Ph1UJcc05A4XCMqu98g26vkz073fyj5wyhqBarqO25TbX0rHa1PNzNj/7E/v
IZKblDWRs4rYJpUW6QsIL4mjxwRWTgt7/hwlXjQRvYLb3mULUvv9ED/3HKjOyjcTQW8gwQlQIUEr
zHf0c0uYimICtk++56Kx9u9eUAv6RBYCQU0kSujTf364Tg1WrPo3ck21Yt3n5AyJj4/3JIgNaqyR
JOqwFRly+0DrvyFe0lfF/9UHLb+EZ0Ek7PwTDzxp4dKUWf1Ooo1Q2C8su1xtLavXZFZD/bVEW98H
KyrRtitixSsnXyP6RKwIt1V7qoC6GHpbEi5w5JjegVtjcVnDolTd0Wd3F4dNPcBZgEUhynQhGqJK
tuoXWer/YY/ILGdBehtv9Q/mWTpcvZHqqApU7QXomT30kGD3p30YMe8QE2WDbgTjqTKp8Q62ugEJ
gPiu4xGWRxEUz9sjhzG/m1HITXpDPKVq0pnqkMbbkYBnfJ1dT0wtZCxi+cqIf3p1K6rfrChsdaCi
cqvzo5ER28CfcRUZhZvc4N8FVQmrp7HaCtQX/A0o1/bMsKOT83MKJmtrB6VuSnOydlrXq1wvV0Z1
FXZRyOAtGk+KcFPnmKWPZP6Cy9Zmj+oKM0Rlme50oTMzAE6FVfMw5ai/31c0lhlavr53iE/9N5gB
u6GEKCOW60ee19BxMSyJzv1UdRxcHCUxXghgNA4QB6Ci21Z9hIfrRNeq/Cp+0tNSysIgXe1l4fa3
x1ayleQI5wx03tnRha4Reqf/SFOfT0YUkyoZBC9fqTGweFnmwkSlZzLUVdc+WvVSAo0SQ681Rohs
tn+axdsDvXPK3e+jLhINBKr2qZ1rwr2clUNnuJv2ze31Rf7I9FZ03JxjTd6OVdeoHY6HXf/j6/4m
HiqTUkIzJ2mjSSJaaN4yvysX5trtq7py7dpwfyXjCtxobK1WTICzHMVD+CvKPTPnHXDgnFFJZ8f8
3BI0NJFIKfHEmP0l0JPOJq5PUt/LtD3u/VFEqeGjg7bGIDShE8+MESjZm2K0P+zLzzw8kMgfwP2s
nAbLKYf2qfZr7NBa89u/Kxc5n8CYXQ0fPLUyOJopTb5ujOXruow2QUOsI1El4g8kJM2A6zKbk5aq
z36okR6r0X5RwwqkT4g8+ZywaaybSmUDhVaMkMTsk0LUGHincN3w/dchmKV30GYuB8H05fgJj0AW
kU1wRlMXRfeVRbD656rmjMBpUB6uGnE1exjcfbV9hIzCYWgufa9q10sH0H11+D+tsr6BTgVcazO5
XG7rv2Jp/sx/OHLBvObvFErT2m3n6NISx6iVNqcth0wLY4O8Fu3eUz2NEfZ1c3RKzBUVTHJ3HF+N
MbVjTlXTwwpGbcCSSJfhKCofdHZvaqLIczb/5idiyurWoDclVRQ61B2cHCXe6GO7eH0M4moZT6XA
XGJO41W8F4IxQu6gGL91L2iUAzoO2rUJ4xLO1B3kpSzxtDLZIZIkl+bgHyFPiLdbodhI/eu6JU99
wSKEyzqHg2osa/8ECVr1XZXwiEvIaUI3YLMn3NjWhiXjoBseHI7mqbqvTMTWRwjlu7wrkXJs1Xds
OuewLtuW5fiiCAHtNKd3WP2yNfNq3xE8DE531+xTX00/3Ri93foAyROpIuQO77r2nDzoXf+wd6Vn
aAzVaeTo8kMNbO/S7Il3LTa/EBydya57Rcajk7r9oyYoZTtGnSv8INvD6yk4sdknUIwhvciCPDSK
4hUKitRt6VusTZHPNfa4MqRNajDH6oNpbpQokWPjA6kAtl+gijFrlOc5oiiLF7gtNCk2AGCfu0da
BW6ByYyWQa13JuZlWQy+zhff6qcSlDcWtHxeIM20jTEEfoFN4Ku7oMCq0IDR7yfC4aUXzAPOANBL
EVhtejfOY8caU38w1m9Vh9MQV7f+KIicHDMmND7zzOMvABL9NoefQi61bExuzdYTom7zCYH5XvBm
dFcK2DUQKjbzw4xUVpiCQiZcd9xpPdomr5xY5Z7nBJOHXVgr21GuchUb1pomi5rqRdywFe10Ayl4
GEMK6vAmgrIUTX0qzRmoyz/WjgO5QNSZY8SQUVUMpAOOcLDJ+iEDtL8yf8eNYQu7bM/KUY/Bn7gF
iSNxTHO4TOAGv41WUtrtl+pLNOv+CUr2Q6vbEN1Y9dO7XBk5K5wvBK5G4PYXHQUp3SviEA5tXpy5
3Sa+vnmLS5Q7O8Vce+RO/GegDtGjcnxhkV03NuO0dv6y/HmYWPB+uKGT7YU95C0oHDAQmgAta66R
SEm0bLaUeBNa5HBQKRlh9MrnV/dONeviLv43+3WhtVCh0LQShpKQm6b7CJ+IlOUNh/LyDIXBVZmV
zsMNz2iFcMssuyBD1c5HmtTtpSDBTCaPVU9IIe7w9HrRWYmiiiucTeq04vY4opTpVfcxW9yPB/ss
0qEW9oyuYexwT+yjotmvx1Y+4kmlMIvVBzSphlFd0rN0N02DonWCF3xTpc/E0jsN2V1vd+7G3Yha
s8ukNfbHgF8SgBBiiNLsa/gHW0ZgXkJviJU2s8+kb2kdQoQs36qKVWsD6974K6ykFcDIV9SRakIg
1/I2hgdJOetRR/C4gex+U5ETawLO0JzLiCowBdbkZLP34W+ACxQE67JqJi1km03wMFiF5s04YzCQ
u9y5G+cF5K68M3ET65joeoMAkNUCjH1jRbHQBcEFoYA+5VR6L5Zsvyp7dstZTA9QUoedoo1mDlIH
dEb5nYXnx4HIkC2Ye+87w1eXnzfuDM6n2jum9eLK9WIb+rCfY3UB4pukv+0TngVydKyRehGJv8C0
DpLmhcBhCSkRgh5Nwzu4z8jQSeSTi5r8jVd1YhTnU5rnvpWEYGONrcY2xdXSW03WGQqV65UaW29x
A3k3BniGdiFJ7A25KYYHro6fzGraKrJA1gr8Y/dRSa5yy7S5f1KJLrbIlIBulr+FU8DGXNsVH0Z0
8kFhkVFm/0SkqBGXS04Mzs0QUvqrDla7brTp/QVjM0p/9WkjrMvRboiPth+oKT6whXPBm2/jzptT
2bvMImExF9eYjcErYavm2zOH9oJKqyFThx/AWXdV8UccvZgua83f1I6qpQaHxaMQT7T0e/cVSJ7p
rVqC9YaHVpeM6fdQ2xC+r+tSaPr2Ovm1cZ/Ykr8BOUGcZCLXd/GqFCtFB3TP8ZqnPMg8FHhE8+PA
/HPrReJ/pjWu6BX5v8AUtjSupcT9fO/eYRAPlUnHg9nZ8Gq/v8nxsU/iArf9TV3bczL4DGDbqDwb
ZxKYLcy8JkzLTKeyWqJc4n6L2wAQPv0bPBi6DQo8OypUxsh66e+eINXK2tSRGeV1xg8qrCpInJfb
0hfLEqFwQ8jf59NM852eb2aggLMBExRf4LeYM24l0erCoEw/I4+uBpajxvRP82+DK5ghPyPQnsIh
Y8xssKYXgJB6X26j5qLTglAvD34QvJHZWuHNZXszvcphDJmWzItvbR3j79qrjw37PQzxhcgRCFgE
VzW/cXMzpPOJ9NXf8UZlRN6pKUIxWW5XLL4kuXVWxSluXdXY+AQO5RdRqtq5UgWtBLX6jgzwaIqB
wZNE4fgeBGeaIVCV1WwkRfiZa0ULR3no6Th96iLwoGxqkMMELmPLhGlOzHxcMcy2VUq4+ymlxxVv
6B/3NTYvW3q9RHuRxj42aZpMv+X8zoBDAlly73vgSxHCkDAZ9cUmo3Hcr9205BuEmV4iL6d20Oe0
FWHcZob8xAeiXwuc80OoYSILLm+oRTV+NxqYM+GghutMJd0d8v8Fo4QC5aEl7fu8t5LeHuUpDC9/
ZsjROtDXJIgFp6lXKPabVeJ7uKIlHsoPreeoSqufLvmWugQw/rzoGP3af+z4kd7kWumKzMPGNz94
ytQmNMMLGIVgnie5ouBHqguWqwUEj9VhixErlkWG4guIJttx/EJ75BsWU8quxrVXf/SKR2gMddum
0DdttdUvkQZycxv0Z3EtAwJW3oXXH0gvkaVnfR6odAflQTAsZsE6KtHA5Qo4mgfZZJLfed042TOG
Fv/LDTff0CGFHTUZEQosBMTLObi62stKbcayKVxWlY5dvV/sg6hsElxdfTjOvfbGoNLgjasnK1i9
mjgPXu/OBc/1F6nw0jPDTrBBeXlUsrVfIoj0f+9vfNb5gdOw/pJDyVrlyLDBmRCDIixZnHldMFgC
eiyFk49ZRx37Zkfdh9hkLeM+VErGp5y+p+QHmdcMZUOK1XsXa1p0jTToZUw92+yX2onrczwhti6O
43vST13BNmPw23c8GyTbtIKUOGtGACWmP+esi1HCjPDgLAQ61PjMPHL3qPe27GEeSjNqKAXrpvOs
LYAEEWsm3Rz9ffkby/OEpokPn5m+YmvN8IKzCJ7Mbl8kbX0AtLrSs+eTbp/nm7OV59T9UDFG/3xq
jy6ffCe55f7uad1TABNgz8mYey5LSPe1ynlTC2xFBFBIWkIra5ucC0MVb4eq1dearxFT2iXbhe+d
1GUPrxP7hvLu5UiqDZAXXrQpxJb+ZEXaCcWuyHO+nsxaP4ags9tCefND8PdN83qCfSNNf88LUbeg
RznBiAmi2pk8bySkTEboT1zo5MmJ3VDYnxPGuguDqkWYuKUieI6zTf5I0QJv2PLrcv8/R4dGT1nD
UCo6BIinJ0b2jeVtLtVuikUqDQBqUpHyEKhS7KH8UGyD1QPVy7mD0x3V5PmIYBYkXxHUZH7mrIbY
7Hx5NbTF+rZNX8Raxj3RVllLiUVG4kOITRsYSOOw/2McPcyP8GWCSX0j93iv0p5qKkxYyBXmpA3E
24GbvnwnYzUewnRczIXu1ZGbjLwl6zZS6f4LPMYN+NY4sdYTqRCyR8Q672EIrA+NNEKAmRA47R+s
hIXvPm3xeaHkIz6Y/Hp+qJmeZD9xuCSv5JW6NYjVsIOftA3V6gIuYFMfVdWrR8IlowQp7vrrqNJI
bzaLwJWZssa17u5+hwOc9t4zcyNy5MuogSFrLhemRvWOw8YZFlfr64/2KIqsPC736P+GYSYMwGlQ
5eq8xxGqh2gnpQuWAdjpqNHO0g9EwXNRejJQ4hjbUEiZLsqy7+EZRYsJ6jMXz+ULRKLgkq/+6mCQ
5jREsJ4eMJfwsWy98iFatN6DeuG0FMrFPqImG/ybR2Tvd8ptfBTuUn5ZBbeTZtHtYtNzOoi7QBEM
Lz2RrfUxQtafOkrcm0W9WADs2W4ojws1TRyjY709UlJhRTKxuh8/IHmdgfHyww47MMahmcI/auow
GRrkP4vmoj3KL2NsBqsrf7kU8wXJNhYQzCITxt8DFY3A0JdOHdJSAzlUk18UDMfPMgrtQWMg+G/p
bVJo0SkncApxrCKWPMtIPuLYPaIE7RJ3C7MQdaHKByXGdpXNHWnnQysHHecz221hhNDQIVXJlTRx
vnBW9MxISawRlIaDRg9xPcwPcz9OT2bmnBugNLeixxXHTyBHTfbJbtQ1NDf47wg4/UarT/VgaMbH
+vh3PKBQmJosfukzkGCp25st4ls3+eSfXAES/jZ5o1XHjzDi+owKtW9Cg3erF+UEdT7nRnA1OBTj
GI/UYOToCXDEJw6z2JAX7hH8OI7+6/NVs14szdC+sjuLQ7BjUMKtcaUBBh70HBQcRtbfQcyNuwtC
b6B42YbOygHHhbvs98RFRX3AUBa4jl4vIfhvvEmDp/6gap1DszP0krHYiEIPmLZOUSMYlpkG8SfH
LBVjVb8BJzjm9TLfsYAWWrdM66sF6QbquL91FY6twCcFlkNem+7gaEeHyPGAvfBsgESM74WVEazc
KhGosWgJecWAaBsk6tVjwIs4NQmpMU1a78stjhV192MH/+o6uACSykvmRiuja9HH4F+rsbofjXwS
bmHlkaJoR4MK+ogfOkEZ0z10xCq8KfHbkVPCM2Fw8iGLQkF4gvMUuyz63JZBhMYAZELFBfoBBwnT
kKOgFcfB7rtG0bLvhUC+BWpMYfrxFfO0tjryf8hXbOMMj7muOYvWH38K+Z2zrhUB5SwjFSSSr+pI
Zgg6RYzr2kGIYWhM7MovFYwLf4I41CO2TYQoVaNAHyjKWQKmojdAGezYoOBUMAIUXBn2TRZBxGNa
NrqrBNxsm55x5+xtsAEVw5uUBIH4GvBBpLef08MDVW5TvSpdWtgSLUxHtsM8aDYyMcoGBVhmIb7n
8s8KmITvb89rcEBObdn5BClVKvJt/StdZ3wdn0UWG/1fJTMn/xp3zfae0p9l6afi4KKjsomXoqWy
/x9xfA4lFwW+0gV3yo7jI6dFcGt7n1vJjq6qrywIFCK7BvaFGNfEQiPXwZN7mDesVGbXpflQ1LM8
3Qq5UI724EQccqsiNuovQTd6EAQcK7+wxhZsgejugam3M1BRCCY0uuBdA0jJjjJRkvhN3SVtKyHX
YESgboEybiCefd9O9ZkZqf6bcb4enC6SH+oFnNhpWgihi+o4fT2nfActc10ARBDZjaNa6E/F34/+
b9oCrjxmtpoDvfuZPO7lv7EoEB03GRjtQoUloM405aInBy/9W81MmUBKOyP0bMrlPmw/a2nMZQs5
p1WAG2pTkZSZpIolTBDLvUtBKYNuDJaQ9HPTFF+b5fcUOPPcoG4L9fbB69hXNcaKs8Sr3nqnLm77
YqXd+vOqOSG4YWviwzxNNdkwk52vSzFptL9G6RicAREjlED0mKV0iJU93RKkCQR+g8FV8zvTeO0+
K2bDdELIcyCWCzwWkKVBuEETE5NJz40zKg3MZsdHjB/sM3YMB7QD76/9vQwTphX0NUuUZO4tCb2G
mP0hU9T/vcFG6TbUAcznvkmMj0Q1vK1FlvDYKpUooI/qaszbLgJ4mRZWu6EqF82PFsBclsB3WX9s
x7fUa02VvO2UfcTzFZVgRQTwO6+bUf/pIQNw6DUgeuK1hAcP7ZwVSpGUc+mXenjIWX9g3QciPlr8
nQS5Ewdkh7Ls8Uc7u/mkWIgtYcYa/b09HKaureQZOuvv9PjnlQ2nWwabmgAtUwB/wmi+3++u0GjZ
5B4pr0r1OPikUpY5IKfrgdqePSwIBrS0DRBR3DDLpg7x54yMgYeN8wN9GcroiHD+fjeyLfywxUt0
wg2XahGVjH9b3USRYEv4c7v9gkL+xzNOB24Ae8HcPst5ATfQV7zZv/yrHfuO7U8jqOmvzshVRD2d
B3AMIq+n73+w5nSrycNUGnqZODLGYxUr9k6/nScBWBaOAB0M9xEntMjCbqoxtXvMb8WN3UBlL1wA
cZY9u1qPg2Gu6sdy7vMF2BFLEwmQrYN65CkSEd5E8IewRbm9mCghChI9woMIPCsmEmizH6csh0Va
1kL9b7Tcp69RXpR2QQlDJxZe3bu/l5OJlLUJLILzymZgXvR+3D6PfwF75RevF/a6fl0M3dwWVTOr
+Ph9enZ+WFe0rIaXGWySdMeDJJ5Zt6zfbplKhpRCzQ6V1OGMV9LWiNJVSIa2DCrNxJoLvd7I/qaA
f2ss0bANumTXwf7HmPcQ1Xbr9RMf8vgIiv9BL8ZKj4Dg/epQZ3jzWweAM44g4MHJdnUrCPYuQ0A4
8VsyxkCSXkdon8UqQbDl90SJS2TEktruhK8hJ6CB0SB8s0S7imsO92qCPA/nNA1fWbsY4MFRxisi
lQQuuROKbiqS/N4t6APPq3ClNnlmEBGaRoHREDX7MMFdNfuUq8RYyXTnRgfd7vb4+lG8VsIKVSuS
gVdpi86Bj3oeD3zQkoIx10ASXeF49jEiPexBiQ7TF61HWTzidP+QWIGajyWaXJHCaAfyVrZrgAWW
i//o+rzbltstrpGdH8J9zishdCgu3BYze+HvHla3xfLs+2xF2LY1fvorsYgW5yQbVf5cQZdNq4h2
7ZrHPdBJ8f24ydsYtMgBhttJogqyA2O+7qrVluQL/tbiZccTF3qX69J1vPDk4JPMP6Y/68wSpGk3
kBHGXDpymC9mF/v2GOX2S8doSBT9MrEHrUhlRmEhXfA9wA/9972VAQrh8Yi5I2dHTJ245ZN/+pW6
I+GPufqubvoT1Nd1c/XbXIkoyoIIjYa/VxedNAbugrx7ctlnpxleriDvyz/v2OrLSP7Tq1lZRQf2
VkKn2ve2/SF7yf53thbbeL6kqbaVTsm1PGfpaoRaXQ4/b7mb+GDXijnaOYxqefPckCGm9b44zx+y
SaCU8x2nOSVHCHB4MUAhj+PH+jQudlv7n5t5NoyK+gojdbVoT24L8ClR8C/NUFP6qZfnXEwK3ple
Ub/lIzCP/ZGc8WDWwvCGUd/mqf+YU2LQaWONdKqSicgZ9hMgjWBxhfk5kSi5CPLlhmzcz2vpCkiy
Ehe0m1kRVdowrKakmbg83hK53NokRBLUbALImqwOzlyQXLuoJsXKwe+JOx5ZMVrm1DjmkSAd5xp7
NjNZxboz1mvfugiwjyzakI0ASaiZxLaOGuxgIbMn6JpVpub0uZWjDUNhM5kUbP481X7bSEUcoKeF
nmbwGQi3ZaeBDpo9aAtjodgfp0nbTM0RZ0z9rj+XKxW7kazRwL8+WIK4vD4ElWVBCOFCdgAldG2O
9NZBQ3zxxevej5qAMjq+fIDVbJLk9NLwacJQbF5XFHRLDlr7Asmpxl0OhN3aGoKrvzC4TdykLwBV
e2qNUU0S9SzVOm7cXsWnQLwKJNx+SdEATO+19tx8JhDF6ESdzaNREJIFvzGLZdWIYGTMXneYpZ8F
HTaxW//67xPYkzaO4MldZofJBZdeV4lhVi0xnPwrDAxC3NsAdYSD/UYuqN3uU+gYxtWkwYb7EBBu
59dO0iKvHzCpoCdBv0DDzQBgY/S9fcpsMO7r4IpZbPqbK7osKzyeho1gY6Rt9bOXc6TIuTg6Hcjw
yZXqCxo1ya+4JF00gk6FqqVoYrPPOkiuS6O8CP0XPQ8LrwyEy/cjHeY5+yY4VNlejo3mwaO0usTe
yjlQo0UGMlCc0DVDmMkrdZudtD9ypMAvQw8dTbbYtVaqxVP7HLC8OPWAt1xi0Rsg/bUg9+aSEyqe
miyRVP2lyeVG2GgaYdaHs72TDhg9ocVHg5vrIvaXnkzmFQJTC1f6MT6FYKkQJMUaDPBXImpk1FLq
YFAuioC2zH3ZWqPnJ//f9+Um3c5qng45EyU6W07HJ9iRAf/HcXC/KQ2nudYg/uXmKG6eSqYlPwES
bod7VOt4LSUzPF6JricMeXNxrJLKIxK64FAxAsZLi5AbeFulJMAcxjuryp8VwsCiOlJPPpUuB0QM
D/0TRNDoDdcwmP1irr0vAcBu8XmFq1EmMEOrAB81LioVOBCyqZ2PMKu0wLjot8fLfLvKQqETbc+G
eTIGcgm+iJNCpbP2ebSTUUQvvCE33KB7BcBby9mlQoY+ytdZRk6joJB9SsBkDQ0kdlZo/30QTuWv
a4Ibk5F/l+tcBuktrBbH+kf0ncZybVATGj/IgepYyd/0xi/VuFPLKwfPoiMtFGBOo/CxNvN9quwJ
qCf3dqX9XYY6dhF4PI4LZM7sFBK2gFvbXiZzf2mxgZWYm+MNOo5Gw3/VaxspYzRopmG0qYXiN0UY
6z97mDc+GlfgQQBPuQ4REDk9OFEV7MYYQyB+90qQkvyI7+dNY2Hbo+js01KI7nwYbjdV6vvV/BLR
EQAXIn3JZkzIBT7fKKUh94NxiipWF81/K7QYSthITCVJL4d6ideqUm9h9HVeMiBpjG56a704iMx1
j7RWy0aMiqfiJJKY+YC3OKF3Yl84o5AQsI/hRNxZSM7IhYwgJ7C9MDJqyyDL1GQG9pcpPPSKdost
8Vi2k0SU85eSMOSkAlhPCbvzigNxY/Hi6yfwkdkmB7WnJdrk8DYmIo5LAMRNifAPbU/ZWemSyKwP
FOSohDv0pfPGVkb3lqxIXdSjBypLr0mMzwdFUQ06Jl64kCt7EAtvfH6A+hVVbuqsnxLHyed17rct
q1QCTvZ/zg0y6NWe6YD9d6zn00E57k5pbm+1zz7qgrZ5oHmrGkYrN+n/oia4lt1rdz4aMBZ6gbN1
CtIPwFh8YLte3FphwkUa8pYgJY1vbnWyCo/mvg9BwlWsxC9sVjTegPUNnJtj1wBtkM1m6g0gL0Gv
psuiokEWhGSZpR9Qvgm7F2TWpooPdVOEX1IyIVz2sJV/4R1EYQHhHOcKY1GMFCOYYs/yakmpq8t4
WHDHCRsa2VNTJerjCuJbdKrjOTIttLfhN281+PcVZEcko7BqXayiKqFm8pqBcBQ39tIQ6UEfr3kE
J8qDua0nI6x0x3nKs2jagCbhJFTapIuTFvdL4gTN8+sDIZE5V2a7ozyS954Weev/IvZBjH7ONAQ+
Ef9GKQ4T8NQmcs6CF3rotL1vAea7afkcEmhZoQ9eXzUR3pkfLpuGzvSiOYzOPqbvxm6NLWNFVrwf
LAwVkMpO4yN5KxWm+z0IrCdLKQ/NerPktl9NP4fa+mZ1VuzPEWUMvylafTpq3qp057/XOAehQrty
1dEpo/qCxwUbl2vuXXi5A5Z6Li7H/Dw1plrjcuhbI4taKaz7ZU5kz+vKC3FjbcRMWK5MNoZudK40
gh+i1tMMQ8dsj4mM8n0Cwgo1hbHWkAk4s8DlBs1FZwZrk+0y1iU5yrEa7qB92m2+N5KCdim22Wuu
R/tKy76UTH09WZNOb7iXCeZpWHVzs3X8tsu2hAd3J7NHP4TuFd8ouVpgwPHEt0ngjOxRXwNjKusS
uaI8PIUjNi+OTpmT2ivld+8cxcgkN6qrJRt12OXd179bCuBckvHAUpZZC3tqoNe62C/LYbiZuEvw
Q8NX2Li9xF2jp6vn/1w51unbO8Yy9EhssAEcFgwuLkN9UgYncxCxknA35/JlImLNae/m3A4CApoQ
PJpI3iMNswiXsknE4c5t4D6ZZHNtb/A2FcyLkXo3LSKAfucsiLIYtTTovSqAw9ovfqDtz+nkPDfW
Y3dYKDltAr9vKc+EGdt/OVsBQe8XaOSp46Gf59REbmjAuTwRb9qupaMI5MOWVk7Il+wsNDobrPMT
zN7tJ8DsRt87d4MVAP2g+eRY8yqhIPIKJREMYxsgzvAszggbJXdsxtmbITpca0W0yzy4FsylblzG
N8DzRAwvB/kvhkEn9uv9JsZyxoKTazadX8g3MLWAt6NhEdpolIHdwSxNXzlckh5QVUEqOEZUW3v7
bVU/lY2IthY4rtIWaLoWPIhX62MInfRWwCstJrcgAWM0aivkCsBlq3O2PTFQgUdnLnhU/n3G8sUR
6JW5f7WAmH7lzrM+vImTNMC+zyTX+TAd4JEOUZSRgwf+n/ev8D2545/PG40ZoRXaiC9I6i+kFrEY
z2wm4Qs4hrEJAfrMGq7q5RTCPBpRB/nrdCQCG6zxwg39I6zB8x2wvCKujwGF2FWpSlJmIcPWZd+5
rnG6ntQVj8pI7EhEk43m/cmS19qGcV+U7SdEx9jlityGNn5r+5KRW+Ukst0HDb6CX7StEf6ple7E
2br8fi7/8r8P7atqRYbww6oxYQ9MGX+eVLwZ1ANlP79jo7F2c/CBxH1/sM4btRdfL/wMv8gM7kNR
ujSDmXfLMih6Tx3lpcZKcRsv5upjOuWdCfpyd8fxgr7d52fzhYLSz1zvXu5PcRxCFJFowsG6SDPZ
86kP57r3nB3fDv3WrK3EVgxdsJ57XXMRnvaNjQK7BxaA6u12lgbO/qPLyspFMO02o9cqb+dmGCvB
ubOymMIw0RwhgqS8ee7l0ga5W3m7L7vXr3HS5Ge1fgfiyHU0TybfQaPxeECSsfIG8dsGazEiynlt
PznSyFk4yHuJHsoF0QO9G8ZzYMUV/4yhzSILbH+QlGB0hxxVzF/4ZToI9WlZmIG6NrLfQ7X1zZqW
eRfrJ8lbPao8/98z9ZErChpHJwFuDPpkei0sNcdILwkkxx8TOebfALoVesG47Gut7qkG2xjihMhq
f+LN/dnPRDMjAV/GBY2xED9X4b4dwQaHW6ydl71SWBxIpbQwGBZdSvMlpTO6N1hGJrrbNjElxV9a
cxB2vbPh+rFCD//25A7MlwPLtmDdStWOqa0awVeWIO3956HO2Gm/p5nsQm2k+jLm7A1IlfpIudO+
sUnqE/l9ONYaV0+oyN6qCE5m/FO84zSHjRumfBDHHPX/xmYAJFtC3dj9bwQJSET/MRAS+ZFzaC9E
a2AQzUviH0R045pUlnTCC/zPe3FcYg5J/i16GRoIY0TcNdJdAYquzG9yxaPrtMmIcrVtk68w3jdg
ACpHvkRhoAUCDdd2Vi3WbM3Lg4OWpEu+bCUmGYooSiL8nGnjIVzpcNsi+zRmdRa1PtvGhkHYLz5v
h00Aa1QuqMABPheAamkV4cghKPQ2jem+04DSstD6cEyZ1tt2r94I8nFpHLQ5/JkallpfajoOI/CQ
qOFKX95ocJY8YpRHPPJ39kWMJiEMiX0fDPKrhDfTywy8L9yVuZcfxnAqB6QhD0myK0c15xoqIeig
Mq1Bgn6pcr3fSX5xo9w6eg/jpw6zBzjGJnz/i14GMhOM0K5u+m8O+h51Eami3S5yWqUUYwEDYr2w
/CVWEWGiLtKoaXrvNDpvCCG8Prg5fysCT3fd5h0q6XXrQXu8XnsVZXhunap64nZUFuvlxvaOdRng
ZrXXwBouPVn0QxT+1QM2NYAsWAOaLPwyzJGq3VI7tN160JDmauPyR9WQ7ip6zOsxlN/+PhZSgl7Z
ndOOsM/Wb+NoECgkDB2edA2Cx8xHz8xlEuoPSl0iJnb0CxOeyG0IoXd+VngLED/aTWYkMpWy1+eI
gX0BYh03pimSfoTpkSc/29yebsrLJz8pIu+gW3udk8QR4vh6M9UUEGCIeGKP+rFMOs6v837rCzN6
lXXk3d7alptu+HIBaUOrE6Bt3ZC616rY0KWoUWjyVYPvS/cLDLrSKHzQO1LMIf/+jydVV98dlXAi
aCg5OTeWc14PPBbcLwFLiA6lb+GqmjW7ElPmvoyMd1bhkfxrv3Hcee4RB6/ntg+sS5h5NbKqBwKr
2dNGNup/+Y7qxCzAmWgZn8vhbcYJtKiJaxj+dCimrnf9YZXmjP+aihonhNPKRx45j7eUtqCQkP27
qIw+AHgBvjWvE7L8B5mSTQP5ShV7zLAIO/mWJXnK2+MQOBgQ19Wrev7JZP7k+wDY6Ej4KNr0w1Xt
SEHEjPys4AFZKSvnmPLodMAVPsYaJyzgnAl1KNEBt65QFbo/qeS1ln8Ocy6OcpC2SDHTvpKv9fpW
cM8d2A1UUUvyEt36qoWan5SNXiruc7fD+bkl5bgV9O58RqK4JKVYPpHz+bhKxvI8LKdJhoWagJqA
rpLCaE9G6wKRQ1lwPNlMz2OLx4xBzEefxYAistCV4oaQh9/Ra0KFlZABAyHkRB/Sg8ttOr0DNKe1
Rl6df1RlIj81tsocrViYz6X0a37IQ0Ah6SfIJv0ubKFK4f6Obn5JPSgLx0xbwd5QA8YQUxwjDJ1S
rJwtIdEXS0mR1G16XpMEw2a1UbGqY7ZWsSb9r2bYOY7/a0ipHvsfWJZHf7YcHdCLNG0HOdeBWawL
UmldVXS8OLi12glZ3jCd2PtQs/gaU5xRGCCrD9/3IW6mHMZRqoo+Bkhx4bBqBezC4GoytIn4XLzS
mQPk5En19w2uLdc6ZIVvXcVRHm8GNdM8tgxPoLmqee2e6o+RiKL9jIFrNTCxjQakAi5AO597OmRj
tZYaC2K5rIK05jzVNYXw+mdSPLrI3gTaJ+EqmZa+ip42sIyUDQwLsIYfejbGLgwZY0cfLq8H+1uO
mjQMcsLbYL0LunrwSnm2mL32cvdebav0CYGFaq3QRRrya/LddjBRR8KCc3iwokGgFl/UUxElHgjr
BkQH+JI1T8diZA703TFGvGOhNMKrCm5Dtr7tVfSJ9p1BZrqAHzWAUtueG//G1/qp6IgT45k4q7qV
+xOaemcsmKm+r2UvYpoVlkTm6BtmyRuTGdGV+f3fPXP3Ck3xZ2zuMO0qODL20gurV3VdNznwuy/g
pInafWFomV5YkPjlBQXqCUoDtJmPPx4j+sf+kLn2WaGQfT6Qjjg6XTMT+fakH/48KQOkvD6bToCU
jk+UO0BKFKd2MWNb6N33IORkYzZZywGgeHPkoD+J8CM8x6qXR+xsNJPLlmeUy8vSBdc+sWjMkmTY
o95NQVpUejv/SDU8YioPkbORywQfRWb6PP/YHv68916kp3TZrTgX6UEFBDvR0x60aloigUlH9ImJ
dHQLUltG1KcWYE+aosK6fwj4nEOjCoNlCo4MfFUcY/+scZEZ0TTmIzZ8bS8920wauAj+iKmH8p4N
wjwXE625oaKoFPEyubdE55U5CbarKNlZUuATkQfd1/JFMnTl1Gg/ZeeNS5AKqumgr2MJ8+eGeLGB
3mm8YLhaOOCwoy3aBK1LG8+sc5GvgsaiWUdTFitBMlbSbM8tgf6oFQUd6sT0nXJnUjbkQjN/pzP0
MKsPdptIQ3jJINrbZ25hx9pCm4/yxM27PzuN4N1q5lzuF3gFLFEldOdEdSaOeUeUbzvcDpcoA3hH
ybnChTTBLlMP6VUB/2GjAtcUVGyU6rss1erf0loA0lO0BhkUXIqEvPDniyE13P36YdJ1mgwKG2Ms
opsCm9ESiughboObBa5pmRxCkwfO4CKmq7sJudkrKdY17i0SaCNXBHDvV4g0mcbO0rLbSaAP1LS3
H4MxcYe5GB1wUQYL7kuORE4uSLoWcZsBEi4VV3NjEPyogFaQoKAw82++rnMXdLAqhMWQoXqhE1b8
ytg24N6Cbkshlhgld5pOe4TDwFlZrnfwKEb2sTO7VxRmWYLuqReRzFGp3FVwTJR9m/Db+IQvsXSy
TsikkXHe3yh+PtOm1N8rA3ML5sNR9HuLWxdk5qXuDttikm0bySXaxtx4P41E4LXLAfsa2A05R+3u
nyT0BLCaqvivvNcYRWkENnEGOpqZvUUzWHg6dlvA7+J8JfuQ7BKUJjzI1JpFgwZUQXozjN1D8cbz
izLa9RW/QfXDu8WBZNtZTnn4fVXN5href0qNglpgyFOFVLMyuOrJBZ38Fcs0WXJsrb7IKn4zqtGH
e/0Dky5g0FPm8ZA3pnidsN0KKbrqKxIgIRPz8d5T1BVVNtknwOAm7VsdLvZKtLPi2OXgFFanTc1Z
wQuQ+VcD0MSTWWLvjO1LsqYZETX2Mb+3vIc/JThOJ+/0uAa1xEkZviAsxwm/86Nv5N3peDOhOLQE
yFoUmKPBxU58e+cG/iTTyJElxYkdu183+w05rZevPhq+jkyrfxKPSVfoqESX/2qR5oXtn3gJ04XJ
D3CXPx1BuohHK3kvEFm/+g7wp+M+XPV0k5z5G9NbPwhbZUSnjKMkTszU0whuI8b7z2vLV2x+jYHI
ogkuO7OgqgJyQB4aB7o2u2KmYp+oZRyT2ZSaJT5B+8WXeD8cyKLEAD9kdncvWd+7x5Jh+gJhDIAg
JlFR6V81iOcOEnz6t0cCO9bgA+/m//M2M5bu6mGF6KwcutnxL7Gi05jhr506bWBfgEAXRqAjgsxJ
kmTwEMsg4j8U0qTj8dVvPNFSW2nkg8GXgcm3GJbefIwQPzPH0uq7D3FKkgP5CqSZYL4uQ4qH7a3/
H/wdUXhzB1HPulJJuiaFCv5MGzlve5nEo6c0TsnpHkl8QSSZCLZgtz3fVWP8DIlLxJhnp3lR7P+m
LMHtrobWGRdwU9j6INmSy1oStJb+hXXq1HDBHgbbh2IhwKs4P98Fs6nsUKiB1kuTEfagldn/C+0j
ZXUQHzvdMwsbXbl56AjL/AS69HQFLisTNUxmuCrLTYvB/xYXnhqwNHYvYpcddy0TWS+Q7RN4m/8F
LYTlq9XzeYipREcmAiU9/8oLdZBugr0FvZHROfoSc7jd2fVR4N+eKpF2Yk5zCuitcuXgIjwo5Bn9
tJyqVDVlYY82wVAvvNjte9TsAQSvMtE4/e+TBDq6s8wXfGdKoTEodPRNzt7g0yhdq69b14E88JGf
0C624Z30sAFpcjIazlId1WTvc+HyeCtlTuS1HLS9YiHRjY9KLcEy+CqIAmFIBe7cb7p/fghTMd36
E6G0pV9MVFhWmOrl+HivLDMBbKKtYymFixoOPdDEEpoDEdQySKaPHZfqZA7ljqkD+WryP7RuhTKC
mlijLKjbQZzyW6/E1aFZvMkFPSjSOnN8JK/u8ib8tafE2o3gTyX6bSWy4mkIvzf0bvEU4oqE9DUX
1XdAWZ8+5eMdIE3jITtyMQxpZrqRquTXBH57PNJlbSN7MVMZfWFJd5kfW+/pVTMrZQ2grheWZof2
aX1/kTldUnh+micXbrSTkd4mXWOgcynZ8fb8Pt2lVpVqJKLkeOnDYDhaS/3VSdplniGDJaI24UrQ
btd10C4mPuBLZw7jPTdo1+JAg7yGv2fPU5gcH8sjsHQSTzwb5Lzpkh1vVyQNS6j3FbZIRStNMB2B
BMKunILfhviJaS5X/wTvhJMhVe4N4noBph0Vsf2vJ1dwnBlOLHsfV8GwMNzSXqxbnV+jWGON4WIN
l/e1CCvJLayiXR302mLg6YcKVvgMOXFDh1B7g1AcDW2JuXPOKpXarLNL2zokrb6O7aKHyzShKJpQ
th8WqceBw9IljRCXfzo6JWupOs5pZFjWZwCAfJ4xj2CtrUpMfSCv1Ov9Y+YkuMNBC6iQchpRQbr7
qDmygZd6Wgtop1Ls8qcAzGxbA4z+1JR9NY06xwGnjw23g2bgHh1JXcjVgDgotS0KzNMw7N6fHphi
NvHXuDZvsy/CtwUcfrEfCk5a3UViHa7D6i9xX9GeuZY1vpH01zPCM7oW8EBm5EqncG1ykOfRXTmd
aAIia45Q8aH8Ebbn806BaCSDCxRyf3Y2z4QUJscR6lZyo+2c/QAsdIIBmcFpjQLwRuGXhwMyMLti
aCNPio+/MqJIUlnkZr89Mq0ugBVaqbUEycNzImi27hbeFQtyNnW3UQwT27tFWRLFDnwVCd7qC2hJ
qq0Q1dGxFmtxdNPCs9Kb+1vAEa6N7LDR4Kar2Bd6Ujjo/eDylJNEccvGyGeFEgiRjboWQLyEKDLH
LjU02I9Z+wmPYvS6slU4tBHf1x2tuPeYI97VDqH9tkNsLpdakezTdQ+6njvCQyT9vcYti27vYpfm
DGgROqboNWIaZlvWeCVAtn/GTtyw8lXJmNwes2UQqn8ifOGJA63DUrEtw6JxYRRPHe6WFgVsz5FR
NKIUL/CaAbsXQEYYnqmntIZVijh6V3FCriI+7Y67a2UvDbDCXzrZds/7QXBDxRaYUxn55tyIafv5
ws63DvAJ4zE+tGXqSyax8tOnembSIqX6jKv8edMZAk3RDPjsyKGtIDenI5Ehw4oesxA9Hk4th7AQ
SHZNDAU9kLOB+JqsRB2enalggp6PRPFg0U7OpegAUcYYZ4PdSHLW+WnhskXAqWiPW+66oZrgy9bX
WvMWVRkUioO8PMJTN6CkXM1lkOvApJljqydacEtFTpGcgNPjycVzBJdQ24Fw+5aMXDupD+P3LQAq
cDQR32XDcIQRpo1DyDe/4v/rdpzulZ3hsDdISZUBetxjN0nG50p2nmfFKKLNH8fsDQjtXBo1mgXG
HAuB8UAUFjIK5ndl2n1fsQfk1nonWvyBBhJtqvhVak+cAyr4Wv7BovGMubk0DnGnwpiXe+uD5mgU
2WSx4VaKmlAlpaxyfGfhzK07rueEIO9codp9ESOb5YlfpRgXh9NPRnAl1fs9bTBEPxaRAKsW5wbu
KFiL3X5q/N3EstJyOgFpEy6Yn/rWBKmyFCKSa2A7lWGinhmmWGR/7VzGubkNOOkryCd1hHH7wazx
3atbNdrdfkVbBs2HdzDJMg1utbKUUgD0wdk+sHPUtARdCW8dp5uVdzFbYcvnjj1jMM7Agsi5LAcv
NyDCjRHhoQ+tiSeO3n04EpbZtXHFs9dpQH/BjxHkG6+RlYCMNg93C3WiSj0z+pGw5suosSvHxDMm
hGfTiBoJPp/j4xFvMyxePa2gIuKCvZAGHn30ztdAQ7znKTo5NV2iyYZKHvHGec8aw+vmz30dL068
7X6tjPHsQEy4N3OWGuRXFvpMafITP7+etayEn+30YfEstuu8W8lWTOh1SEU/nHioso2nZOTVyNPF
1GO+j8sADuZwUAlCREm+3/uYCWULT4klHOUEAUjMqrPfHKOsXzC3WTCmZPqdoAg0TymbsUyoGhFD
gjPnX41fTSXSprFTxMmXQ2njPAGjiSUgL7L2ociGv1A2vpBfagyJ9vvV9PO1yFnOR5l0uUvdfDjU
L0ySu4LqmM8d8mDGl4kqV3kZ7146DaqC4I1o1exSuxS9Du7JfNBMuLH0U2gzl/jABZE26iqNKieF
rMFoo7sBxNQONdYecnVmh7gY/OXqz7t4zlcVZTv5YtHch3ES44l6cbpLoJeD83igrAZEBoJVVW9P
0nucftoY1j7Oh9jCg+thp2BzXF/mEFQurcebEVcJ5zez5iO6cJfcdWBgs4+ThczhnCEkH8g106Wo
8Xm0ICnPHmxmbezzVgFAkVkhkgOq3kOk8+U7DfuRb40sbbv4+IfqksDGtefyOXWYdW1r4UUjNPat
gPd8tKs0aNdnbgzSupu3Aof67StSIt1/IsMRnxYDnP7/6Wbvv474PSHoYfTVf+R165jS+N8/IKuN
W7Gzly7U6W37DTjxk074aAQJXcYdzmoaYBdCMXduTnq5ppcgufP6bjoqqmnuZkOdZBDrTSP2wWC6
ODH5EL0gN4I+PAKuIN9bnZZWsiqc0yojMeFBrHqVq/kb3ktW1sLgR/a0jBhnijV2QuS7A6Y02etg
8DzVtrgvlU0nK51Oop3uW9oXzFXBQ0ngNCB7mR4kpG0UxYZ+iXWrl1x32u2+Q5xeP6i1OGIKMkxW
jc4Mj6c27eO6nwMLiFGPhnJiZ/6S33yzZ9pNhNke2no/80lHsdoo0h8M+kEwOsfvTFK2j9WjQdsB
U3SiaINJJicLkGSBNf7QmnQ1nzecZpxXmjuiXUba/hUVjlSRjvEiWvw9Y8sfVkWFbW0JfXzBSOG8
DObIe2bKmgBfjbWUlnZnfC7kaUwo1XTRmm1ocSj9eg8zq8Smy+EemAvH/MrMJigOpKUeygVnanEH
0dmIVPJVi5WoRUy5pWV3+lPi64IL7w5vuXqVGNhPE5t2KIWrdOCQBDduj0qWVGkEtohI9FflwmfV
ZqqEHmVXgeO9pL/NZa2SbAtxWaMCy8DFUylz03CSA/1llvELABq1xacx/GlfKSc/nOst0Fq5ANqD
2V+Ru3VeYc3TqiCaBBHENmwRCP6iJ7U5vy7lJqj3zv6CkCo2wW9VNRrVXvVZUxBEvRy0pCKWe20u
GQgd+/XMViCxQvGn0+Xtp518Lt+0AF2jmXuPYAyKermgIy5h6XlDuFlS0t6O3GmHeuFaZe58RNay
TGZtuKbKgseu0R/PGIWQ+MWZTXPO8B3C6UMSNj24f5LdVo/OzdzOBDWKL1YJQACOfVMGjyukCw7n
fasSixcy+Nj9IOtGOQL/1Odv1+SMBKZ3kCe4dvnZvOnemwWoBy2ysM82hh/GlW8thuzhOb9HtBfB
fMJB8qwWfM0bTDODbbX22ct/RJ9QZ6f0h1ozHHmEhdMZHWRL2JM7A9I3/F37AeDHNvxUtfoXh7Dc
NgugLrR+/6klpdnHlo/29pcFT1gkL8R5i8oT8EOLbLM6Ew1Nc1BWBvSGDInq+ZAl+A9/0TE3cIl1
ky12KH9GgHtBdAxuWadWwKt+KOOx4SPsVB1nXURwCIWSk1UMRRbAVGiUxWXMP4ypx9fh7ECAt2sE
ZvUS6PXPaKLL1e1JZm8GdZLnvp85olE/TqY/kjpnsNRtwIv/uVTHCBqI7loVXqyW9QA9uW3uHJ3A
9YEtsgZ2CXmcKmn1tygU2XnfPepfBpkt13g3rnRPmtJADPz4Oe6sa3tOkEyfAE/hPd+kQzUJg95x
jTlriLzgwwz3KhwcawAoPhzYFzdSuC3Pr5BWNhtKu5zWiAYVoKaAhs7gl7Sr5iQ/bWKM5Hrm8pLT
tuZdwt8Mux+FqwslCTtyLluljOzQoofJiXLOZ0fAIfJL0EkwF6ToK48IA8PSJpuExPEczHvN0Lmx
RJXuMAFk8yif8SGLBSAfXhqvUlR0FerocX4vYHlNoIRguHjmv3UNAoQKzwlyN08Mk0qHTdZ5hwq+
795VqFuKvpxwJbI0eFt4GiSsSUP6Qu114gCjp2ZX8kkE9qr1YyHUwf1dUZxCiwp9gnTl9NgI4WgZ
RlOTmSM79weSJgPvB5cITcYFl07OtcQaB30BRp9YdyChJGNT+4zC7wZW+6bPktxW66Ndo6/pRl97
vLT2MfnRLDhTT94YM+A4ePuqOXc0nOVUVtJhOhYi7qC2AZQvWeZseTF6d9Aw+LisKON6NAMo/h42
WbGGTqUH8J3xVC9JDeVsNEzyaaBM/mfL9jis6ez8SGTBowu3EEs6WUv8MhvEvxfMlygIXGKO0/6J
jERqbCe7eqbr0+OqZ4v11k7c/GfNZ0F6qXstPdLWwj6jQjIP3tz8JAKJh0aQisRWBU5iXGX4EiHs
xAbQ41Sqtk1CHajQAp6lCAgyNVFPn5m9d0YS2uZVos9WDFNUwy6nU7V4fKZeSTPa82hgxj/2AMWS
UsMclN8K6e9AXPYuO992/AIFyqGa40kvc9aGx3ByjGa8LmgvoC0glyqblgm29CvZS+Je0w+v1y6p
yl/KkyZkDobwoOXbcnEh66kHl/ApLM3PesSxjtAAyenI3WT6jXvZU39RMS9prICM8FU/3unUXnxY
xj4EGfI0izLpwWrfMhS1ZoRReuMYYWUsPZkwtC0qo2q0C4eZLpRRb9URitL4jVDWY9hHUQH9aD7t
G305H8BZ6MpZ2OEbjMdT2lLPzcItF7MmJ9yn3RFcMUeiK1bO6sV4QRRSlahvAWKlG9fZxKSajGpa
AaVuqTOqiRUG/kMs/G2cZDDz/RfvWORsdcnGo/0Wjg6YDHrv7kWUU6vw43GttK0PI3aii+agc0W9
DNVeuGhr317tZbxd1XIujeOkaWfbpIe1yMTzDUIBPMua75vnzPgECZIm9CS8fQKmcsssM1QuyeGs
ugV7IMD1hPLDS6R0L8D+rbNLckyricOdwKjuJu67OCJyNwVtS4Xc7qXR6lFP/0RA3DSLyz5OH6vy
oJ9jSHKwls6F+HjnVlNM6bkMeTDk6EoV2gc73ns1NEkNEYKJnX6w7xtn20cG42Bev7Qy1T5cIwDH
a/K2gJHSIM8QYYmvW2jmbe5ekXYnwfen7Q1iZmI6y0TmDFJSawrMsakMd6tTphUymIqpKREPaXy3
asfbX+6ADU5uVIHeZ3wl1GpxEtyA5DfjRi9x2Da4Ooob+ouL7KGLXeayeALOqGSAwK42sdJ57ZOB
y9/zCw/ApSenucVRm4xF3t6ObpGpcPH2VXuyvc3tRj+ZyUaDweuX9xt9BeK+U3KxP+mTiEsvilBo
jCDlT4jAE2A4Fb0G/UZ6/jtJ4aZgsE7ttz0Drq0DSgjLkUN2F8P+r264CPqCffLo7vGguDUMBGHs
EGhK5lt/72lXw8L7rGmzdcKyzG5+8eXmk8CVr+B+pqIwjdRHvabrytkUtibV3RxF0doD+OFrn93H
LnSUFx0vdQ4GXLnIiGNIvHHvJUi5ugkmeILocHBpqQHk1fftBV2nIDifcSABzxu3RfmvUqngGrFb
6ILn2zgxOb3U2o0IUL3bzK/PTF6POAT0VZa6ldUN2rQqaOPeQ1+b1W5rnoTtvhjXlup3uDSygx4G
G8HrNsZsJyT3rkpmfpV34XCfyTfQZHdB0XI3tntpT6rIsAzUIRwInOZNvsBdXOt3SP0dWEPPiM5p
4VJAkNDiD8c6qfYCWa1UeOl4qHBAuSju7RGAmvnI/0U04FAgacUeWKsoF6NBq5ne//++3s2fH9iF
r+xbOKByRN+ECCz4ohfKgXO1uJmncIimH2oAOk7MDe7qruZbPVBATzmXAcQIXnmebhEN8fOqFcNo
2ncgZgEDUq50u+4NIXFulNvCF4Q/UVuPr5Pz0sPw9C8PbZC7ge0KUuqLoWweYZOL87P1zzL89lQK
94b4UulotKvXGK78T4i8GXkB+RodOVxaA+2Jz24VFPrZsjwBR/gmKq4W5RE8YEHGOfRRmvpV7Qa6
LtQQ4qwklIHeUlVtCdmFmL60WDi+aB6CsbKMwmF+h4NI4QvYFW4EMODh+E+ihxwycVkOwNmEp5HG
UyauxTv3kVRDIS1VGAdIRMdVnN/Tle2J0ED984NOulOfAiaXrk62D96BdfbkhTJrvi9jKvmdPJ5M
bhC2sH6c0w8wmxBJu5tQsgGBdr7kI6xMCQak0q6Xcz8F4RO9nHqYDGOFD0g85kEthQ+X0wKWDwCX
bRH7bchwLNuhgyUtcPMW4b/7eFgcZcrOrUZSHx3cHLFO1sghmRblGGlBwQknhKFKPAGz8Z8zVfE6
s8j0krY3rGfQX5PdntalIyjljahq+y1nJimPdE19yvS8UFXLBPBfA9sCEYmt6/j2ENvBnWo8gmS9
uk6bJa0KK9ocjoNaNWfL37LrUZMG9ZseunrLhAJqMrU0RqmvVBDLrWfVilQ5eIu1D7PI9QmRosue
gvq6hO+3op1nsPm1jXVmV39xCscgQ44DbesaA84Jr3j1qdCrwnrZqixqVTJhQGzVU/+wUOWTRkqM
2x4nlv1XjIUW4PYUe1i3NSY4bkNkLYBguP8HaJiizvXq/YOcquDCJVHYvEf6H3J8SbA/bVMem+Jx
c+pW6A3Jb8NOMOtaHuJ7pdG0tGEUk+v6JbSE2gqcIVhNzsoMdkY8O8vmazN83ACWpCOS7oEZi8Dy
HRLbPWLq02wSZSrUUc8ABozPNdhEd4fG0HKpCQ9wSPzv6irluTUs3K/Xf0CigOrMUsC3ppdPuNRy
Cdn/s1Wcpm3aMw/lCHDYxDW8koZm2GOjimy/jAb/O47Ag4uhDCWBOviGOIC18yM5RGcK2kVFJI/1
gESINV4k1dVHAh01agYqw6Yhmfzv/tXdX1+MtrcRZnC5sGroBP9cqZbCAW/kBN2OukdAPKtATYKc
88LGkW1mdJRlH/y8P/QMJInlbv+ZFWo8INLLOlzpAGMYIjiTYc0R+LmRWvkWwDxxMu4ETJbMoa5k
cyZy75LjyWVooKcxGjzAHY7NB8+Nurv1K2hN7zWB8i9h0XQEovPyxDnj8qcJANgkCfoYlbkGLf98
D93O7rGtmv2mftO+X4AQA5ik31SidiimgTRLK58NSAfCk9Kq8LV0UifhURRWWECWaKYcGNYAF/Bs
PzeWZz+IkMSnV6TS4MP5VqBRnWshcqm1YibLQ+k70icYJGJ+mUMf+M18mrzLgQHDdA8uQk9xFXT0
H4wCYhrqmFdmN2Ung6H7e5C9DAIeA1GQ+jIg4mvbIe2ec47XnVl1iq5dOSvwlQHZWGQxjTxvgRV6
qpdv9+2kEgig2quob4SR0kQRe24pQnqzyCqVdK8tso43ZH5DzEvi2TAin7hlH54TaK9POvGoHLax
GTCFZ9Hs9OGn3j7ULtAfKZKY+UHHr2GmAa9pT1pShyU3ePkKAh3ihczvFxU3OwbiBKmEuhyDxHM9
6UYzvi38Y2PbWyFtmqClymAm5Igkk99254xg9CgR4Wzqw/7FetoH9lo5EZ8pzHJAK43g/F09REBc
bOsGgA4i1CZdtvgwprVFh92ipVh3qgHqrE7NdgdJJHdwyBnJkDnOipuVETXlWUkiXqqdh2RjcT41
oZZWDaw33GKsYM5ukxER89NVgNiYEDEsejFwsrPURtSe6086sJ1Ior9L2UHMigjvVM1r3Cx3Y8qe
N7qruQEyV1KSRjt9bZMoYNcu3cItgIURdb4oJqcvmKBWPqU6c02UE4T+GPW7QHNcZJPIt/27MeJ1
/0Q82IB6tsJWrZJGQUc1yhKB+YVI9tBgJP9+DCgGq5fHwMV6Diu/AaamB8N9cj2R/14d8xMB6rE2
pBUOWwziqMk32qMN84JJFflw09RptVXDC2sQ0rXBRbCRl+wNv+/JUAMYOdww1nneq9xasRo++K0/
ifr4Xvu45FqrKF4E9ujXC1ltXY9bZPdAP5iLEr+tN+EF+IeUFAAGmuKqI06DwdLAGIJ5qy6iln9K
nvvZmO+29LyvY2Yx1xBWU0wKJeV+WyovqVfbytc9NFphkmjr9B8Q9dFbgMsu85g2QNa6FHqw1P6w
gedAGUsDdmhDeblxi3e+SkchjZRmci+XmM+2CisSvXypEiqH5EFGJvlfOIamZsTjPFb65ZSGvSyQ
LIgzhFc+X9zmNDZVhg1AzJu/bI4T2Vb7NvtuNrNDP5xl/XgpNwXhaUpWWBJzOKfeK9lqgiz1d0Ap
TEIvVpH3QgHSTJv8bzNU1/JhnJpY/pK23f8lHZl4O1LfkMXsgg/2erSArOimrkpE/QBmym3PKqiR
5Rve6joCiD0qA4I8knYzlH0qS6ZWDrrIcHdbUE+z4EZ+vAJGSG7i1ICRFhsJhmVVbtBPh/n9l7Iq
2y/lZbOWTJh/amBxuMHVnJ5qaRlkE+1+u05H+wpSqtabt27t+TRTHpV3BIQuU1rV8CAW43Lx0HC8
uGG8N77XBOLPd+dPG53x/FY5wQfombSeu4+M396khi9e3cLuH3XbqD//jUZLCFv4uTko35uatd+f
MZSSd6iVEy+CseP/ms/u6cT3q8w/NG69RpVZ6mg6JzkzH/if3Bke/d6/qvzLpSizg2PRiHzpfcYe
frCEwQTFjDneUQf3Ha79rJx7u6H7SRzU6jNG5yPGLZDdzsOb8kpY5wkkoURQiHEzzyw4vfMIXeIE
gCbx0+QXUeZ97VIh/ISw+ZqHkCx/T3cc98FXvku0C8F0wTBglH7JHj4je/sv4XVZhB4NaQOcNECg
h0hFJXa6ONVgN9dqwD+fz1WK3lcVkmAHZsjU3GSdhQSgsl6HRyypK/V8jrIJdo0mvaRzoIGK5s88
vF6qVgJDbs13EXLXmoUHh3umI6NC4S+W4Y75/ZXXfX4DRpUrfANxZDWnPxyq/qCbFh+Odu0Lgdm5
KdFfAjbSj3soHMlIpmHcZBy6TMURPbkDOKNC5QkpCnTXDoVPJDTZEDUGYulzhT777cJ6oQ13UYbU
jhl8BYf0QfrFmZgHfOWZZrm7yVUqQuVGlRD8wTIKBpOhbHQepVaFOsA1AAkvLwxMBpcemAv0HfJs
t+89TUUVbJZBRt+XeAH3Ieibg2qULadTJdLhiruAge2asog6C96EAbUXxKtmq6mfuo6gvgvrcrd7
1BEVPdMSeFwYUpZdnS6SUnVaitdn5SCNoOmNQH2RpmmXPZljwnSmDANO3lseUCy1032DPnm5ro6L
cJk/4LquMInr9uvDxprwyBGM+zgsOfglRrqm4eTXBTwwVtGt5W7mz7R+cL8Fx55WLCiHJI4CK6Ym
tT6CKID4sJEB1QMCGka+CmupwXviif1TFYYJMrsItzRLDsBkq7r+ZWEaZk6nDIa3fWSIzqcuILc2
6SPKW6F5jy4TlC0MqY1GFhYn2O1WI7HptcFd4pEoLexVX5i/VftipRaCFpUnDkp7KeQRKPKpHSwB
VN0CzwipZ6WYCNKdlEL+y5ETkomQ6LPtdwoUAl63Ab4d42JD18RS0rDsHWTb8tTQfIFVILIUBxV6
HYbfZMA5xsIV+InqAL5mXMNYQgBQ3aWfxpCOGZKvt49v6h2JUIB72yD+Z+mS29tQKn60EmSuVXg/
uqSLY3AEMJfEUsv2Kjqh4iAt3O0cQa23g9SuhJqwjaAPMSIZsCsCN7N3b14WPi0UfbF9UtjfwxUk
u6nMeM88aMQ3HJ+a9qYptFD+6yyrE40yUv6ooRUyGvU56RwQCQcghSMnJOMtoJKlVDtE4sWTbvUM
jZJHil1tMETTERO9jGRIblJ3loWAVqjBtHvDpOAROldFwU7Gx5TuKY3tEpOcfqq8dXydS2BNml7u
kHszuEWGqadyZuc7o5LR5o5Cuu9uDwV/j95hv8WLJvfa/3n2iAzziqlOT7qe4tGC/wqUr/d4+XRO
Bo9o+u1isMT1YOhCRYmmuxvHkS5TDH1GwnYIXFS66BnOMVLY0YmV8ivFzHBqB5H6o/zlRhuqTDZz
E+M0SxzdYCw+8yKjBmEFSr5oIX2tVki59sNvlTxZOsh5M5LeGFsfIcJdfApVyjf+x84GVbiWEW8r
YwoAHseJgkhfjmCFNXVgjUCErVEZ7QMI5EUkWaVmNYaBEp7joIc+8fdYk7phu40yh8ATf0ixmtK0
so1huBAQZGrEuu4pd29AwlBt/3Joh7+aqiZowjYz4+SswSdZZ7VJDa+801RBhJwTgQvRYrjQSC2L
i0oIroVhToPmc11VPuIVkHNavGOY7RNQTrvvDT4ErmePXg0cxgo9P5xvePHC9AGm1LauGGJMCB/O
NftIPRdzpz7xjZXNWA7KDPqvYm87Usr3dxVcXMJNwmIZmHdKkre5SqjWzRbXN1aiz5FSY+ynCSjB
MVyBrF8WmDsssSsWx/s93BavmwRaNUyxChSkqWw+ZAAhDQsYz+zYBz57ZE7q5sezGGYZk7sJUn5K
Lq6ELEQV01XWi+tgPKKGZ9Q3Qu51H3Lk+zqFz6Iej3Piwiq8edPTI7vhi7Blc6e3Wx6yheNwGGNC
q9SuhkcrnB1mySlKHIhjJp/bkSiuPBGtOvUZU2tBq7F9HFmRR+1Q17DW4YdDw/db6ekiD9qWDAz3
9s32HPqw0ePQVQcoonQGiGtvECqpIeYibdU0RD8y1wJLq82HGuE7ZzpqQniaTIZtn5wWi32lDsy3
ON+D/aqOI/BtKtqBdWb/Tt8ZDCQT+lNDDERIivoipNTC473WzFN3FHT6mXaqI+kWnjZZmliGS7fe
Zq8yufoomPrUkZgWegCTmcm1fNFVtbvTwfVS2OUQ3d3JWTHVb2eJdJ9u5HYYesvzcTgSRGSBU8gU
IPD5CPr1omUmEMSSZ1QOgzQyUNwE0nmenzL+4q/Hu5PSGUNy5doX2kRN6Qyn+HpjiuELAl/uRKmY
BKBa2TqBfXw11PVWGamCJ1sBWcCiCwbS4Rg9uk0yTXZvbgHhdKiCIAXt3I69jfL7VOVzGRXGl621
SV1kH7+8lZOTz0hkiFmOBxQaFeUFXijrx5STHN9IxoWbTq/HOj3VIb0c6WNIIq+eXMyAapp8TF29
3rl0STG+Kzc20hJQGQMNck6IKXqFz6OV0Q8lN9UKJ1E55CNnnui6KBy4qpXuFcpd2TxGWJaHNEZp
fxBjd5nxsK5xNhXjKr8fPOQhHiWjard7mqF/k07eO5ur+uEgsIwrjiTZj10H1t8VGL6bplinCJUy
Ownw4stezz3GaS7r/YedQYsJtPUrQ347OnWZIr3J051ioC6GOAoP++rsl99azbIALuOJMzcKMuvc
UpWC3I/IbF1MTvIfTtaLABBX4BXtVCGaCmglqPFPTZnT4+LLam5nKDCyPo4RrxqAZVcW0h8zHqr7
TwH6R5nWeo5KyGrMtKc0jvSK3xMUf/2ajHmrNur5TkXCfuaDcnZ4nfpQ1zR6MhLM+AeaJS+SDvgH
8ut42jE4WpExuxaWo8GxAlXv/IZ4n0Hrl0Nu3f6BgVpRXV1RIPaiB1KnXuXPH5vQS2xg1NW+avBY
hWBlYRd2V/HM9RIuYJ9grVKCHh2FICWXjH43Fsz/tMQpzlWDuuBHqBU7sRkCQls0/gem5+nLfPb6
fctE7zllMMFFv5UX5dlY/F8t3lGgN8XQ4BMEq5S13FpH7HnP+cIhtTvV9avLS2fUpOBv2RrszPh0
xvuyk/u7ZXvDgyXlD7xfoK42hAffRh58pQO7ndX8kgiTOQc5Cs0M2eZnFiYleCt9OvU13+Ce/fId
OPlsJOb5P+joU7maDnBKFT8ZK0MLARJa6HHNGq7+AS7nCuuPNmNFWIo7Okv6IMVMC1Fl1U4qc08O
VByt7EtR9aj1Rd774IVVpWcVe0QZrhDq8q+UU92qsqugE6VBaTt7eOfIs8pLL/FO04TIVOlCO0P8
Lzn+2yTOUSyAC67hKrDSTBbzIOpIE8WFKeF0hKayqEmvDM5kYw8atk9ThZrO5hrPdav7AZpYHTy3
6+SqI4A4irK6Nue0rqCgDNpTmfu5Nd2YE+0qR6tWBjghBtj2dtJhAHY7w1YDZx1rmzRPek/bgnuj
emR+ODb5PC5819GjT0D02UMGGq+IuIvhYlJobQBfMKffLU50JM7IOR0yKSzvVK5DX/8oUJUKK4gy
zYd1KRkLQVbPiDV3CCiKXOF2bGYrLRXc0qiMmuy6ud07WobSY7JuKnJxS2RM6pPXIp1VjnYfPUug
qmPCvhoFaqkk2LnLjfYY3Sk4p4mYZvi9i4EsDuE104kXLLaePxuyajKfhkjXC54DAbwhTPuKXvRz
2pl4BFK9NFv4Ac5PnybhyDCnjcJ+j9Os4fylbzDNZmOxPn8dgvYa8+FlXRPYUf/OD0343whElGYA
mcZwVi2G1Iyk856HlwawpdhM5qTbX8aH5wsaFGLKRXpmHjWCTUz9eU9CvoWGuDXNQbu6JnCNMQl1
B9+N5o7Ausf9R8Iq1k3H5Aeai1kDtpj5VqgIdQV+hMW+0LzEVkWkEB77ISwuvdBc802FyVd3MVnS
hpjIhWdkjPeK7WK5iD34DOsYkd7/qtogArCZ4LGiuDNA/33mr2qX8WcGHiOWQfz+2eHs+RUTI01F
s4wL2KCTiZQaIfpwla4Eo1xCKpgEMxLIx+D6OB3ujtC90AnC9ZrYzdo/uEPBzJlY2n9w4JS7O3+E
ncbHWOrYqkFCE3HdntUuNBohVUcJUxbJJzgc6OikH7PbHM/+5Au1HP6Mno8IciTARCAV0u13mnJb
2uyLK6bm2QBk+c7Q3jiIOZwOASu2Q2+iIXN8LoYSOnCHQW1EYR0LdM5xRiapfwtzrttOmEDwhLNY
sepyBId8ZM+CgePRruCzwd4uj/KdjHo02aceyzL9k3mA72YgF+b0HMDhGWVxVUNlbrmu12tq/Zbd
CUDxwks2p1YqAkVX0Fahws//EfAUTO+0wauSDOFFVPbWINLXlI18rB2aDuxSqyWjrG8PvhTDU/Kj
SK4sx67UBgd4buA+dVNaQzMi9O5BGo8uZ49uD5b5sarJeZa5X1l3ocP5S/johtEsQ4Xcar7sQx3s
FoQsyDx7o+zCrCTTbsa3IliPG+6JIs/F6AlBgMqFXpsJwDn8wqi3EMEx9PWXryaJ5wzyLprIlvrV
FBzcox0sjgG1uN4AJrwzh/wXys7cahtCntbFHtgBZlqXCs0bu+/tI7xcmL8MvutBhiDTIx01Xx/N
s5LdXdSXGQ5PNAKYNM1oHkkgZoFEzkyHnBwWM7o4wzrYcLvHcQ94IS1pmpHuPIPqmsUURTEG+TW2
4UJETRHSCTYfQV8SjHK1rStzdSguTNW2Cs5fx66CbHuV/CDOdT1mr6ZmHZ8rNTO3fShTTGc5C7iE
MBdDo0v/uL77xQryf6Gd3Byu19DEjeDrwPXWGXrmqiKhy4lO/qTx1gmzVYY9m0Y4k4GWmta317kK
060qZOXFiNHVvmbrqjaNiie3/0JgPlDKSLaTm+j7y8deWXc7qzj6LdGnL2QZCHSuMOPUDTTpdVAS
XiDaLgPlnY3YQYrrC0/sfsSAOAUCYmLLIUT2jhf69efu7WxGTv3tKabFTd1tdH8QsFwLK9IEXNN9
NZWDzMx6sJ+kJ8cFHeQumxSzSxxaHzoIMbCEVabmw63uIYFPP1XHdomr4DuECkSVwq7DtZdvD7B9
Fp7gRXTWUImLnBCXwpfTew7AN1/b/hOShCH8QlEQgRrCFZ8wuRYLqmoYoBOa7bCMtzhnLMFqvr4p
lZyNGlWGwOy6dJCQ/iBv3zv79Vo2Tl+Ib8vXowQzDnwH2FO0ZNpEtKYTjo7Tm8EhGJorz4GnVLno
QJHYoKVDUULsCUJMeZ/cbqR9fUu1bpFnx4m4kiewBN/0Z0NHF3m9d8RLV5y34m1Aty4vDwGLHgHm
EPDqjka4yBYeN5hFZ6MeUaD5jzMGu20cLu2HKAd4gs3gz3crYr+PsKBVOkqe6+sWAudSTO3XI2Nj
O1oDyJgtvgHKzGezwDBjNavE1d+14N+bOQiW2MEPNhMP7pdkWVLV12qW+/AjlnyCtpwuop9FFilk
tCOBHHyIBd+wZCkQDEK+/WuzmzvgnjMLZb8Cpr24HfEY+eCJZjn7RNijiTRvp92+quF9TetYWKHe
NNj/Ylh/+MFDdUdjVQAkE42s+fQ409lgiNztvaHotRwlUqYI1QAPCc8vM+l77vOjpYYCu3Mn5hgq
bfOh6iH7e0kaeoJoPRI0Z9P0lQ6Thg6TaXyJhRBLX7WobBjk6Owyi9KxryKehYz+18eLPCcAYWMe
TZAtZCOx3Xf+lTxXiFBdl4ebL3K7drUk1BtzUIgRZZBDCBiFMbTqnaZpAG8jz2DGW97gv1OgNT9z
1QMGtDI0VyYI0wpl8qWr+Pg4aVHhNw+u7qDrRjc52uElaWJoD5dUBioYGfpJVzemrg+FpbLpmT4C
L6iq9YIorKgXSUcYN9yj8UDQtP454TjKSxk8efPCtJUqm4Ywt18tq4me3JyzmELywBD/dE0AfxTx
uhTCXMnlPJkZstuSwmZHWzWOIx1OL7Z6z7Zz1xex8b6hh2jh7HuAWl3TWCWNwiQlFEugwOXuzCKl
fqFbQnrPPmVnneEoCAScNq41IGB0RGrE7119dUOiObUFOSanypee+U+98eQXeK+ywbX81Hha3Z8A
WrW8KJe3KSytx5iIRi7Xp9FTE0p5LC+Wh1l/PhfpqFJgeEtWU7oqILRe+96bL5iQNujlEs0JAKIq
X/LzLANMWaYtNx3PzUMitJMlJCl3zRblI+qxDKNtAOsQhCbVYQkHWiaNyMp5Xj9DtsGTJP497Mh0
GA0xPfTnNU6l30X7xFht8AfaYqKvcnA2b3m+q1j2Ifv9UDnyFjfOU3BcWMwDxPCiw5JlC8FYRI9k
g41KqTM7VRolkAI3Lk7V3/KoN1GSympvmkXI7HqMubvzOsyx+Ig3pot4kcwYdLX4gX5pl9P/Y3lx
r+w8yGlQGzsJCCdxz4Rjp7cW/oUwGkTWqn0hL6H86wT13dEdHHXDkZFNcWzypkj6BNgAEkrwMohc
CmylIDxb1rDaptG3j/D0kG523/iFYkT3LRavar5NyrQeMUp1OFMiOxVLCo0L/8+b8002HWfg39ps
JgZEQA8nbtC1bvLP7XN8YUfYKB0uJ+3zpFAgc6cobUDNEyca0+qqME+Z9s1gxjqWxSBzr0+WqoP3
YUJX1ieHRtxt/ryNpHW1dhOZvbmU1WNj4STXdXe5W5mbudXylZ96DkA95wCgBYdJ96e9TQrYVhVS
GG1SyLu/OR7CD6u9DRbtX75CcJH/rtQR4qvbwdJPSp/ndveWuTckX2yOeXR/9r4r8Ij8q60DZv1o
GUwVmaqnxEknRoyyidYAtV/i1lyIBQYJBJJdp0LCXSHAcAnm1vj8HRHUUjidybhqwCRPHgajMWOv
ti+C0hwMZm5y2FwUfx+G8sXVQAFTHXFwI6Qjqm3Jqx9MuRyjCjiPmVqOIyevmNmIgUCh6D/fZ/R2
vuGUft4dFCx8i0gJ0XJr3ar1L2scye/6EvV6Dw51OUvP7HVGs6HB7VRurRY3g9Qp0CY9mq3+PTgg
aDbXpjCYW8xFyLAhmrBokdCG3o3RsPjdC9X/3jC5e3y7mOZ48Qxa0oVJqgNCoEGFxRXIFlvpJZeT
fqFpRXaTLx6J862JNVcCJZYX6f192yPVXjjlPgDB/UolRH8n+NS6rjeo0IbAKiUWBQK2p9K1bBXS
vzYl9tWXkkE+DHP/FjK04AS5/WaN9yF378voRtK01tlLUcgKXv+/6OFeqCJ2s7bPtBxTBchfQYs2
peHCThG30+YllKW1N+B46sEs33zaTrwZDFOmeOQ5RH2pvBiA4K/vJsyvk9mG5wwNvhyIqhg6tljG
VWw5c9yIwoJr6Vy282OSPFgkZUCtBNgp3RpOOP4fcWAGgEgRIkLjddecrcu320YPfQRLv/yF+kxj
9dC991rf69qZ8JUiW8INYj3DJzDuJ6oYQeJjGEVeAyNy/oezP7/8TNyjqOb3D2tJACtfo5/fKqXn
hiHyDnABMgLE60sO09UdpxGD9YPw2kx5SJPMoXw8H+xY1/zJy20ssJQEfT74Sfc2F+UgGhVk/BXa
nH+jPTw340XEJpTjE9PUrl/BEBRxQsSbS0hgNtPcJExFFmMnZm8fwKmvnim8tM2sX4X6b4KCWf9F
ueR4tkdwlXsLI5mwWzmfxzpcu7QS1I8RCk+9Ykm0X70NRvCGKvTdSlJqa9driCmCg18K+09e9j72
uLnSa6mlaUjn4/Pe2Umo3bMx5glNPSGNVTiJi1c/x9RELBSSl8beJREgTF802nWXH21C7T+8XbEt
yzYS0ytYzjJYO73npj/RDqIOlCfbIpJvqdXMGIv/emxZgz5FCoYFdX7Lue7rrOLR6NCy8X74R8oA
yEmX7tcdBxDRreK+ISh9qnN/Swbh0wMsdOePalmExzHjjHsKRRGvj6H2aWRIqzD1FAmWhC8uhPe8
p6SS6Nz1B0iLO8EugL5IUzM8iIHW5zGuTt3VtyRfFkvpPUmXeM6obSM02+Q3JGcNGnTBBRUR0c3x
aHjw2UtyEic0ztELcLMoag6GQhtssz78ZYL11/+dOLtScNbFWwVrSJfVbDYSsq262s07VLYWWwFN
hXxwfDdCI1uQVMJ6G8D3+iy4SV7Wwqv4rExMOOmUbNYeRiTIjqXJ/UoPC4Vofqd1UuzgNBMsKwAC
Bl2i6DsZG/Y+iNu7uXYRXv+z96E7mVazMqsevALmC6udaIpO7I9nRTeShes7goOmPC8XniJYAS20
xW0gFDyaTFrifLALZVXsc5eFWxdm7Md3iViMCvRN4cJzqVKIY2JWbF+A1jXAM2n/ifeLFiGU7QaB
TxHH3Y1YV1C5EGU+CQnx0HaMRjYj1tTIEfnAcMnkI9XmEADxhQ9gRcZoM1AwGjVxF/d9OlvRc2Qq
liwioCtls89CXzME16+ZaAdUK+Izzhj3YUvVrakVNLI6eVR2QexDEXYRZiKjtDxA+hMmGp6RiDrs
3EQGwi3Z9jR6wJxto/JMPgV4iEjekCL55plzz987Zv594u7kshmiXpfBddFM2/1r7ckzNolx+xM2
4ODwZlQCPQWpN/Ntc00bB7E2SCnG8/X53hqUgUO3p3cSrAQJDnhdvM5M7h7ri/uxTBTJM/nZMxnt
W0QCfs+zZUQ/VQKMVBhfBRmW8Hfc9LTylk9arEhVQPgWR3B9f2JYe6dkVWPD+FTP0GGDkHgP0/iX
uFQW76lhFGqAum0mS6TLqeveN3sxG1jCCeWXnTrkbahdS0SelREA9Hb5qBRM6aBSZLwKp8WidMUi
hRMWLVxUPPhLxI2BfYkE5hfce6pwL/XrJCU/9O7zOnCHCHDxmIVNdSgAcjKhofois8PcavlvtmUt
0c5o4oI8MhsnujVnDunQvpDGgdWfE6km/qBSPKgiR4OHwJza/tvDsu+xkWi8IGejxW93j4SAxJW2
gRTQxUoNyqc7VgmRJKhgeQLnwP2mYB5y15q2b/mgLFbZ/atS1Th/EHCKzfHEFKtlRifq/4qIW6ny
KuTVyK9CNBg4uCdVTfXm4BvV8xYKq8erZ2GawoIy3uRUa0y1NR8Rg47fm6kNWdjuhILNs56JJ8Yo
ltebQiLxvpyGNFfUUSGJZnt+Pn0ZXQZ+Npc8KAjRNYo5GgMhCPiOJqKnfF4cJVnA68IkaYR1Z2yu
euyM0/d1k5KbUx6C05csQvx5oCQb+iA68yKJc3FlJoyyedJ0OQhDgYLdQyTTCBZRbE2NBGwfys6V
t/JTVlmHopMaD6NM9rRnlyTFacTruLop3ALxkfbHLaADNxMppwT1FfGz0yJaEZnpQy37NVaX90cX
6VhX+zE2IUQZGdGBFO4GVodDdZ5CDbhbtpo5j/nrNCqAdZleIglpEC6Wlv3VSU7gb3oeUp+AYP+r
Ma2lJLQlThSTW7zip2A/950368rVUnIBe5pxp2bc0t/ruSLIotL5hckNnM7+jQZQOY50WVhnokHf
9jGZ2xzjjxRQ61PjudqfeT/6Ll1IkEprsRk6YFvmtrXaPhzRcCtKPktKeTMXQch00uF+wlab6BCi
8No21yK26nnY1Z0G4NNvWUCJ2wtzmIygvK5PwhA+CSP3DO2LZhuKB5YaAiz2r3niYPYSH0o2Pa/S
txiJzMYT1wvUxQ1g7rKuN8Qn4k9oNxVa3Q25K/YHy8Kan2E3fratJPa2wF8UaaSEcMG9XwMNLA89
p/h6L3AtlWeMJjQbb/iXr66K33Osjoy/c34VN/Z7HLe5MS1XTngV/8gHP323erGyFzW5q3PvP3j1
3Bp2HCcubKDGNwepvjWJU87JB4LBramvobX1GrmGbGspFYsXC5I2VLWfcPRbCHXjbHLyHTLBy9OY
48yASKuUUKpsKTYRIbExfNyUk7287WpBdvVUtsYO1100k63CKLwqmI0WTK61Ew+lm0DP++uNc+RY
7us+PCweD/SWQWhA4S5701IgPDi7TZppfy5MbVdsswUuleF9oUDk9HnZpaBUrM/LT4YCXtrUq1tG
KlaFMf3DCk1sSLWPC+pddp1J2L7t8DcCq7FGBfBuuyvuRkZT8XXLS9UaVKZ0NRwWYyRctW2fVD8t
VN3vaW53VuJhTcvjYXik/mEPS/L6BqkiTz8KAb9Ze02MVfJ6fXcs6QUfylWyBexpr2okwDmouAdc
otmwMaeBNrO0aThMiqZX9B6JQqDCE14nQ+9hK0W6/9MDeX1dnj6TvMk2VJt91SSd/D45G+ergshJ
wHgytt293w/hMxRFw7vXuVZ3KbRUaMxArIDtMOqxmF2InjaqLBXlEd5RKTVxJwUkd/36Er3q7h6B
0A7YIdjCtroCzL/50MulJ/LKOofMxOZftJxJ3IMGXFBV1WJ1YjedBi+yDhN14495s4Zq6kB6GqRt
NdKPlB62A/tR9HLaHISm19sx2tEzuDt8W8fOwyE1QOjLKzX2clW20isyrh05stIE89vW9Hhv2/se
14/dILSy2oNLQuDzmgMp6qzimG9HE6fzIGv00wAQ4th21EwdMfQDclT9Pj3vZdtdBpIUJ922OJwp
PWcgGTDbaeg7cjcI1hZ3zK1yHT4uFyWROchvp2ZP0eZA6SDPFMEdueqYyiVv/pzkR3N21p7yOVu+
6WaG/g02D2NMkTrqplvQ8206sK9iomITZmcTSN2h7LaGyLibtx/JAchJ+J0fmuajw+zRXJSPMKdl
J8m5mS5tX8P6WXQMdFlB5A+D6EP1TY+PmDMvTdbAMsFEI7HhJVvHtJjDzuagUBr6PvUA36w7de9j
gQyiHZJkm24vIiehlNOw1Z0dAwzgoQQ0NJps+P7Bew3Wfk8Bkp45OmwNT5D+bXaNL18R8MnPQ49b
hDO0RTZ+gSoTaKAh1vh+KgDNJeZaQZ7elEs/m9OgxwJKPbish9kKGoRq1MAQZAPtnhIPU6SgBb3U
HtSAbKJcyC/Pig5N3yROvGvTAG7bdG0k4jVxhTamXN3X8j8Ue1TIVtHpX9iUtVl7A+9HAeiv+8B9
AZGaHvAHjOMDZGSF4KIDEW1P0GSnyCsTUI+s6JdSGEGO7p6raW2LOAVaSjixe5mMNPYMBN7dHi3u
E5w3PYVnMSLHNTb3eik30QZ9ifkwxFYw6Nnvf0wIkS/fX/bFBdJaJXQeE8aKg4jTUbyIbyHJdp6R
WDXS6N1cGSa8k3HZcX64hGzPsfrrJ5P2+YU20m8jAQs12ooKw3x2gUDRAcb0aqAm3uP7qs5U0nyt
woy/1t1WFmiSmYPVEmQGBMldO2x47tpaqxbPyLJsqsAyMZe6Yy5goJH82ksc1ChsCl83acgflV5U
8G0xjYusGTuCo9GS3YUNfrZXEuvnw/ZudAfSryWdXI0IM7sYRKvzSVrQq4F+A+xpmLf7hCvkdyZ5
ehdIS7W5GP5dyiZvoEG9ZEbvGePbh9QKYdHJiyTEqX6pSxHgdKDa1ztlJXUWOM1nna5iz3XYv6+F
EWCCnfJUaIOhXAQWr6qoQXM4wASKh6ULKXoUGygO1HADHX6ZtjOiZ2ootfkenIfM8LQoki9JFUNn
Jh1lgFBmdxX5WITxzTVRwl+KxZpIqlDhTECuG9BDiEq1Tk2VqFx9zUhJS24ddKclSsCm5MpNslXI
U0+rLHuPpm9KzHq3eAA6clRx85Rrz0EPeFhEiE8cUiP1hlF3DQWbp7ejUgX/cbY5BkqWfjo2/4o5
PGePdEmm7YOvXVNMXyO0mVFwaMuwcSaEOOSjRamBMDzFohxZj9cLNMyNE5Yjv8db1jEAelnN9gp6
V72kyopm7/akbh5M4o0nla8aOqSK78Pv/3usha04PRwmenx39vMxdJpnRA82KyJlKF9g0hLBxgHO
ZNsz7Gw8lYw3xNP+FcMJxE+kR+19ShSSfZIZMOSnM9Ws6v7t+Xy3Jk5mCL9P/a275kjXE3rKYTRP
FNNf9nJh1+ctAx+ojqhnHLjHpbaJkrb7aFwA/eBxy14DEXVVnWzeGudIuKHzOgxy+LX5fyO+xQ5n
SUKotGP+6SNy6qi1Yct0vQGf5faB6kaW/7akHPV7KLwxcjtb0EKsojOlCD3anbAcSgX/m1v9CMxw
q9T7q8MaJXZB8cmEwVqbPdZCevPphntvuco2h9EuuBXEAnm9TPLY3UJlyZ5RLcnf4EU3THIFXYMI
Es6TDx72+8iTDo2LITlipp7UiFX2BSl/aJHapUspBr9fbMwC9gIPYfSOk0yDcSAgwfIXoIjREeQi
gKa8w52L2SPh1PFHBiQq+wI3juPK20LDsnn1VG/0n+OryoTvH7nXV6Isd9713/tbM6lcLlByQJCL
+4rGJLsdPGXyHeS9pVmr8VsZ5mfkfvwYb06vRsBdZ4lzPI0qYKoOiRTTQFnp0qH4LiizQFXWlUGk
jFKlI2ZqZQiun+dat4E9su1JU5lpEDPSadQGTLQBGWFpvBdnLV3C3GE8jAMMUSbUd6yyXI3LI6ol
arkFimbV11YgFVGwnxRWj+lHPYffyQ0rwzBVOR+bDnHUZvrpY9Ujf86y/2scbk16vkfrocmJ8utR
+3jq3ocnS4FSRD31iMZGrVmYd0Rni+fdY+CGFkopSym9ye2tQTOzt9hgM8NY7LNgxiWcEdapWD6t
VGU1M5OV/81yZ2FZZGu3hPNKjxTabyA5TH+Ouy1qQejGFK443pdAHvThloOjV57vYi0RU8p7SXZR
ANaLK6RcdEe036ozKByZPE1vFouIATiT+XdrOmknJORc85ne3gu6YYRkoy1/VT2oebXpMtIyhGEU
yJ/gLX/VZMufKtVlicTUeI/G3vH0cdDE8diU1m1evplVfol/QUEVrUEHpEa9llCXBPf9e2Xra0X2
I0JDoXr4kSVRCn9zpzUCMhdlCkho6LIus0nu3TQtBsa+T3rzjyEibXOUHuGXdkR3VnmJAXtAKAoe
42pQAQUeSbJaW+MwdR6GpruVP8RNxWOLV23XUAIt2RaO/BnvU18LHLOIgPCXZezztxqw66gcOdWO
BX5jn94V9pp08Zy43VYcfW53qsVp7SNBn9DiVavUg0hwZDY/NW9TM9CZLs70o3KJAPfJVNHaJwxd
oVmb3tdiJ5GLcp5HB6fIIOTY8jmRwZhKBb4sd2EhiEd7hl9y00xdz1dxBd3dfM/mfly0TJOI+ZQo
RkAy747wneT5YHTvT1HgZyaD2VuNj0CM+Cxk9jgG7gCMfEjUXmkpaqUpIuK6WBbO7j/AJabOI1LV
0qobxkiLmtOKFWw1unfvnpF2CumReHtkUXreP96Orgs/8vKdVBEMB2ohknZ6UAWtXIFXSdGuoHpy
+YGrHxPiW9+Di+SK+0s6yQ9YggWvnnSE8FSYpVC/GvaoTvyJMiODhBJfsx1xMiL4Sj/DzxE29d4H
Zuo88lpjDBxSSI3RRh218wKGKDSExVcAb+H1KtU51nncmGEC8zVgna1oCkn96vbvtk2JFcIticfq
5nL5FEC18fIy3YMERTRNFimhfLgjRsQNVJzyekEGuZwDVDtjU2kYUAUO+MYZbURtIycaXYGoWGsk
VgxBewxoaBNGvOBqPHXy7CCays+YiMQU9p/otOvmdvBVxYnJi7xv5KXKPp2kPtCh+cVQutGdq/Na
89DoEfAPiS0J8JahrEf/4LsR++KIidzhkKaE8gxlL6T83EBkGlZv6fCmlKyZ9PuUrjRcz6KiRgK/
w7155GU5yygmEx6ZtqnhpjB1LwXQLLM6GWoV1ocTW9bsz1gyaEMWGtv6Zu6/jItYPYPbxtl22lMk
/6jBkCy/6GtooNqbKYgcuE2Tiab9jyOUS8lyOA45Hif90zIWfN3qJrFhH2dHs1+WnqoenLamyFdw
TYpGaCyIJlT/MLHrPe0HYyOQz6w7OBfRgWoCcX5G5+SzIhu3qr/F3r+McfrFS7LYSRZI8etPbxBL
KOpo/reZzeP8eRj7DyGADXlJ1mkcNqXF8XfEDILz9vo/p+4EwSACcARuWn79X3vEVqSniPlPpTQp
r9kKn0i2Jy6oAnc0gZD7Q/sWYgP1pUjt7GRtcXMGW9XmF7wwelxG3ufeATiRGJhf24HvlFcFLYIu
d4L5umbUvJGHwzaxD8h9AdnhRG2d+128/rHHK6B9vCOXM7r5qGexRbeqSzMoOWFa8/KqbDy6TwyW
uPjCsmt7yA92lNuH6eM4JtVkRpmCX+OLUCWeKN7mkYwgiYJMefbJcG+cWirr0YLu2yZRQwTY7FZl
oBYaj2Cl6NCO5tL7awQyVwaIm9Q4F2n9qp134kuPfZE+XUtCFitl8MmSLl4oZ+SfnBc5LPtBhmgJ
X0KoNBCNzTq8IxjWkOev9HQxSuZmlo3zUR2PON10i6fEt94P0w8UM5hd878naCd+hfNK/2rrh4bd
Hc1hbWqyZbSYL1TaIJi91sbFA7fLI37H2grr9UdbCWOQzgwH4lEyH2vmIPkqLh1SAiXscy1WfFDO
vguHFfYArL6LV26KENBE1De530hPhsmTz9A/pvFSknAG1XhLPOBKR/TiMwl+aQV4T8hWQwELxTo6
rxUmg8aYCsu48goT5o3QfGIYov0nEwRDpFeubNW2i3KhgpqxvDARTso5A4/BNB5d2hSs+ehFYkEi
k3rHv07xnL1nlK7cbmpDeKpKrzQY3ns164Udy1WPsuiKZft9ilt9kB7zGLbX8HFq85LLMcTXXWVJ
zHt0dTQYsQVxDJoVcYJrwiL1/veGJzzToXKtqncxxz7MqqxWKIyZby9Q5cMVtQnG61X6umWNR4Zn
patUuTSgU0M80Tcht0N2inmm2nd764EAwe+Dn8On+Bbul9qLdnJbR1jlWptjMts70JsZKNjcEJj+
mMpYoyBwPnvJ2vCkazRUYf6bkF3RcBhNbTupXuXvy3C7haoDbZyvIhWkE2Xz6VZuQLDWGhO01RVO
thVv+5+N5qKj1Sq61BH2eYxBEqdUrmh5UO/GrkFRBZWpKqiL+3odp6YNsb2MT2bpMC6fgXKHqCH8
gppyCmK7MNgCqSBVSUb+fFP51ZNmvHon3QHGqJRzWHqhw7ApsalwHYSIUvqbDJgpau5gHUXkB/Cb
0CeaxtP4bIv0jAu+NOJKTNeCqGQQcg82H0ru3n8Q3ecHGT1wNpz7Slod4jdz0cn0G6ftes7Td8UP
6po+tBj+8XBtIhN8Y4T+Wh3F+eLYFHmB8fQVBAEqa/0D3xV/yro7NKMv6enClL+Ax95YOJ3LsgjZ
DUkxB1qaPI9Lo1UJKG08NF+ewEupbuGbrRXuAq4lNM83xG02/toXaEfziclhgaG43FuS9E8ySCbj
TtqlM8oqt4GWVOHKWDTA1qURarsdWFCwk3EKhl7YJ0Z9vAgnP38JOnxIKJd7PSIBGl0miJfhUgLg
Vp80bBJwWz6rhCXPpu82evkwktZ2UN5TE8uX667nnNVYUMuDIZQltISK5qPo6P+r+qJEHAkFdo06
WAyZ0QhwDF8n8b/73n4Ms+HYQUN5Thp2geAXoCErL4z+oxIutem6IUZyI/YulkFj3RfmoBWzpy24
qa32EX0H+V8eZNMP8uoCShRy4LCx1/toM/i0nEPiwwp/7j6o2BonX6gr7SDx8Hy9y1b6Zx0gKWUX
dpTaKDKn2tTaNq6p1JDavNZh1+WkF1QepSdkLH/1dkBzwq2OhOE058XESCEFhKnHgH21EcyV0VvP
6xPkRZeyBLN5aDweD1os8KZpSlwYg/38Gh/ZuSpX2/IkLDPDl7vkW38V5ujJGIPfrLe/8nvonCg1
ms87Fobj7pWT23+Am0Fa0ZFikbwrSogGY6JDk+U4NKA+IgVI8bXYI6B3oUeNAWjvef5efZAJW93I
ObluXbzLALft+Nle0J6zFNlWci/eVbimjIxJoC5xNr9fvWWbBCWpG/arNVyGG/dL07SvRwCswAmO
aSPOkiVBI34v1BfpyUSUO0eOHGn55WAoUc7PULcDnCdaOelDYuNjY4h1ATSbSrPmF+XHI3uQJ93a
zq6atJQL4neAZe6ngGSLLPWWE6AxjT/DCCkbhBRDWhioIksRK4l32pKV9LtwqPnULddp0QcUz0Dl
KLx1klju4WuKM1vu4x0TzHha2nUNha4vxINqvI8cfcKaBuctAtUMZlDozuZmPunGJXqxmw69xgKH
zyNtIZoaJfNivMtAQ5keMgp/s7ZKVIa1jluRCrh6OzOOwlzr2MATYSgH0MNeRkJXhZbqPxADsbbW
Z644lzfckCTaV13oQf6B6FmPiUtDZVAGNxV5RoxWJPnnr4XM6bIWhtRMBa98qgZ70zxGdgmt3YPT
D1Ggwy3s9g5Mi4iN+FBafUeE+5cfauGdMx+SwvSl9veWlba2kxHsyNpzQkarTUMHxxzs8KQySkrN
QxdKJEczCFGqKc3dpV2zKHXVZPDxNuUOWSKIJ2uBsEbLOclaAYTgbw8QYqLotBy6Ccmviz2UmOAk
VaGWg3pgeVryavIKTf5fW9+kukwtLNmqZgm4m/0axTN+ikVh1AaJ6jM4RBEicI8H7An4EEBWpKcg
Od65fSEkJYTnq6LwarU4jMkFCWm74JxDJhI6AYseiPivjzM1Jdk5CXL1iPXXXAIpcJo1baaR8Dke
lVst6xnxEMiUpucBWOpFxibI2GBKouquPaOaIKC5A/1N5GzStJ4+dveRe6pg6VF2rj+/004MRWdn
IJEyl31xRKbCDF/et4ADgFo/lKDqt+WqBYyjXexTSxQCCIJmfedUOIndXvuQMGci4QB+Chg/XANa
yq19ykc3MvpLbBxDQtRvBbLzzxQ4foVfXmsGe5UABuPLkwkHu4ad+q0oGbyY0cr0vqIAw/dk9tOB
Tg02saeAHLg3ykqhWEZRhg/zUFv8HHXIseE7LVOb4Zunv3rC+NT/E/ZkaWUEoD7lDHGoL0wEWdyI
cMqsyLZOCMEtG5EFWsueEeGKr31wGlcwkZBs5uKGFY2rb9IFTEiO8BcorME1Ocag+S7kK40jqZrZ
axyhcMEWCtfmJ7Y563J5Q5ilNVU3BshJRPnHU5G0L0mSuYL2imOYtRwpAO0BuUiBYiRZF72YMhLY
HIcER5oPGd9kCmtPJTmUvzrdpYiBaB4vpFBNVflrrgaT6TVk9JjUrr6Xo3w5U9ecjRN7p1fRPvvL
IbVXJj+Y+BAxj8J54ZGvy+Tx+edzKzeDKo45O9BmOuvYenD5lNZdyYLdw9sOkw5SEV6fgjv/UTVC
GsI5owNZPWVMYu9wnRYrrLjPwA5pDwVDZXWumk7CHDWvPmVCBIPp9ch5Ax0s9cc3BTnokyAXb61Q
QT/KnKDX68ajZUAj+Moxd+BKlwi2ox79qFdU9lBUc84B5gUJCrqYF1hlzxp3SiPWvmPX4ytQ7ehn
nS/C9onxn7YOatDU4havHQ/oEEyaskGthGR+wnwn/NlnT8x6cpD3HTei09Ge90Fb//IA66hCHmKo
f6Oa+mg5bwQ+fHkzk+cEE+JAuHPBhgcJC7Cq2HwmGSYPbv4NUXUPg9a+uAnvA9e9S1fsml3/kW/Q
xziARM0tk9OwKvOhXkFcbU/ODcpnNvYzfqKGfG9tlN+oaLdVpYKsVjoeJjDJYI5q33Qc+g5lWoAJ
uefvJ/QqGY3riAzQiyRS7bG1vY3pRd1CLYXw456coOh5LLC9SQEhKM953xz0kMNfCwGbAUuPm3i3
szyvGIVWEYcjKpfJsZ4LEcOWPXMrfzip7i7c56jdB1iRRnMoSfeJt2QKnjvF5jsCyXjbYIb3Lh/8
jzzP2gRItMxQZ4yCyhRKA8lP7NX13V/cIsfOQy/+g7lpz2AulVqjzE7DhvCi5WOPY0HWPHepF7KQ
/4S8bx4Mo2upvDfUf3zf+leWNapTsjWPbABZ5QafZEGW7UIFNFbOF6uj1S3GgUX/pRRsjJRInQTY
BCAQTPF/qUyuFdqP5rkJ+3L5/H1z7NFnAfltX3+fyQbrH4JOPmFFVsrN8livqqROoZXMvNloeX3w
pjhwfJ/dnLc+Mbrl70QuZZMSbcyM90oWCnLbTTmIl08Mgz9tvi17h2x5HAdoeKR85QgENkUwzEky
MQuole/6AkSZJA9lx1u2NSb6p4e7/pvKs6zmPudr55vohBYmm0QSvRoNd+daB63Cb37qZT+Y79+X
OMdi5OnvsN1JtzwU30KyScBEMzBdqwPwAhnpdXlI0/Qi2sa2lSmpe9CXWcEmUxNGuYL3vAdDLQ/D
ErIKljv+md++tb6HdmmD5ZO/sSJLjPjSr6op/oJbiue4y8GfcUHb+MMjKzqk5hG3/mGI+exKxVhz
SuMJf5nrHwf43YCa9S4cPq1MbdNd8UyLk/OFmaanGYQ1DRs8rOscBQklFAdldSzTROUeQQMglU11
uk50sA8IETd2S4ck1oNK473pf77Myrp3NHRKsqGYItdzw5oltXvlWiAAPkbEX4al0JMKPN+rJJTF
rMRb++/V9S41VekAeZ7biB2yUiz5lL7tAr5uAJ4F4y1DrV6m5i115t2bKTtuOLtLwV5/poLWlcKQ
Nsm4UXxwhRaBXPEgPHT/9dIhqYcTp0NbGvua2JDz5/sUkY7NdsQU0ZUZvJd03x+zdo5WfkPuO04v
PJ8UDsSgZOhxQEU/SUEuZMVqN5gN1OU2LAVPzzz/fjMc8DuxhZ9UFJ/l7KVTI78sUv58ycUto6lS
dupav6n7SGbO3xrcGqqwi3SF74FpZ1V4LXaFxvm++bCU34FRaffAgW7zKFk+I2DbyNhltu8k8HCI
XMW0+SEz8Kwz0ioyYamhQwhtWxhuYHagNrwuOKJsyPcO7uUuoe2G6kr2bSFelIiOJtWa30qA/6Gx
bKnUOBsa58+NG5ohTCQJTtMh1BQkPI9l8BcJNv0oVDeoB9Q0xge0aFjW7bQkW7zwxnDVvNfMblOI
Vp/3zmYqO4XiGXakRhHFwnKXTdaiV+lTIf1ZZ5jfKoV19JiUMF+nyr5xcjx4e6yY59qn2ROgO+ng
BWGQbycdAxOEwoWLEWSp9eZBNEkmi7Btfd0G6E7gxn4EQYz6lGdLofsNOs/f+ZIQJBDf0g/TmrhS
hR666Pj5r/6Vc8HwIw7EMIwg3Vx+wyoDsSMlJUS21yRkVu1OZVubuheOHMlzOP/ddlhPIICYvM0g
43ANlC9YAP8DM2zRr7QCfrIbcT220EQElJHqP2qtT0Ovinx1YGqmFTQCfonJmz8D4weob/tX5IFv
yR3PPAAnLwA9j4URjEpnFFpTS1HX06QVlvaGi1ytuqX54ywPVlW4At0eaJL0hvAY3ECkj9B9q5bd
eODg8zYCkUImyEvBafmN0vG6AkmQ9CXXl8LaGRC0WO6QGwnBtxFHg6BWz8wHK92w7YwQYY1h/C6i
QeBLPr4+ZjblkelhZz7PVm4VCoxaVy1VGac6Xwb+2zwQsNPKAIW/TmcF925YtAcgWw0W2aXj++w7
mEOx0Bf63tUJVEyTjHQYv8SiG0RPpSpRMLj4/c0i5sPzrXuuUnf/6daFaUvUrRq+PCJn1oDOKZJ8
bL0yFkYqdLfVtBNLSEfsPR5XmH/l9Yi38ipmXFJ7ltJWta/mqUKefbj9sfsJmScQiLDXpXYF8pY0
bJU6QpONDYmvNXOf3L7bsiObwGbIsJp2okXuPqikmtGHGt3M7DNdDT7e4fEFkkZOLVPZsLK2bu4K
QjgynTHOi/hya4krAg6koL2OZhoC1Rr/W7+V1wTB9AXgbSl/JjYyYu5INTeTIM9Cz8Ze0nVzS0Uz
P8H0Jweg6g8PW22dZbbyUw84Mk8OPZmktaLf3LeRzJl4Ehat3R629FRxE+UeWc/rrQZqYat/VYnF
4Lp+ep0/XK7TT/NF13WOD6QF+P9dkFkp06bzInNKtLYJlZsLpfdWuErrlGhxa1R7aALBrL49a7ka
7DO5Wi9aCjsnB+EFkuMtMN/yZA+X1tkq9qJSEIV69Ja7dlVoecfz0nz1FvunVPuN+Wh5Vp2hWJpy
4kXCmmvweMnhLoz+Jq6/PaTCrOVi/6OjvujZwv3xEPAghn635bejYyc3BKEz1wPep5Fg4NoavBUh
0LILG5HBe7DkO1fOoi2BJxutRcAi4JKiEbxt1fKpEZbfjYmHLuMBPPgV1VrUK0u2jYot96ZVwyv+
EpIQ54uZ6RjHjbEo3oXFR5VOCvMK60xmVDv2H+HXryfrIBQyz+6B5kXnrp+pAaVO/9wbdsWpwABY
q2lOxFrpSipzsC1wVK7Jirgpy3nLRGmtt8uJSvjzTPpR1yzpkeSYPluCw9qy42PSQcP+DZHEsS+0
bKUUJEtK30TosZXeSHLVIOTCM9j3FBRkNenmQteBRGjW9sQlgVzYT0OCb9MaN6/8mAWPZamUhKg3
sx6bHjTVU58Lp+MJsPUP5GLR1FlfMCIzRnJ3GA5NiWLThfeKqrVgHi8Ewybwu73LQFfoZjoeDvRa
85QEPNBrE9UBn787jC/A3s9by22fZqtynJ6dgT3ssplV8UIAad3/HU/aS+v8EaKDszn6orLBnLhv
b0VxfNzpXpJ/scDNoFCZzKHs6NygV5wBwMucIJliZvH0W69RvbVS4T8Nef6xWi7K7jYA+kDJUnoo
l5hngFnl6aP1dhLeYuhCFtPVU3octzKpZ3oHPGqLgd+q1t+Bn8mCbM9cMs2Z7insCS4YOky7OIhs
pDSBuZ9bQdfw/GJHDNJqfT4zMO5fXAyLigImzUy1pQbUp4vo87gOrdIMC+6NvyDOvOFzqLAdn2U/
OpNCKNXNacQaOuOSpQwbOX0XkYbnD/NAphr5frDxEupQnZGPPDtqXiW2nKKMTbNLU3+T0swCw5rM
vSGK6VaMxvHPus7dVjgka7prYSOEXHxwNVMElyYzXduVHzPP+XE4wx/9f8astxlLBwNznvFcymTN
SgVYPG32C6YF3gna8TqQxHzptTdatDQIPfVbAoykhQLr+dUL4zE1WFRD6C2FjpwxyERkeNKsSiuU
hYRAvNn7khe085pOcYG6v+hWOyxnAM5+jcUJKwAhREa0pWUZbzwyG9676VwuJmNoZB2RA44+4A5+
rqWzTRVop0MByQUy7+qyPO7Kja9HhrY/e121wNvOhKhJ6IlJ6F7oKY14oTuxrgWWFduwtsBXhgQc
jwNZ+cwtbQlvvh2d8M9zel4yvXKmqeYshXoo5Xo8phfEAXNugz/1xbVibF1NK1xDf/DTf88igYA8
cjrwlq7dzzNzrV2yWAAqQSRijhDFDeJbmJk/xZb+3pfW1pYxseBptBQkOZ6USVpW4gPM+tK68R8b
Htt82kVsjQIvSQmRWnqxbd/+d1AADuW9h6BxzgGSEJXKjA+V3RKKDerr/NiwtbF5ELeuUOdu8cbs
Pfu4HkgTMY9r5zGgxPJTB2eyiepSJRMxPY2j+xqGXhRyMFWXbZ/WeIJXSnIpD6gIZ+G3rw3dNeDO
c1ji5TiHv59LNuHgQywFyv843M6OTQ9tiumo9OgMNf8+ebCsShxCXCtOuyWFzCWXY8+P2z2rzGCD
9TlBn20Bc6d/9sCiDeEZBHXei+Pza5CTccy2Y6dgAnP45kphMkJgz/2bjHOJ8KfRFpNYkV/yqnZE
iedMw3e0U/bHR+fwOHolNL7iN6HYSj6/0/BXfP/ZA4u/EzmOuGHzlLcsFH08SAi1Khu7N91AyJCL
P/rPxtpZDBxyI/73NWwhmpyRQkY2dDNhjR2siBpOkNJz81+vixTYagoCz3tu9pXryDBrRYY5jpMO
ErBKxFCsEwKc8rjOs0sx9DP3DtxNZ9QFH1BaMVRFHzs33p7wP9+6BKUOMbCI5bgbAxOFg0bT+JzL
w05RWHgK7qbeEszbgWgRiekhaXn7zj10I056yLoLj94ChKBER+ITg+hQIopOsi6DEA2LShPzuUIK
eL84q/PdCj3c02M6V01GvgdgaQq/xLEmT70WFK/irmAPxxXiKUc+oxwdUtSN0TxSDn2pzXiQEqRk
ymoyYN4tsl5nyxSO/H5Cx6jNdcqdn7Av6rVM2VnuaASXGl+SHRqxKMiQWI1xcocgWsYhJKtNj2qq
fblLX+VEdVndjDr/cqYK9ote6epxIJ8nPo1H65frND1FfuPa6pX61FXABVyTYXCocP4W8IhaHAID
Vz4AopzcWnsXuCgqhxd7wKaztkr4VfznassK0XxlbScwkV2qnYvoBeg9ht262dpdcZDnytYgBtgt
A5tkAt2Atn4J1bHt22bFlHqNB6qzH/UX4+L95hT6y/67ZQBIw3hVuBNBjKcEawVsetbcI2oB4Zez
EVBrj9UlOpJFJTpPHVSM1/APwjEPAY3ZFNcD2FlnpuobdepiMEqB/BYJcx7QcFBvm7qPsMhJNCSw
fHs0ABp0qmKNy2/ktLJYv9Yu2zMnfW2Ayg6J0vO0+uWOl3l+AUlyOOtaIIvMm//4SifKIj+J6Q3u
oY+6JusrsaOlEkfApovIMuEqqtyToXYshtOyo0J1tN8fBHRYh2eB4w0U9/PH4cPMVy1u6L/a1EuN
fZSAjz4nPFU1WYnNfI5UDo/AzLxH5xcUPuPwow9cqVs0uCFwNBS7xTLY7mpwj4XFE52U/fUg+gr+
bZZ6HE8liA6jWvjvcraK6ynYVW+qyJDC4c+66yau9+dNj2YNBrG+neyvQ6KPPF5Nuapg+fpDGAcD
ODrpUmBmQxJotaw0pFfixyEIOvav11PymiKeTx2law5LBDA7LRnSyccHfSKete1W16n9Yc4FLkmD
eYQzAyjyJw+vWKc/o4pSJGLOMu+ifPXiU7tY3lhdgEJYdPdMSC45zVEOFOSfXQ7yi77lsVKegf3E
+tINGH6+LQKoKFHP04UWr/XspRqqNwEs5H8MlgBp72zSTR7ZHQ4+zdHTCWmMjAJGK8A8ST0pmgsk
I4FgcXZnGGu5lv37qMlmuxeMLfp1OoPf51u1ACklTwq/V2qUc4gAykC0zTFXjnLlxstqMWsjGiJN
ZHcEhhDbQ3frFrDLSw5IHYWGW1+UI0fIOV6I5c7iUD20ELnAaHBa+fl98uimz82sfmEv9K3Fwcdp
CSOohcGVP5yf00hLJMOz+htwRrApNjM6WY2hQthsFoOR5XgntYh3guMW2yoy2qaedq5DHu0Oi3bB
1vbSmqVP1CIR+jT+VLYdqHP/FkufjuVTJl1TnkpUufKTUkMvtLVc80dPjwroSxKbezKqek4jy5Ys
SGmuuz6VhxW1aO2Rauir0sZJ9ePzovOmMznDEm6NeEYZLGtItcT/1mI7pmFb6FLjuERyqEM+jim2
Ypo/XEYNtoR7n8AMjzZZtqWCEgBT3S93Cj7PMeDqwMTSfp4Vd+YZKNUXNuy0uqEDNhyPDSTj/BR3
ZmOQhNXu5d0ElX/WQAT7ZzTpYBPOS0RUXCF34FExnFmB0RMnhsPq434ZtvQCQePX8l+H3/VGEQLJ
OI7ipHQ1oEXKgFo1uT5opKpSp8/oCedLC6CFrB9pSmHn6gdEZ6rFkMEtcw6PgxwjLg/LujytwxUq
Dy+g5C1kaDaDPEaT7hS+Hvlb6NyQN8f11A4ZSVK1aV+qry43McpMGIg2koaKDNHA1z4j0T1+/9cr
Dk4JSpyZiJ5cpKpDAwsaTJyj99nQraoD4LOMv5XYhqiHN47ImEigfDeJuXlLFqKcWzPyfL2OD/vv
SLvfq/IWpQcw34weQ2oaVUMLkHlz3xfvQzzFpdQsJV8gD4XSo3NN/aReUs4fK3XvuJa3vhQTqjfe
VeKDdO+LljpD/VWyBThDHUv5T2YAbnEHvmq5YXJc4j/hqFVwiyDDuPlsab0g3YaNQbVm6LfYB7vn
R1k8weflJng999T/76LFItQ+zMrr68J5xlasveJekFFns9mNrSel+byE29piHbiCkeZt5xa+2INA
MgNxQEwyImfN6ggRht88GZKUEKN48JHJDL+YewCoDaf8I0dt4ZFa9qLPvBMpVtR9DZ//osb/CXhy
nMre/w2yzCsXMLZOBiWiSX1w5F4J+mbFLSGvp9LCqPxxeC5Y5/CcRgyi0646DOS8DWEGA2/1vuM+
GZ5qp5VaFURjpIZXI+Y2tJMl4UZs0UNJq1+XwYfKyi9eLFK2X0r1OoFxluTn2uvd0+e58sTgopoV
qapZQ29Zckt/ak0HgfICJdQo1RPqS8K9C1uueytV8bi7+LXA8YAj6y4l8AE3PhI9WztHubEaTP5v
eH4cC6CQ96o+jqGKCx/VQmt/BtRkKnAtP8NzuJmqlHxX/EJUjUyyXEI+QUcqgdkhdfOPSbVCnEss
BlC2L5G9QNOFs1ZWgsTfU6XiXVUNcmlvnFbWWCp7AlLf4FRk4xFJbhFgmLDLbAgNRWsA2oq3zXI/
Z35UExCitZLbGTBiDmwQnMgUhaoK9e5yfR2/NiZ9Rj+SMg7OPp+k3fuhbxnlEnLxO5Ahgo8npOfv
+/XELSMZg4jml1bbTJPiOC8H1EYbVtJNlX70ilbcPn/uQ8XOHN3pBq2nJrZa3iuJP/G9r0EXs8MO
/opqH318khLrG2I4AHRmmIYYWNZTMknZg6Q+iO3GeTvQMuZ/IFVSB/d7gPlua11xjsiM1MDSLmQ5
pqh2eTTOpsaYB1nLhTVbCQDn8Xk/oEuAdZYr+lehSnrvbekDhFlnNPWmWAvkimd0HtI+mzCLqvdz
crAnoH3eSbEV7yErMKHFbSqbVQiNeWKjLjnP/J8WPiUAoF+mR6duKJ32la30EtJbqksBS5vm2mR0
9k4AhzU50oo92Ol/6lu886y4R9fn/tk80Pv4f1UnAFKYScfL1iam41yLjnfuH6SETVTB4N/A4Rx4
kAiKczSSvdazpMYWlwGWKyY6AfB4mDu1bJBCrqx7eJN0de7wEgvJ5zRhF5Jz35YI2OrpLBjvAReS
1xMiEGSsLqGeOpK94ncF7Nx4ftJh4fCoYDQkB/Kb6A9J6MRfA6erFqxzAjEPHXrHfxZ7T2d8aDjZ
+cuDMB9WmXlB90DAKU1eEOODJwp+fPyBfZivuj/jV5uEAb5ejGaN21ey+35SaUDoZsgIFx7F1zdt
rrvMmk3IrI5QK8o7QvWV+wYIj8PE65cIf6ac0U8GWhT0k7XLwUCj71EzB1GSISMwmszVPdHINDB9
dglNXqxGyXyyIC/dlXstuxwNr1BOYnoGpbg4fUiWkh9Cgk9bwl8em6k4YRXYGAO8D6jSwBcxBECH
SutnxXdPtqEJCvNby4XAKzGc/qAlz8unlbJEyl+go1iMF6nAiIgddOL/TydAzZ0rO3/gOPAjQXL0
RXJInIZKxVWlaedSZ8u1f64Zz2qekod5zgrOM8I3apfTcvCwEm6Z0N7m5UCzBrLMey7t8ZpVMwAp
FUJ/aax13mgV5E0NLSR48Z2D+Y6LWVji8B7bQ1K4riMjpPhMycOvj1ifE30mW5GykPSR+SnJXYXa
jKYA9jvcZMRV0ghZ/Kidy/6uvFhyw1OjpKWYgE5i0wkxH632r9lAIf6AYzHp3ExBny5tovHUpfsV
ZF/WZzuAfBXQUM0kuptXWDT1dMJZON22QahYlwZAEeQ8yPQsIGRmDYmTzIyngTfmatqFDbks9mRe
q+GtOcKlwzoWkYPRpHco95fgKEPCq17ckl9lrLpuxO/j/q6W9/9r+ax1+1LTkMsHjGCdeRJ2TVsB
JjFsKEpJuGkscqa4Rg3x24QMOW0Lx4BXYGy58dMFXCQJcP4+NKyNEk1td9jXNbgbEIVdb5EXJjqP
k/2AB337nlwz9+NEyb0eOHZ0FnBtANoE1Ylap9IVGsoHfZ33JZzzcWnp/vxhhFnfTqcX5geA2vm1
FTdvTaiOFJSNEligmzyo3TrHrs7cS3Bwbxkly7UGnrFoHiUH64APmJsooKmRJorB+IyLmhaR5EvW
07cwO2++IJ6c/85A74vKyYsY1CeZ69AfnqDc3niurWw8EaPtRr8NJdrpxJebD3WixOI2HvfkyvLu
cTmB8gVeWknFHWHqUeADhvTgNbw5l9rx18Oo/djLulaKJXAAL7tAuXhG43/ttBEO9D1CnUTszp6d
Ewct9y4q/7599jzbVfbiubaLqCsa9fGPYc3rQGfh4GS29hYzz3bmNhcre97gh6Sehx94KdYiXtmM
z+vknYtniqLBqScqQQoYswTHjFXwPDsAMceG7aLSzAroSaQMoHDmcvVipBVhpOOVpdXPIgPknk1b
TlKTsxk+jWlL9A9UaD4XKT26UdwSL2dBVD7BKTQT0EBlhwGVn8Jdnc4pWH5nzXqUg4Z8DB1oM57S
lqNMqtn/FIO0838JGw3+PSwZyzIQzvmWYsfY+NAqoP4T6e6OrCNc9zVlus09VecEz+dKlRJjygpC
ELrwAavF1mH4YEJnB6+QOENhBmidkxS0vtw8uC3aaxT8Hnr4yjRRmvZ9PHGBiL/LcY+RsRg7MmM3
QX9pcUwy1EIXH/q/LxFQST7qcZLvIDCy87aMimHhl/2Mi6mdriawujccPrLA6hXb3TdtBVvN0I9i
yxEwLkQdyYqx+X9473Oipk77Gq2pC4yu+WzWVSMSGeCsqiYlxw4aWBThY/Oow58veLnygaftSPNr
Xu+q2AVpRuo4B/NAbfaHwtmhHw74uMGm8y9pryjMaHO4hFjep5aR0l4rGgxcRXC+0hO5X21xsYl1
unKvwdYUCoTe35IIdi6ham7TxOlhN8LWU60INRLvckcMtV5ywwoNgURV35UPU9yhN2mnmBv6zE4c
l+ImaJvMyw3retCowMVP/h3HZ0Owc7FQsZWGMFKKPkrJxhpoJxRaC1Un9AqjB0eQb8A2AxVxADzV
sbFd7nJyJ0aWsmH7cWC59QYu0FlpGg/nyMOg6G5eluTht9DjQcquwPaUXVr8f4OOkozhv1K7RUdO
qR82Ki+QPCBznkWH+gj4u75yazZGmrM3a0L+uDxRaHR8A2X9dpugnuL2BEb3gm6mQkWc5d6OuXin
1JrroGNMtNZDDEJzwn31LGvI9y/AlqhD5L3f5yoj7ZU6omgP/5yrrsjm8KoTCEFDX/XfNaQR477u
8wZqIvWmHfoGD3jFzBha/k3N42AGlLr7npXwTJ8h0lpf0FIyOPhk0SsA65qvihYmGETGLThEQL+N
8Ke2ZXcqPeZ/MroGzGaoLw7DnOfr0tz1pSzuK7eEZg6908lbUXqZW/Sv0niMBHXPNgyIc/kIdrm2
HKTVFW/LTff3UzXAltVblP9cEQ5pv0GrDOdW5ZbBKzkMPJ5PjRWGD5mjXioaE3f/vcR4STzNYTbM
tQGki02ybZl+Q249FNtcig6rYXKKrMP5X5aH1BlUq5hkAwbCG+3X49ElDwSWu4mhS1ke7XEdURjI
N+ILx5ZPtJRWbSaBm1AUEov8w3fy0xgxrydwuEcERVq2YPsA53Pyn19nMSk8qh9OQeQKQZohG71p
MooSafQaww4vcmBJymymEouPCB1ntPJqCO8oubFO/fMtHfbYG0/VWtCh8CMABWjuezQwseXGicsS
I1Xo7sMEI1pvIcxQDlo031pqcwKIc3+SDSZCDU/WaqQVKBvkXipINEHbMV9cUPHIBV43LBXStZ6b
JXEesW3CIpa1n8JW2nrlqAQFWNpOuh+KUYEUC4zuCMyknQGmkIwfL8kwJWhISEkGNxKqoiRPdeml
yPM01m0HKkkNVx1uyJxJhY1Z0aTLmiOJm7ftohA4igYczFUF3dFGJSWJR7gEbuqONAbYG3y51drF
I6SqXtkiE/Mqfbrl6ADD0hCjgqHpfXk9fmE8EJ/joIG+dGAjLu7YBbwm7wglVVD/0IMQZUQLNR0b
lJYy/CKMHTIjm/nRtg3w0IPUjWICa5xoBP5mKwplPZGX21r7mXAqI8pgn8YrFBvKMg8zgmppUVLv
grP7hbu8j4UvqjdGAUJ7rGuCJCTtfvATWSXlD5MpGYqKgAOlqGWZf6Z/G9lhdRrWLqEDpEXFt6yB
1Ub4pUrN9CPLhW9r94FA9iLfALZgPfMrOZKDOQwM9cRB9/ETzeuSUnywTzugNQKhM9HXagRRymDO
8kSLydpLLaL2Yjd4ztRoFzmQRzqjVhrHufyfKMYUlEeb29AYJHBJCYbOAMyS4q3l89sKeScNiyvR
0Tk//Ld4obe/c1aQeZ98AXdyaBOocMRkz6WClvwsGxVrpq1nD1nZhbFQ9QmI32dGWr1nlV4hRkgr
G53tKIp/znTeM2cAZmk3SGQe5UbARaVADuIlEy4raiXfOFE6J6SzUJxxRvUtZfnEiNZLWfzQJTf+
DXSTTo5yZ3h8MVuHSO9e9Zb7+/Wl1MKysG2uM3EYxFIxQdSa3hnAgX/38AzWPrqPfXicTz8px5sN
qLCYTbtKK2NYHqx0RskLti2mE/APZfXtrcnPXbr/z40O0CyhmuxrHWTWTDLUGTxKDIBeDhmYlF+b
6iXbQezXCftFCh/qgjoIgfdM8p3najyMXhKC4SHjJ+d2QebGxXQLqZvG4y+qsWKps2HZtCDU20I3
aVqhXffEyyvcWow05L6Sr4SH9LjeMWE1/pb24u7zj1RlugjZlkHwCqDIsSiQvGPiua3OvKdgHgym
upRIIk4ovRfgPX/BD85++2ULeoW6wVhx1hCgZE741oRkpHEQsUMtS6siAsIbtmuYas0UJjM9Zfml
yScTAJRA905634iRXtWCoLewvWfXQBw647Qi7uJVjlgk10YwDvxWs4vN9qZM/p018Ug1VdhuWyKq
rZZ/V7P9fdJ1xtISsBYu9dFkSmxVgZ5s8SBTbRkWu9bv0MHLO2U0TMuriwsKJhxKlbqUBr9pJvDt
jmg2Km96Mu87rQvqVxZRR9gTR598hOrSuhwxl+GJOG0JHwIujGhNHZpi+F6vh5R/azdgH0JoF3HI
qcrd6lSdmyKzc7yq/CoA7WoFZWRtGwmjrTBLUBxtLrTKX2eD1gtCuz4CmkTc6g5wM3Bpq5ZBzOpI
y+7eiuOYBBHPhgUfp3rbTQyNdDOqfwxB7NFk6PnFpgucJxE+t8z596K7VaNRAGSSv9qyrkNqr8dU
7iynMtnRTlqFVdpcJeEWYXpObOGaj/9mpSQh4BfcWleySOnhcIkjFtAX0BcY7OyY4SdZze/CBg31
iJEY0HlthXoh8X/1ytKhrwVC4Es/8As4j6HKzH69aXt0UE5SSQegx9kP26+UVvI+5exAT38ezaC/
KgRKYVFXsCQ6elaT11Si+SANRNem9CbJY5pwgTNaaWtIBQZFGe5PfXMRSWtcdSlQkN8YGGuNeQ/p
yCSVwtubdT/bTBgopS0LaiUGqVkfKp/tKfLZIHlbOsY+Id+LxqEQK6RGm5GxGzY0EDSVDEAhuVBd
qWnuizt0IlxxAhSjmujQXDcFqogn/OOvT0YxD6RSxMxuKXD46HAPe2G3LcJRVRABKuuwZG2Cckpb
JgzQlV6140J3KudsaElnb/tAFMlj4P1nbv3CqTpZftYGeuBJ0V2oa9iBfkeHwuLpmv1uHuVHS2MN
B0oVYNJ2XEBs+HzRPoC2/Y8+RzZ96V0+mMi3kvX52QdPv2QISzDaEcB1I6G+ZIdUxvWIvzAFapo+
LLh9PhYNxOWjq8uTw/Saa5dvd/BGkH9fuyc7+VBpWN8z2ThvSYl4VKnWN9FhRKjR1nSN33NU8gtk
g1Zmqy+xoK+aE55Tm57Ti5+bvl+q1u0EPSsBh1sILwWSeaxFbpmFqyQtL68ZRKNoZ8wQc+ozyCnN
l4QwtAveM4IOAX0CEUiMhNaUCwdL16gThVsxPDAuUcAtLxDPPlLtz6HIIPn5ZQgXVyy1zvEl8r5p
GnGUnNEANMOlhrzb2FsqzNlqa2jletY3mWa29zJ1E1jRYiClUVFeYRnj+Ttum3WktRxGKtq5vXlc
V/4xLHTuJvW8mqrteYc+8uzPJWa4NUhKsu4RCefgIjPBqJk1wrqwKiixCWmP+YZGBx+FQTn+Rg6W
l6AuTMaSU2Pg7wP23WL8LIxnQJnibfrkk80cFSt8yNOPrFIHkVMOJTsXDReJddq+5pvAQ1/lqbAf
7+1/dK/bedGqUq6HdHH79/67kPtoWSDCMENUcY23sXo+B43iUTjJHfKKZaI+kmV1NBoDIHi3WPYB
DJfRF1+3ezZZNgXSk4DyY4IWGG5Hp5nz5j1EpKGBvpyUuxRYAS7pxlqFVIfX/2qF4v6zKnXYIwAA
ioD00uUx6fhjFUpcvBwFqs6rrYZFVBbai7Y1mMm1QAn1gsRMVFhkrhaOTV8dtJjd5cRRzIpPWr4B
fRVowuc7HDM2nJNwfC4cttImeqC/8VAY17i8ajiCfSkYMaKPc3e293J1bCeIEl5NPf+nZbzxL1hx
YnRVk96nnn+xb0S6g6BKxKG6zQWVUStn0SNDHWOfmvcsgah92QBfr1vwcP7m8vSmDMUfBCVXKvL4
LEz9WNmH+r1qu2BLN0xTRxQY6T5UdSyFhzlIhj8Nc7dv57a8nlcSk7JGyLgpg8uVJFdktXVYkMNu
F69tKsM/RJJfMxaOqFHy99WG8EZSTUZ/c18l6eVlOo5mQzxeVq/ySiuD+FWlz3QDECQQ/X9GtCHw
z3TCD3Va8QC5PgVMdWhIDjqngElzS66QKgqIbYI7NWWechya7orj/t59NaLiXusX9Jri6WOblSQY
IVkdMVSmE4TdFuTQ7pLQ3uqNEX/GI417ec2yyodaW8/y+8BsQ+SqwjE/aXMaxikJVNurTgGhIT9u
nvlM++cdzL/PQE3bWlJcopgkL9NeOdS3tV4D6SDAdYBQDr0pTn++JkkIIxahwplUuBBHSUhUOdJN
5lV/i90bbpF45FTcJ2+op6TRS40Cfw3k1bQXEJoV/OxH/hrrL6CobgLpirw/l1AxDtvu1Sseafon
xfxHC20mykYqYz5E+XkRDgiFdEE03NWVfqBwtb8qA7s8Oy0/a9a4yLj9ovtRI4ou4+uJotKNvkOC
W3KzWg+4HGFB4ccwajcVoHIF7/itLpFaxdMX5ZrViDH1PDlIcDyQRcGbXPW7FPC0Z3qNgP3JMKC6
B+0BH5czsyD1yG6WWMq7l7OCjF2yZVq6+fHvxN61yyt66zIpCs41dLfOWNzr9ha1Yoh9nS3oMm9M
Ye3vdAAhGMaAlAvlG/+H0sUt7XLUNBumMckHGr6i7XXOcd5xzfYC9BBocwqSk65MvHNnTVkgOQ8e
XEnb/imLRXleNqztChyJ1ZGvpvE5MVwnh+rPAMbZti7eloW/bNW8hcoORxcQa8hpwWrmsf1Wh4CT
leMNjVuyvyyS6duwO+vAGDgAfs7Incl3RWepsdSmvL171lcrPmAlGJ4kJGxdUVoD/l/WWNxxx6ow
15h67bAPO7qkaMrJPnUh2qp6U3CTbj9dJG7vJcRspPeRl/XCnwb6cvI385xz9HHqkVleqc1GsLtU
FydOUsAlPzjWM0xT0JcwEkPHEHt95xKBPVxhkkUwewaoI72JD6PVi6Ncx9f973zG/W++45olgSHg
ZictMGbFN/ss4i9tZOl9wDEdTbELILKUiZPT8hQLSx9KFnY5zqZatbok3ikIQK9aIeSy4RI1wvJB
SG0fF0+3BgJgL0YUXB04eXBqs5Q+NKC5PocsrM7z309ihxEU3dcj9uv2RaBRmdta6cqImeGxcfnl
J2aHukqmsjAMRy5ks+GL4rb5ZecY/+n0EkWNP6EjDuIarCrB/dujwoWVHhi61EmK04oDJY8X1KmG
IBbNQhlBn2+bVCgDHAyO2Vmk+mnuZ+PdafVX2StugIBIklsgF6h6ThhDO4k0enS1jwFdGZhHa/M3
+C06sXbqn8U/Yf6nA1cATF5BxrnYMTAjMOPfeqCcLkACFLsi1UE0699PKqoVA4g2jFQNHX7LqJ6E
3zKfOgvKkMfNG4XwVMhRQoLPKMdBkJhcCz4kmgvMoHBSwCHa2SbB/anaVsMUmLSzVtoBrLJAC1J7
UZCQyh9J95bBaI/jCedVfi32Q8A97YZV8+EYcLo/dU5/Hkh9seM4+EDymehKgUwnZXC2EkgmYPid
PidiCmPEO1aSaVg7+GCeYowmVi1jodJ8lncddXcnPDNHeCKBovGechBDODRiC5FZSNB5X+bVFeSq
iHxSiPDkW8hdAnRAfzuyS26Op77GedwbXnC/d1WkZIYQ9D3cLFQ3mEgvyJqZJgilCeefuB2lQBk0
J0M8aDIxiwO6WVn44s5iYukMpnTNIJIPqU4Q9tLWDsgGpLxXO5fb3F5QKgrpEZNoswgZ9/UuzB7p
Khz3aJAYiVBXH/45UWSXqaNqNCb2L8kcW0ApSi1kDqNHFXIv0CTJCqcJWrgM41xWqsmPI3X06mXE
Y7iO/VTgSti4bJGUwuJlM7/l1f8PggyRhAcb7e1wMHfXnvvHoulTrQNFDPJOUGvlBFGNMDJQRHyy
NF0IzC22XAof8NDWF9W5/bPyInoAWV+Uz2TCVEmYRkbphKMHZj8WLg/mU3HKYb8FLQSwht7feWmF
rogmZgij3+idAbHxrHc5OzwE33DjP/NIk0GsotDEaeHSVyP6/mVZhl/zYNwuQnN9irttMFV6Cojt
35hVHrn60Ou7y6mJO09gkWOapfY9WSNnBB09Uf0tzPoyddchG39fYyAduReIOyos36lnEe2cC5w5
9TyRW8z+mDakoyaRl7XJp78HlvCCRRN3il93kTtf6GoXkrnR6+tfZaAF/QTaR0yXE+OfFzHL0fWW
qpfcjb+khWs+hNP9Ffp3s/LC9y3DASGQ9kumFpbYzQrhekoVCHNHLaTlq8MI3Jt01d6ElrFtwdUL
DwzzBg+M4VyJbdFL4XyAXjF8BUvwBws/vZbTTIiEUH9S2OBZJGCu7klzQj2ojNN9yBs+reyoy2dU
GB6gJK9+j2DVg0WqDYz5baQ8Ine3UXOobwJLwkNAHiQNkCF7bLHAU6pFYySOBlmrBU1vCI7nkkQE
lsxQqL5pZ5PZORjjZykLBZJnU4GSsVc8NRyBhSplODhBGZA5qj1fyqzt2xGnILbhiBN53GSUVVL+
zgy8jkTkS4PwWhmV7CGPGY5urNbQG/0P6Hv74Xj+EBTfZdrW70LiW4z2aFvxF9RlHgy94PDDlvBa
A3TYrRzLmcU9mCn29qcR98BJv6Sw0m0/pZUvce8u22hqVB3Qyb4sphA4hCecEfkRMWwi9gWdONVy
pdylVBxy5nnf21lSKo3kl+BRuT2JzA33DKNDyoMqBO9I+I/4EfYheJfzqmWE9QcWVa5/wWnMLWuS
X7PgWgb/PTIgEpPtBjL9R4TADKyYX6LSpj+VBZO7LxtUcLv5n+5U9SF5bdoSCytDAlsp64zh9KB0
cyuKQ3H/g3srCgoDo/anCFZxIiyPlpiLszA7Heoyu07b+pyf3yNwLw1p+SPo6JL4WjwbFi4O9lG3
vh0Otgc//hHzHXHSNC2DMpBZ61rYG6M0hAxCnpkLeZ4ZUxxkgSYEV1MvrPu0mFhSvcNrGKieRAXM
FR0U+wa5aFF9Rqjapi3AvuGSPT9F9S5Ee9LuWpM9NDooANWHwhSmwQPfuLG0epVLqHGGM286JcGL
NZ8q/Cbx0bOzJMqbgCLFPl7ju5U7+2Dcb+PaY3LtKfSMKlF1+U3IfGGxjY+x/nLf0WJmeKTImnuP
VXJuXEq5YscZdUBzJPXtUPDB4REMsH2WO8DM8QAb43oon3FjKvf89K1ZCGKZySRCf2ikF8F5L8Aw
FbLOuKcEjdebl0d3+kS+BM6G6TWOurq282nCkUlgH75Y2hEPmRYEQ2iKo9JZavdQSg8sPI0vH7vY
9ChnA2q5YpUwaelSR4EFauRg3xXMnn8tqjV8GzjZpatoexHzrUZybxCboACBr9pQY7XU8NYQxxTw
PfwRJTgnS2087jpdvmO2VOHHdHNwbuOknrAM4luoNPAM2exntuLPn9NyG6R+1HJ4i28O9tnOAGOW
RNVMHHF834/qWqjSw7tCR1lyr7JX95UzBHEBxzm7xFTwZlhQce/K86aYIgOcPD5Fdfz1VNkHKjT/
QNHzeN6cvcj72pPXNJp8oj6qn9c8ylkYxNHSdHb25XcHqTuR1iPRrYR2DtzcvELa1VNuprBR2TJY
zg49fo9uSJlJT9VDw5o/IEdO/LLv9byqVZ4UK534PMeQmp8e6nrbqqmybnIBvn6tY5gmmqIaeuwb
1ZZeaAz/FeC1FR73mrr3xubmF3+yCb/6nxB2HkZrJjXywH6VD8TktyX472HNvbbekc+KWIFfwZS1
L/MFsyRPMv6hgK0gyQTHzr663SHWttVKRSRgvRUoU0hbrU/VmcQQHL/0E8xEgmC7WyzR8QEIEbPF
2fQx0h2A21sQefLD98x5mUk6Tl3pYf+UnVio5OsN1nBOdCK4Cp41nAJs1qr2M+Xq5bylLoEwkIc0
/WGCIx1cQw4sspGvDL5rwlBKPt2LxXLcB49ZwzM3NvYDIBBKgecX7Pe3rpA55vjiIcggUXNuMgWr
ZtguAlsh7ODiUq+Swc+zwxC4oQa6vbyXevfUl7ACxEDC1/gcX5bU/9eVPP+Z/dS5FkL3jUw6gHV3
AuB7pNEZMSwhRa8jpPfzvU80iB5qXe88MKiQ2riT4bINLEsygFPt9xhGDDiC/E3qtQuZHcMXDSAX
QVUv4+5wjgsm+ATAnMEE8mJYoXan4k/PeMz+EVQmw7MyApVDxH3HtbCCinm9PGW9IkpiANUGpHUi
paSlq0hvKIx6LuAkbtp4pd4EeD2PU7BaohLDWjA8mKoMmnGp0fKyHH46NGu+gbjc/95ycTcIna1b
wYJQqoNY6k185owRlbXacUla0Vj3o2XXG374FlbXocVUaxKKKmXr+/VwJGrz3hW9knFaSPn3qYxw
zvu8v3oCQeX4jOUlkgN8S5KgIHYzA+RsuytRM8lvrq4K2+3gC1y/Gh2SmE/gNfxDyAtcTcp2Urvj
FyLS/uBhkNcn4QtoRxQdPKrysW2JPJLnzcJSbjyBLaz13LG7k/AM6GgQ0QXeO3Kiw6P3sUfJTAp1
BBgpND71+8kQq4gF3RaJocYmhaCTOOOtPynchLteTI1DM2GgJcI5AbKErhb7BMCtCz/Sp9xWmB0T
5wn1vFvBBgWc3K9Xkmx6U88+3mMI13NuOdEKXXMI+nx/AcHo4sRcpVexGflw2UsJyvSLJgpZaR0k
LXsfjirGTjL/tu4x99e07E2xaz77VwcUiUVXSvxM5R17ONb683eqUTFWAx0ybPbUG6Z4r5rSZsya
UjGdg7Ty4kNoaoeInuX4HTy9j+fKyCwbu6us7I4OucMTrQrMB1ZhBSGiUuC80jlXSEtaaS4p/CB6
XPjPlZzAjpgvvChpYE320hcVM4pJLkEM/Nm43LZuqYiVlTspzi1JHMDOhP2BeoWHum/dUFFf/V4q
7n/ZHP/xkEBYf5zxPqn+1vQRGPkWtUdygTdKw6Z0jtLxh1BmcUGyPoSnlWuR7ZenGaGbX5X63R19
8JJifcWs4uPwj9fy8TXD+nOr1wR2RuVSFTqRJ88X2Zizd6aHwYWWhxT14DYsI0jJxKrCkz1rtibm
cjiHhmMvOU6dfyQxjhh89NR571DqKXMvZo8pM3cfpaRam1d5/4eoWVys/QSQ+2jnqAZraDdzsSKx
DK8or+6dbvbRS53qPq02Pyu9VDHAUOxTl4IsuydXu2EcylY5XrI2MQUNF8qdxkGX+ig/u2UJLRd1
vmAR8imqV0lp1toXIEbm5yFOKsRzjM1VRzocwuGq9LadFvi31w7tgZjVqvGSxIHkbWAu6rTHx4lq
SjED2W5yHzXjUgGg29nqFaRwUQ3JyNho0fIx4V4i+0cI9hhtKoPkiN2nBukCXTbhDsUZ4rUSkWZX
1zq5Z1z1kU+1DbwOHAybLYF0bJ/jfAiApskNlOuJVbP0nP1B46ss6KfixCxb69aF8dQfwq/nQp6n
qSamt5NF/FoNaz+46FksYEyGwtiv9RHJplaPiQUmfjrI6+y7ECvAhjUWwDTyrq5Ioo6x5/sSv29Q
ZUkR+zzabzekqPe1AlUtFcUvsDgkWa0KcMyZPxs4aMp1O9q28HMzwIIaTeUDFysRgmG9V62BinsD
Hf4PkjiMktlJUlHJFomYaLEnI/ofb7wYno3eTYYHJYPVUcuHUW6NZPluFfMYSw5gRtWePGccK8qb
xYSz5M/x13YcwC5O5rPoOlQVp66cLDEpqw6L68DGzDI7cv+NDHay1Vcg0mWdMYW8ZbKTTTTNy67C
f5vE1ICAw1ttwYrS0eRcx9Cbm9VUmSldYLytTIveLO7mF45QYW1tq43vQG05RAMXwysQUHmvTCvw
cdqxI/AC4Dmhb07aD4khoMuD1ZW4oQPQJ46UVUqkkZb4Je3Nm6j78oIj4yfu0QW2GKkid4z2yzGs
7PWYkmX29e3+f20rTefxPpMIcZXiMr0Sd1L7dUWF3LfQSpHQQcF2gCCMTSJqG9py8ZVI9HvsRi7I
OdliB8SpeHWoQQnEHfhnWU5zMf68bKAImNyyDtdgYtfsCOGJ/vQ6rTmVAXbEP2gBiMSt72gq4IJ/
oKPRN5E2nSamPY1EfEffJMktzwmbifIC1Ja3Mz1ugOA8IcHu+NLT6+TP/T3FoyXu6nOtBttuQEc8
X8wTxSoflmJZZ4eQ28VfFKyZzB+lFbV+fDGtKYXmdgqN0eCEqNWdmsRKIEPtFkS3XgShFw9IZv5Q
LO/kJzHcVHF2GsljTTRI0HUVSlvUKZgY4FWie8DTaOjgAzg2YKAeV79wgSymgDF/1+z2pbKM/1BI
JvUWtS30EgKyvgAdG2g4XUuD5XNr7Rnk7ScynCsSKGaJo8RXuJfU270WeDuwDa/i7STI6cXvOiWD
WsxlryBK2EEe8Rd7sqTJjWE/iNbBKSr8BrCYAe/WyAq5IfVqnQdEW5eyqQ8/bF0aLdOWAl3kml9S
GKRjnshNgkYO/2qGhZMYhuy+tzTKXy0egwDpVfkYq5igHMv8Y2Qo6unweyDffiFTQ4JzrEJbstAA
g/jfU8NaPkeRDU7WCClTr+mG97iTjS7GKgbAXZabo42MGeBrTtA1j4hf9owlDTupw+M+tr/y6xIA
9K/0anQzCl2JhhkE+JDGooWJHMQ2q4qaGAb+kjbbn2gwaC4vM5ikBr/0AbQVtWFEFE5tb6HGsnNE
O/fSFwL46rv19WjdTy2YdNQhiy0pcr3rSggvwvvFN9eg6DWyOZgZYibfw572LSWxeOASOQKygzK/
KqXp27KhQ9M+P6jBLg8JCdMN3aJip6HughynKatRjiKWRwhOj1dKcZX3L5S3qRwRlH/eglVWvdI5
wpvcXCkRucNrRfi0IkPYX5bGEdt/aIgaO5fxFMVd3dSWV2hLEm5xPMjW8emDDJuXKhNB2RYTLX0w
IO9kxbJ310cJ4/uYWHFIJx6IuTIg3pgBBJXpx9mEtdjUx/l85zl6fVTDXfOyDVyUAn6foN+4fTQ0
V0KPs6sDH8AbjNxUCjWO8dkX58WBL5lNTuRIPczCxVmTC3JPQozQUDG1GKcbP4Qq6iODuNqHoyJN
NCsha3XlEI8MAgLZj3iToT8HuQK1+7Jl+9UjxeBFXq9ntgYzJjzJfiwQVRPrTcQzEUUtox1DqZ6R
U63UvjNcB2SP3x5GgRhKYa43vGMoYBKsFf6cjuZDODcx8BxHHUs1cZV/Vzhe6D03IPkF2VmvorgU
k5WWiuK3ta3nkbS/mRtdhdNs7kI1UB5OL11s+Vx9uFVZOXr+oGYLBhtkPQa/k9qXGzDqKCzOFwSD
2Ocb/Hiep2zvAY4CyFHzZqncEW1XGDAuniJLE0tl+0/ZeVSEeIOu3S/Ymrsp/iD7wRH6jG3bT5kg
/Mt7SxvWR1dYvtSSQwmR5P7LN+LytiwzRm/350xfjp7ZPaWAolArScE7iQNnn7nWLTZfUYp1Xguq
pRdqgTjZl5HeNjPK22e+N8kkovDtSABjSJPwtMJ+8VEHetrhUTohOBIj1TPGpdP6fJLGuHWpEVZY
NBG1VOAUiJy5qLWeqk8lLlJbz2OuU2F1QASqGy4Bp+5RBrvDT2hMLFr9vYGk2/ObYG7JDjWx1we0
NaiFmuX/sN+QsfvZOuY0Da6eM/RDRtWcVFWOqelJIM1nNq21KHq9uE8BdTkyuRimVrx2tmszv36f
FvB3YEb6VF03XELjy4BA+1iyWDhv/v5WvgRu5HOO4HgZbHQnueV/+ws581L57iEzXzw6SsSYkbJ6
gqzM+cF1lbxdvsvWfzSSk9kxsStXCIEKQ7A0DfT4dXPD4vr2OKQc1tumqlCrj4l1+blRIwrQUI9e
pzH3iCNrh1xj8ds2wq+MsV90LWhuoDYVODetqsfZ8jkXMt6SlFCyUm4BFbWCJm4tmarpNI2C1uiS
M1teS0aMp5ydMfCyUVONXHEpZzBJ64geKs5k2rVM2HxiLiW3E3l9iCgeyEAPXTUA334EqmxzXFai
1sBHMCpl+BQWxlRMyT8uiQtEg7HgHSpXxt2ooaobTR046y5ZvPvU3gdHNLJU19eyVLT1HtyJEq6c
s+kHZ6zdzeW1khDwlJ1si4mz8R8nvVcnRci6WNI4cVqZaCk7ahRnuKGh2chUfXaqjNuoi1NG0R/7
qtbN9/aKJArhlk35ntUrwAGNIpqF+K7T6ott0t9Ft4NlUFWUcuK0zDdDUJ8QaygDz9bOHpMKV9fH
cfC8P8wXWyd+j520/a7TEpdHjDnBglPmZcgc1bcDMpuG3lBZKM0iSt7WAWCZSzcFFuOi/i/NlnUX
9gPDx8ltyifT7Rv28M23ekt50BBgr5iWpKOkN9SmUZlC0xyNuQWlXy4LaDI2G6wfh1n/slJ+BU3d
4eAWqw/5TqKRGYoLjsA4S6saVNxexwjUn6Iez3h+I6LTn5cbVJw9x9g/eI99Rb6w7NUkz5F31AJ8
Ju7QrwFohwUsv8Ru623A2Nn64i5oV+ZLUrez/7mFlHoQGCLE6tf4GnubeSNTJNIXYurJgqSdsoGs
ZH4CCvhAO5X5M8ZAT97SWY2uIhAD9tjd6M7mJHYFKsyTjE7RQpECWgSzvJyOWOxLZ+QV4vWp+Dn7
7peSj6g7fcJ8q8EaFHow+S7bDxSTtg7+KBRz5ZFG74xkP99AITojzGMO9uqswg8PD65+HPETQhEP
Lcy+eyRL28Vz4nzZtMybQPudlgX6mg+Pi5JMKFq6Kt+i6IIAvkeqvvJP5uPu7LhflyOqKX04v7ey
HzW9ZCATUMCQmuNiagVHBgREP/7CLtdSANZvyyUrf866yx/eYK37LankMXG5cpHsfxDTtjTmg8W0
qOzzf26xtWic71+0fcuXVu/os7L3lF7SnooY436RyL/PGbXPdVg3d/DYNN9whyDoDzBLG/JstbnN
xqo09tj+z/Ci709TnzwtkJfZlfw2W1NKUXcgi1sNmF3B/852CFz8m0IZreiwF3ruExFmxBz8IATe
U8OXv9mGfm4ZK/Gea/43tHrTSOjGedIq71BR+BfAIsBMQe7JnRHqylzcPxASSIZmUlwhePynARuA
yvuXSG1kGKcnc4FfKlBE8KdQIe7Y0CbmnPfX69Blmy3Hlxubmxogvz8u1ZF+FM2JRB3KBylqY8C8
lbR/PBXIY3KCjjF1vjanOhmRFLkTDhrGqbvML4lsJfDSgM9V0ru/ikeqZBg467OuSG6j8o3vRm6K
MWjjKmQFT0557/BcPD6NZ3oh1NGb3PXtQvlq4bOUITzW4B72bKp56z/OApRwynvW9valXNtAPQvG
VmTvIiviDeOvz5KQ1VGeaff5dhV+YOscr+dL8yudjD/k8E7t5Ky+oA2g/g6h6SSWsOsMEBNFzC8E
HRGRQan04LI4J5qmwuKQxV0JPEYcfy3vzpXPHtyphMd0EwlA1gR8RRXiLt35LTIL4CcYSPmoVokr
76Ft1K7yA2mljvf3SnkPhkWGNMWsRSK9JuDn/tsj5mWRib8c50QEie8umNFtPPLqs+aR5oJiIslh
ghShm796kUswg65fAFA1zKmyGuQTMk5/PkkrrRLNDLErC0Hl9Ecjq+AwtzILbVUszjDZ3UUOAVgb
09EzhLcrtI9R/NznuC1/7IbjEkK5VkY6F7fv0JE0263XUALaQKBlRRjNvbURjZE98nd65TWdiPuz
Vz0ScmX2/V27TA8bEYZCvVUOsSXqvu75UHyh0+YOcSTLy8oKFsfqZgHpDj6pJGbkTf3newmo8WBX
u7mKRsngTDXbLx5eCTR2Y/EwH+OB/azYbdkRYK9g0oqnL3ZN3f7Ju+t8LqZAT7PkfPB4ae2S9OZT
nQQut6RBaBt4avPUvj5S+K5nyT9sMvOVBEqNSFok9zPvpbxw/iqSwdGwZMFshZixF1amJWyIzN1G
zwodTBij7UWfVzB5Ns0r2f4xvZ/gnwzkwE8L/XKW6v0JTnsve863qi89Tq93FTR6AkCjOpHjCfG5
sXXHpTGGeA5k7WtIIn4Pmx5RdvYH4y/pPcHUoFmeZzPOaU2sX2B4Fh0MsxeelxKUFaiebsN2XePg
1jACFkgm6a/ZpHkJywG8Xe/Iigarc6glRviN0RPhUiz2dOw8Ki1mdEBuzq5toLo+1t91rPZ+SJRG
t4m9KJ5T6yFwcPuMj3IP0aDWAtZyUENNAt/pOE1X4A7cA/mLnallHDBs1I1UnkXLfcQulaubR22e
i5fEOb3I/a+OAnSe87x7PgBcGfL8/70r0mJNXn6OwdAnqqcdO0pXdFcseDhKLZV1b6tbXhniaZMB
H4FVmU2++jtURiPio793JnMHsC7YyG/4sy8ucyV+j1ToSb9PTzqrCjgpcCkZ+UFXHerkG5yOmexz
LySjfNzy89XIxIbXIkH1jg//qQHsZq1HYZde05B+X3EtFPep043iLGzQ5o6eVUpG9Oks9ebgFhsh
GhwJdPxd69rfZgsxbzKkX1VuzK5wX0fPS63NbWMHPrg0ECn69XSxrElxjM7nAjheo5F5n1GayQKT
EzhGPcf0It8gaYbu9sqvVtL/Q/dSmwtwplN11zuVFm3VR7h9Z7kWFN9uasF6IHIY8uqZYSMmMyNu
xOxZr355SGnrw2oZ8r/WdqdZBpfntkb7OdZ+fRbhCXutdubqf43FinstRhOnGwTvRJ6nRPfVrKlO
npB1CNwTkBBYXRlB5swP40GlH+rD7gZ0gFpGsxFXQ6SQKb2+ICGfeR0ImetvV/5viA9mLpWIBbyg
0s00tKeNK8xUnmEwXJ7IKDMZPl0BbOxJfs6slfWK+5/RqKfZe4KMKj5sKHp1GM3s62BvI00g222y
jXIfzsyfO5yYBio6Vm1U60uMbprPkuF1dV4fAfoFA8OiTeqo9ojgVZ9exSgn0fAMDHFWZnvcrEV7
t48sJYg43u6wb6nD+YWTZjkabOk82cRXU9Sq4EVTgKBTHlynliWpZ9Bj8s79kC8CKXa8vEqeYrge
B2iqlRCDwZoVzwNRmork2RwTLukrTtsEI2Q/BOVPkmzJzw5GKUp9Buf1sTtmA8pbnUjyWjaMUJfP
gcYsppEiXCVY0NdyiQvykoO0+wfuYm2QywI1zxQHA5p4ggGiaP851rThcKGTCtIayxfahjEANuEd
AYbi54NsPTCfmyUwyyygIjV0GC9rilyQzUUUv6zTld/Qk/Cg/R9sQpc5n1HC4Lmb900q1hU6mtY0
0J5AaV5jEXsZke2EDWna0tLRJoScnywObstw4SbksKUZg3LYNchweF0Y1ZIrhDcv5yuT7wwax6Ns
Slmwg96YKG2bOKRu8EJOvzXOqMCxTUcM3e6ujWwEr58Z9YZUsfPrbSGpMN//UBWabdj+qcd8KGqu
tfWMNcFoXmcwYftLx6PCkzaO8g0LfPFDOpJBS9wbdqONfbIRp/zkMJ5oZo2/qLACgMFBxs76QVvK
N1QqmtZzdkB0WeGbsEfA53EpHazP1w8x2k9SmKBWOXdz6THJXBJAv5vjXiu5X7xdiHywFdFIrvM6
oWYt3Fy/QmpUcP0Va9qjITGhuUbThuhyneAXDoNaeLuvUpKw3iF1TAyITyO63eAqTbcWcSLl8y17
AXkosXAcPzYWHcoi3U83IyyJuQ5lHIwP86s+kNWJlsfnJZeWwVd7ejj+HnEuHwm/3Ej4e/Nv0VDY
l4wixVrNNAh82VWagVAWI6fmkGQ7HwCLeTAME93AFhIFSaVH8AUhqvt1hZmYd/8T/LwoBJAyqiOz
v4hUmAOob2bXO/yoLvFRJk/z+5//ZHssEQfuxmsWOmS681k64EuseZuESjdBTIMdjC3cXHPIXT+r
17hSUSykTg8NEmuo66ZOQQJH3oN1EA0D/vr3I+iUWEffVARv/+TN3+UuAUIQYirE+A4T87qNnEWR
D2/fGle1UaQPNMt9hpjRv4X+Z6FnH2JZHAn+i5yzJ50hcM1HNfyGJOiuul2NnoRvZepGIlVCMwXC
WfKhBP8els82h2UGjp9VeQ3F3S2O/yMq5Kc2MPCx7PXMji2eDWUnEUyrRh6ZVdcbIm3j2flp3qks
MGBckgzW2g84iELKUuc71nykTvOkKcciB20MGGTisqP656yUeMcql5y+MnWxalmymf6uQMtnO/M0
l74iEk+tbj/TNErdiwIRLsVd65xkbfaka7RS34mlIb2uGDk7t9gxO6OzI1XYQgFi16IQSN2sQ55k
ruOgl0WU5+qBvMj2WdKK6r6GcyNDeLQPThjKlKsARJn2H8Cx8JPLQC+qqYghln67OjQ/V314ynkM
yIkH7Try1xGAck/+Vp+wMUHuN34Zgh07X1Hfte9MhyZLF37L3NxriJ+Z8CRBDVRM92qDYZNcXUmL
O636zU0KUupfs14d2DRZTzuMkIPAi+adzrad7w31j02pbg/l7140OPl262pfDISNTUwISSOsOLXv
8fC6vop7qUW2zZ8C4mu3HzA/RNmooFajxMgGC8LtEPZLdgSMSLzm244O34qgpHA1rTcMWZd7Kq88
GQonOA5yrELrvDa3SUF/Tdvk8y3f0tmDywFZl8mmM94uuZHA7Tp9IKpYDlNxZdU6IuoxbhuaiZna
D2qqMlPQ6mIS6srbaCmvfBlr7MkqOpXOZ3akAZ0GqrZnU3brIz/apsGnwraP7DiHT3E1Q/IwvCE2
Xc5tVeucSmupLKEcEwyabNmvO/Wm7zE9afj9whlSZ3PAxQQNtjEMAlAiTJivaYkNW84HrKr/Rr8/
hyOSrckJK9NksEyXwanCeyfOemCApxQWVxBambY/mJ7Ae2oA1TaBdbdxh8jPtZE9d7ppt7QC9mD9
lApaSgPFCnL5wR3GXurQNL5nlRHkCTBwewrNYkfcMC2G/GPNS+uPt2ztOtd3/4PIJUaKtyi0QyQ0
VzmBJOS/ZxTT+GBb4cVbA1p1M00ldgumZhjnPoJLLESBww0FEYlB/BYW4N93eTwhEjrKKca7Vf98
CxJi1WdLH7Ac41mzA1reyElkxxrYylHcSCyzqbrtDJdnS4Ai7nZy2r0KmLcgjiUyidDnd/NkSRHl
XvwnMg+e8D5S19B0QZ7SX9+adjC1+feTltt+hK917G8vQoN0/Ah78bPhjCcm6Qk/E7H72zxMctEv
egtvwJfiYIvg9Jg3YqiLr/oqxYM7OyzhzqFGZ4UPI7CKrnOrM7cMrOG5FESFJYWrdQ5+QGM6Wgdd
yy0S+AUtQoBMg+yv79VDnslxmAbpSY+EYwFopc95oN+F+4HZ4nBJeP3HEA/wJzZFSb6bLbmOpqvQ
PoYdPNIESfrjE2eg9Mmmur7ZPZGnzdfAzHEXtwPXguNpjXWSRQlopOs/lADpFyHRE/P1+O1KNDM1
hyBfC5mE+W5sY3+riR6sqMKi/mEWB2Cmx1E+7H/EM329IgbvqlfZmYXONIgL3dlIYcLK25rCsz4v
oluedyd8p7gDnsxBDqzghujR2V2XgaOyWsJ3+Nqp6Qw2VLBxot/sB10u+mtDGU5Pf38vvfGf3qGz
6/I2t0BDG2oNvc1P8xXaQWJrnjB8lr7BjefjqjIuJ8NEZO8pR1eDrlRIjbcmDvrX0+ohLX4jJ1Uv
/AkFUt8xKbXPFk2tJvqGUZDd9NiUYCWxxGYz37bKST9WV5lUXHb891a+uleStk6eXBQgOizzee6Y
twwPH/GxI2AHX70eI2npwkKZ+qiBijactcyxPiLP5rHyfyfZ4AC/BW1hzpRC2lWaWhk247ow5SRj
1TptO68Njhk6/iH+xgI+JTnq7wRd8CwV2YEVVF4cStxLyLQxOAnr+aY4/FmIQugz+5kIg7CeOYWU
aybIHg8IB/ckXHb1sVyGDYvuXe3V+EnjG6GL+lSekbJDdc+Yjr/CmIv7trkPH8lrlVPcgwtm76Sn
73CEqLIOd/bFATiwsjgCKuCjjPz40aHYhV6bQqMy3fKtMtGS4bVqXvRVFEvkEwfGShA7Eb0l+KyC
vgUA3wktY7fos3XwiRV/Rd0gTFXSX8B+e6f4fWUC6D39hczdJ/C3/fTK4IUQ+ONqGGgC12NtzUZh
kYyL0d5iEparyg3JMydoNzaqgibj8JVqFe2b6dk+SA1EFbv3qlDu0rjH8fzcE4ZA/7YtEWK3/TC4
6/Y/weHLrsd/GxIQrgpSasWbSC+ohG1i8ilXGqJY8IuwwpDddM/cZRlp01sCVFmnr31SAkuywb9S
WsN4VIsshavkYVjLY+xJ5GPRD7DQkzZtY275YrWgE4RErjEmbvz2LcuR59Ff3tIAsy2ZkbAxNuVQ
cm3HY6k7wQ3X7oYM6z39YBhxavoLa30zBTVuvnGPK9yiKYvRfrQvo90YwGlaXP26ch7aiA836PQ4
5GzWexxGGnh5cDDimMR6aKfk6myGCZG6Ewih9wxSU1vQ3d99yf3KceVSJRI23sAwYYs7SDKwGj0H
cd9zTNoPdSUVayKmZzKBa1tGT/oBFWjKgh4zhnKUvVeGigKl6CKwyb/HRfTgjjvq4J7Kn04wGwaa
clm7OTE71KcxMQpULc0p+1+PY1gX7+Ro68Dx4eYbnFNBuNvC8zAuH09G8anf7Jykf5gYvbxOaPK5
66AhVS9ayyOoJFQEqiEsMi9Y5rdb8lTGGAuxECepvyL5kGIfyyCRkSqVrxle9CZauhRfzlZ7QSDV
7vH4gEuaIWqpYkKJ7D03vMmbDbN43Xgxg9nCRnX8IGYuddI+tJy2Id5bsp2UmGWtu+oTX5nbbGEk
4TFld024uXE8VOh5/Tj0q6SrmZ5lDm6eJc/ZeMn7s70scaTCqPpLiHFmUkypKG4WFXuaz6CzHmNq
8bCpbMzZO0R9AMhgFR1ttASZtPn7hp/qQ+UbbiE4/nIOyHwbKufcQ87x9WBVve22eOIvBL1GSpwk
L0wWpeZ7s0syYFeKSQCi8DsGRV5sXipQzHswjYgBgaziprAPPAkvRc2udDlRpl25KlzDzt8pfw/c
4+rjweJLWvHDf2qLK1vOJkiLUqUNk4zpWrtuk90AA0DpVBjW+IOKTj3YN/bNwzeXwE0WkEI77glM
Ohqx+nmntEfSwPmEy3lFoBH8EBgjw+mrG0lQrd5ZXmbs1ssHjZu9TVF+i237+JZTFybUkQV6GDes
yAM5syeXMUGBxVNmiy3fVKxF3rMqrXtpMr161Al0uLTC0l6PPj7Dy8yeF+NhDuYBYeEgsTRsLBQs
FxrdgEx1gQdlLljmf2Pn5U1hsF5PoBlzwxS4Y1efwm4g43J/y0WIPc/G613SehCE0PMYMvEqrMQA
5MoKV7STWUTC4cP72jZOvHWggdIS6XhHfdal7tLPbA5clVIQtbM2R4IyOFM3t1pH9CS0bk4WY2dY
PmAMLAGw2rypxhYVJABDjqc7nJm9RJYFRxZqmQiaWfwXgfVsL36PLTZmTNklvq6voem5aNS+2459
fONvIUlddXJvLDiTuzbk+3jvxFCyT07+24FH9TONAJ5feUGkyZDptasLO2bKpGY1EupjWPxG3CyI
PhLMWyGXWZSo2yOjj4eaz0Q/GEZ1XK2S/aU0qzttGfE/SLTp6jMgFePpEkD6XsFO/JjnVAGZ+Rir
fqBOJauB20FvAmcQr3kC5E3UKfDOGAZxENFCSdpfzoQ62PRG0cGtlqDHbWHfumNpGSfwOj+MVuw2
Y4qSED7dwa3aimrCUQdH5BCwjsaLCcFvmXXlb5WLlcN4MfOfpqL39xUGAguytBnZwKi+Nt90eqFj
zLmwCpsQATwoqHGOYgepc3t3xg7z2GqRB2u5E6OQ8ND1ccryi4dSNfOUe6TjUwvOjHSSV4HymFAb
dZC9h33O8zf8xL0DzdQmbenxcWWiMJ8nCl2P37ZI9GtDf+v0u8GtRpbU9+UPddHHgn31ROBp5NhD
cEAkWO1+chW58YuPuuHOmNN0MEsVd0i0Hgnu0CE+/k8mzTYkhD2U6c37Xbn6ZmhR+dc2a68a+IO6
nD4mqTP1r1HB58O7aCDdYbKPus+cejv3bTUAVBqkfFBPw1KcNVDr5d7bf5XAOUm8D8s1G8n/TSli
T5FCVJjF9heorlJnzvTgwfdRskzWSQenLiRgnfvtM55Xe0dv4bERjLINeXVlcmccrPWLyQn0t3Ah
PCRy/kSV+URSI9FzM26t4zJ633ldITsF/+ST5ojI2JRIOvHPu7FKBS0jSMw+3r/U+rTSJu93U56V
ECXTV4wBK4sR+ehBdiKq9xMuVyhKVM6Xwt6kD3eV/5XYF4nPGTCR6v9nZlnVRsECShxegyEP9/nt
AcIUd1B/8hmNqO9bq0YWDapPvq+SFw/H6aEO1BXgyjVmMNXjF4nQ/5fnN+ZX16R38Kyywkv7CHLL
WOUVsWHzKw2FLvfNULl0drpp5AMjlwscsuJdEzRSpo25aqdRLI6pu7kWuXgkBN6y+5F6pszWeaBW
q5k2T8LSDX4RqYyf6+Fjo1xpd3CVQF0tRzhFX4oPgk9HSgPhBdv4LNZgoC5K7JFM1y4jFQZ5Ofbg
zOmlYjAMMyeoEj1V8PW+ngHXmGp1/dM1dgeuyDtYpkVIumKoezTiCo1aBxWVDWzkQDFJygzLoqhl
Tb83tVTPhhKQAjmLQecw7i90+RW4GL11lkl8VG3qAc1aEKsjh0rfEZPVtopqqwWA47IG0NgE5VsN
yp9LOqBbxxVo3iV3PtHLlz/rKQXXjYZggz1c/Q/QxReoL9gi+Ry0ir3mQySYt2YOBVH3ktu+D0IH
2FUHOxp+kj3Ppv1HssMiCoM6Wb0WYG6UkeOwe6KWgYt05KB+TTk7oxT0XA/1pu22Ef3tuQYBi6ya
K+0EFgIWIjji4c2CjifrrHl6hh02iO4miVe+AeIP4krro5V1r9IcPeopuNlE40y28HBbf57IwYZ6
Qri2WZBvn+Xm1tEZscdNbTw02zi/0dPWdpKH/Ua4SKwXOWM/O/NCrNuIHxQ1DAzn7WxsvfMROA2T
zrzo6p5VwgXzYT7nM/RukdE4N+NlXp8TEZRBqypDyjvMlbmvChd4LoQCuTPgmDTFtqAwtVNve/qS
oTIHeYQ061laNO79Zzzfx9eT5YOUUkor+zYMc9+6vgvrilgKjfw3cCI5OqZLb3Xj3ctzOPA4FQue
aVU0ceObI8IgJ9BrYUbSQbOt7IRZ5OQ79+rmTnbM497lN+YtkBp2n0+3NofCVAh+8/7MT4/Rzx0I
Th14+kpjBAdPcbeC/Hql9UWvaoUHjbWfNP4WlNdwhdR3KH8h7sIlvt/WCYYosB+VwfuszTyiF3AA
4CVjzAov+OpRzyx8D6zK7jcBrIqRhFuP2dycrjlKmfkfCLiLE0BjYiTErmyowMkgFp997G25B5UM
4ocJT0priYJsYXbCzm3bZEVz1/d2ASXCIUpT2gDtmEzZBCGcyVwtL6jmpEkmM5u9ef+KCYbR26Fe
ymWW/b2nJ3udlfnzvtY0m+28dQT27FH9nZUFLpDERtxrNX2r186TBe5BSUXVloeGv/BaFB5shrYW
LxcPzNIFSrvOVJ+kR9YjdJuhihpGCCv4/lILapIhnnuRa3khwCSiE99h1MYVWHJAQ2u9Y1+Be5yg
8JWXFv/PJUL2VeyDC5F8bFu60ApHu5OFJ2vDeTnm4vNhaEgdXgSwK+5Ie91fWR2nnvcsklFbL88E
aPhCDTWxbOyS3iuXsf7aHTbTOgfyp06BbGGmP2iCujZSd0h699LaBtjzUEhlWRpHF788MqI78NzO
JNLsnLJE5bylnpr5MR4bvMsW5lI6bSHcwuQryz9XWlzgmj8/CDFIMIYeG7hdxKsqtVcBx2v4WI2T
/Z11PqQeXkrr3SI0Gkq6kemv+d9Wn9JTjha4jgA971QljH3hi73oMDiOrRlYdoN0mSPtzxs5LeaS
A34ANtAfH4VhDOW7MI4QlOBG7dA7OICoJkUsQ7s9Jx5H3m1VEKnEHdH6RCff2tBvNKYU6n/oPHS5
xXJWdMGuq4aytcCVyemNIf8bU1FWOr39sfLcm8HUiRDlxGVSc9L5VLGX8328QKH+UVLaHZS78CdL
WNsyQKsajWg1wQH5Ba0SWZsgaOurFaYgrisTiotZtxdHqE4YXqC/efVGxyRiOaIVz1v0jiC2i9nv
c0fIJ8tOQmH43BOQJkZnJcP2UU7ltlYsV1onvBAd2ymI+dfKunY3ti2Pjn0EXRzDPcK9K1kCqJor
BEyTludrNJnqfns6daEsqepNNLlFFhlA/zSgKdPBel9MI8XvjW6KhNk6dRpdA4eEKkqOd7vd4Wj3
Box1uxtM+kdpQ2Z8+JldSYafxpODmHuSn270vlawHbg0IZdTx4nPGrq/DWvHHKQADSdcIq8aPXCx
tB2crUDzVt4qsKu1A/7a4Y78EaiSNDTTY8z8OkJx0FTD4qSw4LwPwsNxORjWJfVYuQ6AGG3JyGYh
HQyz5B3zy1Myjo5tAPor97AY5nig5Aho7knmDOv9AJN5dKah7/Cl6nmJaVnLqUWaCVChibtzGFUs
CwHrNpbXA2D8wIrYkQYchDODKGYWNiB2odvZU3xzT34ztqD22ITagJOYB7ApZfe7/eMp7FPIEgfn
xjiJJvVnBSsy8RA2wNO+ORGecNMyL7F5KMG8qfyyhXtESWn4ldpvSk/nxC+9wkkQx9ZPwnYUoV0W
vtbupPc10MbsrF2e7xPeBy1diHl1opqm9tPwu5DUN1Hu4Mfh4Iz6tdrDUoWGbyXI8gtGUBQkn33D
51bv3BotYAkjVC2Pj/5WiRaoTHu1Cdqeqzrk0MdVTsl+giCiZE+BM03f367HCQdJBz3KLYb2jEgi
Xaiow7KaE5nnLTTmOyJAA5eVI0zekMkmExCUj8iohnmaXwdGXMhULxSASFPel0WzX2/UF5AW9iRo
jrv0ey3jj9kkwOMXZPliADZJxso1W4mdBVw3du5XzXfN7SfSrkECG8azCxlCkGOaMkk0Xbajblgl
Tw84v4++rxd8FjXP2QLVpaSvFsVLdqxI7wi93goE7xp3IkXHDIPsaBsSSGqRQaObGJnMbx7jyW8E
euGcrBFb0ovbf5Fhh+cGH0NqlPcnkZUqgbg6iWYKu0CS8aU0f0ZxAezFv3KNJ55eQNDw94TFTyEc
GMBhiIt5QewsMbfcXPlothXO+pNvxoAMHLoc/kwwb8KQFy3Yh/QRI8987QWkU1UXT16H2e6+wMyZ
jSWf191QAX0t0YPo8NM1XrXgnGX+IdHt0iPRBJiV52KpFTWxJX+cjjsD49qU/nP0j37EYqSCjnvE
/4zmPJeuU8bM2uGMWFJdB8/fb5UxfuQ9ZKtrPC+YgrfRhBACe8fxQJ0s1+pGYhmkBxyV0uucmT8U
nmF+12EpIWBAlqgJLLKt8dsSA4k1b0z6FwSQJwUsQ4JQ7AfzoCm4LboW3bNxLPGTSI4Y7JisWX7y
SZkB2GZzqc7jmf+7sRfeupt1Ms9bSe/SY11iPBIinfvJIxKoEWbJy//G7/NeI6ryNQao9FcdDBau
ZDIGH9TW8236ud+nZ9dp0qU1FCMmpW5fAhYAHFet8EP2c8jzWA3dxFl3OmGmoYa59y+d3reguvRd
bZgl0cOKf6lesyz4T+NYF1zeMES8uBDLB7eJL2R6xSDBII/w4gqP3OguQ49KhLTtJOwsqU4oChZ7
oF1fqJV6g+1Cf4PwFeZDiimNKj/+QivxKe2lS80EwatTfqLXsHpSjbCGa2F6eCBU+uUHgvm7fyc5
RdCgVEIK7JUS15j47IbLQAfkO2URDmJnt97aTHL4TYfyfSACKtSytgm619OifMpgJSE4CoR4a/WO
DS4uEZeklX9O7kUZghYTY95jkLOvIXGiRZbnqap8T0OgoHzESa9Aw+6GRKcQgVyUXOE84QHs5Wp2
sCLUPI2tsNhwr6TozOwEIVqbgZLhcv1NWn7NONBPkv6E2uVE//Zd6bH5olzwa25G0BTyrWppTZ0a
clDDUb0cvQvSzt4lmtidByB8C6lDyUsqvbV3a7Q75VdTyS18qqcToXnvzfWnB7zEiM7lLFzKcFcp
a3r6dIpiKUqYeSAfMAaUMK9MspObRV3DNYj5eYWecMB5ZXRIBhUbmkeLGW4PLeTuz+RLHWGpJFDF
X05hTv9vEH62JBHw8kMJK8ZdsWMuC8WH71+aDLY1Utk09jzmwbvIBV3pfQodMoSpW0RppPluLeC2
gyH0nvPLEIe1ISehLuVtHo/+aAa1nOruvpcS3889UBjum2c8m7XpmhENKlYbcGNepVmckVnbkN0I
VHKb3IWXpisyzlG3ivEKi2wXtpaEF3Cqpzt/4VnofqT7tDn2hD81xvxZ11OGo5yhKMTvq/Otwe3e
YbLW+2zlXyCfph1MFuIT4E0O3EsSq2RpzLTgzLNov9uAHAmRxHkBo15HAaNYHrb86hxXs5QhMCH7
1Dh+qltp8NTHi/rroN3zEOhoDj5Bp9YLpn8tmj0wGzAkh1agEl8uIkAe9Ic+xpFgmUiTEOT0gvMN
y93+vl3II3eIUNhyCtvXKqPre9iT8j2ZDa50QS40IIHryi0Czfwz1AA/lYyolBIJydL5fQfyvNo7
ypSLy6yHQNAXEnt8NHZVXL1UH09rZCp9BbLmGyge/IvjRm2am26ghXsiGCHgZ/TjcxlUHOhBpOMz
tj63LMVs1b1cezATXRnR3wsdVLSfucYot/BfxzgyUfBLia+uMc1pKpOxNyn1BZFqXd/ZZssv0PTx
Us52aJ9FD/sKH7Nmdk0Pv/7QgSeijAS7V3X2dEZ141S0MDmLIFbDTRyAMXAgg2Nlu6BQSSUI/nH7
V+1nXh76bemXmmdpT2eH63qEt9xgu/mo58vDMbimdoCV4NwOVccUdJcLPpWTFZkrGPJHVLbpYmM+
2Wo5WFjdyFbVEstsRZM7GubhN0RvdztNSMLY5cpvJFKUZ8OvDwR6J/EoKRnTdWqPCgbDKGlwdEdU
8tiGUkh4kD6jlY5vglBXXkVoxLE7Du+ocjSlpqyCGrtQ8nFDzsf3wrZ2aE1/Lu2j5RrihUuF1Qfb
bTwyEJvPaRN3wVp/RmQEEw9eK/SqRo+QpSU9FUUjwO9FuHH6GGR+U6MW3780+5HRWNASr823MHZr
gjgvuJe/dkZQB2MeQjaz2ynoWwf8F0TcN8wG375jmQmjLA5cSsbHpwNhRQDoY2WEOT/xHWGOcK/1
lz+VX0jHORm4uo8PMuccSPiFtXQbSpHilZcrsVDMMqgojXhrU9PJ2scysZ8YP11xUbDy7Y6K75sX
vOnN+qsrmo+wCJG2mamwV2shJObUDHpXMSL7J0CJVZyQflBBpHwze0VYkvfWg0lQoWSNniCcI/CE
07mOltd1ar+SVTpPwLXvwxUNTND9OJCMl8PKqXfKTd8c97BZvVmCOfXbCPtuOmSBbzA0FMubO9kF
fz5wfU1GjwoAoFP9C3R9hJAHk6lY0ZzcOi6ctpQY4d9a6rBAkRoe2Gz+gncJP1A0MrDmM1x8M7Rt
vYrQ57HzDhZ2dFBiWnTKA0ZILCHumc8pbFGSDS66xcRGvedtGGxHV4OrotvnB8h18luO3nlHgo26
WlPBZSWEB29T6nDl2Xq5lTAM5w4clbz4kUKDoe+dzt4eKZcalpphWQUYQXtYVRFpihDIw0l9tA7a
K4GjGJvo4FLuh1Na70BXWJvw8060MV/80bOHr7YeSio2ROGBW4Ny3GKYqutG3DO/ujkaANstld7Y
EaqMwK1qaG1Sg6mkOoCuCzdIxupuKoK6x+L/jTh2Wqap0ZJryZd9mde6GYwE6ajHBjHlvhyYapCJ
xq8j9GajKFimIKZWaYGYwluInFyDtLlovAKJ8OwYZf+aHrpQNqSaivHI7iPPAGYNPMJUjHsSm6+a
0T4Bt8jXr/Uj6mbnONK72sKTbKntqK19YlzEOZEdiXr9bssUQuSrPKEho1VsLzX592lCt2GSemcT
Z6p0FjD407vSCFmjMwPtMM6eFu/IosYtoC0ktARdXMR827G0g52RVgriqgd0xFkQr2rMIqnqQu8s
o3z5o+pauP0hDgugijaTSqIQL1h1uV7/uc8coSmPYb0YMrt+yQdPrBtS61tLh7W2161IxCTBsqsu
0Ul3OKUCn2mV5E0GHRiEWao/eV3s0Zes8cvWcfIBwijqglwlKt6dkiJyAisYhYA8scGG9yhe7J8f
AztkBhN4yAczsMe3h94H7mYBRmyvKswkEB8n1f7+3XHlqqpsFhuTBCputTMAOcbVAFK86LQNZVhm
vgLrHrVR0UdbkdWL13KHdPa+QiqBBWMmm4IQfxGB5s+yIEDvwh6sqWbcdG70J3riLIsLuLF3eyG6
AEaFZ1qqS6EHHCE8v93a9DvDG8HqEJTE0vJWDPe3hw3JX97wkJesYwuaQDNb8Lw6mIO9kRGZQQ0X
KrRdqBOC+hXqhsSJEpWGuwEfTbMgeGpTPDzMyxDKpZ9+lhfN/AzXj6WX0UKq+ZtXi+AkJyzbfgUw
/hJ0Z+A836Us5epvIEyHznbdFpwANOrHPJCwvLtRoc2VRxNyhgFUrAi7UXvgQN1aiiVny6Nawg/g
5FpGqqsnmRLmuTOgY2m80sQ6dljvWwo8upLd5hPZPhGumKMbhzdZNHvJG/w5kZQLadynRnM/RVsV
fn/EgFJwP7vKHJXN34IcouCGB+bdbSZm7kWwNzjUzlxAOPq0oyA66sbpF9EZUipWfoMIlVzyyeAr
/uVLp3F9ixiSCiqI+JCyZMgRUhQB58PUxkjEZAroNAh6Dmp4+jjz/dGVe2f35cLw4EHc1V4hpREo
L4BIbtO1YYLXcPSJCFYQCh/3sRaWgivKGezSfC5ZHUitBcnkxU7xo7jH13lJEaiOVyxWC/L5tpur
aFaJCbMJ8eXHh+4QNEEIqVu0yMOuU1zd47N6cER6CSU0ULpKoaZuVJ/NTgSYyXPqWlGhQzO0sAce
kWGxHLKRznyoPmBMEspprsrRuP9AeGC9l9VjMfyAq2/d4fmc+VsyMkac8O58/F+hh/1QL9b1k56U
NVEtak78eU3jojVsYFPguhLMdzTcdQWw5vECOa+sU2X+sVCvykFyhJkC4I7If6FDhUcqNLL/swPm
3GOpuAno5TCu/hh8OPX0vWOOI2jPXbTtTs6bekbLwN5Ogga3fVBvtkgZeXEfMRV+dBEu6uS2ETrb
KIwjvBQsMu3bq3e6seNPY7wVHlx9qEcXneb2ZdShWEJCTGNZv0iHJL6/xGZa4LhUUMJ/t0H7GOZE
FNyNDSaiVxn9Dp5KV91raVZS/CzpgoHEPnTzph4QTWPAb4nqbhNUqD8W61EtscBukWvc2uF7HBVG
YhGld8Rf/ZwSCet8Cp6Rx2GUBeqQpUtF+8CCSOmRIeT2IzJQ/mLv3NhfiSuxXEshMmWrOhLfl8+N
o1SVpd58Thysdlgy/q8mS+4nceCiWFTmo/TyGlozsRGkPgNFMEPrt2JaT5KI0je18Ke3K2yHpprW
lepg7Mzis2sbLVQzgrsYiJJPwutmoK76H+S+zrfdHXz9vgXqozPbPbL5L3jsPnil2U1fsUrsFnDY
3p5MJ6OrxNGHNn9tNxEqpcMYL7gqz+CWrxebvJwNAWO1Y3krjt0rkC+yAi/yaFgTIlDVET8x8nuF
q4ezMdUlmO96THzqLfwKoI3DnLnDQDLjO1W88h882A1SD4wN2VEq/5/vRj5d6PH8ElPID5GYJZwX
/ypK8r+qvRCBA3wzKySgzv4C69yT1xuXSK9znZzcnkzB0tLczREsjOlWOBQiZRUdiDm0XsB21EBb
z/YbZiVCrGJ8jIr2pfz14VYjaQqF9znHwyGbIjc8mZ9xIKpyNhh/o2l4WqR/EozTKokcL/dFCpKa
os1FXx2JUz30NSnCVdKBfbnnPiJb0GdCPwO9QGP3Ew0KQz5ggS5N1sNpOvCssvyIYM0ohEiaFNdL
tf0C+V2cMK2V4BfHxBh47+Yv8tA3FBFIreyytn9fzATkUSDBHAJqvtJwI/pRtNZXLmB1mzvqqWdA
yxcnpsCei/lBiIv6l/xGVX9hfAAnFf1kWPt/voCI+zUKU3SLvipSAqPDqvKenCg+d7Faf15yfTqJ
c7PkpkoW6/h9pjYNvG8PkAJ+lPfk8M36AgtKAkKdRS3M39fthTH9psUdUD6vh405vsTz+4s0Mlbr
gGRAeazTNcoC2oymHy5MOT6Umfjg2Y+piyjU8kPAw4ZPuQlaL92pxIuNZmL3Fw3ffkQGTdOsLagq
7jQhQcWbSgyw2jIJle/j27kV1Vgp5bfggMI+vff+RqE5SuC1fOS+sphc11PNRD7nc0ACQhRseDas
9feWKjwEipcuzTVWJv/p4k+YZLWHtJF4VhjIzz7x9XttIYznN445jG8vXvcGUx5AnWDYahJvl+Fy
KzaSFLdeEYQ9s4LF0shF5m4Fj8ZoNo0GAAM2PbEs4zp/TES+W8JUaysWmhnGln9S13ss2FfW8uxg
yerGPyna/NW2eq9EEHFRFCWdYtNEBB+DdvS1MkPRP4aCsH7Ypc6XBeS7Y59iGtGAJ9bqhzuvrQXl
naHc/Fz8JVmzDWpAScDqh9kk+Gu+ss70P+mtoT/RJ+KeoWXhuBgOoJK93yOiFI1/M7FgMIekhqux
WFmMTwkUJgLhskZn1TgJNvCFkSDg3gEk6qA+Z/S1Gk3SGO3flg5vonvatA1CH1v5c7mkcSn8ltFN
27Tq9PhDLxyuGr1piI3C9Cho7x59Mq/e87P0w05VJ2WpD3JpuisWeVzcMF5HvXYh/FGYeo9PTbyh
Dct5evp99CJENTqt8mB2Z59GGZyv0zDy7tOGh+rvjwGo59AHo1empswnRSkldZclRSttUgIVBfMO
X0OOezDm0AgMlhTRenQflPLuYK0rI0u6Hcf6QOunyvyIIJHireccM5HNVGOR+Js62mEmpdB7vZsV
oH5T27KdDfmnjBpVQNW1oFbmZCmVZNnvFdhkizkcmSk8zaIc8LKhZ+2x2LdTT7sVLM632OJEYQQ2
9nZ9Vk9VdAboVdgrO2ySXxHcatuDLMQusg6ZqNwgtYoqaGl1fsxIihI/nMmVmxpUqWx5ic+iw9Ls
gVLpQQxxVhZQFexKcaClfyd3AhJrYL5VDeA08gcH5hTjXerHOnnfEgNN+HSPPfEm+LgltEzWfK4k
R0U+MbZuHK9A3N7SclbCQ5tqano9GZQKYIFIcLu6VIr+Fh+4YnDs4hnlvUpvghBLj3xvZCMFAZbk
ch0h+vhlUjOTrmZ+9Tc+IozCkDmXyomYsFNduYhxD3kmuHLaRWi+1892QA15ROxIsWmkk0IhPZKq
2/43C8TQunnnDj4VpWLTRZvgyUc+k84xfz/j+cQAzXUiHBPRF/bLhTF7pOyVVWRhX3VaQytTSvpP
jyIkYf3rdg0VZrS8rhGaubxwStkbT9Un88zEwfL0U19EHwkWYfMQeSmzB4vHJMAF3rDatyQnb0ln
PhhF8q2l/tz9HvSW1Xg8EhnJcasKAQtTbyx3FGVqhW+ovHfPIttiCgcn7ggZfvGZoN3CDipIXP57
SCDk7Q1U0Gzpz0qt6zwbw4jDLy75/4FbY6jLbgYgkgRxwl/7grfQtRMO/Dq9sgJEm1zBLaFlBodW
sX2wIGatzzaZDA6hGRanLlyzBv+OAL0lLFqWWMdvRz9ceDSk3/uI0+1dw5ST1t9mDxAueZk1dBu1
g8ZkU9QbW6VqOnkTmHFYHjywhoGSjJ9rg1ZAsvOKYPbA6vhlw6+NOeOuc4xu2vfPPBRVGzZJazg8
88K565vmmNcNeuqCiqzPKDejNNuxCVMx3QbH+9ocVHm1TO8tyvKLuEZm4y24QR0adKBRmd2FHcgj
1zPfsPgZ6B+qKdUfLu7482Zvv2R3TCvFycnawAS69jBvi9xzXRbJZ4B7+ZkBlmKXdrKhtWbeUF06
N/SnoH4eNdvyBVrl0k8LI6Zmn9D80RfOGgYh4u4L7H0dMs06MS3yAXkNQm2FT1BxYq94cpyCNphV
NqFt/LRE7C312PqHMq+Tzq1TDgGks6i8va6YU2aIXh3EkD2NVuVbL+6W4mM7wa0WTe63jR33IChI
l/KsNIFcmck6rataWr+JtiHWuaM/nBSz+S5cAzmD6L0YRghZ4oXY6x5l6IK1WbKs+bfD9FluQNIh
/n2wKdmQAdh5StLvjRTZfYGxoHcEnd91NEgvnE8yzz8PzE/BOAG+dgjG7RjOqA6M3XnRWDDCcEoe
5+YVubb5YbO8vxzv023z8eX1NemhR8Exwu4BCW4kEUcglw0VZJxv8HmCnwgEUrK96C5c6SW27iWV
IYD9uXDbAvq9rVjsuke21QBGDx2Aaa67MOElO7jnmx3bdWKUjEYJN1YjVf1RY8+Tretf82dqrfpo
TJiW5rjsfKo1J1wpUgpHhuR9ceDPLQqKNN3dbhXTg9NGeLU7BSeGvW+ie/tehtZibJ43Laiu7I17
VPCG/Ug54g2nzqx7Xk7RCTZMN1pxrDtGkvInVeRN/BlN3ihEozCiv7HqCp0avEalXjBTo1Kx7VNo
ZPLdTyUBCtxW5T5r0JKz2Wb6CJ8DO/Z+FclSL+E3UsAiKkcR6N59xymhvdowi1d2SyB08KTapxw+
UE6UiIP4IfqJEr/CoJsp6Zhgeez6KCprrLjk1AFKMcj/qBTZgvKfhw866M8EzbVUpZffKyY9S44J
k2DD6lVDGFDLubYT908dQ8jD12c58asEvrzqyO6rWV7AVBa6DqgMwGi72Gyipj0WWRioHZWWWEBs
JHQbm/Zf6rjpOf9ljZ2UyATqzaduZxyM1T/AsRfKfNi3H3JTFD97EoFYfysPyOnIiTON+RPojpqE
p5NiIa3Y0EwgZa+47jkZP0laD9dyHqMtRrmKk+dZkQpsi3TmGU20IHPpYWCdkCuqBfDhfVpe9rne
oaPkip0e4FrvB8xc+EFY/LwFdcaJZpzX6SQZBoNSRnlpFuGtw7i0f/432OLZer8zAqPWPfqLrYGV
A5MN+9kpgKLhYLdv009/FxbLWw/53huQFyULZIeUOIDNti13drfJVrnJDtOfvHFgIyNaKaU+Xq1z
rjzOn/Vm8Jjs7N7O4xn2VoaOhQ2pkI3PLr3GT2pxJdNsfIRCCQeRJJ4QRjzCgI1pRXwGufDJiXog
HaI1qr9ma4egwPaR5izzshD8zz/oqm71VvEzDuXk9v6eROxR3t0oPmgC42O0bJfR2SsnDX1uwbey
vDDlPr1fgHtQ2NLZOVKmfbzaH3/6ii1GmY5p6AXu/5HkpFgeyd6SqGvEdamVPsMKZAldq9ZfhMXk
7oGLuMf96vDJt0tHEALqRbL+abqyguW8eh556CjWi9AUxHTDaekn6S38DkFmvWqrKmpTzBU82JKC
zU9MD/VZhhcEp5yUVbyZmfQtulHcXF8/yqOKL6mCqTD4axmm/Tkji0tY/S/SJxM5b30Pjg5ve7UP
/gDKjC5sKdVtkP22qvKm3Dkdm8VAeGOb4MMof77UzyN4o6XLI7AOYac6JpsqIjmN5mO7a7cIGqa+
NqBP94Bh/jR1oAwFuZnCb8JjwMqvGfGFCN7yi/1AETpe5VqZbFWbd0xmsF8Xh/wsl+HIaVGyiFtF
Bv/BFmv4wUXLbZQ0jzX8loQFYTEUO8PrjDgoqQiK1YGwSmOdTg1su1R4Z0DcRZlKQf0gGfqyS+bG
2vOP7ApUtDfTKC/coHWFpp5fKSWUe6OsCNMkC0n/C559lIYJ3ivpmGStz6WufsWYILaMci64+W84
ye+doSNmQEfd/wZAFjCPpCCD2Cx93dIpZ3e8h+pucLrr/z/Re/9REu12Q+Enu8+MpukGsAhJ9364
Pja54tOoM7K9B8Yvx0Tqkr3u/qWo2NJm+BPR3D3mpfvbVyF3wWoYMPPYnwalz1QWjcSuI7Il2ytC
HV+y2u8Vu+72JKjTjYOSw+GrLXgM4Fh/09lYSs7kFaXx6AtvSrimEZ0auFAg9vAdvLNHViVGUmC2
LdIqIUBG6ZW318wL6uYHJy9u9s7dzaguFIWUm4Pd9Y6qrALkuCE0PqysdkkPxYjsQF1VD8oWR/P4
GxRhQlWgHcQqYEy9IqeCReABfLmszTT0I497DEvs9pU4vz55P+n+Wdb4xqWtTcNorakNzCukbfJ/
eF3h/qDh2n8fn2tTOjR+dq8B3VCrnGKU3oUdd3AQk3QnGV7q9hGvKiu5KE5Jmu41E/Nka9Mh4lpa
NVlCp2d8aXwFbLz4ECMjrbiCL78ihLRpFc1m/xZ26a3ARm1D8RqIgd/mInrzJX2xtj1CfZ9SL/As
hyMnmDHULQRqTQacTFQnLwfIp3qWrV7RqtPiEgW1rb8wKWZVZbJLQ6I69C2J1j2rLJHIiktGcpSq
ku0NnquYVevBOVWxTv6QO9BeDMhWdVQMH5mzgO2ckvlYd92NQ5Q+ABx37MivtrR+WQoURZU2ogqF
t6JJvtiKWT2qnjwSCrd8deuEldDHXJNvNWKij5raLPI1JgaCNuqyIff9JOGHFCc5tQ5UMHrJEgI5
nW9FrVKfPuP5/Dpznk3wjF2szGBTTmhitOQZZkIMg8p2PbQlPOMX67ADoRDrp2Kke343/ZjmC7Vb
4t7jKJpPswXZp0Iv2d9BKPNm1N0XGBWH/BfpD4dnTB8eh+Ov5iEjBTQjp/ONJCJkbmAwiyK3kMTW
Jr7A5bLA4cE4kqZJtPyixY3FFleU/gxQDz+J/ku/uLJEcI9HIQojvrOKULDPr+lyzsadrBAByaWZ
vcyGJYZqwy7G6VSWHJ4635GnvRcm4N+DCUjk+I2gxaNadKjnBVGr917DzoIwFNOH94CM0gXlAeZ6
aL7rJg3d1XqC4f9VTKmZTRIDSQhLfVLPs/YQJo6E/2JgBGrrPAriTN6/HGWho05JxYQLi6FtwGC1
TqQyyNYOy55bW+viU5PR6py7/Hqzur3SLEfPoXDypO9Vd5gBvGiP4sRVkXLFwWnmRoobNKcWD69V
9NEsAKlhqccYtAbFalNwrYH/TsLWnSPVAbc3ErwRuppr492iB2UqFktRR8B+8F7VdVbe6sfOLXGs
s7jz2jMua2nkyXP0IcpHC1jBx1btVM9cbehdOrH43H7HTMVfc9jslwgFAN+D6r1IAxWv56oTcTAg
zIrylxAjRy1tqIc7RqsTWsiVm+jaCJVoBVvVzDZJck9/WPpL7maelJI/V1EY5KfsgzYW0ZPT1RKW
WSPv3D8sq3bzQpU5+xyHIcTGtNyZRHXXXoYDluPrWawt98bJNWh7qLHfYE5VG9EOyxTfGVIZXw8h
0Mpq7NUaW6/r0Hw3TMa1TFAjvKvyWosdxQmfouARDQvqwNm0wvxwW/OEo/eDif7gZUA4DCQQ+rU4
Rul7n/FYZH7oFUOw5jOGrWUihClv7a5ytrKYfqnkzSnpflI2r2IkEx26IlOJxj/siMCItATFzmzW
x4bebHh0OIYov39G/2qCcBjtuWbGnIXPRmEbbV/EeJHr84yQ2B6F6ymkMVSVB+7ZLDiHJj39vZsK
Km7egddDzyrSeafReRzbgZxfC/k2X10pkhm5GKHifqNJZc+Lr0LU7PswL0GgERThEq2tQFyo08YN
i3BCwiN/Bh2LV2NwAypw0kbo8XOkfHZ2qwVNYzVkhASYtlx4XGUwBBlnQNTX5ceLVxs1E39MSUTP
KsQjv3X8A1lCckuEq/PNAV6km0wY8CWBvwvO1feK4pIvIQGAza6nDVe3pIWqjPy9ZGB0DyQud4VF
edIlgbC20zY0++PmYWVxJesrxoibWEhVH2YI92KnIu1K10SVeVfSlPh7P/m8YCvkJUS4LpI3w+Jy
OXBwzu/E7t4TCGlc9D5lZ460Emn49j7n5aJxBrVXT6a2Y461pJg8kU/jwx/fU+JTkVpVQyKDvlWX
sX8xHiGFnjd3WvcgETipuXw8rE4KPM8DZRVNRqJXOwpqIeh3yfhGnXeHRD4FwyypS7ctqyxkYc6+
p30JHGNXlOPFGYohNcTEUHV+YHFbaN9IijBTy2HGcepQ4nnD9t9TSqx5zHr1gJB7r+Z7iL/2W0Mu
IrH9YVTm5f7Rd4aasxNAAbn8MHNPoCZg1QtKw1Abx4E/DfwFOhChX3Bip+xZ8dh9ukTdMJsRwEzz
fCMRUD0NNG+QlJP3lsrVqGtg8cyrwfxPwjE7J/g/w7JERZsBXOzASoLTJ/YruVLUvDPDSzgt9KeY
ncURyRCPsdyNm8wHyVLsZj1SQ3FEHKsBg0ZG+1oaZIxJ0lv+ZnhHOvtDC/qHy5sV69a6yWekCyg+
Rz5i2cEcvtEsb5DOMgaapNFIBwL8MtHOatY4O/q73AoJG6z+xLekXo6XyUzmU2b9VQPh9M4wAuwG
FAyBQvk30HLa936c9J0RkQyvXGOJAsjQLpUI9WhaUJ1RzToISFfQIyxwOzM22tpHpNyO8P8XJyQ8
n+BYoKgysfUOInoSGSSUpX7U18+SxflSgRCdlhAf++LtIH24IRwpGpZjyBB9q9K3GFdp1GjZuYtk
n0sFlfJGi8QBjJvQPvX4JRUXZh1O8LkCMHrRBmrjsGC+pfcdRAlCQVKHftm2vEk8huZ1T18lrqmQ
usdTGPnbnt5fdyrviUpBrRbSQq4FTeArRZDmUUq6ZqhtUi2DYODGNfoBRSes6FN+HBRst3I7HTye
kEr8WrGgH9s7oSPPBnnpTmSW/caUHkuaiS6PzY0htNc6drSumUIyqEZ4vMWC0RWi3Q74ImI6I8p5
8g3GUtREJ2ez5y2uH18f6n+5hKW/wD23cqYw1KzuU8XEyE03YtqmHu0Ou7ulDQFeAol2dV6BKweh
TATOq09AM3JECY9lloALep8lbGDJUEpSeVNgB/tahAhhs8KpJZiKHV/SGGdE9yJXdprFxXhUARft
z3+8d+LlCrDRgVTLjQGBMuYETJe711H/fh3Va+TQuukG5ilR7xYROOI/QprEhKCb0Ugm/7nP1OJh
LAidp1TD5tl6RCfipvuv3G/HVBDJ6ha0RvEGEh24/mCD2JHrR7sk40DkUhwQFwPj9Kebl9MUBXjM
yLtVgX73x5Ha5zHjSOpjtRunVG+eJe9+xyZeEceHNlTxHWT8D9YUA/cj2ZcYvfDQAimQlQFAE8jv
4UK3AzKt/i2vPtREqSep4hZSBMvZdxqhFP2ANdH6kWPpRW13lazjNter9LxwllCbsQIJJy+DOtoa
MkMV2rZ4Fwset/LpRJ6bwPVCjVqWqATACO/gUB7s4IXJwZNSnSk051FMOEvLTld+9BXyOVYyvkef
9N7kdgbCqmo/eWPvB2hdPAOnN9OJ4GTZdbwEAKFvO+8LygsAUMA0iM9SQSddrNg1j6k+OsPxqAWQ
10X82Jqx+mRWXgRwETDYDlrhtNoF1DFKF4ci8GPmNr55TeJfdPhtDGrkUDbtBFUU76y+1LKa0Wa3
BgFDW6nAFdw4lCqDtQkSJnUx30LGAyQQHmRvYGUjrtd0T2D4z9SCFjf6R8pXEqUM9rzSPG8UoEb1
WZk/y+SEvTgZVvrIahlMrj/HXDvLehDbHFwW6q4EWDZxj25aN9ffLnscZS2IPLc4LOQtGK0BVNMF
N+fk+kGqlZVcAAK6f8ntvpNbJ/cJU8fBwiXy3FeOu8PI8nOIk58lUwPDDaHxRPYTlVybvayUkibD
Rh8pIcF9gQ2x84q6eXYkbkqj296m3i1Ww4E/+zmYr+pbrBBP+2NIS1UYdlHG4xX8vJK7DUJYHO8y
JBHJN2Z3TifQplluxFQwo9G3QWzuqaEzkeTEUi4K4HjOkJ8WcwKRJGkICwQyLUIcDBdgh/C6ui7f
/NkWsGy3fyzGCVdimsaDhnJnqothKV4ETrx7o8CCjs3bWMbHhnHnRtPZjDGv9YXk+70UVAnfCP94
Eb2AVnzZPDie6qY6BwYRArILVjYlrx9k2Myeqgup5KeP4NcDgvQyWpCCXbDNocT+ImnnTUpCtYE9
c+S3uUlubM8hmvymRRFgVHQVp/mPJfzQdQULmBZoYcl6KH3sl7QqSo8PXxAAHLqDuKwJggt4Pbtd
Y/5jdgzyIl4Ovllk/S9hm98O2H1qNZJfOSCa7AGFYITPQiF9D+mmVYeltbAVqH898I4aVh6JjYfa
mDQ+RLedAsXa1rL6hZgHxpYhGzlQrZo+guecBlPqxjxa0NMX7LKBV87vQUXVeVR1updccH/Gp4Ms
LPY5UOmtRWm4ZRYFbNW+KmiYwre/t6QKMSQnMjIr9AKWtJRyBe0P38k7v++2NZ5zdCE6JeIkkico
ntO95lPFtXmjyQFpbmh+7YhSmoNNJs83A0JFX2vULSPlSwj263XIbJl9A8FxU5gZfHDCrM3VunZZ
IixrN7pxGZ7nfX3X0ECeux34XX5OadoQplI5d5EL9H514K+gVTs2byDQ5BRNSbl4Oy/72ywti5Q+
SFyicAqFdfeZFtQeE6vQuM6ZVRfFDJ23B+0xL9ZXoB7ONBG8yDSuEfJubD6f8UEZ9RUYGyGwO0cE
NNhhzPkp+1/9LRPv9RYnuiH14DlyCMu+YEdM0jN4KT7DNiFBT5Lr24oyb1a0bcR7RsMQoRS7qbGv
2ApiSiEWEFFNOKIWAyuItLNdQNfBAbCp6Rbeoudt5bCejoQwq3y//He8d9jd5Z5gYusacFiJCgcJ
uornrNvkEJJckS03qr4ntNzccncmBKc71ZFhL7REiYw+B0b8mLEcMozlDrRiEoqU+VE5KnUe70sX
qHIVc3SmErC/Xe5du3y+qyKzcUkLYZc9g82zYz02T6oVToA11npz8WYngtqMm+mxAlhXlNOZ8P92
MBaPppE6W2fH2RDEpSFueD3tyqVWBv8r6WEDQ+TH/TJXk5w7HwECbRBtrw1M4DIEs0A+auR/9tBe
QRR3fgKGaBrZ2MtJWyMxM5ZLa+Q8qO8JYOew6QkxNLnzyFmCzih0gKodPnkqym6n37AzKi5yFHSy
V/yUB8eRIMIEz37MEPm9+hFDUylBRBCCtav2BvSTfnXzpoTYBEwPiVo988ZIpDcd3WuK3ABF+U24
uWNmQAh+lL6aLpFPQVfq+u7gvh3N5zxA5HcoG/hGL8Od0N0Wq0vZ98Lysso4BkZfyEm1OP6VkMGF
8CtpKSrfBMXqhAs+PQgRQwdjxEwUl0SA38DwhXTGWmMPICdW/XxCxYWZo/gwNzVE2m15Wja8HF/V
lzvvAgmEepije0M8Qb6wlFBaIUVwd/qzE+jVn9j+UZRpmlAvOt4LBtmPcVz+y4dHYRGZvxSgaF6G
M4T3LnZeKlui6iCyuX7TPYe6S5jyXCpJiLJP5kced7glzSZkMdcACZhULp1yxiT97RnWsrJU9a7r
JM0phb8HHY+1pKNCtWcx6PHZmDGAU+bkyez7ZkrLSiNd1KZ6d8NS9G6C2UzbM3xZnPo1Sk09VijF
fQFu64mFsxxw7fW6DiPAlfzgL8gOwnaEl/4VO5ol8cOYi7aH9L2U7jH9h9b+gmOfXoTWxYhgSmOy
tzgER3YnZABt87LwbbPEgEkQH3rFPsY9hV+6XqARtboTqPASQB0XxsjaOuI2DmHKsbuZn6jJzjyA
tnNzslpvVMjJNOVLu4Wk2Aa+jjPpaLErokaEZQ5i2OsNfM+dQXOq0kZ3ER0ZlNKYC8cQxVKO4zPw
MKCgRhRAAU2kW/j6AZ1bhlKMjEAdE2S+zNb+OkJ7Bi3NUwvaspV81Yq7SM3dC/tLH2fgt+4NTHHB
XkMxVCBzEMB0hkJ4YSjOlEZes1vVvhdsUBLkzhKudMaZyBC6m7sFHBUr1myWWsOSDXpPKMXpZd1H
pshZIbv+cD+P5yGtQgQR1V6PeQfTTVGq5VWwlPjImdKJNAVAblVOD+u41uPYt2RZ0fqFPqgA2BN+
2IxEXIOQAWqiKHrDId6C+qOzWZ3oUW8sYgSZOQtEBKZiJFxtJzlcVfFenLqJpzThoJa21t9RegSp
RpqITIgOQgQi+6QJjhQn+I+E4spkFPlrrqzpIu+XYaBdYG8T99GB/pW1pwRqb0Hb0nyy0VvGJm30
IpxhW8dgEWGJuUrGFrraJ22WQ4eac4Sn84kGb0th75CRJ6bYZrW8NnaXImkQFWFdIYhi7jJKD5pO
Spz6UniL4NLEP05SgbbmofIgYSLcG8ArIA17QGreq0yW3AyVrYUl/l12RlEN9VajAEwhWOUZOt3s
4+nlPSpTj+8O2dn/Rgm5DldbA8YEQ1PAQ7M9+WflMY1OWAkT0iolBAIu/KSs4E5myTWqGmMfISnf
EvRXzX5wv/0knapEyRpQoPlNSOWlVVkr/JG7y4XUhTF5isZBb6dXYmXZoxT6Y3sHzM6yBgw34m/o
CXbqpJ0JBYvrQx9ZM0SoBYNafJ1Xd47S7F6y5YIJBbk1wpq6XPQWxFw4RwZe5jaVdlXjcNhKetB9
HOzWEqnVZcgsFE2srJf3EHdPkFcAEos3fRIjN5LRBItCAGdX0cECS8RAt0zmOCPC+kAvOnlhh1bW
qFPDHGIrwhRAXzyhWhpIiwFO+rB0EZldzOJI28Lha7tFAAy4kBtxbj1E+D5iQ9LZgiMcMuGgbCvv
l+Q+nKuAvXy5MSisACF9Vjozp/iQqz12N2jiLCg0XNGZuUxd6XnCRFow9LIOWS9Uk15PVwEe8RMB
XD8g5qSX/aogaVz6ktYd5mEGAcZ4dBygJJpX2TU3BawytG+WIfRE74oNEJLxBPhM0loPbk2SgKvX
xN8m73UdgYNZBIMWiMuzXvdSgsCeTrB4EV0wfi75XJxf1OOWrWm0zwTc0fh92rGQmHYSfKVzC/+F
SGPAlI8ZwQLDYStUP/TGXA31eO+o2lwgVVwbcOIinUZPP3Ya1I/CkrVMyZv6181VEIbVc/la0Mps
+iIlV0gVpljzhV0knPbSa6M5T/vb38ef4M+zDqaijBWmcFSYALmKYzu9VKNBF3ei2bO0CFTF/TzR
+HMUcJhFX7kv9EqHCOqOPxCYxHY0zqL9H72jw3CzLdsNoN9FUzLEHAGovz4i3NVr/wjvFR5VHTPW
2xCLm1hkHzLGv0rtpnnSZyQGSca002rg+wHn7O7MfO56WpMH9wlXpY4ZUJqC/YVu9va1IXsSVxE6
TFyoCMKWmTWhs/CFksBvnBMHhRQJiTu++7Z6NunCAHVdYXA5Nxaz4bg8RS2MCoAYj460D62aRChQ
5sYxmtlh1+v4gpm0u8bPfvEGId3sNDWZwEA30hTaa3f2a6EycgizpEWTC7IupGdlkEu/6tZIRTUQ
+Qd3zQ09Ema4VubW8asMF6E6Pg/QEfiLShJpiObSJFqVf3P7yAEwUWuwuq2MUheTTOAbMOEByRvW
0rZ3S6zokqui4Z11uB2MUbUD56KQQ4T+X3bn3HsPYZfMcU2yTmWxJ6fqxZ8oCxY49NTSjwBuO0CX
WRKtkhJm56J0URZU/sxDffm3GNQlgWpIzImNc7NoAmXfeo/HxhYVX04rNeZLj5KFHYQVSfv1DD4Z
82DcebbGw4Ei03KPdHwy49vOay7kogmAYc6lMv7VOoUfKl84LKWFHJ9+Sc2Y/oaT3V4hKj/aEG/q
Lsscx8VEwI+JAs7GGBY+w2a6+4LI30hwwC3XHYfIAQrAOL55kvHi2ijbv5TA0mIIjSww6vLhs4Iz
1YutIBVG/GI67aK52qOdk/9iYrPJwEmqbPxpVVvGvmGYogMVQ0bsbbK5m4RN4hc7k8TLe+5qUUP7
wU85mkYoIv7PMwJYAMHiog5aQ0hcXTNjqEEgAVTk35IYDZHA+QaEK17UV6Abok5V/y57XQXjoh30
TRfrXxdu23ya6Zsf+AOX+x021cEsweYoqn6jgev2gAixc8vMyv9YeQSncYApJ37Q8lt5hVNCD9Ox
sCoyDi7yJRqGiOz37LC4l9AIIXkkk+XPBX8buBvDjDruhP+LGRtrEh1TmKygGyP6uXPlDhFJh2aS
pYam4itEqEpQq8nFHxtNqnCg+IA85xvaAFZe40+97APrhlfNTZMaIwKizrdbE3drh6tvaynZ5XpN
L+X7epNHucsfSmTY3G50RE/xeEqHwBa8fAEyx0ATapY4Z4xDiQ1mrB+aKKwYDVNpY8VSWi3mkJf9
2fPjI47bBwf3NwgDq1FOXscdAJZNA42NqbZUWFjxPsOWFqJ/f7tN+V0AwsxosU9JpDDbor2RtIQk
AI7CVnIzLy99+dc7BfLEgyPlKg8UMs+0SQlPduczSl367Ogx49SPm4bWrosJ19Jbjk3DH5B8vrV4
VsfRytD5cKgHzAoNy48QX3pe7zbRag+0omesJ9cgrjAtNLlECvbB8z0NJ/7fBPKXhsdKTFMR+2AE
xXpLp/6FzFhRYAdBH7eEllgUsXmjKVchMjNhSSxbJa1/LsPMVYcpXF+y4bOSaHKgbFtf3g3YDsue
LDUS1iTha/XsfDAzC019tt0/6i/ecVrWXuVbPyVsWfTAl12XNzGfsIa1tCILZLH/+icbP8xssWum
bNrB3kpeJFCr4+TS8Axvaic4KyRhgzz7pOS/L174SlKu7Qgu4Dc4GVAxUPPoM6mJ7LFI+fH4JJA0
AgVN9zkNfQT0FfSyp1IXEtHt9kqXhSAFV1PcWE4SAEtAHK03w5lKJmkBhDH8E8qUqHY6k+qV4bUc
4LI/dATmx1uAqOVZdgrlyPweUqNyDL6e49Qw2GIvRY6Ca9nX/SeVg/JfEWGtbtu8fIhqrofgFcCi
KLImjrjP9EJIB/Ia8G6CSHFRmyW/yc2C/ek3N6vJ9ECxDT+W1ntnBu/35nhAIXd8FdSPL5t/4n5Q
3BuEb7hrBBGmAJ9zLrYJu/K5Ewf4dd2eyWRU+AQBddNaY4wMFQuTFZNiPwh39yQBDogL+i/NdInW
1Yq31T13R82UpfQNlK3Fx+XmohvEZpd0nhebBmXqVRSCWCMO6CobSS/rr6Tww1uC58nf4ixghZ0I
0zdV3wC1ZiElGkWvjVDmRk5A7TqZOUWMVtqVnSQrM2dyOeAiIGz8W/n4lsIEdIgse9kImwnlqHVH
bYqjDqgPXVqv0O8VTPF7XpiRVK5p+2lfgg60l81NHr1TECdMl/9OrE+Byko1GbjWJR/Dp+FkeJ+v
dy7q96Zg8V70jdibXvndq7O/GsMZHDJiy/ezdLaemWC4xI3fEM7E8KoafEjV3DdppwlZjbyVyHu2
NQdAl62+tW0s2nVWzXMdUUem8Pr/5vmtwxgrJWx3qyinEy2X52Jgmhe12Fah5m0jm8FLHb5yMOct
iOJt99CVbLciElNVYUMQ9Qg+O3gbMHao//ISjzdfAvBv92o44owN3us2OOU78DfZ/WCS7qqRMdGA
3pD/E3esizQOiW9+ChCu4hQnEBWOvHS5DymeDKlkWV5tFJKZQua4/yy8vQNspgGlhfRreHNkSomR
v2tPlT8Q2WIBLCEsr1qALwm0GG2RJI1GWP7tQTV5wVW8Ypkb/oTn2TEknQHq2yyi96Gj4XKy4XQp
9pOH8dgGDVPewCXmEwxNLrP/+LKtzDrcCSVDb14NXqc/D8RlQQascdvmzU63r9tvgoquoCNmFfS7
gDCgwruOpvCq41Kt8UNKsFG8wbgXXiR+7iDtk1jR+bWmehaR87LvH4Plhl+Fow9ifPkfHxzsh52a
twca4pVqInA+rZRYlYSzx0yLKxS+8mt4IxFXzRlRe1L2eHXf5FOLzCyJaLZkRhg1ijYmXkKTXAM0
t5fkQIp5LwK9zxvEgWoLmDyU8X7FS7GZxZEy/WtKrq/C0Qtspe8FM4PHoPG4jDNPH3csGE5wElg9
oI4GVWIZJildtDI3gTHU9k4W+PV4CL/5FpTLXBGYPKO4OqNVUtjwZvGoJ9PaKBi6xwwvcAkcJwxs
Wbs07CiXuXC04IFYC1Yofn0AG1F+nq9RSYBobtuaw1j9UUQMszcJXjckdto4eSb+V2CvMPmkpqas
tu8rKOd+Hcv+wylTCuAcjVYvMAoDy2V9WDg7oQvMUEbRgqkGkrtApeUNBXiWZWeRF3J+99JlKhcJ
/3o2f3kDCYcZo3uDgyK0u0brvxEfYeUFN6FloKBZ8BvnWSJ/jst/CMbm82X/8eqXBC4/c0l5qVVx
0s1JTB2bbGRdp0RKajsVrd63vfhOEUJ1nVEPmYBTUyqbIP8nBojWYC66vK/uUsIR2x1XptRVxfL8
mqIzzXrPwq2CBYF0FhO0RS7vaUgIeOaqpfy1j97WbkF83N5fB+SG+LFGmJEwNIZymukcISMSW3Lk
Stw049wQvrP4ObbjmelN38UhHOS+A0z58zExOQEPnCdLm1Ix1/wL6gLg0CrVWco7q31fOmQd58Bs
RQI2JacBpIuEW+IbnoXnp+lYmfwXXeJ7QcjU3dQVAUgum+DhsE2l1+I/R6TZ4BIySj5xZWoeJoPm
JttG5d4KPUA8PK6HSogvic6ZHGISgy7rC9qJMdQ2dbPzUUWJIhchI9RxlNlZBFETlUO62DpxIdFk
novkRXIKPz6UKns1rmWibxh5Yxrbx8bkGyEDkciVy6BGO7MlZA+Zf9YtyrmnXc1HfMBYvD20gezf
xwRLjDN33V9g8zA1Cf58vydoIFi5ykmV0nhODCYpYy98zFGzaj1GdJVkOkp2D1+ipgUVnnWzTwYE
FuHx8aaJ+4lHVy4EvNKqayiD0w43EMex2iqUQjLbiyGxHBEvVMwzOqLNvhENUQhXVTe1cZ8/+13T
JVaeiY7ETM8FaYoydNIuXvtQUrmco6QjWNsNz5EDGFGzkaK3crlGv3LrCN7/hJb8XxEA6BJduurE
Zv4hqOSt6MkhzFxlERPz8QITS5bGoOTVvUfgfLD+/6IIySmjre7Ooi6PRgOLYBVxjFASBh0pGK4k
QW1ugFSL3umISS5tOcdzxGcHyz/dlgqnwIc/uROo7S6oXqmtlpcLFn9Omx3/e/KHHCkhfADAs/1p
SarPoGZuyTRH9nwPjpNhx1KH1utK1JIpj5gE2VC+4XafmzepyAzmMeSiaC5MoSak7wdb4FGPhoi8
xMvSy/Lr5/4TAmyyeJMo+tNzKzWjyWjSFPL32Rqd6o+Z3gL8cjXYz9JdywtH/p1VVfJj14LXKdjo
Q607CsEVE2LEZImYnREdwXfNFg+vvqtQhQ20fr2XkxrfVdzZtXj5OSEi+4KCvAaI5kimYFTxyg9N
fddWCh/uQAPgtYewGg3YIWofhaHwCn5O3w3fsu1fkZedi9A7uT9MfDYRtKAZQ39srHZXuWdfQ69Z
yynleIm3Ogs7tPZMlI8Y9qIV7RhXBCfTCAKfQPUXXkiO1zscRbbqyKx8QOXAD4GETN8I/0Vou+uR
/t+i3CtcbeCbyE3sP/rPFuWCUHwU6XccrC9/kIe0YQYxaRnB5IN8jLiH+7567SnhYa66D1DjXXpK
xXlT7wE6+sdKjVDAjQgnkvpYyYcxr+haaWX950kPO/BmxkOD+MZ7VeXQDooiT2vPlg76OWEdRDOP
wkyUjApgSOch2ajVaR4mxzDPmbVD6IPZxcauLNlT5MmZw15a4BLSLbeG1DzdsmfyvtQq6hzwG3vV
Tl0tkJh+3S1HXubv/HhLlqzEKaV9y4hHaNwzxvV0dvsIrLjgUGVvLADUDnFtnjFSCILsAAsqm9GW
Wcb4d7KEsJD7MC0EIdXfDXYdCJ229jjnZmBlyeAnV4YyROlTUXaqX8N4cswRgfyQYVLAI5zt63ca
7LkwdiQidcUHKevE49aZmy+xHVQBzMrdp0UJwk3Nw068J8BsIcFyU8OyWOcC8GLn5mGF0B8gMtkf
8MUID4MBW0qCbjcDZdtzm42GnrZ7kIWYWr2cSYpn/Ymt//tnBBZpZmXGg49o/RnAX22Z8DbTjgOP
6bFiziwQ/1jzn2J6s8yDYzaujv8LB26i0YYEolQZW9Aejoh2IaUF2onA5HD2SP4+r1xZncMI6lsS
cQGpkTJ/a8tUuPjHXL35nvnaSjUeb4aSac9Wvr1LmUjHAvCJV2NeXdVC/WHNd3zi6+v72pvRtpWA
se2qJ8CcE91LttQWkqEBtRD2/IkbX4ywhH6M74RyIrfjF3XsM+BLLIZhqVnaYDTKBNg8tHByTS3N
5Rxc4N8WxwZJ7VmJ8LFeApBOj9brUswSfRAIfwT4N9UkR3kOZrFdZQbnKGD24XfvSU9FdbRH+NYl
BRiMdCBE9eOdqtGi4WxL7bls7ypqvYhfpqU+EEkfp5D1WOXXmetkGgoI2SwQw7woyCZ6EG5/nqTw
12oboC6+2GnlUG6O/hDJomjls3qcOYjvbcr7y4C/zx9L8AGGmucq8XXibdkTS+7RPg/Cx9bV5Ccn
5gYFoq4AlWqZ1B7K1VICZ8AfcT4eHEzaa8Y/ut0zBOBRO+7nFVVbZMx5ALXiBSYvs/FJC4uyWFvS
kR3z9TklquFnT/OaTxy/2vo3LQ2l9WI69vnTL2ApgSpfF6/0Zi/cUguv5YWkR1N8lRtIulhnhINN
UguIq9bGWi0IqKMqgcLEPP1IUEumx9GyBkbGdO/PcJ9h7PkN47Ox/bRGNbY8WVxGXZNI34bFMw6Z
qWdalcePCXDfxuDbME2j9503feqqjI0g9kRIy1sQQgXexOaOLDdKgyxykvrbaMSDoCZLgKSXP3dX
dFtANSetjoN86sBctSW0sByuXvWrTf6QFglr6jGRj/Xt4T1RUSeglfJl015ufk8VDR7sTAzeUDZQ
br+hnWjjJ1kPmHP2WYqHwgpEQA7Hyp8Av6X9SA4P7N8NSKE/2PTriKVpilJggXXV8laZhJRcHQRm
pQPFYV8HUNzEX0AWJ2ftYfAFdrp6lVt3FDVlrJWejqnfOLgxFXjAq2/kShaTDnVQVZj0pHWIa35v
NUZiG2qNiAy+tNkl31D3RY10Si5KFH2U7lRRKDciCipEjtDvDg7XTiXWX796+mx9UE8h6Hd1vEP9
f2B8sm07jBC83X4Pyg7P2/hB0R7WCAmMBQdRzWPa5sBhbuLpDqP82Q76FLcNqtQ1DhB6xfydaxQG
roXo7RHKfh7jiG1QHVgHfgAXDqSa812lxDKKixrHesJbBAfQ2/+vIjTgpvlzUuxhduHcEvlsnuXo
PcDwlG0xtm46BFQzuCHOT408QvjgpjRB2B9WYE3CnSD5ndaePNmU/GTMA7r81gwu+CM+1gEI1uH9
zt5iYwn4V5cOeM69CsNHho/CLdxWRE3QwItHR573Gzzm108yKQV775bgfRMzSNBWr8Qgr6X19u4K
FAFN2TJfP0GjSb0OeriG/p3mxgPJS5NXSrfp77CcjSGQO13cI8oUVDSubYwl4PYo5Ly0XtHXX2YE
ghRUb9N7PgTeH28cnafGkNTCiSLLTmzBJ4Ybd+LSOEB40C45x0wF/6d9QyyBoNXwxUQAMQQU6lec
73Lhy/gSW2HCIYgNL485QNKdaPrR028KFHBKzFCpKYYUULVLpPoC1jfdHXTXFCD9t5ezNuYnXGXg
g3Eb+yYBgKjsVz98ATiYIuStqe82nPakgtvmNtiDlscqM0BklfhNaySFdyvgcYZjUS1UMmBGGj4E
GZUUim+/v5xJwsMhuV2N77s/7PHwujOKV63hJcsLCscw/bYp0DVnLzjSifnc57UofBUMVLvM5xsi
gFbGcKrKo/DWoq9+TUHiesEm1bOYEsWSNLWmU2K4u4WvVk9HkP8oFu5x9AA7fwBeYEEMxz1S6UXB
qkld745wrAtHMtKouW0W3Y03m+AEq/zas0x2XDg2s0bQO5CWUnOgHbaheJsD8sGUeg28pj4RT43F
ADmVctqCyVQoI8UTOhNo5J8+kEeWKytAjVST/1bH8GOGVAgv9/PeatphQTlspsZMg7BoJ0Fb9DfY
ynTaiJfJ0wVEOdni054158Mj8qWRrL6mBrMOqXpe5FYR4QzLrUhq75XB1JW1c8SjFSFm5jkxpSLr
KgZ90A2/qNB/43YR+XPnZ7rSv5jFDvcx7Da9l0E4GvOr6O+GJ5ETxgA5GpiuR/A1h/Sa2fbeA4CS
Fq6YJ0IU4H1At1YdlF1xSUQ0eYp8pexiCz85KzgM80nHlVga4TMV7kN7NMsiydbMuFg1J2z4r7/I
4X2Rmi9OWW5o/P+t2+4H3qOGwcPvBcRLwI0BnBS78sawrlPyB5RWnpWhI1BM7dmI9mZ268+M5dth
BGVlyUAiHowFD7ueix3hMVAzZo2pb2tLJCUEWRWmDLPzhQMB297nVl7WQX5mqrOCKbeUJmoMojj7
k/yep3hx7TMTJNlaJn/IMHZWDo2n+S36LMTHpGwNGFP2saGbGW3psZrVoo69avBxnIMj5s4rzWCI
RNLOAxZxGExan3NF5bAwYGAf9VLUD1vKfO43mrx7pQZrjuvqawXRLLISK91CMooDrCpE2JZpT7Zp
bNoyFcxGBRChE3WeC3fyYnKTjyCTSnimVV4YjCAvOT8c4fU0f1zFnD2GhriMSzXxa2+upu61pwI9
ccdobi8t/LwA3VgXzZtbptY12SpPF7Kyrzmlm9R2zIhlLPZEJ9WXWELEpTZa/Eq4s7v/T7USIvnB
2AQDiYJ3LXBWQKn5y7IEWI1oeIo1UR2dGQ333uidNvzWj5Y0kkE/zdC0A4lko6tuKHdUVuUp7BqU
eb8TIMVdXqHRB8kJ2FxVgDwirGTsdlLQvAqHekiOnx1tqu/z+NradB34imHgFCn7ucLu2BgtSNts
Bbz0jMu1ZQbiTw32MO0/iYjDnYt+aZ1RVynm8XS4wgaCUwnz0Ok6YW2vbRDqWQDvM/Z9QLNEZKyM
AW4XUXzYS4dIgc5BzGnxGXRRvcH5etpwNDYa0ytlhMeFCXVbjCNFU1NY8Xu5dB1fVVfhiDYAKDzg
W3fidSJNCxVbbxgDOOLwsgt6Q8r3vdRAHAHUpHTLF9+KXTWbFH8hyUYwMjq0iSjX605HSjPSGTu0
IbUhe4ASTj0OEuYecd3w8UK7t5mQu3l6Dm6tPaY4AaAFB4bzrv4/tkY7D7MK3w4BA4HakTSFnxei
SXwZo8Q/9/0M0bhJ3DFePwWgbtJDDSjfKcERX91cpbAsiHE9PtXIoCI0K/w/uLZOEWsPkSSkUTJx
8LLTG0pxEvt5Ay6magGhZXP+uRw3X9pMaX8/8zxGEButgc8KYiCfeWx5NYAc7KqYqkyLKsk3sqOP
UCDqMZ3CqxBK1hucqF75rkZs4I4dM2TwlfMrVIL3sq70MPtk3KbJFk5Yes7M0eE0jn5NRzdBmRVp
mANTe63HAcmaYcVQm9bvUc+lgyMatowMYlq2e0CXH8UrUYVfrBDl1DXaGT4sjb9kEtq0p1sMYdE8
59cXSp1mncpsR7YJWe2V4o237OqtLIjZ0Aq3J9gdLAyfVr9dvZ080ZK7mViawjj+a+1/qNW9rbDP
LzVwxlRYTP2FBKQk39fQI0EGPgLtoWiB47Vo1HMPra4cD302iU4ey5lSk3NBG1sXZVNDIElAbf0U
q/ma7cGKHMs1wSgAN//FoES2hECtQQ5H1TqYe/hBDhU3d5XStjkqCU/noUEZYRD6LvegyVB/vf5s
bioHOUIiB6cctKvovBAltQXo4MmJjDSNcBZ6IMhR4mj8mXX9qhw58fcRdDX2Nsxi9MQzV5Hp3Z2v
os0nnOr1MUbe4u1283dk6PYRvqLfOSsb4n3dgJeZh6cfcYTdk/86m0jcnq6upGLrqyYWgED/7mH/
aTxJdt31dmTV/9wKzvNQNFemxJh/0kNu6pwhPbdSFGw2dX9RWVN7xYk9E9aJs5eZlHJsL7Jq5KkR
Ii7jib/h0kX1CelBvrAniI6NeoabNf/30pRAVRIL8UASjTw3kHJRF+E48oDA3JYkswCXo4wPUhOh
vbxN5/v1PWYXcm0n2M+FRaQcrbFSM0GNwmRN6YnUZ6KgiCrMLrelGVX0nB0/nmXC4SlUht+1xwIz
tHjkRRJhzCKIDPttKZqc/PneXYg1NY0C0Es1VEVixplRSniGiamIftASLe4A3b8w9ohdOX+VqF9z
0kWc7vWT2x8wdyl5fsWPN5b1u9mwN/ZgeZ3zL5TcOzUPGZF85KR5Yl1RXL0WQdLPkf53VVwUg99J
JOFSGd1XAxfocVuQEC30ASAMMBECN0oGWR0aI3QmtWU5NyCzBOFoPjYoKniDTlBJ8yJnN/NeqL1C
rPhGJoMT7jRpIjrGjjhwmhE2Z7ZxrTs+iPwesLcjzDDb2cuUovLyXpZuNqgydFre+0CpFhot3n/x
AojlRy7VyU1plo4lT5JArJ7ZcWhxuPsZPYZCaGLAdRv2/P0Y+qroD42ixhAK7IswB2xESyNlKiL+
8/MRZ32XICrESQcpg7NWqhHnfzPZFk+W8nLF7D6Cnu5JViG39GvHK+seXFwGGmtrpn94ihtjo9Jm
rd13VwmQAxJe0d9JNAEvWEgH53V6cUf6wW8mWo0uujIdPTsXwPgqYBOE/0xWSeiphGE3HAb8SwVM
fbM1JmO4ysiM5nNIhZ1FW+BjdA+ChhnIZnlDiJ18eqXUvwJJKbCg3gFZ7oRb66JgaJBLEF+YAho5
eQFBTtMLOcRo4gE14zXEh96OB+jI0FDXV5opUJ/jDQ1TV5k7gTaSSdRf4Ou1AbgVcYuU9xuudrqB
Y+MHu1UsUvw1IJ/zUkbIDMI6XF+i/ugHjxSqTIyqh9ko7W0C8eSS0Z0gMKkj4He1NDurfchgcIfU
zkMJJAmyviwJFBjoV7KJkB3S7IBtyj/3Vb3HQhxdVPz8Zw5w/YnitYRVja4LqCpkrlfgGITTGheI
QqUe0X2Y14A67/N6KpgWVrGJ3hZGtZgRo0/zH6vY9+SfrgoTEQFJBIS9xeRoXwa08zpG/a79ZXP7
qPh9cmor1Be2wKE1ux+RmDn/Q5KQy4JNzzvtJzV1NJqO7t39GUi1naDsncBucofXr49WxXJaUl7K
F+ecW8ScdDEF0YcCL5OEgyhrntyB0j5P9gdWXEmtvjoFL3d8oNkoKxIWtDjFObT27v8Ql2sOJUMe
q+N9Dvbtud+SeHhD94BU0lH45ypLDCMGjo9V+/IXZGKIAARXCH/vpGNNrSv/fwhm3G541ZBI/mRb
XhXK3KSyh5XkHafoOc6zHQ+9TiyRMxrtlm9k17L+ufsEyaUtuOXlzEIlCSK/e7vyfMZCMkrsEQ6x
NPKHYiWZvIDp9qDf3xTz7qKbFRxSj3/bd3i5MkGD5jeZd4shKRkocBATK6u2kDreFP/BmgHEZQPY
UBuRoBHKTXWCwRccndooTNqhCTvrLrE04wDl9J6JyYJv2B4/ePJZhTsnzCnJ07AVX7+k1Q8Xpmot
TwEQqugPabxI7NV9mZSOvDCGloZw2OKHtUiMhHoCJcjCYVnN/8GILPUUrUTSZ6h9/qEMIUXZoIsN
VuMMzNCnsiAaRNiiysxGNlplSH6nz0fKLw6EO7XjcwtLgK33rzHJRPeyHZh8zssYJQJoW2hkrkwi
HSA7B9VozsshViYGZ0JKgdTZbBBYd2SD1DflT2XocTxX4UNBtRHH/kIArzJk3z7WvuBqrVaki6mM
8BMbhXkQ5WOZCbnxreV4a07ejB9qYQh4zfqNgUNc05zZrnQfctPFHn377vWxSDvwQJ/t9YNbKnci
5qZzmhByJyKvO0CA2AZbPX7GaXUpTtGId7cHGch8zeMqcTPGtUsun9KKnfK7++eTEoOi6Dx1HBzy
ryWPlUJymVMshadRxwgwWlY7SahlwvRH8KvNEIHsQzbkloIXjdtgvJP9VzUZ5oUyaYN7FO5erbEK
IgrAB2+m80N57kThiohe91UWYbx7KZxjDI4/9BjcI8KgyRKzwsXy/jJ/Cm/C5Hh3K6uhfp8ELejI
TGNdklYFIr8nVd0JGCtIUILx1PlFPVBEQ2rppsvNhUnEBbjLBKENmaB079Jx3/j19XIcWPxiTX2I
LboG/GI8KYxqGPZTLXtdQF8HwzfjTXdoQ7Q8G1S1WVqc1W99xRNMGp5rDOlcy2aDI0mzUFBH4ZVz
mDiTXP1K+yHdTks8PlxltHwJW+N8gbMxnfgQMUvmuxHAqsF1xzAy/mc5cZZN3t/lRvkhBOEvT8RY
xkvrv88b+dnTgM6SP1xgyWh6sGJmnB+q0vPpQKavD8YQMAjxOk0XlVHcfwXg02lswEU0pDVNAYb6
SFEs96CO+AO8/dBbCv87mCT1YbedhfoEA42tQvr9Fv5RbP/coL0amq2FEOi5swo8q/Na9/4/PDrd
+0c+6mRZAxBwlXy70lJenLwENl62Pk3MLORoqGkoWCtdmdGMM8NtopXEPu3/geOjAgffyzkOzut0
j7LW7143xYVbI6lRnAvq6vGUELYoRqQTNBdkES9ccxoWXcUIgOG3Xd0VjtWcYhycoyDBeECKh8Hj
VL8vkeSESh/uhB1FrTfStw2YhoIg0AHyQDINbov+fXZ7leGKTzoeVmMMWwRv/EXSDHlkrRrHwGpZ
cPhpJirm5sqJyCjKpQc08oUraTyGxGYZKUHGwe89agWM5nCrbsz77kF8s22KQS6qRTtsDabieRyp
lGVtB18/GJXrTVoLxuIDlCKOtYvw16BeTRdCd6fory0NObGJxLFrW3ufF0WZ9ay3oqQo7dv71ETI
J7zVka8aMyEttLL4I4SqEvGpLmfKORur/bTtddzmNyhYFpO1Dn42Cri/iIwBEgcgM5EbzsUIJddG
FkOzSglQ/krCSjaLpNOGQoPYxwHshP/6T5pbGVFU3iUNuIvOLjMK21rMI1pib3JwGaLLoKrZxKJ5
xUPCwd9l0i/0BHueU0tdUmOgv/IUSPR6nWlUR57o3iRRZyYsuYMTyvtha/0XQv25bI3TiyklrCCn
6LbCdN6dTgbE0ZVC/2YaPjTinaGenD4AdNLhekmdwUDkvl54Qvt0OeVqp6e9Sb1yrXJKWG23mo2N
c5QR4GuuaJTbOqxxX955nx7rtZDh38pVx465bVc4JFo816I5na0l4aeSOBN991x3YP3Jewe6jDU3
z32potPmC6C9nDbDtIQwtiRGpCFpfaBSlxfxXkptyutBzHv6CBW3cN89Xie48EFT/OWdkRCLPDv+
bgqAAWpUVyCxgHXSXDQ3DQ3TRHcwAGQr99PZC2cBwFspl7XtB6/eABDLe85T6FomOUxfUzmQC5HV
2GfIhPR4uDR7IFo8l1NNHfkHQX4ayPlTMRF2IecXaO1vc0Em02Sq23EdXEClXBad0GAuAA27euB4
4hPBC9pMy3cZUvaiJIC5apUR+CsppbjMHadcgOuVpVA6HsN1y/WZeQZmBg7z4TxLxQ88PNgJBvuv
6izuDE5okn4uIMBKhIZH1jzNx1wYccKfQccTLJhZXHE5bBR+jjHgxBMjiXZ2dylcB8O6+35d8WS2
0J40adpLZ7YR+wG0uU9ZTLkfDxICAncfTxCO/QfQVL67MATWwPzQXpYfWUtXVh5HBOKki78JuX74
FyJ3PxpzJ4Rea6vf7zU4hVhbbmZ7P27cwQFQQ2fA+QtlSMl5lwXNQi3ugsG9/l/gDnxPqy3klIY4
az715rzy9m7TRwj2niXt5wautrcriWcyH4tWQpiBAyxFp33lTyQYw4idUVBWIdAqvZZVK3e344DS
visTfz5f/PoM1sgf8wGQ+1ujzmD/vga2pV3ighYmZLArhyacIaUDuXCWj6FKnXRMXS1e1tUkFfaf
y5BWCZ6gkcaP2vRjoxce8H4yEj4EDr2Mb8psfTviUC/aZDEjT1ILXuk4LNbkJtoMng8k4mzPoEbe
aIr3OcG20tHqrWgLaU9zitcUVYmDz5a7T41Nt77kOjY4GG+5KHHeNL7ah0G+4009xUGjl5pyH6en
uODGpwkgeZa+Be9DPjNbd1MFxwLdfCZUFdVcrsGVKQj/OD5MafsJdKpDaW9ahXzubRnxF13A41qH
7wy3fX476n/G2W2xVYVkes9PHb7BTAZF5z36XIKljSLOdGp5TizaAiLAOpsBSsl8IxxHyCNv1PqG
DI0+9OrFjD5Ljj46dp582o/IZ0NxOsoSbgx1yU4hJoY+ezmaAdr2H4l4JO2SQ7PNgB2O2KIjUMdd
AIJ6K+Bmdo6uWELVZ66VwqCDTAhJs83EIrvWEwAimMPSrCgnD2ETw2uP8Q238h8EJAsxHbp6smXe
IX4LVSzgr620zRe6l57eptqwlNMllkpbCvZEfwIkBr4aAbaAW8LHWzwYdKdXCl0l9mHZ733kUPs8
fgfy3/+tFgpsQY5AKSt5dNjlcROle1ajhvjl4skyRWx3ilre9Rt0e3q6acV4IKby/3A3fM7YrZN4
0RyL+O+h7lvBuY/TIf2snc0SDEd+h1e5sWUMT+PL/3pfYU4KPpHNrNTOhIWCQkdRgiMqM0pbtjby
lkMQ1H6s92lakbupzKNjMf/qWMNPc7cjgHukK1RC9YUuWWoKDKJ93j7ozx2n2cjja77cbGrElqFB
Vw+6ZWdpS1dJ/5dkCj8kyy21P6jJW1HTZSDYAw3r0UuitSmVnHaLdGd/Ume0h5dgPNV1iY7cQsP2
qzO9LWzzhKJXyT712RD1Rgf4w6C3DQy+D320eOnHCy4OFTXVPoaFUWwAHev7Oikc+pyPWQt21rZX
jU81zuvD+hMENqz8HCDwDfGkL6ZSWprqNeT7avMEvAwB0lJr6OSoyBcOMbjjll+q8PSw/5PTNwjK
DOhY2nJbJI6IZCM8EMIj7YwdNdhF582O9bL7bIX3SOAVsVNusUd/+UxzM8UGH4EJdNQwnQwmrruL
ohHHbU0secUjWeCCFrvxO/hrFiIzMUt6Ax/4WPindqeVHEsCjT2ftSpchJVEktbNBfiYu4C2J0OG
9ySuZd0jVENDl9UVpZVvCRmrwoZv1FP4naB1I3M+l0e563loQyvkEfuuzI7cOQYoL0tTcHTl3JSB
SK4XGD4aQrL3pFens1zelLv0r+EUoqYaJvhFsL1+/ovoas7WwwNQeexOjwZ1YZ0ve6jraYuxssl4
3wBkKUduzXoMrggPPl0vdg33fgFYWLzZajFpv1gRYgQmxMW9lQxaHiXwX6fjhdgHHF/Vw5wF5uJe
K2hy2UC/LdO1FRfZy/lWhRSlyCc8SbMPXw+IcZDlvHlBxF6nuCu2uGe8tBlKEImFAZJp+zE4aw4q
Eepr5CbO68F1K5EKWBRFqgA9d4klfUYZfv0IL1VsNQ2y4cHzlATazs9f0QyHdGRnLVXG0JeW1M8m
wpHm3ojEmp4lPtV1lr2ceuEZIfLeZz36INFhyeaYtssKtI1/vDj+Ls5fZfwQBOhmwBvTykzBrjS4
fUyIhG9PF0z+jf/oyeT2vwcxyMaGdTxLmdtpLMOjZcetNcKjxPQoijnv6WHejuSfPtfUjfUMuDNG
TLNZO0QZt9HMG+SfgZzBdd6t1OgiYJY//PryYEoq7AXwdig4lMvWhOcMswVKPhmVsU1WlDBXgCVy
awZU4IpJ8IbxxHsWEEgb0/a4XqPw+2EFqMZ7bVi3tSA7Jp1AnxaJo4yzVi5SsM1Ryq74BsNjVNNr
0uUv2jjSxe3jbowtRyOnoU4u/D3DI/8f8Q6z0Fr8ZXee5o4z7GFvLdfYoUUJM3i/Do7xzHf7iyNl
+ujszbTYdDUwxdziT/NNRJ9G/ICH1c42Wz90KsinL3/LmnbmS21Y1b0iizJFUkOe5frBTcFUZ7dg
q01lbneVTyra5nz/KqQdPYay42PTuVAGje5UlPz0LEZtLL4r9TD4BOcaR1uSAZowVRXCpwF7Ks4P
3hr9ojUveInldpWKxnXttEghn2gfV1LDw+mz+RUiUM5NfLCayFM+gNhFymuHd72nDrr8RMdg+oku
BXVZpB1l9Wn4pb5IJAxDirBu/dmybnpgJrlWVPJiANZfjPcrKu8kQLquG+FCn5d+GhHlg9FKpl7N
0yP5KJ/gW5+RWAFWgfoaFfN8EZK8bKebIeZzK5Lia7pm5wNS3tbT16RP/qgXgkUZiJR/ldo7BK1A
qXBflm4YFlXunA0EqVxhFjDG5vVXxXhcFhhxBKm0qfI3wuFro1cfHhra2tbt2j7HNnUNMHXzgvkD
sGcQ/OLt0DXmtjrShnfE8M1YaL4FMEtaal+s5XUlDw68jq3iIui8yZyG30DbW9FYEjIaJNZ7kxNg
++DZYvlch+3ZDvHmaWY7j6/4qOGAyk+iWXuJsfR1+pUipG622WcBsI2Jr+awmurHydVAsY3hfrYI
2PUHIqqTsWW/WMU8XhNFc+jvAhZs3aRHY7gzyWObNWYG70xCI/mNU9oJx3UEZd01kDDHQgBLvv0M
k9CodzB7c6MAi0C6rfl5+4z4TScEBCcI8bFXjelL77lFECRv36SbYn5wMqTKtGAhelObrFgOGni7
DJSzprPtn3T4bE/yg63HAhRNNDKOGNNwtiQ4uqnHKfdddefBoBTBZTosBcrWIjk23XGpK6eqeY/W
DA0vriR15XxIExXZ2nO+jVeYa4/zqETnGH77DdgeDZPgrmSZ0rCMVxxzPbdwic4mPPirkGNerZBt
/YPreodynwsb4uZYUvugdpd82vKCklzFwY7e1AafJkWcqGuMz0TqemPxGjATllg08kDXTRaBFAc7
yohO+g5y3NWdY7qtp8iabVxxU5hOxWJtrIDWahhIA1FUWqBrU5DS5t1iDB7B4zWxzcLc2demPDVK
A8XSWckb2gBWFAsh7Yzw0BGgpDQiHqEu5eJN+Al6QxHQlMSmshYgZG0RIPRCHQjQYfrQWmxhAAQm
jgKih2Ykv/4KnBZ09qfA9XnF5qPEzQWb0kqM3+2BH45/PgJyB9q1QO9MWa7laT74oK9XIhitnASg
wv3md1NIq/m3wMJi0DRCsnI/zBWGQ3L0wdOvZa7SuFBGkmIicclsertBHf4EwwWWNFuniTCIoTUm
bojeRvw0+BqU2FeoWJasE1sbhB0l2wer4LIrdMZSRhFukY4nmpEA3y4QdYJZMTxXvlKPsaDl4fSf
3bGGJ+hofAjjFIZpLAOfp7/4qtU3RhvlY2C3Ay1p5zaAfulnQs3AdhWKoJMIfI+vGo5etTnxnQog
iW8J8GxPQmbhEc6GuJQP/Z4x5zjk+g41/Kp2bB+ocwYuoHT6PV7x5zAwkIiZSYqXu1LZGtWXkCyd
yq81AjHjHIMg3hnQEkkxPBbzOdngulqhclcjEFTGYj933ken5G3lfmWEj1buVOvAxUvZtpSO/VFm
c8IslRNBfgttG1Ar+cvHGx2pJO7jPj1MkVe9zgvk8YpxBRKHOkFCLyqWr7tSIZQ557eUAWPMr9qm
Mat3VraXkSVLCfsiX5JrmVGVrmES6aQYnAo2o8uu1qyuXp59i7Akxz1NmFRZGI5pH7N3ZNpTllib
JsQd6K+xvjUsFZtfHzZsorw1waJPGMWNJbRa2E5vgVP1p/8cnlEokBVBMyer4I+dhcuilwXttcoH
zjpPAeep4ffHTjqnBVI23v3A4eSi7lNGACsZgYBBtgsstjtbcWpYZtAs67DL8Q6138CyEKb/U+eH
maOei3ePQWZuhbsSrNFk+47BPVch/U1XEnzswIr7ksr5emWXkgpfxUnR/yzMqlKUqaxAGUWsyhep
mubPJfbP8vSIm7E6R+cz5LAQ99c9ru1I+jgb0aV7+QgyIo17MXDxzSRX33oENdqcFrGuoC7CEsLu
pdkR8ztDzoBlOPOA2c7d3SqaSIJ20l71ZHpXwrPVMON/QaYwBdSb9x6QIfDi33mvM/eZE9SP+CqR
gpUuZ/JmAmHG7un2b226PxfI6y5+1ywSrX7T729wXP20oRM3HmrHnijF+PIFBeEGmz/eC9dWwkpk
rxopoCr0liQ+MyXCq4GOCWL1f/AkGSxjK3YKNnQygSImQHNplqgc0aPne86oZu2jw54wk2PxvfY6
HFTXDICMrzMDvpkA4DKJOViVE4yyP90yM6yj7UmPAK/fr4gAdsiNt6ka4LN8hlzwLlobZVKy44Xc
NUuicFUz3KJLzdD5U8VIyoZbYkAxVLIsMHebiuL995/A0fIYkMw+LfkyQmPd4fvX3RlJM57z1qi2
7yDDUoyfrCsxUIeJdibaoebetcw2wK1Q4UttauvijY8tlRb2H0fnm1UjAbamI6a5omTVLitSr99+
jo38yhn1tPemiVlCikFjMrAHMXhuCBk4iNeSDxkzyI1iuAR9UgqIbzjeAoJOOFN6mlscYakMwiR+
SiqXdAMgmNN4AR0t178G1U2vhZX/tVDvTW8iMYzx9zice+XQcbja/bvHDNb4AVuzVSnmD4HryjGW
JxAIRqyQcAeszZTJi0OExGisXHh4HLpPuWDv/u3wgPB1Z/x+gBqmVjKaHc89TEz74M0GlhMGIFBc
jA+CnZ2mkL6S8EaAK80KkTO02up+7mZXP3+DZ4379n4aleWLX86PRPfpOMsbL5yxqGXWZVLDMGpj
XRXXx9lSQUZz3algpG23Aaz8nn97v2eQmdkVe/Xbf30fY24E6BTPoorwvG09Dh0LTbY7yVJGPMCB
dmnbIidmUgGct96asPatAYAz5TcO0wCnRC/S8638CVrxPSDYH1ESO+BZKes5wAU4syvoAohy4hb7
qM3Gyml57E+OSKbC0rxfLtVskzroLLvjLJ1EYhoO/WBTxLuWTpfkfJqWYDMnTA7qzcOrfCTD7s+o
xpleDSAYzAkQiiGpY4auTt9DIgyncoy8cg7pq6N6DOPGKKL5P/bfdM1a5t/vYRQbpJuH2KsTLGP/
QNGH8gD6FFx7t0wyQDDTRMDZzOFeUKMQQHFzz3dQMdMjEBAFXhAYiaCQPyouSsVXEZmka31S9zSX
3FjguMc2of4K3P1wM8VyBXWQuG2oVOIuMZCVn82RtcDnljUeHf+DM4LNdgIRaZ0wd5lnATueN3bK
JfX95Pisb2uwfs6b0IviDIgv9Cep33V9M6JR3zzCqusBaYJV+V9wO5ovX42Z/ZznDy1dNuoa6tVD
4VquWkPGViEtKvMI+krbPvbpCiCV77N2soPohKk7L7umYhDd9w3FkkS/iZw58px7LrcNQLXc7dnC
vSyoR13KCHNVuBeE+VC4dv8MbYwxjMWEHYSw2Zha/rwhDVYvlrxqDi79iiIi1Vo9E5DvEoUTgPHV
dIbdGsBcgiUSKp3vF90Ej0n9ZhZtSFBJqlK91xdMQE5cninIFjXqh7WlnxTSd8M15A7RAGR/xA3c
hw1TKzmMszGnelhkgPEyctzGDTy2HUi2hf1YirXC8nIDz53ysBtdTW7q5vdZ/IIQWNn9AAGShxHx
sNvCu3C7cvs6g5713B78B05hhFEUjZ8d6dpEi9BX/L2DwerELiVTNFEWWfUphwI/IeQilH2XQLcd
ZCcNwUCjxIU94oDG+BdiABdEc/1yR/MlpHv3ESms+Tfylb2xt0EL7qh5kWGuuirFW5qVo9ZsVdQJ
SOK1vQqtgDvXnbc3MYx4afE6cR0RqdifhQkZRHYpUJEEtLE+tfLrS2vztFaJRhI7i/a03+NllHuw
PIIbzZVWmzGGTt/wYVYHEK1fgCb7ot5qxp/vyeTscCFmgPbQu83SXeiRrzRPQ1EuuOWFaFJujKNF
0XkYqPOyZ0W4vHYg5nKtN2Vq3e9+7gJspaI0wIMg06GWnsafd//g2EH16MmHFxkWAKpvgLfG2e1O
7U3IpJrwNQeg8j0V1wwcuJ1fb4r12uFyizSWkAGAvSMYXPev/DWDQ2NKbbsWMMGKDAirgo94xUYL
Nv2HMSuP64dIMw7x7EW0yKoGI3uAr11SyRRes8O2wE41Yaaj6pSVoI7A1ZgOCPI4UwvsFwDWtnQL
cbTXjyUihXn1zUxJRi1h1vIRwCxcj9zpxsEuHVfehClRWava9dobgnzMczpMQNbC1KyYJqygQ4XC
Yu2nvc2E17HOgi0bIIAlMwH2mzIfdVJ5QXYt/ye2bySV94XnLrszRxTC5CmPnUEEfh52MkLGOUxr
4YMAFX6Nk2iL1HIc7INs1RpRQQPoisfRF4SNg0OWBRjhgXBDoeu2X/J2Xvknrdd50J/J+OsqQFjQ
kT0I/g5AEWu4G+q3F1D15aQGPUND56Tqs9Lsaueg1+tO7bVXxRyvQKQYusCGX1aZsUm/hjDqeEIA
L2DIH/P467bqq8D8FyBdY7StzPTol+d+E6Pc8JqRRbCYbp99zAhPTN4wBy3DBFgMj7vah0ktkHM1
cTm8vxxgQhcPqm8QKOXldinxnO4kq5XZQlqiA8Ex4gac7jOe6UtMn0D3JO0+snZFRaS+CW1Pah3M
z8mBW51Euh679Hx0nS4wlpxRU2hkv6Bidzq5MxAssNbrnaQ1CJUcDCZYwAGzSli2LkdLzgViVAWf
Mq+pozMakeJB3gymkqvwktekx1enrOX5QCcQ+XkP1x7VECLwu2y2zteGiR6479sx2O/hE3SRU6+O
gnZKPaT9vlTPC1dIxsjmUrdvx+KeDvrOdZQpRey5KaZFVnuRpEZgDCbqL9muWvF24YqHudruRJ9a
e1KABCCNPRRJ6SOl8muSwEP2YooR8YXLpRwpl25vxdC6S+kgJZduBthCwM2Gl8jcLVgUMrZfKJ9+
6DvJHMl9zTFH9PslL73hq/9xO2wmpMQJl98/ih/+HCZaL63Vn84NINc8IHbiGv+5tuA6Loyl2je1
QBUp3rZx0C8a+cWNlvDF52gWWYyFzTfLHuVL4cYL5TMM7c7MW8fctBLRfaDKsA566tIFel+RWl44
kzS7w6bImS8Ou6pXtAB2yDmQtD/54huqcIS6WeNzN6OckY9GNqNaTwLPbYbRtSC0RkL7r6p3KWis
OV55RR1elyrl1Pt+QwXh8s8OCsTmeiKMc/9sPNX4Huu9jFHMtuIdMilaLzdA3ZUMYONTqkhgTNPe
Fobq5OfmW01g4UTNo88gtMUfLrIHX3udCuvK10ALgjwztZ9nqyZ2Dwpcf3QPZFzLsJvzo5KfGp2Z
etiu+F3Pgq677dKAQi+zV29gHiEhQl5PIeLEEitrU76oeXNcyk7Bm28XqJUumH5Q0cGLMHh+WJAM
gF/JWFu0toXQ4Dqkjoqygtobhrhl0WneykSWpK/yP0XEyZRWG2SfAIyvOKgYKnHIvoxQi7WadPlY
bHQNoG1lZZc65FMhC5p2meb6FOrWHU5I9YKCscPnIlP2EFkbxGhouSbcIGs5vM8n673pB2UayywG
uYPrBB8Pr4KN3dNdEwwZ+huaXx4s3gzzpYhRlJdbik83ctt6suFFUmYAcONnRfc1IOTmZVpkjBEr
g8E0+w6zob7ehW5F03tchH0xhpeneq39X9zaAOhHFv1lpjNBrnnUKYZuivWofhu+WV4A30rHXikY
SKN8FHQndTHNgsxCklF1hTxjvJUBwHiQR6snDt4X5rIRYlG+5+Cb79tcsYotig/mRDcp1/HsTd8c
t0jnt9hMKwE5njhaLQbm/nGLfA+P/eGBv7AA2S7uBdmm6J45yR3pd8uibLAT5ZzEBf4wN5b3Ly3i
u+gqpZSmDE6L3FkW8edeRTI4qcRWzO/c4eqwcBtt7NDRxVTIcWa3LXJDryD+IDqwXCKCtTE6Yl8u
xpPoobV3JJtMNG7OQ/1HLSf+u52i9su8rnGdjZB79J4Ewojf4/P0FJWQrWCy6zCarkpHftbwrYej
E1K/4rujpYWF4ix3451s9YjmHix0kKXaPg4/u8TGI4R8AHTYSzVB20N8S7uU/5gp5wAohvqRJasi
CcG/31A0cuMYoTsuszpuFdC6Q0K4uWvx7NP/10pht4n1WbtGKwaJk0Z+iKGdRv1/667A1i4TEHxl
UrOyHc9mdZ5tVi3J2FOLWfF+t1Dzlz3KJwlJEZUCLCFyRz09pHgLJv+IHj3on1gW05m524hx0keP
DncyjH4etqo5CG3Vs4r4p5voffd0hhGxUmGyN06oKrmd5N1MCiv3TRwZJw/BNEjNbncZt4KgeLUB
1FeswmDbcUi8DDNJzpZ7ZO4p5KRFzMl926i3wmudHD/GMExhzLXh53GEo5pPIGQmzCeRTivlRpzS
X3lvlIa5Mf0cCwOxucKybCQymriIYw8xRRF/4Wi4DeKmR4JhEg6JWb8uR5I4jhnapgNuqV6LuubA
vITFtxBhd0d70FwQi+LBbBXlGOElEoJswkgBJIn77u04BDk6eB4WS7mDJu+a4U00zBWgwh9qRc7f
Uvg2lj63+B5vLzcJPmRHp5li/oU+bDPZg15NR/hzcpzkKed5tdWINoMonSmJ0VCRB+K/o+gjK/O0
fPFSgnu7pbo1e/0jPyef82jtZbdIAlBf8pXtoVXOOgLeq6442sM1/e6vQP4k/s51FASGumekRZeW
o/4XOHaOF2/vrQ+gQPYUGTHACVi7MufGJ32/mT76/iNe1EZNTSPXUaU3C+7a72pT1KIkFaRIIY68
uyVg5o4Xs2LreBL/+yqu2J9pEPzsZIt2FvVO7nB7ihhtlgFYKwqoeQTuoQTtjPzWcf3ipkgF4UEc
0tYkm7xVnYc2ALrmB3X7I8EwDBjMWDs93RoZh/a8Bg6bHF2xHfY9ZbpZXvYq2PekgnNWdEnRjnnb
7gA4uVyaJr3lIG7JROpt+fi+qTO2rOUboOf8wf+SNxexqyL6B4XwdX5ewdyAo2tkQVrHF0wWiVFS
rancWdvW82KZJzhR2sJIHkLgtvTugg9hu4NGv/knWEHEWkrQMP0LOrr122oLg0LC4iRVkjj80DUD
cdJnOznDfoBpHQZK7eH/TJ+xePaqDReyz5gNV+tnzzuAeb95a8aOSkkVRJS4RrypYfvqVqHwv4sT
BBEPB2V3r5qbKKewTVDfqrE+FdOEXaMP3nqlDuGHuzDVBb8h6jQt9CJH7PW+gPeLosViTXs3R/5G
BgRHaiPdD/ut53FZVEeOJMMIuNmHMrC1Qh7+PLQCvI1x3VGemBdQQ0oUbPIxo9+HC0pTnLTmIpiX
cJdxDgUFIMoJgtKKtd37AGlA3E5Y+SeZZPMF19UYoTe36KgrSlL5tGFd5dvY8S/O0v6a34lxWlJm
MyabKo6x1gtvEjxJ08KvLUZHVjV9punlu8taN71UYA27d3jCn8cQGW6s9T6AkIwhMq8sAhQcsA/b
91bhq6ugEdmCC/Ph9Cuj+nezDUpBoBU7chHOBeJaHzPvRf8LomtvoljPjyxv0dB0NRCn3/IzKliP
cWp1Kk68u+TiBSN6mnfv4tsmZWlwzaXFPhFPpwp1aoBPZV2dqMU5Vk+5EQ8LQttkbL1TFUYcQrBw
+QbxHDfGOlIkEeYbyPgQ1SlKrTzLc7XdN0G5wMDPXhbUj7+dRxsm5QJXzMefSSrJLCalWVMHdgnZ
usv42LJRxOl87TNDa38s9jj1/9Mn58rP8D7hDlBOAipGsgnyut30pK9jkgOlNYFjAOSivC1n/dC4
c+ju0oXDjblC55m/XyOP1goXxU6kX43vJSFjOHuRXFajjcObNnDV4Ic5GhKxQDVlDaahuJm6n7pk
9LFxB0K15cZVwKeBgrZN5ws7WZw13ygABPP6pqzHpC+wlnx8m5s3hbcD9pTKOCprHnX9X9XFHACY
M03i05BkRX9XuKa0COKoUlXxPYVXFna1sSV6rL8h+M6dUd33F/Wgr89aMhGs2dldQ6EWbX6/nUvN
+0paQ64jRvmKq4hulFmQW06m9qOzPv3EXAYzi0zHDmxMQYLRP8+YIqXh/rFmmYMwbPgFhPj5AtCV
hOTDjQ/ZwjRg3JITkBt1yo/MhfIrYDSz4/6yqZD/t9Sj0N9u3IKU47mLTHgLHwQIQuNOV1cezOJE
bzWjgtDmt7EsHJLesX1miw2M+lGkN5vOWTgPrWkyhIJ6P8uh2mjWi1XZkDUUV/jYqXWOg2PQjdx/
MwD7HgXMGLSWgoLj0MYEMP5iEALhkVnS1fCV4C3/MKismyER88198Mz01ovF4NRaRp3R4oJ+NuoJ
jatx8IA9/L7CI2XAhozbneK6lEfbMopGFTRgCTajyZp0SjJG9T8J48hSgsRJrBv2Jv2ocOsM6k3U
PO+gVKc/p2jDFBxqggLBbQUw/ph81ejE/bbuCO72zhLzfhl5E8B/UlY8sL3MwgLOgQzb+N+q6KTg
X0nyOkB+RKw7bCuYFZdlJ+KJ4AHFYm/gGbf/9JZXDrr+ZLHBfrBC/RGs+1jtLQuBw3/hOTYvkCsi
Ge7mv3MKA0ALkDThiDszDtuBR6+z/C+zjZNxEQgVd08oVHPSPss8FHWdJf9xhQvQWF3Q1je4Zvmh
ryPwgeMt6uuwapu8Nqs0QqigpQTddDTYUUkQFqUcUD8/F/Ad3MjpL1nXfmi4fKXAuQD06m/wNSl3
GYIdPZaS5hbXvDAM4Q2e8RaYhTHtN1O9D8DaYRWG4A8NXlkuYqt88sPxDWBKFOefnJ2DFs8NthCh
aVkHfVVXgN5ZxS7YU8qnlHz/q/4A6rcAKZbg28e5ai5WRyLDxotp6OjKHce2en9t2H8GTQEbXwJ0
mIOY1iQ8LdVSWllJzqTfBp1dGWsL6oomjvVY48wqyWJ9kkTwU+vKA+NXXCcXMKifBMq1MYE4mEr+
aySzJoJUV392Bij1VPXZL9Qg1bjQXRmsh/VBt579LXi57R79xTBR2mC2TiHqiQkPaMU5icw2XvGY
FHMOpUup+AeMmYSZsUAfffa40Y3AUyBMV+1Lcpgm7JxwSX8rHiu9LWcmcTUa0PApIEAtVxmN+cnQ
58OrkeNN2CmEJpuOs+bD5uYI/wWH5Sv+DDYTvi0MqxInbZoSBpO1lfOOXTBBabZRWQ8CliK1oXiZ
csouNuZYaNUe8KXESeaTBman981hUMvM1vi9S8VIOLl4U4rymmMjY/Rrwwwhem6gGe61St1IHsRN
rePx2QidSf0AqoZr8g2zkKygaEDYKVblLyD1WYCV6Tix81Z8vFhitza8IjhJ3lm5zCgW5SafWQMw
/WHUvtuJVUyHTpS1uLZ+owIyqq05LgseKpFmko4b5h6CqSibqSEKKzlVufo5R0M09qNZD52LchTC
ze6maNSo14mKNjwv7Q4S9LUduPPazDBKHVzZPuy3x7LpcBQT7+jCfij3uBt1ZcN9BA4WWJfaiLAm
vxhZr6p2+ah9MehdhOlY6ZU6e+JhiiqSXl9g1TEO9M2Ia3DPyNEjPC61/PjOIhrrVjfoS/qFdVJl
GXQ1o9e7LJbtMFYEAbR0pJFhjJQjtDZjKF1wyT+Myi4p/G45xmXSyssecjyGUwLLOfXtONpMayJg
j7Ka0gZjMDI9gC5VPcr3hmM5d9Dd+xnA9dYncv6p6cFd+du+Zsi1AjToSMV9qRQOF5VWqJ6IEBdw
xlxRj4c34TIla71a/vyYqq7M8L13p4ew3+R7C95Hq4Bcuri3LS2k3UgYOVze4a+9Tf4RgJ/uXdJd
Zrz4bIDxmMHiNhBC0ck6go/922H9epgr+gKqMuHISP3iGLAHAF1YvEvaE9y05UP2lWAONCC8scyq
Bs8rFg1qDQqI/7UtHZq+rM1AR+r/tNcA/GTGd+6K1RYIVJ84IBXz+mYr1mBMCBPmdNDtRgEudGUV
EdUKWBe0TwskbNl1RSBxSXUcyd29+oxl8ihAzYPqkvuoUGqRzN2n7WaWnF6TSJpGBbxwxBvA1JAE
/Nh7XmWdDGiru91q+NRSv0utq/QD5KkGVgGx+qXZBYijhsfukaHOuTCpFZQ/w2FKqOU/bJ1n7bZm
lO7dvZV8KtBF9eSOoeNRsHJFmrNCTi6TW+MxMDg4zPNYGJPlj/TJnshHg2ih4K2iRiIU+nRt/I3O
4brQZz6lkODxXuOBRiiGYRClbJF7FYAss1QyDkR0/MVYze5kfv16VpBHq4upU6lI7JxUOtiaD3Ey
0y0AYyEVjSTtd/bxdqF2Ye2vioLzMhKO2aLsbnmLpaxCJ3IYXywXRSav+Z0dU5J8IyO0oOVn/8Rw
NfZjn5Ls4fzAEiILAyYAxRgwqdvFJ3f7pLQr02dBvbN1zPaqf+htSpS8mmrldFBzQAMUMfmktwdP
on1Lp+VnGjElTW/wEdNeKSUJApkduCninyFq7qhAoDaZvlwYlSHD+6QdrNhZPuPiIW7QRdW3ZWYm
R72JP83nNr8LwycJPilEntBATRcjuVRb4KEobpUTOHfrNAHpus18dWyZKGWLoUrXIUvR5ue+EF6w
NDkgqAYI3pBEoYEAxN6kmK4Wn4izF5ib1tCptWt8mAleRRT+aC4qSbv8D2RFXK9UdFKy3mNo75yx
8oC38vYkjqgpglznCnhv8bTqjJkXOWzNC28K2hQUmWmzxm4qf1tagK+I1bgGnBT1hvhd3zBeexb9
qOjm/f9CJoXmyaxYtX2j07aYHHfs9tSWM9hhkXKK3ir8LiRiP1CbzutJC4RRLjiBATGdFQ1Ow7Ey
7eu38KSPX98ikJ/K5CNN80rgbXqdjnGbMoN8HyiRiwKMhmn5TLsAtchin3Gh/F6HU7o9eFaZvKTE
s3YZoenDFPUO0k5NrWI0YrW9AcUnWv3RLiZc8SACwlqUsgCCkh4WdlwsM2U6XEC8P/T5WKtT4DtC
T7ZJt8IoSu0RkZ7WzPTGbfUEO2vJ4EKGQFIlevlBQ8wmYLc5TAzhQtAtsRNgl/v4mjJdtKXNs3Hb
P/ws5vedygPOBh+v+2uaImiYkpzGhyuyw0FUwfMBJtT0HlnpBpcXEfTu8xxWjSzH1fQNEV9o768w
d0qKWnM0+FL8iAP2S8PnTiO/bON/fTSPp3IlF1vp//Agp73TZm6MU4TWCK5Zj20KqE4KJ91aCRJm
5K4VGNsM6S0PY87b6FXwMnpRP8wYlJRBrVS7425dZn2SDLvs13J27CvLjhPPzW0zakwZTChKgk4I
fhbnlACfWm3dOY6S2tBsnc5O8molzC3LSsVIc3oC9WRikKhX1cAvsMWRv8r3g+7oQYAi0NbRfC48
hEFvC52B/Sj2ECpSNVyJ0tlwTN7MXNOImVFAQfNrNQAniRb0yESeol3LoDqAIrNGlzdOz7H8P0MO
3yls5aJ7Dkv0ETOTIlcmap6c9P+HP4NkIrp/KKvrp2SUBf2/K+ICaJ724beCe4G6lIj6xYuwYnV8
sQNgdOq264VWDQ1kpSv8TNB8X02LImI4Es1zlp4YqpQAig2Fct03EYkl7AaHMwxGTnySDI+9erWX
YwQ6A0f4okDfNTMsO2SmMYYdKr7tnpspj0xYSmY5++Czd7xVjwqk6L57DLqzp+wNFeD8TcAsfnTV
bdnSYEh54eTQaITv8YOtAlMJKMlHGXEu7294vNvDiv6+uokCGwnAn6XN2+DNrLlP8cU0032tXlAC
xC+kfNNvixDWeDb49F8Ra9hzyqmhpx2hxXGoNb3eDIh0EdC1wNFB3rcWqUHpKoYrqCop+ykPp1iI
avWbX4q8oisOLV2MDZbMRQAIiMNxWX+KtTeZMj/fPDgqYXZBG8TO4N6FWWdFPLu0lev+5wh9wi9T
fiIzvbxuJlQXdRRpKOeGWwXz24XAfaVj5soxzaA1YXpQg6keE74Psuy3aF7dGZjvsqs+aaBwir/o
/ZErGcHdpGC35TcZOmnCtxISpu5a3G9N4IDydzTNf3yY1IW/GIit7o7VBFP9Nw1imUhfzqwtYGPC
H7i47DVUfz3jkWST0C3e9qxcmlXR3Ixw9RkhroXOLCW0RypSkgFuU2F/TKuRaj8SUnwK3IhAH9gn
uBqsXVBFszmrob9lDInJ1sY03k1K81lf/yhQU2r+pubSaIILojMmciMc0rCcZig7zKfmr9vZpRYf
lpFyUJtop0hykNUFSHwa0SsMfVutHGggDV1BZ3Ej3voCfvChQay3cwU6YhMhhVAtGFktXj6XDhf/
ADHw7snIS4Te1TvGsCpV6f1V0CE7OHDjOmUBtRNkr+KXylSMcxTg+XKvCls/3CbsnImy9bYVe0HJ
ITA+TH5VBQFFUv5hSOlDWD8BHLS8cjE0eciOTmp/ZrWGndhEGavTAeGieh3Df6wK1rdB/AsarJZK
JyflvP4YleuVNoD8oM2rdZfuP/lf8rwfZUzfaHqXIGpnQPbr+/7J8GsI5IveFn6THeJqpfr0if/p
lKT8iYGZ3u8D4vbyMqrJsj4cl2ySYv3lxOANefmR9HMtOQOk+dI3N3CEu7jio9CClrzktdkzO/re
wg44KQyZ93+3RcB08CsEfNQYa53L4fVjLiI+xnXo4yk7WTF6I8omnRZWIr6Wp1aQnRxnhMHnxguT
SK06cFl9A2hRE5sOFFoKMqWc+IxOjTrv2JuM7VPqKu4skKb40ccI9JpQmtD8XoksjMd929ZGOmeb
5R+ojaQxd6HSMnQROYauQsC0R+4+6D5xd4ysPPA2ehrdbihiK20UbRBY0Hipt3wa30yn7wpq86qJ
pjgY4EP2Fa8KZaMLAlANql3BcdnZIFoR8t0LKBLTBKSifgZ/30F4XjbUxPrfliScnP67/hlW/9UU
fM8RtBEEuM65rbgN4xgeQ4KYM8t0uVM5AB/rhoxS1uPo6EvzLvrnFFtozuHlv1TQKbhKCEU42dJh
Qb1slRJzJIedub59iKMgRGPkBCS3dVkB8rzq3veFvJgVO+6d7UkX4DPqPRko1ykwLxNZ+u62vruY
Co2W0GqzZIiZ0CIEPtwPMhDVKaiFRZ5SZAlbQsmuwuZnYhYNTdnnok02LX5FtVikU78P3o1W4duU
pIjjhw2gxDXlhaXZ7ZDX+U/QHuILZPHoCY9epo872kB+TG49sh+YyjPuUDCQ50pyQV7/Q25Goeeb
S1N26scdzhjXd0Un8i3jKhH7scEMr1ww2EllxKMe7bCQKNiBoJ4kVTKdgauIh5Hq1iMLS//i36At
bbMxIUWcLENFbvgRHiGU20mhCCl910a9A3oK5Awe5Ek/PDtvNQmLIKfFsAp4c2mksRYTVrxjghQV
GOalEjwGuKT3ydEpJRt4ge4hi+GuGWgirGfnCNE//XyCn52+S06m3FXTO/b6eD+bEx6j2f0UVmUB
lz4UkLJespfaDtVlc8nIr53Rc83yzc7M4t0JMdI6ZpskJzurZg6Vcb+X2SAj6d/cOG6E6a5O+mAT
Fku0lZjbyLUW51wI/sg77akh4mLlEhnuqqHYl+p4Q/WoivHawLxYbouICuEWyg5qyIw6SP/MCSyp
d7iFvOfpiK3GM2N79gOSTrgwYQixS0psw89NYgj5u9LfZ4ubfbnGbKfm8a50oHwZv4VRI/x4BbN0
Sojv/ndxdhEWBKArTS6h8hbQvvFDUhnbWoFXfXr9HPtX9Uy8sj835bKaxGJ4djajJBmHWXUBYK3e
2dZStm8xkBSqw645r/Do5Y/azSDiZr9KotdTMkvPYtkUJ7elwpu45wXjW4rJl7cUVLMn8QeB1XE7
6log2fCwmRbv+jaULl5bmP3itx5Cd1d4d3Nj2T4/9yOT3anJmM1hh1Srl1/q1wHrAqOvfhjtOA+t
kZ9QXCx0f636pkBTDFRZIaJd3LU80EVakOTHOoasvsdeQIu4Mheps1PlKg88ISpb91xbpcJMxBQx
QfXDEjulJq1OEZhNDl1FyAeAOEH3Wc2taAkusHjvhh3B0DKKwLPG7iaBGC81DzvmDA0LK9q0on6h
vasDe61wkN65z33uqfK/zjPsOgdUfxjPd0OphBTUP2QadPKogrDCV0p6hO9VJDMkR/jPBZ1h9jUT
NL8xY2FvZziT6+WtwalHaf3HL5mN+53vScH1ocikpaYR0F4n4NVEUaL4v7JoYrtIr+VxIxEXBOyG
vWwoHeMGqTL+UmHx8YAO2aWtoCOdytSsQS/x9s3G6dhO82KatD70maAxHkZoXK1cfG0wO7hSRbH4
o8eJWUj3J5BglMUOzbinU/inDPuojbJtIJHfCJ1g2/eDipIF1BfOTbBU7rFYQ3pVihz+UhxtDMhr
D7T6+RnJTt51xHIyqxA37enSdZuH5X7+/z3KhKUHutaEb5l7tTX6qKD9nuVt8U/DvMATW4snyGBj
zSDWgslGClus38RuA1J43TX/xOKJefJj1m8+gMZCrCOuXBhgj7k8Fie+nOiQn0fnCCVUVhpibx0L
D/eDA3f92W0DkZ6WFKKVlOUMev6vDeJnhIybZFw7Rb0vGm7GJS3FQrmRpGc3vg/Q95zoQvsrEE8J
kOPMMS/3lWeYHlR2sAyNPVKoIf90yU8VZ1hALvf11VMwjVzLIGcAHS2hlaZpDMEm7XRru/bwBm5U
HTcdh0IhwEiSRJySw4DCqACTqq/rYy+G7Z1/sSIj/4VOlX84svnMKT7XWc25+cfUpRy6EZfqBwRD
Fed0RPMxqiVhkYrfPmKfegqlj7Y9YT16LJ2rYA739AONnF27nZRImwDkiB+NZuGQbXwJ0dl6SZuO
ik7ACMLFfARAJGuLtZPF6VBzZntWd6se9di9DnCyncgSjVzJ3nQ3DBGH0APb16QN+TPTW9JEypcJ
CrppBTvn5UeuEJUgWc9RNLv0hxDSyQGxYF2iWJAiRJktln/LVcquW1ycqqgaFkUpzAEd7GAzSBx4
SxmmwvZOg8Yza+RCCdoUuT+Lb9FssZ5NaKjpGP63nna7cK5VVPaxZ/rqd/DnZfVH9iKhP0D7h+9B
z+L8roYDHC0GawExb4TdsHwjeYuAZQrN8xEfmrDwNYV4kpqFd7eMQcQDY8YYu1DR5X8Kus/RdIrQ
feoV/hQtUjh/0dzn/+Fi/1Z3vCePxuqZNyPVzNwbAx6lNiIO7RyiQHQdwUkyP9koDFgzTEg0laO4
cMsuM6LAT7oRinzKEciF//u/UPHuaOkJGpxZiMYM61bQf1zHDC2JZ0Ykfe2NH+688UmeDCJu9ZZ2
bdHkvt2Q+K5Ep/2Wl5gFm8vache1h5R6aseGOQ946eLhsx2jznXIku2TP7yUCaTY97hpcNF165EA
i7NbbTm5HDlIbOuaaEfBWsaTtuItOuBFk13ragaAhw4cpnXI/gU6uYlyH/jfSoOoh7XyjGJKjWYE
xqmYr2z+ki0bW0ZSNrIF9WBZxtRIcramIXPDdnpquMc/+QWN3wXhtjUP+0ThoyT4x2QctAmmnC8v
M7guJ7G1385nSGjbTO3eVpNaMekUNlcmxghbHl6Psy957TcXB9442PqQ3+n+SYYoAVUNcF72Y3+l
a8GDwXCOuYdeb721OmyrhnytHkGQXO5dqrE29W4pFDatkIFi6E/LHxfe8nB+vRJfpgfgXB/324Em
kbo4PYZqFjt6k8zrtCkKy5ovQ8JOQzGyyxtbH0qGnEAfAd7/9GMuqrAkD3gXpMJ1zrJr3sqikkiO
3L49E2jb6agx68S8aHvM3KGV492LZ4vaKNhEPxFiF+KTqLsjf7fa1RSKF9mUimW2B3L9J+M5rAeB
VdsvI9FpyJ1DSbarTwJnYvy9eKEdNJm5WPaC+wCnzPfOi4afeLUPh1Jq0AZaWgGZxGwreAAbdxrL
CJGbaPlzMaXl0SXJGeJzMVhH2EgVipRBRPZw/15VmS0QSqEcvXEoXMLDrECEx83CfpNeNrPwD4v5
T2nBQ719mCdr1J24OrIkSv+I21YzdqNMRWS2oWQ3/3k/FybjKYCpbguaEb/Qe2P0UzN7L7YIea1s
yxNhNzBKOXdU4Y2PSQXi2elpMuE8pJqZGNfC44dT+kmqimNqJrclgNznlZI8c2aReK/TO9jVOG8V
xeVGrMkhsg9WrRgNKdMWIdey8b0XNLSLj8CklOBMOqQ4wnsIkPLuw6WcL1tah/Lh36ZvhHkxgvqJ
Nkogd5HA6tbfy4YRCix+tziG2U1HlihaMX9iA3PpiXx1s03qeyTKd5lEC2bakowXDRy+eQGrAjXq
iEwoW6Gf+cC1GcE5M1vJWKgBRLMlgIYqTHgjb+x2UUOvUkZt8hwpHgYky2tjte3hFwPTbrOsVZmk
ldOXS4mQpUiDmypiGPXTY4l5YLrc/ZeBh1Hdfk3ds9xZITDWLk8J/Q8O5XK11enYWkZce0oz8KLF
+bAoBstIyiSXGnYZo6uN4aalu6WBskwQQTqNcgogpkLtSQtfuEUWaMW9hecYPj2eaju7t883ZJjC
5GgYSZJ05fItC+IjHkuy8k2+V5dUoXnS/RBDvLPi47SrvwLFCz2nC5baP1d7Oajgfkz8TmBQ8M1Z
9nUbq4Vp0T37ODUZJG/oK6EHam9q2U6W5TLybkbPaMFvoPjMaFQew6n1jJWM0RiowRUejhEojsWP
oBwscnaRn0Bv3LvSAnBQlNcgNSLC44Gb4TAhUFpVFb6zYPsDCAIeV5L8FPOByhKiwXbMJ7pWBFSu
SU2dhdPN++dhFp48vCnK0MhXxSwOk6gyZIvOhgBZiFljd+iud03q2EA1e4hZBFua85otV5tBRsGK
rn2Y31tb3boORXWJ9obA6Uo1dcr/yPj02wDBxM2/RFcZb1pAeQK1o+w840Ums8mjwCd7Oavr7GCV
y0Zw3SHixK1W+J3xKwlRRBRvHZMT15JsQhrBDnRuNlP5KjtsCj6vLIhvM+2YZ5apAh0blP7gWTBB
L48lK6fKkqEBH30a0As11s8WkjrjiAnI9QJvvt7ANk6OLCkFxlNtZ3TKTl9afTmlWv/0Nw1wqbVm
6jdk6dbDFnt9rCEYvPfdSQega6HbwbU8QSESTFSdFvWwBnsnVXcy5i1j4YDr1nkl75CtG3dusBsv
6Dx2a+ij96VV3Aj+AHUyCPOkzpUbMyBc9+8PGaYhWFtwkv/EiNUEvp7CcbmuOhSkD0wXpmLeFg/K
uAj8LBq7Adfn6Jzlw5BmyXIJYPnEbQ7ozJYSd3DE51uRzBS52/quyWyU4IbuQa/H6SOIfQmOpLrz
yEkV3Tqyrnsa1pGhk4zThqqb4GEuoxLC1PXo/v/BhIY2U531RNVk04DE8/5K94nSnnwrDpDxrPiW
F8S6l+FjABQzTIWM1fcudz/ndpChwqy0wVatdyXxPnY+2OOWgRDfFiCmShs+GLH6/VBT2xrKRxUG
JvG+3xU4pTioCnQvBPofroa+ec3Ft3a1ZoK1GcpnXAIL4URoi1x+MBHorxSnRhbLF3ApB3Q/njKW
v8MZ63Zoyma61cFuCMg3WYiErgMZbm54vLjzL2en5VaKSBN0CY/HonohYh44Dy4ULElQ8UXNq57a
FZ89D28nQhqP9XKTz09vyHzpHggoGEMfW0gMc+GCdE4numW5AUvRrisAFRgxb4u1zlAaNb5tZCCb
CPKF70dMzHTIv6qxg+2lz0TzT7fL1uYHBR3Hsa1dZcwZD6R46mRSUQ6ozV+PKzDYW+tDldIZpGPJ
sszcqsPbiSd83JVO64lSLbzckiDlEToGDvS4vEd1EtkU1WJTtBytJS/uD0LKeoHYHBuQ9It6Bnie
16c3icxhy9wiMKlnypXf0yBXhQLqlHivFWVMe6UkTQXLqEos5+RV5Z28L/xx4GQN+O/Vv6HXYpwc
y78zvlkkPv1Mbsvv4LIHxdyGkwgoHTDNvbLRWMVD+A1Lvm8LzOKJZ5hzIgJGBnJ0TYQ2xDAX/ou0
q83X2XTjpquudcKEEbmZ3TbMEkzuNYQWE87B/CxTn0PfLgpx9O/ZivTSW6s5MRBwysU/bj88Kwsq
Qo3P4HQz7gvaTGjX1ttwe0h3B1aFJC3j0mrJ8OKDNw7A1oW6QYewm00GnBDED051tQxOGUPIYBT6
lRDUbd9pYhZO/oRmqaNVJUAN6buOWB6kSZa4fvKkeMJpPj2Q9mGAU26xqOnyUL86T0OdY157Sx+q
KILruxMxh42jxaZwyAXunOCph8/bU0jqQyzMbaM397e4yiHL/jCz0t2I2dgUNnNX81UlnmX2Uorq
HgtEpV2ZJHVisBnRYeEX1hUTImHmznD9Ou6m+2HLKnpHVaxMtKGgUDXJtnNOnAZ7Fn9CwEWpoNK9
ReI6umrkiRxGRnUUfdeEzidAGJVinNt83rJjZr7RTNdNxw2MOFopiumGH3YkLDUl1VClkF34dXBB
ZZVs7/xPWyywceoRrQOeycJZhJzxPi3+PFqWxAntmmcV/K4cBD9BT9+nVeRZviH/x+YsRcf2z/cV
JeicuLq0HXLGspNeY2xUXTtKlhGZx7hGy9bejUGG3+20jVlFGlCsE5Flq6mvr9ENaTJFHV2UnRYk
kc7xKlGFBZiw/6cfgF9VoCunZbORX1sYa6Wb18wUkinIJcSoZiuVu0K4zJ81jJGJ9QDiEpRAK7W6
1fMUQ1ITa6CUXhVyVMl4aj/LXtJ8m0KUnvqXxxBd6RSj5owYwOChnlkEexkC6dBRPVo4/L5mFzce
H0o35qy1LqCuJ20DtimUtCKqm6RHGJLNUGor6Pold9WAuFyoVw3iBvmsF/oL9+kpIvaR1QZ53dFi
NgL7cWnR/HxOryzPpanLMAQG5rJWiZp1eq57PucSKPVRDdfzUUo6A3+HZkzxmRQdHNJWQP8lqO80
JHzQElcmKJuMSAD+iEd10tpkjhFvrGsL5P2M7oJFH+hzViPEzA/Y85wv6rtCg4E5ubMI8UrYPSpP
N3xUwkiCCSNvfv1JQk4XbkRzvZ9pLJv4sPPHPwdbFOMW1mOf7p75RNXlXKIWJ+OXCHmouVOJyaQj
vGyUoPD3LwCPZc4emDpDtk7dwaz15diDd9CbD2M1/9bvwenyWXzqaXcOKhY8BrWhHC1KXS9nEMSw
vR2fQQzf1a8iS4fl7RzwdGMZVno2sszzKrajn+vijIfqdgO6EJkJhQW+zsq6hsQuFTVwXLH5xP99
bI+e+RL1l6jjVHcdxzfyenZ5WIMvvFPUn4UKPx5rVAvYB5IqkhIOl6EktGDvuSS7APP6sliog2le
LS+106xP1/Iv+dggIqtMz72jH1AcyCt1GFKO61l+ceYXzYRpeWCaXwsuUzpPaDI4G3mjDS2ppGt2
GEoRTpH0H2yCfwMTv6IDv/+t7s4MALBnLMRRQ94yX9U7NWlntsghbSILqbfmrirn9uVKyTITv8r2
KWe8+h10AnRdl+yeUHgWLu3At5VOM37Dc549GxtBHD+LZaXB/BFmQLnpPJb9kP+dXf98wKE27U6q
ueyROyofvKfaTieqfEa71ytabpnQRG7WTF9t1TOXZh2lY7d4zZ6ZBbQ8ZY3l9Vlwz/DunsPBuosf
aZtEFTGsO5fHssnhHqfeNhRdPe8ac5MMpwLkbH1ng3a06H84VkkCwLaMegEudbnQ7EpfX278RGvM
XsKm675HTBED5AsyEOnQsh4UC9GgXGZz95Wx/W1LKhyW1UUG4BDhmXCZRBRsGoTnFfNNciOV2vD4
Spq5vFO1Ek/XPOmsbToB12smUqXz/BhASW02wO1Oz6TUgp6zi1Srcl24ZRyFkuHHxid3eXLF+YjO
F/LLl1ApP8MQztwmvkDsRWF6yxU9ytWgsFrDRAb+GhBgeVaKlstK+//MWfxHSAa1Bv+2padJtjp5
dn7jAr8dIE9Bui3LRSEL7sFHIFehNi1QDjynhd7FukFRIRx/nXgFh7RqBmV5+d4qT8rAOy+4nKyz
a4d+s0ZktDeBr3ahawMSGTDK4itBADw/65mDblSMtsuyKwhUQYf17kHAqobt6tA1jriRoBR1uona
SPOWS9T4um8WiACgGNIq/goqT5MQm3P1ccT6x07oepIiz6Nnn1o+CYdo05N3RQv0OAMkR7Q8HJoA
CvAu84GdAiYTxWCQ4dqWFNyWq2JRAbVbouCADMfVe2pnH8HI1xs6AHL/FkzinvaFdC7KKV5JBqOD
okXQxmYFyjud92lv+EAL6x8TY6m5wKFuNouAcEDRh2E1VtwvfvEPxFfyGJ9EGwt2hE8eOa/gWNwv
N+Vsx3iodzDsXMe5KcuGe5K7GhMLMxFxShtp9CNmJ36hEmMFit1z9brUiWyW6O7NNEWCDkh9nP4B
L9h53ua37YWDJKjWPRwUtWTxqztWALRiXB4kBwHQd0Q+GJkEml2HtI7Kd62mpW5uimRuaumi/qEx
jsDyTmBv6iw+7+2xiwp/RUTwdIgQhDv97u76+vnRF8ogfPorXqWdkTilvS5fV6FMdWk1Qyamh48u
SPcw/892zS8MgYDj0eqaD8tllIudlLhIy+Cj08MTEsroNgmsv+5Z84pfiGpOIUJIlQmMPEIo8YdV
yI3Ht0bxw4C2ESvd8QRClOgzOOCk+z/EX+SG61fcqRGXzATxOknq5yIjtom27z/kceGWfwoyF2UU
sLBw9M5w4MALxR6VjkElbICXzCJjGFF9JTpIaJMoIKsB5RNBTmKhU8iFxWewP33dhdH+lj9rAohG
XTP8sT/tyjqaZOBn/SbSCM1v/8DyZgx/tzrXd2T2GfF2NhMJcMOwLE6cnA19zM1UCJ2xkk81GzXm
v6sbmHoC0O8JFlF3Ay+AX1DiVOGvyBYACT99Q/MR5sOedNEFa9DwUVNq0SDoSnXGpI9L+m4s5k0/
rfVuHLtiCRldbk+n4kvl4vJ17F5gQ1H8Pjwy2K2zXHp8n67qLtd7YU430ggh3+F7Kph8+fSCmRc7
emyqOU2SuK+VQYdC1R8vIlbo9tT8zDd0dZ4ezxAlJ5a0NI8OVpOAH5abSD5ylZJXY0dPXz4ro1dm
vgdPQbu57GnZh7AGYtx0NtX1YJ2xmcyfwpf1Oi35HzBqV1gvw8bMbzT5YW6wmZmMGqZg/3Vf9VGA
MaOeCXEJut97P9VD5prcXmNBybYnkwWBG8pY3Td1YzdDP3CmqGHKoS+ygTLNbnvJld0FGDvz+VGO
FrFC1FCjzxuKZITL9TUX0mBOTg/LoTrquzKNNlZywolP49qD0xEspL7FZMidO6O9VACY/3ph4DQz
Rs3sc47JyEK/BXgjnQA5yZ3GTNr71as4R9tNLJlArvJT0Mzx3SpiCMxveVhfVfPh0PMXmVQX6f9g
wDIGPHYaaE9RMo8sshCCHyqMMlPTBaRyLs8BKdDVGmhCmB7YMgnX7T52KWQf3lu6b3jRahMg9Otn
yRu7YA5VdRP7BPFs1xYqBdGWgay4HlEkel2ZscSDwYamBVILtmDO03PfocOlldl7oltKsXR7o/qm
43Rq715M7dwgSYxrVGyNC/1ZblLhbz+YQTn1tlCy2Q84qlz2iOL/KZwrdk33OY9j3vYgirP+hihJ
wGdyoqGdqv6ewwVDQI+kfhrU0YqOnLCFq0vXjoerV7PkGgkj19T0zT9Z6LU6n3LQhhL/6g1kdcce
rh+gJu4l033R6KrG05zlesUI9QbwABvEd0voHKQHXFZxmRYmJLjbEwwMrUAlgmDtfy+jWyKH4/kO
+g0Zutmijsm64Nk2TbqLlbZomKa42wr0kp+BU/2hb4xNqXzxJtva9Ly1zW3d98m+7qImVT0iDZ51
KyzLAiJbnnp4L189r2FhUclKytfghI85wsh5QD1GhjRR4FrG5uLTt8S6uSxWj6jyErJKxrGwYDzB
JlSCIfj5NAIHs8VbYyCeZxNkiluKkuP2Fyp7M03FeZA1pc2AxLQBlSHSJySHHS+Ttnk3dPdRSAsl
kDbS6HrhWmH9JrwmAksNLIaeP4ScFweoXu2dcza+KEcuPT4LI5osjem9ox1CTIEMrP+pNSlmvpfF
eovMgqOHRNhyWACZ17d2gL0AkyyRZaY76OoNr8JryIza+qyMGSNhyNZGNT+qAjX0RzmSnzilTFLY
14E6LT6HdJ+V8vmZcUGcnZw0Y4luUQ4YB2sSfxUA9wBgF+uOyGe+Ipkszyu8R/6wY3NkxHgVptaL
m27Z77EOdslBCGxp8csQ6hsKfXNDvjhRwGO0T5ZFioRC/+lW9ckSTY7nEKCHi3eN6/lOXftHb/Sd
cnM2MoTXprVjnVocilojn3vyXWd48j9c81kgyGyK+SZ9wEzQBxaS45yHSBwofOCw2Igl1VfQ4nPJ
9BBXGsVHQSIdVLL5X0FObTld0xFnriWhXLr+lu4bTKHwpiKBQBvzB4FfOqcIXOFnacm+pmLit6+E
d2wfgKvPLqVehwpd5y7rXFMKYY5W/CMBj4uwR7uC99ZDxtQWlCu6htIzPW6KxPLQ47gwXiukgGTR
2vLYvaynwEUzzY2CwujVCLGT5oWkAghcGy1wkBhU9s/er3RZQn+/pXEnUqyPF5GZ6Wvn1OrSWJcg
R+Kg960MCOjmrzBTuUDf3RrLvMtsFHKbJEeXLzifvx5Wmd/Zc/H4doJmohgUjXoBJO9VaJpcd77f
fMuk3wS8pRLakFdIaWkmSUC/sr9NQNmv2GRCGoCjmXzBT44GHgkG2q4B798md3xngR1MizK95cDM
4uJ/hkE9K+a7VnosWb4XxwLUrcM4xuma3eBXi5uCLWiY/qe0JsWGE4h2lexMo+mFWn6RXeWtE+NR
qZI895rLYF7r0kTxGHBGY4L/pwY/+59RWMc/YLajdbaOmcRaMGjir1MT7T850i/9ZeQyYG5rtFk7
kwh5kTudGwP4pZjz/CsQ7DS0p5Ha4ut0Cd2z1ryqLzJvD5+hQlmT7I0FrpBasRjqGnOIS63DqRA/
cFC1hf7KJP+ThMDKKJrDsTc9eL6hW2UFI0WNs6Foyi+AuAJPge0XSVJamJnN8v0QFGtN4UjORqRM
uzjTZKyx4nbSDxKP3ViBhki0jWeDinbV04M+0Q3gM4+XbTPIaqSH1RQasun6EN0htDsT8Dxz1vUX
kF+vMX2QavlmLTgUJ5tRTOhpFQOPrK0s2lFVHYxMtRnCxmOx4Obcuo/l2yRTFeUpe9knNiDIGglk
zDjAofW8x8rxGLlE5k1P+M5HJ3ZQMPijPrh25vtVFZ7Rg+KvCgQoHfsu35e7rhmiD5fb40DFKceQ
r1qvMP5uUqHJfYf9kLzdct2eSJoBCNpbFxTbcYZRMUdmYqPFha70uIwkpI7BuwM+V5W1psd5rh9L
NG8bEzc4JdyheTUQgAkKYDkjx8sXtyFAYU6O0hDAFDEPMmzmVwK2buxN2M2WWAMer0t6VkLu55IJ
3aoK7D1pJyT4SMBZIQsEude0a5eQy6/ravbVBrwa7upfKtKqdgvhJtLflpYdUOXvvbWDTW4u8QXr
D3uQDtkDbLkHFHhdIS5aJbEy/+AFbotu6blyIqNehgmUjUnKwcQ9ESiofbn+1bZ0XSPWJv5jlxSj
VQt5gtl9KpgEWxXB4ioinOeORpXyfK5Lt2jvxd9ab0V5c4ggzZuL/iP5zV4XGdXVHVG60mi4zTUx
VjmHfo0PhhkxtIVfD08/FIzXmjRvwiSU1Sml9Vb0XQHMypzddOWJT9mFjUjAsOICq7J3ceypRWRu
UCmIwJzm2OfbQXctJjTrnbmtFlTyGlTgWur4kpW4dzNEfytmbdQ9NaBvRtjFBTjTtPEtvDY0vz+f
OIm2WIMpKXpZ/UO4AjLIDmilz3dT9v/jD4AWPe8qNiSThWUNXQ3wJWzOSn+RdHuuLvtwYwN8scg1
zFK5SzyL0j7i5g8Lk3sbBWyyejhi8mHvUB2rZvrUBWwiw6Puic+XsCxHhh6/PSoB+Kood44/U9hA
5rxhmtLhH7ySOk/pskox9vm/BpaIBb+1WSnbOy18LSZMoPdlHMZb9Q+LQYlkRtz2aMno6YUPK1jt
a815tVraCj+77H7nW4samcp/KwdrJK3/dSIugYVZQTM6e7Hs1N12Eit4H6DJ2u+r7Um7usvIHyYs
k5kAY5goHkhHEYzB1SBvW8ob/4nUmYEfM9e7voG+8kgyM4Xu1XGPz/HYZXexusP0mu2vDbn/hiUf
Q+wfYqMBM3p806lKdKPXwxCvqGHTwvEpy5tXqjMXhe7ZtCsRHdyUoXvqaU3kPSelIv6U1gk6ZooB
dxgTDBuTEJToPUbo19s5O2BldVU3QYypACfY/u5H1H/CHk+6HMrtAWSAv6UDLmgvsK+2esFTrtpH
0PjzsQKpzSzpMBDVlRCn/x+2hSeIpShHYupZGXqpEUnlIva3jr2IZNkdx2xzlbpSgl5Vj76qY4C1
XBZ3afxkWTwCAfL1SsQBHdVcn8054CINPRr0r23GoSNC98aaZn1jvag5hhkXUd+Cokvt1B+vBER5
zbF9kX9Nw4nRJwnvVTx6a7dl2CbDrETgNM3mQgYMDhibPnHsZGjgWQQNPsHEcVLzuZeWnA0veU2W
Ye1vEUAT4JzygJafU+IzbxQRLrUZV2q/rYatFqaD93tvcuyRkASwpdlF1sgzBShtvIO0mw6AKYqt
rDf1BYPiyA+6X69ZpNPTwF1Fz474h/J0jtN5kbFs7AM1nNHCNQCCDYHmfuvaWmXI47QFbqowzvhu
KyhVEj7jRY+fm34wumu9l5fSIkgTcV65VmfeJZlmzIchmdWDOi0ldNfFw4OlKtvDGrJS0ufD5bDw
Rxk2tuxF8GIb7Vc12QG6d+x41q4odzVnDGxsiBtadwYCVVzULW9uWak6uXd/Y7tIQsRQ5BtnqSq8
rSnz36fhK+GPhU5aNVrzdFFuoyZeoVXUFRlcZWDXaG1tFIluuF5clOfHld0zHwLIXVzpvnfURT+P
MsEOKWFNTYZTOhNIjjibqwtsmlHwVsiqN8jAONddnbc0aqTIjpYuFuXAf64hPNCKYyqpvBlw4Fo4
kdmVTAdyu0Jz88N81mpCkA5MLR01YS7sBL1sJOwvsjP2MaIqJ6T7dKyUxscOGdPMxApnlKIXG/ux
BraET9XtnrBNrXo/RlKhA6czPN1XIAe2G2fAOxPgKNf4CznOBCekPSUf96sQ40uqxOX8bl0lJWci
w2P0v3+P9jhcO7lHnNxZi8n0Mo2uMtI7KQuUWO6X5XrggV5+rC22QBeKpt5E+JgJUcQPFdV9EJiA
uuVUCbyPE/jOR00yzus+x5A5m3gmMmsxKGEBQOofJhahnjN0z+gap5C3Mwi3sVxMrxx/cVz0ari1
csU41L1Au1RNv32suy5OKo/tJfdJhen0UaqWnGwmGQQEgcnRFsa8ASCeoODZTUgfZR1/ONpInRWL
nBcXFz5iU4+9Yf6gcNS0oaUz9HINo4K75cz1LGfFjzPsZnBUaRjbsI8Y3c12Wa0UxIm2ti7HRWaF
PcHrgf7J7UJwE7K7VAR2X9U9QLWRVMW7lfcf+OYNpAtmnMlHGVdCIYkkCnkAMejwp4hF6fk4yXZn
YJ1lwrxWNbPxN/AvvbfMN/1rVppyu8owVyfG6GC98Zm0ilSBWgZ4HzIZYMwfr7tnIEpFJ8DxVsQk
o9tpp2NcIzjMQrCo/r7hOxcuVCNL70V1taNV5WX61yE2F+OR8pfBH8srNjaiLXr+VHeN60Ki8B96
tstnuNgr2CrQVXZEZ/Koa8mY18Y0kT+AimcNNsKxxBIIvPuytqW0r5K0vBDvSFlhX/NypexXQHiY
oMUeUdoPtOY+y0rKrxKLXWkZgBoG55THRgwRTAlyU2+hQv1tmKsOy9bIGq/Nyizm++Cp2+VsJfNB
RMHTgkyndeKTQbM6ymlJWiXwqplCgtIS+LSBgbMr8Pt6dkD0Hd7/5Cx3hy8Dr8nwRAgjovmOsIja
/yhlzCd1PYWFTwVWYTRsFIhrIV+/fLr3J/ru1znao/Flvrek3UlZZTnG6L2N9vOmQv/LbM2C5ZCu
fa5LZLg25fhxGb091J0OxYQYGrjbUNvhzOeSt/K7HWruX3PCKFvAAtjpq053817P268mpaxjHa8t
qJy1Qs9Gh+JH4MNhTt1l8nk3lFsVcptZLwqfG+tp8PDex24SREAxIEqpU6gt3HvfK+91cYO47D9i
r3AxdtJ98Jor6x6e2fSYzt7qbB+KNg+UduLocN+9wkbZ2YJmBF1dC2XhtW56IcKQoQltv0wLXL04
hHuldDnxSOkXdcnbizZkJEs27N03FjVZJyI61LNx47UH6MWhpBPRkeXF9CJqHGyclDcppUG6IuqX
NzhXqIGz8hj0mEuTHrF5mhV3/hcVX6E+rhWqfVAPPQ6es1QFc9Bkyw5IQOmfCa76Pa/J0Hr0o5LM
jN4S6y+XLBc8WjPwH0krp6QZVdbejG+fXoqxpLTEtDM8SGUUQkeFbxwi/hNMEtctvYsaiZG/xzEV
eqGvRWneGOdB1CbixHw+SR6aT0lNb7v3EKzXjjRM4fRqZEDi/MwigdfVPL7HO7AjGbG/gCqpzkuG
N6Fj1qgZW1zODR4qsAjQzGSHPIVwm6MxC/mkBj2RRQGBUiUD0e2g0iAjOhDILDW+Nnvkfjbz1LsY
A5zGoreB+lYVJy0op7i7gNXHxkhki+XVMPAmxKQlfSNPRDuvCL4ZCwkpZCYMuQSpsfbKd2epTCaO
Hs33vNZOEHiAWFgXYpyCxG6GZfDlII8IGuAgFclNRi4aahyJk4icQx/1/i94mYmImI0Weq9IOIVC
1xE509+adhbnbh6UXi3tyeYY1OLWtEEO5vLL2utyOBwcCUX10Tu+qbIeDapRKyizRrDec6iLRGom
wkjkNGUTQ3asZG2yYB8tsCJXOJj/ouZUStbCF3lcXXrQvvKhz4DD3HkPR1PBuTeLwsGKltITOU/M
PhXqY5drlycx3HfqIrs3zVVthc8WBdZlqJjiM6xyvBsVjZVOMOfoo8lGHLoVRUbgeaGQLs2oQpEF
xcaPPWeIBtZFjAHekDGYH0Aa1orwCg+swX0sdbnnauhMpx5iZ2pnbPHAot4NHtJVQgu7nfNJ/6RR
ilLUW+m3fshCWj4bbFWMZuSHfEU1wC67dOCTMliZpv+5aKnAMyyhqACYAkFLnFQqJ+RNweDdokj2
N2JrxPRWK9Ts+TiF+neFaOhgpoTYO9zjuDu5a56xt8ZmsKSmhfgWsgHlEacMN/ex53rFenDEpFLM
cRsMbh8Oln6JcmJgJJ92/v1kISYel6kzBLD2jMweKtX9BjAfPyzzpCc/P+JENmjf4+reCjtWqooj
UoNBDk4A7xEbBMFSDEhnSFXWNzlrpCTyJ7QcyiFU2XknPqkgJTH2ftaLfgNvd4oBVPB0i/oUIH94
+FZbbv/R20EKRk+IOy2UeqopfbMkoteAqawXNiQ//Cc1TkOohoylQmIHREmA5DSH8jbviKi/inc5
4SVGvSLSeu+m25cw4+sDqQ/ILST4DS8MygD2Q6NOhCibLiH+iNObYyBGrCDFhAQEAnmPZUxv37BX
otpXFmnqSd1skBURihZCT5CBtj0lwzgZLeHVmUBAWjipATps6L90d4RlAZhA+xuIq2/Cf2A3whau
ej5ZfXdtUTojsdx2Wg+m+uOHywuDnekvgnZ1e8BjBd/EWbICUchKzWE2qgCLZUMkDHrtsV3P3Zm0
6rqtiFyQzTBrXE2kMns7hR9yPF15ql6vrhwxGumLZr5+l1uVJ+GFJCbPvncJsTyfVRzxXqbJVa2M
F4l0RQ8XYmOblZNzXnQITZeCtuByIMVRBxi4le7ikb23CgN3y8fGZ5la2CVNu4fUljFKWR1Y1sZc
ryrAwdrt7rNuIsTgstaMUAQDQiqmtbrCYaZ0H9mUgAme6KRHfFh6ONyqkgYg/vqWY8E5m9k5gf0B
Ox3xcwqjpYjERPDuzn0z2toBv7gSXlVIClELKZ6ybV2Y8iFUzLgE1cxHOQtgYU99g+mH3J8JBucT
/JFYZJ1EImYezCDrLIAfR3EPI3pcyTB0E6bRBZXF0MSBSZjLKODzBZov1x4GqBiIG5rUD8AT6LLj
db4VOXwugA2lJiXciEvdULdJVV+jHl8tHEO5GvNsIIXzWGw8Tr9s0ly5fCK3ubVK2BlKlJQwU6cM
kaC2ZD+ZvBu3Vpi+ecpNGSVrENzTwm85rrROFYuYAyAn/+kYd1KAkOYVjShAUlAY89MjlG3PGWeJ
lCW83XKk1d816Qhb2DrXKyuvMOydca2+KarUTuHX1RhcxtdLn34x39+J7KOEsVziLH37aUrz/X/U
OW0oUw+WmJN3+tDXP62vuRyqHJIu4BGBpXmBKeFKde2Pg6p0Nz3ZDvm5dyNCDqTUJkgvXiE4bY5b
pJ7rBUIErvulsPfZ+Wr5BZAVqEqRKzoRsg6NtK78FeArSXySRkTqp4tAtL7+CE7Iz2cdDDgNvSxn
ZKaJWbFcL/C81o3JZtStAEqQs0Uwh9tCi4dasXHFnee0BvBCBH77y1vPz34EypOg0qegwn5BIqku
B8JBZ3siS38lsZ6Zj057pJUEa0DwTjfAEroi1Tgy9ldBl71Mk8fRP0EmN31Qslnh5Fh3YahuErz0
U34hNjq7l4HvyYBatVb/Gw7EaCSfDCKyxeCBoNU8xAxmASdJFU0ShwNecsZWRZROrTbfJyjLLkUq
zSiOIAcQaT/nwKqNc1L0Fk71dhQoXEf+fojK0jVD17vAYD8HuRzYS2xv49BmMvJrXWGXV6oSG1oT
fqme5P6OmD6SJ+1QfQTqttsuvfY7IolMcTMcKbfn80Q4Uv/UmzjLZCbuyhYKEy4Be58kJMszdFef
I+20yoPHbJLaCve8LREHKjkDpANZivCMUtye221qj4Cbi41jGKeR0Cc2koIuGx3nzdBoORHvJH1B
Y4G5jvClMvE+/xPnQPeGZIIXcXduL1V9VOzlFAc+QbqjpIXlYmQgwKSjlCoM5yHwRlXRwjUS7A20
qNs/jcnwmZSJfgM0b8kSflq+VV/RmSj5X3iNDaGDjmkQHUeSHKRFhjmS0W1n/NRQHK4GPeiKWMwb
agrhde5nFJqfFmeKlql5mGpAReJtVURKiM5S9Ez82XuEyB7K50KHDeNPwsgPRhFhKMNVbBeCXNHL
pg0rCBSLhbIg7Qr/5ndJ1uy+gd7X4INqdrXm6T7OLElCMQz7qyOctJQbpQUWfwBmXNu7u8avNVM+
HD3oDpEnErfCdbYFPoMYHt7ShRKeGCA1iigVSs7dS/o8o4J1rdt0TQKtLSyYCxqkLiJT1RZ5Xxip
f6qJuS3nJ4XO6raaZPiYDvSe3R8jo131MqIfAh/FPzBCTd9e06dxGqEucjRuQi8QthdQgNhn8Qj9
N5yVQT2/I5DEx5Ki0Pi+BZe2bOdyNFA7AUnM1GnPb8Pl5DX8qNmPQYQJos4iS95T7iwK3QjDJkLs
DyiwO3IwtpaWc9uBltxThcPVEggF4VKoGTmVCRjr5ZzsQ+23Lcv2AGQ7uhJgw5h5yK00SfMmKtF2
/IwbfBO3/rG8BcsOfMum6D/bnQFslTVyH+KHDxPoZEy2n9Po/nNoOUXZs4M8ThWQhDZEVY/kI+bd
JpXdmIvCo4U7E9Ch9nzFMJwrSblztioDgBiiycD0o17SXd/z4Q7NCHpe87f9EaeDP1yfQBNJYk0b
pTXI3G5PkAjf2NzBqRIhFeblP1cd3b/VX+y0F5aRc1BmrXk6LW8XO8R5PIug0b/n4hujHYKBW2hL
Iagbi71lMsbbZbD4HtRdo3J3iyMIaAFh3ZFPKiflGBCm8CdUoSHNkJj396HpKGFYnAhgxqg3Ooqz
YeY8k8//GL2XjyOmCz3bNXK8rPKhWC1UdD0tTlD2YP9hkUSeoPikfeKB4Pq8nln5VJkFiv1ku36V
ifaJTyKYG66zEYppj3mAxK0H0jibq1DekiepcIiocv1BDV6RxeJ9axZBl4NxQ0ssPrMm8p1JP94j
42FCjWDjO6E6KR3ZIcOxca/+QUCigMiD315Gp09EY7+UScuuxEnyrH6u5fbhbMVk+q5l/TCsh5X5
VbhOAxVDDZk3VHHgeVpGuBH8SxQAru5aoQYcQlCn85V3fS4EneJpWLX7kRbqFnjbyeyTR8RCWZNn
VMs9BriHiT87o8n6fuqMSD/GKW8kbXv9CmHfC0tEBsyd+3Y8yxLqs9ssiDrPTmalAe3G7paBE5TW
JQoK+l1N3ijAmsidW/j/TKwDlXIeBEvfiVlrbkjJlF7y7ZxZuMWT/dItkE0tWcj3U92aRIwyK9/w
m5sFipJ7GzV6IZOOZFJoT3SKDJFrTHj0S84r0HLdLOTM8hw2BN554j2Koxgv5WJLmaDdjIxbkszt
Tu4VLFDbtG5qRFUlWB7wlDd51u7SCqA9kRccQG7dPPAa/hmUYzl8X0x8iinLEBD5o+iwhambz6sX
F2hhNg0tfqM/MU37xfLb11tZ/bCVEm8ashlYxyG/3FO/2fx2O7jG7Ggj+W2x75Nfg/h+9/N27+T0
oY3RfDfQ3Hkm3sbQkcHz4Pt4XmgMo6s103mcyWZ4v2QT4+jhX4c/TlKv05i13JH1+3HKUpzEX9ct
b4QY8pDV2343neR5zqCAA6j/ywlvwJUd3w2WfZIodUZHk2ndrwqTdX+N163FmsMxG4ateTx0/F3w
FhjXXocQg3O34QPm2HDHOk5sapM+4hbUWPSFs1qINMv1KbUbjvodWfWKy0aifDzbHjSMG6CJzJC5
PudGdYAB+cP+JXoSCITpEwt4ESai/vN787OZkjSMuRbIvTK+jq0PfsuhbDpVLK/DQAzuWhpV2OCQ
AZJRVziA7sku0Tus9ZA3669sunX6eOImFn+LvCOEm39Ip5SdDr8TByTTR/eQLp78aLchCGKSAQQH
GBAhiFOgaJzOQgAstkXRZtji/ejHnRCYKJqYNSMpHsZ7t8IXUyLVL2q0cj3B7VdomV4lwD1uQT3k
xN6E7bbnwjW35oREM866RUR70453Pgg/AjbsDniwDm+YLfXrJfDlOKHlxUANtaaxqrZEZE7azty4
uD3FbWOGgkU/Di9LOD9N1hCNw4jJ1clj5jWJ2G9HMjZfCkgMrAXZvFKHLE7o9BxfaQNCgOPWTh1I
j8dQvJo7bn1HN4oqJyu/zUBfXMWnVtxI5Q/uZA6IkiDslZOVf/j3KgKKSo+01SRykv7Fd5rpNo4k
ysPppc2YplWoEsDcFZwnFvSH3BFCghpVlSctZmO1APWE4cO4ZFm8SWpXdput93a7g090sd4Tr0Sh
B+dj210daEq91cOCAYbybAWckqukd8rTW1E9FHgdz4UaT7BBWB5bCiZUdMJcPf13b3EH0xHBDPOF
Ycq2sfTKL0fmn27SKHR0lC1j3DFVHiYTly1MKObSxpiKLdCqK6Ds2W+Ci0BmWYHVwr+uAmlCCKNS
W4OiSSj/+6E+r18PSMiggraZtRMPl0fXAeteEDNT8QVNjXhSY9s0/V5Ew7hXs0njSVg83KVLfJr2
JfQPit+JXfNImpIBoQQnyWDWmCkZZysVReF5yumD1DA3x2W8NLKHz4gqu/G7f+tKdUPXYiU7OhAD
qAShUTz6fEkiayWUbMePF/ZEmC43Ad/D0GpiC0q5umwdH4IH2jsnO+iyzCfmfdHgVyn9LHNW2C/z
mlKE2wgo/HoybYcyhXdp18kziimOZJQsSvCMouNCaBY/doH7nnC1MOK/ej4JK7zEwR3XcVPGccjo
a3P+omKZZiwiEJAtfmC6gedRu2/k+/nqAZecgOhByO7RShYdCbcEFqYmh4a3jxKYAXsnDUT0sTbM
bbVPgQRlarzrO3iHaHPM50p5RER2fZXDGuIcpWQZ28QXw4223bFJjpBcvwn3IVhZZ1OJYjjQe11m
v26zIqQzlgByXCyOHLWLCwA96bUMA4PVsZW4oqNrsTxdjDkE2ueKRQNn44aA59VSVdc3erORm9F4
3pgwpDQ7sRxn/uLvPDQ8J/STfWBiUrAS1zTobE9ELDg7aeiETRStY8f27lZoEFy66ixodi96GSt9
e2DO5QQ+3rZXspfycWz8gVWqbh2YpqdlkilbCsrvnamZTCBnhFOyZ5/CtFXeQuwU0w8u/JNH3F8n
r/WaiFzQ4ccvFquYuvYK7n2VXR1002ak1OYlkYypdb3ynBPTF7M3TkEJYoh9MAa7qrRQptHalS6F
qoZ3Sj+DOJoA7tiTVJNVhlJL9GixuZHgjmZhmlCLN6aedxd7+T/UYdFmpZLFk+H17Ai8jqLWZtSG
LAZ49igW/Y7sDnYz0gSylZHPnemUQhFcS9XHMwnjo7j6A2o2D9georxdWUXub5YJc4DOn1Ks3FZS
YFyxsxsHd8PPlyDJ+TbWNUOgqGXodbNJKrl+8cXo7Y/DszLc9mnjbBUStawPeElGBHlEpXvdydPy
MrtOMZYera9wT0ujBe9bfqv9eNKoX6IZu0v9bwPIb0zH/8IoeyFrDRVoym8pBxOf7XF9kj3QzKKe
T3w23jsQFPzipr/SWcHXbh4Xp0hevbODfch7joopi0N3YqQC+jtTce/LN2whoQZDr9+ZHHQ02E2a
KEc+us34/naHAQ51w97LlcNeb0smBMa1wOB0uTTON/N4PKZUWyuyTBs4BtAalhA5rp+wLf34LK57
woeMULVlrHhcNd3XZXHnxOhxz618y5IyQRrVeXm1Juo2n6xOYxJDgTUjPAbkqoabrMSNbMfXa7/S
LDGfp9ve/77OGnUFMBsRt56iAKsvxvb6joK50977ZYUQCLVNOr8si96qivJGDZS2+yw8veZAx1qJ
5qsIEd+v8UWoXkFcw3HIB8n5dg2J5rWG64DfcACk/i2AKa2HjJGy2eHwuJmGp6KFhlNPxGqwOL5G
lXF+NIS14s8SKVCjjE42OSmUeCoWf4oqXqP0+RMInR0YfdpKgjOdTRfbxpA+U5fyS6suYxrF5eJk
6hDhMqfGveAGFSSQ436yxo+OK4WtIu93lyYS9wDXi31JGey0RoUPV8+ieCWE0Yv01pJ0Z/hf+DYa
81tsxpQFc6Djga8KR+Z6W0J3ii5j6x0FX1mqgrpNe4dkX7m+aZj9Vyr2DljO/25Lv0zFsTFEe5mx
KOkkl2pnt5myKM1XD7BI4LwAHFPO7GlUKp5gCOQck2KJ1i9/0JCpH5mJyKnPZ0sQt2XfUuRahq9W
ulKd5THeICrbKziN4iKQDMjSE9hC7YPdodAoBLMMMUNA8tdD7Otj+FramYCctsWXW0MsBd2CRWv4
Xqw06Q+q0ze/cYWA6WvqGbN1S5ui/zXgJLJSefwCvSIQh/At9MZSewny13qMlqIqDxd2cDo/J2yb
Xc2Djs5j/Ts57N3iCatRCRmSXWi2F5Ss/FlmfKCoZ+OBX4BwNVBcUQQr5vxpdz2ByTLfCkt+YDJ5
y9mGbZxCjU7AK7Lfg4aEs/DKGa0lb5ESsj+5gkfJz46t02+TRO4L+lW5W3t/9mczgeroBasAwUUB
Lg2j6YbfDoC/cAoFLWKEs29Ycg1S6lJbE0qOgFYnrzF2xEFk0Hudtt8TFnCoQjh1x0StFC1wuhWk
PdpHTz+hq5vV35VLS3pxSEVy3apEzDo7UA7ZLnZybBTbPJit4DWyAk8t0a6izrBOgmFRreiCkse8
Ur7CNevfGGwJe8XdeRQ6he0bY3+0V6aD+JHAsm6nnSvD5SGGVxZ74QxHhwrjcVSRuTAcSVAEXndB
SXhwJBpFhNVvEIYtt92pE7RQfqy3GX2rARg2tnN0d+Lpno5Ie0KcPR/x5CbioiItBv5zybVqprpo
T5e4zpXHGMYzwyCGPVvkoIXx5mhRZehKdu2uvr3D/X9Bf/zzbkXMREU1NxljbKgtmIPgJ8Xk6DUM
r3K6LZmRTaOfwpvFFCrhyoiPK8W6TnV4y3BuQNf+1TGLY6SYNN3oJZjXU/OL9ORrEb/IN1K5AvMY
wj0gQgQ8IsHNmsyhbePAfs2agan/GfNgU+JP3uyC7nvuTJ7UvjPdWhIZhQK3SqP6yYXXtQaBjns4
GNHXUd3Rmbv2CijOG2QNQyispS3O2SIRlvEuL8MLlxNI0Ds1D9vW8A96BSvz7n+AjpVriyXwoQIq
62CU5Q8m5LbmRZBWGZX6eESxgNetCGHjoXN6yUiRVXaEdGEVbQoWqqSYf3EftLEox21bWY/oz3Gj
4P7VmVvad95U+/EBYla8ni2FOnsgpp3n47p0j6ahS+qsrouidf0n8bF58l7UCy7gg7sfbUoMc9gS
sRy5l7vB1g2jdmWJcc0L0ExKx1SopfB8Duh5gG0pUUTj4vUH0HWI+8shtai6hpxIefvF3AuFTN5Z
6ASCynWSpz19zNDbpfdfXAY/4Lhlc8ii3OaRKeKS8XjpLHbN3tJEQ+Mma2Lwjp2+JIeBOgdXlp3s
vScrpwOi1TLL9eP3wkVC7orvoUcY9STUVnTl2RIzsdBrSzb2twl1E9G4F8S/d+MmlG+nqYo+FxSF
Q4sFe7wy4KVU5KSEPTxhj1hCODIPDCq6mwucGFbIhTvZpG3hXVa03xXRZ4nc3dZizhaF4g5LO8pz
X192iSbmc7UB3per9hNz33vkDavBfGiwstItyBxcgshBxgUgeG61v5MrUOjeiyDRy+LNKY8DBr/+
XJUN+qNxpcXSXdT4AOW/OJFZ9ZWWXM+4nroW8jAKPbhzDBc/Hr7kB34V8zODnmekDoO5i1Svz5Mv
PQbo5ccpZEj1e7AXAOCA4nSet8+A9bU2C/QxE9pAM2f9Ad8vQH7p8Ma6HCrlKM4skgMdVlOPsuDf
Hzgz0O4wZqMVE0aO6D1kD7qGXWRv9Cx1y6WTBFEoUawPtqs28wCMEUuEWpdg//oJkmy3zr9kR1Gp
CsLk7goKrC6cJlmph+M34CIpqdQALIDDXR96OJAHExhve10dqFdiCKbPIWggBW/jXKcNX4hOuOd9
TS60/qTBmc/RPLUbQ/rWREoW4z88heTQvVHAKmv4G6Aop5JGukWYhDznFupNKUJR51M6TKcz2YwS
4T1Gilq7k2kYn0TIUYemYMu6uew/Vu8k07dnQg3P8+ZNUnxRSGGgAXlqEHG5IVKzVM7Wrl9ymnBp
Lyfg0+SDu97kV9nC1FVF8iIKllmkgU1vgEsk/zv6iBC0vpkY7kwVenJleqByWogHqB2Yj7HkVdGv
lH3/lYjACedkLDU3RdExTHaQxraK3g4976D/ViNypaMbuDHkVaH3TiUGPVo9lSB9PNLl8MGqjTpd
H1mUV9M4ql86lV0L1Ou9FuA9fzIdQuwImMsTH1DVjBq7xQ6JRfMX5NIt78OBnBaG+eJqfNaYdlQx
QSpBvX9z42siggrkgxrrHj+oy6NiKB7VW3Xkyx0v6b5E+1K1rqJylEz96lc+QdLMSAVl2d+mt82r
MZ9UHZc0sPpDqYvg+R71G54TlYZhEli5Lj6wqv2Wg3BzAtG9SZpslVtb+iTCw+/tk7V4pm2bdQJw
EfGvma1zaLOr0qVq7CTNQVv7bLASVzhDsjz3YBl0HGaqdD2UvNFMN5qehJBcYFHFUoWW/vOu/eDR
VkdRkfZPKBT/+wpHij9GW58w0xq5i1QijktNm6NHOneNDAX1aLYDNRhxDL7DPYucFqkoKBR+g4a4
pwb5ffbll9VleW0LYq4xRD9U+rxPOl29OSP6AJW7OFn+S3z45iLzneC2OK3EbxX9FavqQWsecBuG
L/kHGM4SsEWEYBQnnN122aR7XwfK4282yyW5j2GQoHZ3YN41OcwJXlR83lvbHl64sw9S7RSzPqDk
tP8i2e3Y98kE1rSauWs8dBJfP5P3+cfJI4VmgiAw1Dj/9jnBWf5ZFZ4dR+N8AWD/l3p7Op7mtP81
RLt05ajuOH+pKvPoGYWyYaP0MiSr3MiDrnezBNx+ZNBSEo8g3N5dyTJLZSC5EPNZjXBiuxH/hpTD
hDjn3TV5xjtwJEsR6J274GP7lIRgtOVHQjCPXO2DieBlWW8hPWZWbAkAChP7d4X8RmMuu3+r3mVn
q2wV48UDiBnoxF3IKcCXnFvnKyuVd+XRpVUrxmcDznP5WvNKXZ8dmSOx3HLUI+P7Vn6AEue3cI3v
UmNm9n7Y+2GwM3XI4ktUa/g0WoCg3i5hColdBIbu62+ki3qv/ckUiQ3Ga6NTX5sbjcn1MxXVB5ie
DlkT9W3dI6cv1KkxhkKmM/TkpbMcVVYxkGWgCPbpfV88McQGDWAMc7E/+60Z2Xy70V4C0rstTlBN
MTucqI4xoeVUEtlFIlYqqawkl7VXsCTXWFFPJ4Ja+dpVZTP6eEd3YdPLfS05HMe6JxQglgZl0XNh
BBuGnbWsWG5oV2OHbYczaz60zfR+cFFzutZwzhWRI/WHBBZOrYfjly8oStMIxTdI4w7dsXQsLjX/
cSehlRfT2soggR/ewxPdLI+Web2jLgA/0TAOsxG6gOj8d8QFR/QvastftKr1OMp343wNdMJSg5n6
HRgHm/pqCJ0IHsO/mZ+8JRsDPuYGXc2ZeXdzOcUa/9fJydA1SmS1QZTSdiRoqdVLkZF9F86Yt/fX
Ny8YqxYt4Wj4WdrrmqZt50hnQzOh1vTnwEN0jxMzwY6QUWVEngqBmxv0FD5i5+8ItBh3LNUbosJO
pONQ+BJ5DP5YupiLGezO7Ys37MPDiIFIttj/B/zEK8N5yGFqxx3YYS8PRDinc3R2K7ESRk+rDqc7
Ehvf5OmoZBLGLuPOptWsuRKMYkrfKvqehl8Swp3l1gWjy7krteDenlTgdq6DbMKUD1ciakkuWu/7
FK/Wx/UFAYggKlxEIsIETX/vrXVDkuII0jeRCj4xKUOYMCXFpQbkMLIbd8vOGhMwnY60m/kpjC8M
CFpzNMwxIqX9KXXEqX0083+KeD97OaWM2MpHtx3EobGs6DZu/E8eIemieWCFL8T/dK93v6tBjXZO
V/+EVD2rqODKLP3dBkkm559ZSsLwxsUR6Glvr895VCUxKuZWPQ1pDz4BC4ul+oWaxFgPLcefwPDy
c+z8N6obpMpiH2jGKIKyQTGsNkcF2oGl/24X4opxRzhMsxX7AdRrxfQq0AJxjdbdsKOZjBZ0YxKA
yca2rkB2//347iCeqQl1Ddev/mUEvX8mMy3AKeRb7n7RWbefgOT/Jo+ehzfM9fUfv5E5zKcEkKwi
yPNCjCC2k73sL6kop4P2AeDPcks23x/qbtsZslbQ6WQwn3o15qmtkQfiimi/j4D8FLO6H212WRNu
GayVmk08dEcFO1WErMkY7pOuS3M8EocW+nyijXUIGK+4wI0Ae9KTxul4LpacsnBWLc7VX5cKf99C
uhu9IQVX288mooeieeWuoaNkNvc1rCdq0lkmOXaJvPMTzDO9Lh1bTewVYfzSb3EZm0l41KSBxWNF
KtqAWwf/vx04Sm3Agw7AB5BHat2TkK0QpkS5h2yAXm4Sxl7fKcwYRjK1BVqqabrDDnP6if6CKX/P
s7GiZ+6Z2QTjXVCCjzUYOc6Rxz4zlq7VLx7qCgZpA9uXLVQmNuCOug8PMqpXqtv0FL/ezptihn6j
mp/c8PRTaCBCHVyF/AXLx2agx+IU1q0g780Trhtki2VHKITyy3B5Crnu5gAp88nZi2zrcV3pP1uj
iv25VIAVlfN9b4yQsD4ZvRpFfHahuraXZydjiQxUkRDKXnBuYxvwWBrTewTDGxD8O/xjFiQS41Z+
XaxZ1J2i3nlujRrODHteOfa/6qtZIEY8FJypH7J6IuVnFzrrEVMuZ4h79d7Q0JOaEVwvKu0MZ9FW
OLh2vMVc0yyS40JvilS6lUEEpXperOLfKNYYePtfF2otE5RTX8tHOlU9vEt7kvyATZxLIkPYTPC8
JosILbVbCWO1Xn+VwdMYnLFm4giPS1NcwgdSf0+noJZ8hNhSe9i7JtEXUh8IJCibSYKrtjRdZq1P
4u/VecPQkuAdOcJ4AVoa+D8k/GkZYmTbP10OfkneuWaq65k8HpOHDFhYxfp+tVTot4e8yV6LdErx
i/m9iBVRSVCKmsCn1V9UNhUCQ7g4eMgFP0pJ+Km0QC9M54+BMTJEgmjJeRPG32cy/wPYlfHpIxNH
JcY6yndO4ewbU4eZS6cp5AIzlBeaBBHomIyCZy96bTuWIuEOQkKVNVURV9TVNsfWVIQLeQD9suSm
Ev9Jth4eIOtr/AZ3aK07eUetzTQWN+ZtNRmVk/GtE34ImQ8TyBCt5pssrI3bHevLtyBWZhWjd0uu
VJPckKfkzLVYHYxpWO2j6EPkDkQDwXXdEUI43Kb37DWmlWGnxGzK0Si3nqrx0isb/W5iY8n6HXRO
Ung9IOXO5rC5nFaHLZSs+7CWWGG/GUSn2ikBnqpiWhNuux7QA+1gRBLQ0xdijZpvAEcqi5yNluqE
Agwd5qzYM3UcwDsJu7sn6WzRJMuInawqj7yHfkiDZT0BsbxUMDgeyqJcb7ckJmoxbG44rLBq70NZ
P0G4DHEb2wXIyjPxK2KKIaTrnRlkDA4XflkDd2yjZB5LmVFYr5+dTOBQibvjFUExHEEvjE11SPIy
Lxmo/n14e4Dqq2CCAfW22l8bWc+2RHxkm6u4zKNr5q9ptANJFhr5VNgRTRx80O/uPsxMEuQyoGH3
Pk+aVtxTpG4d6qZZxf62Leyczqkuyq1svpLSROTF7HAFqli8w5KKoqoT9RfKDTbfO4gwVwj0yRWE
7x4TyKwma/ysRFRZmvg0CCf70r9tFoSlnKTKgayy2p7vUCER4KOsEYwZhOoEkN+FgPP6uNzRtFkV
1jiGdr0ACe4lvo19TFGu8NEoqWA4BcDhzrcU7XjOSJd7hU0OfMlJPl7GBQ4c/glCfyG6zCwfdo8B
85b74vRf4CwkMd6SaTI1DI6U94E/ajN8en7KfN1Vj+gzAMYBCygGwii1nBjnukMw/fYY/AQj87kD
ajPWjlHULAu3iSA5HouIiHMP44nP7A4FtGRGqZX8vXzPi3JdLYK4hj2tk29XEzV4NGXYn5+JKBRD
4VxnLBpT97cX5xLg4VnRzPSspyEzKyO7Wg+kwBSRekaqjOvaStdi10v7HKGErwZHMpEXfPRN5plU
S7JuEnTY5lCnF+mRnmJc0RWO6+KdZvnTyW3bQNd6s6mUTJdDXjfxaioCOLF+6Am7BwsqXrc+4cR6
AlXwJpTf1ZDnN0EMMaVaE5fqV/IWFb0oIAQLDUdOnD1Hct+1R0iAV/Cj5nxazrrBVQB8rpUlMu9u
dhEcihX+stEExdnZpR7jC9IXAsfEF6bbO5Sbp6Su1LRXl+IUcYDkz29jLgg1S4v6DBwp0CpaS0+1
80vQg2IuXQ98T7dOIzYdOjB7vFpe9yBbp5EHfI/QVlPmWWoGBO6GltBxDhe3UBpfzfdjTTjgI2le
PFT5psHn/PysdcEGm7UCrAiu/DIFaTFmw/IXBlZGFwCUTrCI1FZeo63vWkMpDGvaAg/+7ckCXaJy
zjUc0uRk6LJiGfjQn4z0UB+uMcbIeTrdZxlCjiJMflu3CWQeVB1/JwBQmT2aC1fotN2s7zN/rI+z
PajlyRH+Jseuk39FUyHVUiIZyBeTLNHxXiw9zm057+urqmMqpSM6i3YjwgxcBiG2jL5rXzhCZ9eK
5LOR7E3TsrXYGzcWyFSyFmmprPJVwz5VFHT+eq0LLB5SHicGwiIEIDKStjoN1T8iIYsL7aqeiTb1
w2i8tllMV/csgZ5jDjM6vkLxb4cjEio4yLXHIyFysu1FqolVHSgxInIszMaERH3tl98w9m9wWma4
dB6zwAaPbgdptFJlTBFZHb/AJbo4O8KxvuzeFrAprV9uBKOgIOuT34eeVskWO4Y0OkWjHPkj8L8e
diIT7H8s/TYfjvKRI3mKVcDW98ViuagqfUIVfCSjcWiUd08Tmrtdo5FeItx78RgxQOo6oEt1v1TN
cmjWOn2wuQtMQjKgDt3bsZIK3V2aVyOZBovOPkX8DNObi5dXumc1y5LMq3315/ZHHAEExPMpJNv5
WMvhbudIiZqbORE/f7EIxaJBnhAQn399/qutbgn8FXAK/73PhIDj1YraLeJLe1BsaWLBzW5sQaGH
JJWBqLFlv7NcgNd9Kz09luEUJByUAMpypPUYHVLjGcA7foZLKYYKjfDfz/vRqSmVkAmDCfwuaZe5
9/1U++06gZwMvg+m1m8euzxVBP6QqMT4S542rEIcYDeiHbMyd/t4bSb5eG2Ezb5Jjytp1Ze0cqot
6pm8VWyASb+T5jPFcwkJnw5pbYfLd4dluXd8nE1ZYDlfDT3Kzosm0FJwhePRUdA3hZ90FY7OxL3K
AXgWXFvyQBd/8Kt4zhIofDOaN4jv2w/1CyLa7h5a/fb6MqOOmAJvomCNRh/VeHit+M2Z2pYgxI3G
CDF6PFRqnKaxLLqIeUzNPML3/tJ7KdOmY6NC9i58yhRZO5J86NXBkIPwIB+m10jSj6JU8Q741Ubm
K3XjUKK/LhnJTjpq+Qu9iDU7uFvulxuy15CcIh5jgqjBwclPY2ia9eeEX4INhtTaK5zdbkaF5m5m
lok/JNzUyCvy6ezwocGOTWk7Ont+uzKhusWzNgZ0BBKfIHYom1uxKScVq/anyJxYvQPzS7L7s1Un
glXg9uJLTHSm7kt5WU+IZ6P98O88QnF/l4tRHYSMuF4Q2Gd1gKuxKihgfO521Da/Ozg6TQ3Zu/mD
m0YW58atRGoW8WZGuYBPit/RMQEPYz1UUnmRFlP6/jek6M4ho1teLmfUj4m18ro4D336UuyeWAn/
VrBUZBlZ64W1lJdD7fnThqOHIv1lYZ0ls0f73hoznEo3O8LajNjhlU6G4vkX5jxoyyOtBJWo4sl8
nbSt0smu9ORdXn0oB1IRB2qomftd1nbdICA2D5H13BJQkCYkYoArBe4iVCPzez3uWWdY8hJOiGrT
nKvaLqFS38O14SujXK+NgDe+PT4qLI7HQaADm4LWghesuaQgwjUL+hPwNPYA6lq4tPOU/lhgBKBi
UuiShVN1ec06Qyd6FMsWMiba7uBdPDblnOFmzVINjAT7SvEWscYwWjDpiBMBBk9bxa2jt+ouktvT
XIDQAW+PvDjFFiuNpkyxImz9fHhE5Dmu52u3rn6qBCoJJWxhVhVYhVIt0zf91JCGPjaiCbWhku/j
vQHMgvQuMj8vxXJBEW/5ac6mXjDf8watipyzMwebZBKg7SK7rB18wQyffm5rwBbUwG1qcUaUDPMc
UvBYryokfjyM1Rc5ZPg2h8VWevj/zAnBzZ0HWX120H9YMm54AZD5CNCLEuhGRpZ8mnLbUlxVXSwB
eHitX3IHYktvX7+NW4n2YjrW77Pmi5DwsMTj4aGPq2K38xk/U2vuf4ZdQTabh1pljS//vb34X9LM
a5drFGNDWuBCmsImIoUcixqjzo//umaOWz/vOV6tdlcq4Md79ikFx0ULuj5iRlfVUEHUSS9kYs13
sUukMTsb114ffeWagqI7GMK/vnNDswIrMpDbkHB2A9hPMXCtByjbXjwnJ0B5mfxHeoEVJT5I7uwN
ZC7XPCme7VkS7kH+rlDWiYVYeeVxmdLbcSkM2iHSMUpnpwDwvjD0DDCQi6QHDTTdhk5URL3W4FcK
UGHbu/ABmeoWzAypr5JAXwHUA956wiDdtjK1EajVsU8pfjtiJ6PDbjPPtGsXStq3RdxKiDiUxfjZ
IH3mxN1Ux+ATDp3zeO2Ef6uhhHj7phF+LBtKsCm4XL0aXcplpWEYTOaewyX+EZ9g4Hj8e806d5u6
kFPiVfNT5gqkIBEwxIGtsnZmYcnh11LIDo5bDK7+tyHxa5GOCJSPX59VtlQRKVwhcJN+lzHHHkk2
NpbX8ssxtzJdk21sgJpQytNwTsMWN6kyNn5bMHQEsoiUeXfi67G/CdjX7/wv5aTvk2gMcL2NX2ZY
BmzcGNwVeQ/Z5295ARpZ1KLqfU9lWA3Z6gw6dgctyWfejX6VsXk5Mo4YOs5bhBif25VyGyTgslww
pOnO8MpN3T1gZuc2ioHhnrUXXfFViqI1oaVMT6B8WFppcG4PPlwxBruQW4E094cRGNNaz2weGNbM
Sag9JfVKXF8mDp5TZHyfkdJXq4r6vmt5Hfgdk108yed/UAEsK5s7t1wQfRR7ZtxapD7n99nCnegR
OguiaAMhoNA9bjfXb9rhZAIPZCsquc71RSfbGXobTYYrgrebqcSOzdtiw4+Zrv1qz6X7VTOluJpa
LVGhspfGHc9VvTDMa8g/CG85RwuJoNtzpKH8MrN1QkCEsEJSiIm9n3dwBHL2jAD+10yV04usorLe
62nMKhKd4LKrkDoeipEoilSszoK+4ZUns7igV/zA+PkipLxUiixrd5EJxMitTz1yvPIqUvTHSsTh
8jHxJkILrHdWAIC9XHSCcYskxzXaib1LviJHmWe307vaRbLTJ1fLXSh1z4/AUYkpNBJi10sQqg92
hsxJYfu/abs9ydECxZUIvpNNXkYlX8b7V096+RFlJoj/d+sAt6j+rUm0JqteU0hlyCfNEivW4WSF
5ImLPR1jMJCvrifkSdDHuZ4O1yfAONi+9e0P3noRWeX7e/7O6vrhPvOY+/a7M1di8pIVeH7cMu64
WP1jIlZoHv3UE8bFQMDSnwU4M0tWWoZQaukVJ/EYb8TFyfJziFg7VxXhpGT4c8bg9I4av7vFXidc
BVLQVgjZwOc2X8/6+3jG3O4bcglVyvADIqHEVs0Bu9Q+d6QvnGYQXbEL+17EgGlzwlkzZdA0mKfC
DHg1o/QoB+HHisXK3LC70PlftVAqPzOzAKHU3OSlKsL8tr5UPxs7rbMhnThTknTHv8NeafXBcuSz
qE/NKk6r+gUi2KbMVBlH9HhG/o1dfkTE5jU5QqDdZhp7VFinrURZkVGC+o0ci25FOxYlfA+F5MtP
lYF8+3D4ALlJfmUJBovFfaHBUq64wPCY7NyDFCs6kYYi1UNvofyXRjA2647OVF0pr+Kp1iPzR6C6
lJuXhuO9Djwfr78c6dA7GGMU8/KDNm3HfqfrYhNgfKovDeYFzAKeYR1b6EkUwKMsK2/QtZU/aBX3
gZNaZ3GXzjiop69toO1rVy8X7/KduvgFKBvja254Q/KhW6b7SrbytC0IUJKm6xhbXKoJczRVUZal
2N9qSBUZ+AdmixftKff1C/8xypljI7TYOvFcCSZMMwSBl5DS9x5twNnaaK819YjJ+bnF9lK4vbgT
90ob0g06I0d6u0sI+bJPo0y7sNI6Idoj7BX3a5Au7bY7+DyFHsPTECj2uG/0giihskbllrwDezPs
3CIAcOBZhEWX68CF0EKf8JTsb8D9Pk4BK5WdZ4g1a5aDHVDynNo+oj1Psw6IJZg4LM/Sg2ELFoHw
mgWXMCUjQJ5jytecs/hGIAhlSdYSybeBD/nWMWAsdWTvgdeejZWEjqN2uxlbbcH6f8JvXxtz23+p
pzQi5NsOp6zhtJi1rVixptPE6Le//5OejJf0NQqBfV3S6W0AFcE1635PCIfQU/mZnexVu9TSCfvI
ogpe/6u4sk/wFGXkgDy+9xK6O7Ru4xlUGZ7QY/OMazGipNX9L/4cDyqzwZjb9MWc0T8dsWktkPzU
w4KkJD9OGAVorO9vsEFFQqD1av9yQYEFC36k9V1FzXHJzlrY6LsU33m+tGOC95AyYvrCXp/R/aD0
JXZmNbdnMj1/RnCxPpfs951VZKnC1dN1ie3yxbX0Lg/+ktqUsO/AaP8+VaUNSH4Tc/+DUJ1GvoZL
rXSEOhvEd5oCweTW9HTijKqf2Krz3hD7TBNAXNQ+oA3BNiHIl+omd7tT5H/MzenPKx+6q9UtvK8t
3GeiNiHLq9D1olFnroM87m5i+Tm5H5HqFNOGagU6vJy2cYB70w7QekrcHO4U0AwHguuMwSyhimLc
8wCT6nBzLKDngRaY56Ao8aKPMmNZTE8Az/QkZesWzzZFwYotYf5xyCUTqH3An5/4KvkEnVwj1EFU
WPUOsdKfjx0Z1vUGLahmcgiphxuXu9a71CCGCmAJ9qtGYPCvZH3uFuycO15wpVey6gbV0bW9WYAP
PCF5k2wMhuKEzQEDohEIniXCb7txoAbgCG6Ro8d9C97rUk3IPFDN7Ef7TKL910kwZq+3UxmHjY4O
gJ1hd6bqvCjRU7eLVxipoh7s5v8HZd++kMjy3x7MsBh0l8kdcCnLyeck978Jgc0o3gKMvwxHYRQ3
bDMEaGNf/6+f0hXSpzOXw5lBQZlCFkjlkP+nNkt64KbxeVFcFVX3w5gOikbbRqpv0UZHx5v2ymBO
rmLkUI90Q8SJA4E0Fua+97btcOPRdix1BM+UGP/OeVzHGqVobPwIgOY2uwy5wJIOBoFG21g8/5NW
GOmWsY10uEM4Cnsj4sFW1hfpcuoelUH7NW5GmkAZ5nBD7vkX4q5g+DivWZJq9ELvCRI6JiPDtlIi
1ez4+2mW7w5q2n9olAW+R/B8T5A+i7AqL3mpTN5/gJinYcpMOgb85ekKEyGogRrxF8HR3AA3IPiz
krSYaOjGAbIdW3xfO8LH0t1Re1pXwbaJEoyInRinBstzjQWg1+RV0stc2Ti2ZCR7FNjRS20oxJRK
um4t9xwu5z12p6PZWzczCcl9QGYlgnBowq8yn3GDv42RIAcYXQvWMq6K8Tw69oJOJ012H5Do8EGd
eGAwTA9l9QNEzMIbwGzevk874JgIyoBpBTePoZaxt26ZITShIDyy438sbNJG6MCEtIAXBO0Ai5iH
kJTWP2c0PoVUEoLNZ1Hk+sYTIkqkT8nOwrmhSrP+r8xLIiz6kFbehLbE+I17e1QHrLEWlqNVZl4Q
35muYH7bITFqPl53Pt/4n0pbuOO+XVyncaKzcdP3VAcD9aAnPmSqImnaKwFSOi+cX68vhGjGeeA+
/l1sEZoj2OS11OLBEA9A6cRJp1KHaYTH6yhYfjEBAycDgBnUqBG/9+nJGWZRp8KQtyas2mwEyTO4
BTFj+uDbYVSa7al1e5PlIi/+b4EaQU7Km+pubFZZ4Yy1hAeZmo0jhRW1GndyY7QVD6Uxma03Jfac
TTXFnh6BZESUIy2wyctuYgdnabnFl8C/jylxgaAEzI1OQ8YsuA23v1FWx/qSCbD2FxfSgC/2DZ9F
ZKkyqcWobNiLN4DfzIGrsXWTbgG+QTP99HZnCJ7srlENy8QTdONb7mM9ZgKiL46oVewKPPes2xeg
CFG3NHI95YqNZbyyiY/OtlXU/tpvJJN5OolDImVLWT6Wn6ex33qYQQdw31P/7len7OjQazFhE0Ci
iZV9RlS4h3VS/Lvdr/0IV39Oasgy3UGnyO9v4QdlkxJiE0v8N/MxFPgZAs9ODanyUB1LwY7eBOmI
sEdEDLM7sci91nEwKpzukowveVAS2LMV2joauLjOsipu3iVboefRdEiFZHKSAJLUV78qoJJtUpIS
9F97xpaWsdQ/G8i++LMKYchQCOyf9nwX0bppVAPrs3mRjV5j19x0vsv45952ZjVHFXH9Mu+15Q+T
p0eKuTpidHhRYYrY7kZDGkuQilMbVLKz/8qSktTWblV2/8woJsIZeXBUoo9bQYL3VD7Y5yzAG/4C
gg0gTSPgKI081huMcfIm371DwLpWLwo5ex2OYLrBE6K8L5BUa4QCYHrom9m1fPQdg0ELlBGTEE+S
iRG/opMdbv02akuz50laeRGJcbGv/7VOORe+hbhHUW6oija/qzuiBk9Bihbu1mp3gdNa2iUBs2/o
TvJu0eoSISR4/nv8J95aCl+Rt3hY7W8K1j4NEOWIt5XOabJ0CNSnGjzVb8vhCHsWW6El/vkw6cfm
XX3rjGlh3MC6y37egLt/G1kh4yNb0ksrHA9bdk3+73fIC/b77rgRJDUJa1UEGRwSNJnkYaBgSGeB
Wy/V/D40tp5p+jO7/IjKRHtvqszOxVJUjK085V9i5gFVN8d4wc+bXnYzdOJcyobnlIMDqho16+56
Q2MVIEDbpVP3O96EvAWtNahV+bdVAT/I1oEZc01lHzot+Ds2eQnu1P4mGOUeflpuiG6iJzKns2wZ
kKiSHpiV9eZL1hg+At3GGKx2ZEdNVR78Ns1gQ99b4wswz96njh4HoqxDSaZr89L/o7sL0xrmYOLp
K+B+29c9lJbOKRxII7Gql49Z1ZPnpeYzzHku6uU1IIIJAZsdGMbqonTrfkHzsi11/ErlrhZsXZHr
V1xzxVHnisEic8kwSNnK/NcAOUBoj0WMe/JyBV73a8LAJe9s70+XM5QntLy/3wS/ONOxOI6XDZ5M
X747XzttIMkrpEjlI/IJEip9cYMpwF4l82lvKlgShoOaziytuxoohTR8BYX45+mxjOtTAZ02Rfo2
INhHacRsnBPaNxZMEshtaga/s26orcd+Tw4HvxhS4Q/4DxkSsU2HZzg2GJcttYrPIIUid959TDLo
C7uY5HdH44ZzyoUTK1Rn/4R+oOt3LZ1xsG/rgLR4fVIVZGU0AX7ORT4XepQDifg0im88rTEPLMDA
BtLIiumZjqZ4dnJX7m7vN0Baw4ViCFObKxn2GOcoRErc4720r2ti3JJAB3I7LnIUcsmP0BgQpJwF
LYPhYdML1m/yFfilQLwyXdBrE0uuEGZppzoQK4ljkiKWBWa6DQV+L4Zz40dsB0yi0m0MzpcDV+GI
GAyuDawFWlNvx7+rPdmXgBE+wwNUtdylXQ7HaaVrOIEps3jCcrrsf0F9JGl4inoeToD+U7CPFWKC
EUnbgzbE2WhzSoKAoq6iN67A9JmoUI9XFEzhllK+fW3R7bqWMyfp3oY3NP7LF3p7l7ir2XESmkf9
uX7KdfEU3qL59VjlcuG21dy9MOyzrGdpHpv+g/BKt02yEseExdm9t3FYbS5XjdMDKXQ8Ukb8SoCj
U+mGQsfrYIS/zJ4r5VvOqQhdZH7Gmhe7hyyZBxY126JYwPb6AUX1x42AVVOP+ZxLk/7MTOIaa8ec
ovnDqjMV0JqLvxY6r3148rUQEMUCGo+AOtP9yFd5cXxopQi9sachKT5YrqpJ9qm2D/aub5Lhv/x+
xmkP9H6g2vNDvYkAa0oJGNAtJ7O6EDBqkXo32sSac8a9BXrFD3AbIoTHIWmUkv/xmtoMtsmQ7v0Q
eujKY9knU5vT6RYl0el7MjGDM767gVZ4g4b69IgkRKci1Y35h2b1kAjbEmrqQLSK9kNwJPyPlZmo
gASL7SzDUMcYzAFuEpGBHF+KuW0qk1E6G+j/YyScyy0br1TAOM0g/LsMmIgclYLOS94VOgS4lPPD
HNx/4VEUeLfQPL5f8OPRCgTs/H8wAqYrWyptUtovdz+wQ8AyBpoxh4RXaW238LzyF5i80m+Hg5bF
OXzjF1takQ9ztki5TQu4PsQVizIuWQKqqkrhEjJN6Y5dEzImi7GT9QKQq8SH7S+zVTHTb4GtwmTG
TVjNoqb9SwfZbHrJO6pAf1F1RuACz85TLmzFNkHcD1Z84A12/uONDsafBm6QiHzerQW+aTpC1Mmq
taEHUk0Qt8O+wjF/KhMcuGYlX18DOY1lyv1523CyV5cdA21kscpajGE+J9CpnX2WBellmdVaAfMu
JSWPfhfOSkBv35ndMa3oFWsVky59eJ54sJbM8nF6XpXguIwF2/8ApnZxMfq3J3R1O/juFAIbPvxw
v6hRU2JWos403+p5QPl49vBTY1vfYACPeqAoVhV/QqQFFamWtbnT4m+A7UADZeZt1SNhPwnTzMo4
Bzg/20yQC54BY6G0dwSzXYzMY3YqdZYeiN3QBFUmRg17BdUItfou3oBldgp16TJHOVENbihSm33B
dS0OOvMc2I0qxjm3FF0g4MDabif9dcGccIcR2PcwruLaWaz8LWKNHIa/g9eNlvcOTxYWQ3+IeNTf
YBFOQWK7HA0BKNXs+EGhOTatsAROKu8YYwLdEZthXqPVF5rS6B0jaFXffCnown6PFo2JqWv3Jq+7
43lsluwBELEYYFHp72JzhbMOk2vdAb4qAuAmaXrz0P5l70+idhsPsaiyESFnNAZl0USijLIGR8yC
ZiqX3Tqm+PSGu4zgYQFaigMW0TaA9mEBAeY0vQiRzojyHy0IkJ46hjTeJnByCjWENcNYRxsT0haM
xSh4gpRdg+NXefJY5G/+Lzpb80iRL3L57XLFmtBzIeyZKHcLZYwQ4FNAADMcEl50rZESmbuYEt/7
j97L2wEF9KN8ae83u4jv+sxnOCvueSOSv2B9oLpJhV31ai6rcATLrWnzXJbL6aoViYTDUyxtu0tQ
41lqDtfHMvpMh7RwlhG19zdunzgXaWFgnzRloMZTQbYcNCDNxtg4eXFb230iUhLPEBoiHe0+a1MC
bkoS4+TfxHkrv+phNYMOb7gwRiGEIb+i3UOYYJE/jWR7XQKJbHlCg7HQkPAqRK2SNIu64JWx0aCB
YrNrPtXZKSpve2CMA+BYbnFZeFnxye3lH0Gv6KCjZzgB++5Q9vsGIr2MhLoxirOuvslJoYZhXY3A
d9k9L3veUyq1N9ockHcVwKodTYo6WeZnbRo9C2UiNx3BlbZ7JPpBZk7HU2WIuIeJFMlRygXRDLSA
qvvPj7MQrt+SvKq3Zus6YQGsQJKAN0EtahqRhaOjVqZrdXvap0kN5n8GmrZy9SpKt5gbw/hwReof
sJ77MrfOn9eDostba8ADBPpwcsA60jsljITxqYDMHGhTKEDDGCXlhf8GMf/rpo4hfbIGvS0OCjvw
cOwPpIhySQx29wrWMiKzIkWYIThb9fXZhgi7dF7/QlLafpgb9PSZc6DuJH2ZY+iWnekgmiTQd/Xl
DTNJTLEsm60n3WmXgBCOQ5/m6iaA41YHoTCI3rO/0bilHqYMemVH9mrwnShDlaQ2Fw8l0fhpvdZT
pkL/PRbasNY42m8iJcH5umLpx6P7X3jMyPGKCKQ6dUhOGMKG49wCm2+3m4L64wqTznbA/JUZsIqG
n9Rxn/caBoay00y2c8xyzJmMEYTECkQCa0wZjwOGO+sEGu7mt5LT1+pO+tx7BQmfn41Dhde1Wi8F
F0bmXpjs9mJOnzAe5XN9R85FhCpKmXizCNpS/HjZ/OQh5OL6d/4zUEjel/BBvXzrq+9LhWznPs8q
GcDnAC2IeeR07WxM0OOTRw0XbVZcRU5Bdo8xjuj0iQmXYCehD58YhbSrZT4G4Z3rWuPoyl9unpgC
wKaHNmXaBatYQ7HZgKH17DlJEGmVR8+jlvb+/xszWsm630Q7GMbkk+lFTcrSswRV2ebpGfzC44La
rsPwl7FimjRxKZBII3SVrPcEjOlAjr5EH2uEg2R5uF48KyZYI5vFFASh2wxk8SLyV/EdDey0yLgS
Kx+e6MEwmfr9/2r0mmxqXz29XeVs2RvhIcz8p/W0FNtQ+4inS+Hjgw66z62PpgUhuqnsip9gxsxW
HzCU3S6yTVcLV2FV0YAnP63+Ww9t+Z5u4hkPteDK8k0w1y8if3iIBa2iyK8XBwUTjwMV1lyeaVdL
3IJPiiFGAZqF400nmIZn0tXswGYbTBH0pjDd6haaqlC4BCWD+hxd3ui9gZpTdh02XzDv9KItXzj+
vpozDIFgrKzqq1CQeFjI+rxsvYmSHG2bBaIrvo8JmpXvxs+2BKY4ityN6YSPMwHOVBNBLSEDFvGZ
IfZRCIutJQTZnwx8BP39WD3eU+efGgc1xuDdY17G2CuOT9rdmR4MMvyLlbnIwF1GccmUuKRfUiKd
sbXeJCDBK/1IdkjJObIhKaHneDBV6EhZhLc9sFQU0pB6Tn+wUt6hn+9iGEP41nj93Wjtfqnu5oXW
q4pzlyZ8FH9xOnEgRa5JL3aRd3EUcMyBb4RQ7hfReZPVKfE5CFqJRlEa/61OvjnfQR3tBf+X9eay
hDzAF8XBm1gicENUq6KCgpx/Yompy3/R9HZ3nP2gD8Xk3InbJmgJOdvn+qS+g+DVAiAxMpvplUWz
JrGCQzU+EUj0F1c+oQZ+iDQQQ6C5FAuKVV8ZMfuXiHvCrRE2J8q2kV1GhjCjVDuphlWQFHfWz7f+
u0YhJ2KojCIlwTrDOoggZuYA9DmXzlcDwi24WQCEM+oCrkRq1tPfNtZq0MGPk4kTjNwxj2TFa7VV
SzgoXTdVbeOgekgFvAAtP+EfJR1ykGxB2tPPkKWLjOG+Ss5G6XUjGY9GRs8eY7iu3cYaZm9OgWAq
2CL5yzg591Q8aqZeSPxF6UYzsNNNOQ6a5KW5OqFC35X6mxWk/mv26oqFxiYNzcpJemVeDXsFhNkc
oGjd8eaxkDNN6L8Hf+Anf2985aJnnTUyoTkFHrzR6OL+TTejsvEJ4pMbm29Zo3xjZDoIpkghe9xs
khC6y1oex+Ov9RlVqVjseOkierXsFKashz1Qy7xYoKbiLAgkF5+Bbb85BAlf+QOjCLM76lzLOZ0N
4QrQ9G8ZoiXX4et7daxkn14GKbhzg8AAdFa5rclT76CsL4HZORTN+G50VSqmg81rBvIoSkoJzI4q
fTtonV6v7LNKj3arbQiNEgtGWjcgLter1jeElRej+WKCtiRnsAfHVaqtsH29u2Wy9mSGD4+Ed7WL
wxnp+cE1AVwrJArmimOipQEMf8Nrv1hQwzgh8wkuTeuFIIwybfErDkk20eABm3ltVQRH2c/ZEu3j
BtFiHxtnplan2nLTApNTbdheh7ECy0kG6w/NofisNcEd7XMG65Yu6JSz5jkJCp5DgaInsmlm135N
5Dw2Vhh0rGORy8PKkk54bjJFcJtQeSjUPZyeYqvaWsn2DuibyZHmbLyTv4QxzBpGBTsf5wIuWYKV
bAqeVa01TXtdlnErtbogF2EFaMWSGnviy+xoVqlZ+pc7A0f5BP7JpPd8YOSmvIgbaDBJ3vGHSF1w
n67ZCu2uI9F7Sxi27y1J1uCgYOJN6T3k3AldVwsdpa6Wc6SLkByDv/9dpbUGQQkyo0cLtG+6xpEL
7KGyG7MinbowSkEJV7WTGVhL1TXnHBagXD48z7aGizNKM9JPINyjHOeFywqjEwr+vap3tm9DRcYW
MD+JqeQt22Uf3j0/Rb7jnTrhuLL21pd/SZKq+y0g5g01jE4CgqTRdoMjDVuM/hnnVMVULF1I71Ld
8QRO8lAZdd4zve6kL4Bm3whrFsxS7sdCM7P/p3jeVmtITeMZLiz9EwQi+sUUEnN0o2jZw+00XGq4
VppNWZ1K3qUmnoTZaABKBBwdafsPZyIDhdgriNe1pItRAuzPzpFQLOnriomF0oacoO4XCKyceDlr
0y8T47DW+7xXjadUiQqM9h56fFV1Dw5Sumdvs3NBUDIvCf8UcyvABnU8FO4LUaic2y6lGGDO9zju
05RXVpw1EARJhWXes9qJgnd805VLQTt/tqpdgDA6mmovtYotwUk0qmZSliXSbevyTz2HKEkfEpUI
zb4BEvJXQrKasuC/lBfjIAspdOYqS0G0YWDz7OH8Scy6T/DMy8DZX/VrMjCiio2qyBVCoVJxgGOF
KcsQekA4zU3xCYH6vK99y5GJRdPRwX+L7qNcDgFtMdq0GN1UCEJYp8NjgwCaCRHMqJuu8aDGIeXN
T21Lf40ItBHs1LqxSuLC8n6im8HfZeCuW/4aa+Wv/qFUTj6ataTw6PL2T6J4EYsCV9BmdyNT83un
N4bjPCucJnDZLaG813btDuLVfpnsxlA0txTq6v5FWoOmpISQtBnIdsWiuF10ym9nFP0KbwcwMf9k
5ob0myGAW9BFlu6mVZvGHL46aHtmazbjlCAoAroFim2qeE9XsrCAjYoWCpRW3UkeFW9h831vn95S
a9+mUm1wm8omdwTD5NXkoP7SI094g9015UIRp1Kb071Up5QuNhgpRjwMB86Mrnze2VKn+cwxNwso
1YSP2hb7wALh2DXwpMEK+1mGZrdXt2mYUforbFvafRWOfp+XcTrbPvkGYVP4+FJIdNznWysqyhYp
EoMlp5/H3Vx/PDCaidbY9uK5frQSxKpVd7mKyCxDMlhuOd3MrUAdGJMOuBjSFc+SOa6uiXAGLux/
Qe+NwmevmrA2d/U/6UITe06W6jGSH5/IYc/CGPc+8iYaTUG3FWzs23F9DpC6LrCO0rpLYYcUflJP
W9wUDnO0oboT/L3Gmlr6dliygfyXV/0Ry+CLmGuhvfv/BwF/xkFs/2dZ0OVIjBj1/HcIeCuJ05w+
YWrG0jvc32ZTK4PQN2oo/8NGgZtWadxnONQMZj4yXtvU4dgXhFccIl1u6k5R0YQarZ5g0dVpc/yk
eBBH5P13U7niXIkGfat4oRANFmElFDhhYU/jSCumUyZ46Bv0J5kKYJHBD0avj38jwC7kqeD6kNcD
Qql4HBVlyFmJrTexucarpwhGSE4v3yIVxq9X5pCmyht8ezb2xfEZyC/p5hBSVzvwk6BBsaRExaVy
/dABTLerT447H4VzE5Aqr3Qh4w+L2LjfwvfC1no0LvSCgcC+O1boyONWxA4nu6Fwb9FAkkdph8B5
uma/y9t/y0+WplC6JC44K2oq3PuJOyHjb/DwM7uDdjZYvAVmbVHz6CO2YTyK7cBP1SY5Nt3Xgf5d
gALlyaHDyVjVakQOEsSuwRsAc450MxUYw6TZ/mKZ4AZN1MKB+puM27hnHTTblh6gCeqPfNi18916
YdjgeFbw7tHTQsDvZubxcrbhFwIbcIyTgNgNKyd/LJCFZV6lJLcQuuiqDzBtw4PHxbhfyg2lHbcO
UdqLCU3Gm4H2zM5ym/NrKT0nvaP0WmEaGLTf5tF1ggH+qva8Vte5wiqInWR7PzV9MATVRtwPmRNH
kgI1bmm4QnXa58XL0KzdNoN0Kh4WWd02CkG1cv+0QkOV1lJcR/N+SyP59tLZ8silZspaiSC9CPoi
HTet/hneGgP0kqI2fgGo/wxcHwYFQ/2qyM7rhyUzPIURjeVeclwfNBZuTGlPuZX+/aU+m1fqYjSm
LN3E9j+dFAqNsva1VLaeP1JMHUKaiOylKiA7TgwTCrSlHGKjEplPoYry6Cy+fETrUt2N58wKgc9h
mv8Q7VE6oGUQauVdMu8odhOceILRJhLHmGv1AZrFE6QYjSf6usKQKhPNqQ2b7fEF+7Jare9srq3e
SSidFVlpXEMCWIY4ac1A7I/M+H73ojssx21PNhhXaEnJVpbsYtrR6Cmpwb+HJrfdReuco80MYkNX
NRAgTYOzWb9GBt4+9/zuijTMOzN5+RmYdAjRzNorEovDo+waVxGJD0pD2pmHiXI193Im5qpESp7H
NnPfiP1Ke/2ckpck732yMoYZTy1unwACdZH7m/dK0W1MeV9YkT4zAyszRj697wgps1S+xaP+wM1N
jFXIOZs16yzGggFdRTWIjJZXifSdCZ9osoWrzt9WLpczevcrYp5QN6k21KSZzrMtVVFwA42EniGs
kqb9MOO9gXbtwX8TBc5jwebiknZcoAq6G2L5hPEoDOhXk8MeEeIgCsV6mmFgAf0CZLr2EZUd1v0S
sBQhkRmMUyy0HASf1HcAF4sZgK3JDmT08Y3RAza70LMCQkPIk5wuu/a3Sj7QwOcAt/D9RFTMQAij
E38YOV2+uzLsYnDBMJITb7wDnpQHNAdb6+l20zIfSsYGkH8k6vhJV2YNGbI16dMT96tMPpO7xcNt
GrXb/Re8J1YwDss3McPUb4LOCskHGDE5gzGUFC2s7f3QJZMSO8tzq0YjJT7ceaKSJfUkAB0O8W2A
sdb017Nfx/FkrXeZQBQwoM1Zj/CTgOTVphoHZf96TkstfxPCNxPaN9BvdigbR+ePjAgDSbSwvzSH
sRKQa+6P0j8qhPAiVqINOuOTUhsWruhHh7vI+Zujiy1QQ1r3Xk8ogrMaOpXO9cacQeRDqs5O3vPj
ZgxLK/IooRfTOOXFgCqxc4KQKXkgqqbBS8eTM4QQKln7KZZzRgOqg26/3fbYCTR4n/U74nxqnA6v
AKMP8GVd/WzC4b+BG4Y/8wI2YBlWLfGMYrLwLQsawD4uYQ5EzN8yWxCtZG6Sx+vknp0BVnsrXDdt
p6smdZQJxNqGuaBmHjhEoLfBm27R6W3nGbtDUbANvEp55NOwh2RYKvLg5Kuz6cl/Mx/1dPTv7IAH
8vT865+DJsvpGBCLt9yR4dNuIKwj8HdrasTSArBj1y1bNv9ksMdMuSMtePeg8ihqpMYb0JTFFBVB
mYm4gR7/YFucNEu+OzcLS1tAodvzsMPxQOL7XhclbZEMujCxIKIs5JsoloTN+qx5XwsKMwwugVjN
5uLpd4DdssXGXdCSHeUbshej3Gxfv95/5qKBx9B8IYAgkIYwf5BqzcnVzWtGddvMYCTIPE8/9TI7
XSjevNsZLrinFqv6q8BITvrd/Ys89JaZGKY00U1YZQl8LGT8sU7Qy3Z8TnxRJPULoDoFmt33w5Dc
VfthBKhlEL86EzKrBclR8dXPXod3K5y/u3HWhryAlVuc0rFv6NgX5CbvRBRCjMDPMaaf39XgbrcL
d/QWwemvclWAjvp6CGRhxjy/5gkp0EFDDu/Xq1hGhq+msICnCtShq2a1P1iNAIMB/TqMRyQ/EIVX
uAgmV9T2yFMTx2sCKmtca0Q5X/btT/6r5tsHa/qtidayzOVCzNCdLPYc7Rj26X/1ZMx+6ZRIvjVe
FhpeFVfhCZZLKnxK+tG5rSg8kUCRb3EQ6OQmT1QMd9+gY7Ys89Q5VpadsVx2qGt/k0zhZuPFz1FV
Rg7efOCpzckgq9IBTMZ1JsphcFZmrGvKTc9Z4NK+V/GifMBU1Oy7BCMjWBRXuEn48UOHV1a4hk/e
0saS/UCXZCmjTuA46hHtIqrldUMjdjsTc/luL5Klf2ju1DC05EmJ10Fe5lWdUKHyrjA8Fuboy+Zc
Yo1504nj3Fb25SfP7PxfBJI9vN9NGIXn8inP8Okxnl6LjC8dAd8qS9uL4wJnUZ1Z/w89FOMFEYk8
CXP7kQZA1SHYX5t3zTocD13bEGRO3Vw3LEJ4pN4T+NGZsunUHLqqp5alaIqYtfliL1UPyamCLW1+
tQ2xCjZXahMIyPD9jNQSb1BVikASoU/C0kR5klpDC4gT9c0wNn61JOaKxJXRwbXIGt+p5gXUeq0v
dDCCjSDK7WQ/NfZ4hXeQEntLvAL4pSrSBMC7htUENfW3vOFPvRy9T92h0ciDeDXIH8lAZnI+ym5S
E9PfV3buGws2NxNiACUV4tlSpfwUnf+BbbFAA0fW7DXEn2BMKd1KFPk8BIsQSVW+KqUpzby0bqLp
PY5QSDTLlpUZMjrPBJimag5wyJKrpFCPbUzVokFwt3dTkEthsnOBXNeYLtGEzRvk+fU4cjxb12qj
bVAwAkSANvUMZ5ewR1RFiTPY1sdzjf8SwTQ1tegTIh2t3wmIqr0RHiVbVat44JufgTyX4FGOC+NK
5/bVAWUeJRiTCXvGX0czLGfPNtaa3yCZJJKNNtM9AH1GyYa8on0r3wKg4XQsOuLYMJBiE7MjnRJ2
UROGWSFqEwFI7yjWiAlHdTGn4peHvPdyYLRJzme2A/oXrZefQijyW5xvKkJaum1Jf6Ue08h3tIBI
09wxuT8DmeIXcDZfWS8zIznZQYoPKtK0c5uuVCzTisd64kHE7W7zk7hjKVYVdDSBar2oHlmvUzLQ
b8lt6aQLaVRIQHVZm80CzdC+AboKusqC6cWkjBHQyvwTvZ3NLtLVQLKAAYAYpqoN27tzc+n4C6Kx
7DU0GDI3N3B6U3h5BsuyldHru13WQKe57rHObpykfoOcm3imhy6xK4fYu7rZZhrL6CpH85iEXENL
4DccoDlI6DPdbPwAiuVucWg7N8ecmPz3/r4lbRQhEwCJjYLm1jwRKkc+uFdZa3u/+BHgYGXAT7h1
RkE9JPVSDRE0kTVKwq6i7bhFmbCvAwb6AdWUWAViAPJqkSdqV7Fj1zW76tQ6vOglDRbIRaF/oSYs
EaiTmvJacX3E9RZZrhrrsQslGq/9L4b1BKmkqgRA2g2l6eTcJ6c5a4S2L28V4e7m+a9E74lsqXzD
UufrfgaPxLWFvKXS2I60ChfzDNfLhOsQp5RxdMgSk/lXwX5m/P/lj0knb6U7q488hnf9gvzzvtsp
ERIabUlpSmqtnHsRUXevzHhGYeiPM8+ieFc3bRL8ANtH2+sUL9oI32WFe2EnGBaZGRsIH2QmZtFh
ku9gktn1uaa9QTmLvSSAxabBBQbi63LQ8/VPkuDd/exbHCflx53KV2WaGG8qVWvIGYjVUNSiIo/6
KYXexPQmCUh0SOxWiwPmOV5BAW65nNt69ZPFB8sdD1QjYADqGbc5A3LUifdD5aQYdXarW2wv+Xm5
8ozXOX0ccYi+8Tl01qYu4KqSp77//LSymAYBW0Ago9Nw9iGEalHnk8UV7noIPVCiWd+eRvgzBVAy
Zw+vT+r2mEO/WqIybaYFvlfgW51oIXrlHpNZK30USyj0ESG6TU7PzkVhC8pzITxKJyc3RY8MLg8H
3t9fMDe2gijwcVHHtl1MdeI7lLU293FwNR8jkvvH6klDw6n5qvzja6nncBXLv7KeyEEBBR7SqKzm
61kFflMEYFAvO4X83i1GAINxlU31vCQsY+Jw8jVckGMbhnojxPg4BQ1yp9m1oyEJ3KupAFLcwPzh
DI7q0Jh2WHprvQ7t+mSf1vsAgTKnc3SPzhLlGtnz9GO+mOtNTeBLWnVWk7mUE8tEC3k+qeQf5GHn
DKj+zMdjgiMCh8X4iv+6OE1cDw0UsOoWQQEizMGrSIHa1CUsHh7YjJ0ZbhhOWyZLjJHUCkY4Y1US
bKUZcJ0WIXon8CS98lENDyHTpWn8x4nTUXm+hdUuMJsWBTLZj4kTaovI/fM79PaOj4J4SKGtk5kv
rZtFxD+/XWaey3bk0Z4KlsXDUA/g3E7nSsCuZaZWY473dTXCT/n1rAYSo87vum6cr4LHx4frNv8P
hO961MXki8iuMw2+Nuuy0Y1vr5jX4uO+5H/UjIyAVptZMbwVjuAbIWsbYDPK/n8ZtpSFRmnp1UOb
149nFeLLz1+4WvjJ7FQOc2fDHV9ndhrsdNKNUXwIklYvBeY01FIHnhX+xUtJUCQ10/v6l7KTFAba
QSg3Wv8FDFVG0unEAPoj9DLdShPQu1dYv+PWwI9q3VZuqdD5KO3GR1g6Ue2N05kPheVEfiNc/Eix
b6tve8s/x4fJkQtwwi/oDDj2JTmRkm5W5WwFjYP/goV3TjhW+5GnabX19iXpg6yBeZ2bTU2Tqzhj
MGxfUJyUhLmFLe68tzBlvEJRhbYJsbB6UP00q8VJKE1xQFOr+51tmFA1ENAmdPuxTeo/k8Lx6h1O
u4AOouYb98+8lluiakEFQ3pJOaCdlk+2MFuyjqECgptYoYT7JQHcIgf/k9hPYx6hLRGY1QZHFymh
ChGWUdauqaCnG8aTK4kKh8oJieo/kp3Fnnq5sYGQyET7d1KyFf6oLRwyuzIP/VR6vzwkCCovWZKR
gd54xwqRxJYwp7QOfngVt+HuKTURxczPbpSXbLs8qsp/cMzg3SjV6fkKxycna+3nfmb4EYp1Uqnh
CHPebIKMvMOQBfS5IeUFoZS1QwLeU29+FHnjVEsENzZt1bGoBVK9quRO5/uViIuGWOiNceUUZGy4
Y0AlLSPbDg4bjGqeOHiKd3LmKrYIJS/8UrSAxd/Z51BacSA1YG3ugdD4ur0bb1bKNu55LxYavAS9
URtFPHRMht1g1hswPAvYuD1VwJFIB8OktUpf0A9dwl6GexaNF2dHH3RzhwbqJkB3d9KmVZViMNkN
gjY5vN3juvqXe4S7k+YE7zC7Ts1WGG5QDZEJ06AfnRmlLfpc6KhqpRfKVEKrLYC0uwhUaXeIqDbn
dNd/otJduXa/K/hxgHnMBIGuDUDV6u0gbwXIp0sp71GYj8MSUNER3l19NlP70GlMDsaLjcL5FRgd
0Rwp5z5YleqXjJ+GantzL4218tHl9NNSGk0ZMyNpLctRsiokhMafVEklvLwraonTLDfRY/8yZ62h
O/b11pgUxcBlCq/UbFc7erV07w+1zhIFnf47liMjZsjT1YSkncg8mruzYaMtN9D22Hf06y1A9faB
8FncnL+jG67TvYopMDVpKclAH/B4hdwLd4dhvD4mJXj7ENWY8sYv88hK5FUdxt2W1TKb2z8E6d9l
zZqLoGabttzIF3xKy3SpwWQxOyFRRwMvNmPSozyBxioumJK8I9xOXzV5Lxlj+IfCRkAYspr1wwMJ
Kak+LPTVo12L+WQ/LPr+ST3Bw7v/wGcMaLcLeZOCcT1BcjpvJP9Q8+XX7uL3q0WbjjQZAUqSYJ67
xkx19//PafSwIJ1hSkCKYg4ZQrqbnCE0wgGHY0H0ZdczT6AOMxnObRTVkSZTmDAqYr9cg9jivI5+
xvRtKbzm565j6a4zrYtXq1pUU+Da+JXYQsKNxeukFOzytjYgOc4EKc468Y3fYjT8o1z63sqTGxwK
5fOrnDCEr5goGxyDmxhQas5zfJd4qiAow/VXNjHpyClswlkHoDwNNIfSp9vMyyxEJEoDxw4PPE4i
mFkX4s92TQc+rx/YxBD/Xo5q/wg4oIj1TVy1BnWWv7e7LUTcxc1Y/m7Wj9CZ8jDH4eObrO8t6/BC
+9Lr9qEctTXWEs3lVFrZeRKaUXbXeVMU2Dnez3ikAwRFuaisz3+ro40QiOT9n+7axwkMllj25oHx
pT4HlFLvjH8hajOSn59MMeMmkMlz/nmDYuNUajOtpl/0aTYfspZalmTbb3eSIKYKQgm/iYLC7Xnw
kt4Ke5lYR8CFKBPyEKhwnPEtiOpNyIFjV0VPRmLQuRpT83JMXul8cPI1XHY2vp8bVjkWYgrBb6la
SESdW+TYlanbpu2RBZQqOufAQ+oxMjcRcZSYQq6tn3cH4Hm9iIGJlxUrARCQ8hQATvoMThcHqV3t
IJY4gWXHPlVVmeNVirhhKwiUUrJqnFAsvQ92u5QpxKmv8A3pwQCJDtKuXafSQrReqxMu+PGeLeYv
0ETSwA9ktk1RvpbgU7uXS6SWw/m2zgVc9cm1YDT3habEoFoahIdtvk6i/z5ERRB1FZDOeTNO7icj
Nh+iXzlEM7KYkCT3fzM68B6SL6vCMXvE5pMVwA0KiZ+G41pghjBuZIVjF24XBaNEwK0djiQMqlpf
C8sX7HsDM4AihcZ3g+YlH6HzkLpftBgR6GjevuUpiLtEvc7njzgG94ttldQ6i2b0fkjT83fXjocY
b8kk0hOBncebh4rLv7oum+uxBIyyCPei4wmliAkihOvlhO3ckTH/sQINVEUU8tJLotxjmnhCyY+a
yd0fqHs8Mb77RkXKOdyX5XPgVgC+RRYY1GWgLsKPSCpcavCF5XlU5A0RZNAMWLWyfLGFIK85LODR
Fa1SEMDtBZRSybnflaJeNZsUXiFBtDYpVc9JMG1c8pyqAS1CLP5jIfncc2bY0IlQxqZymcg8O8WH
ss92HxfTkMdq07rrRUREVbzYiljEzkJM90N9mbLjxErQG3z7XG71aRnZKKZHJm0u3roGZDpeitRj
eWGZSNM39MS3AjeXWDqFNqszw9eMxVgIxjsBopGycmnN5VR43aMtXYdDpDNdQsj/vdiIi/XDKJS/
uXUHFyqGI2l6ULl9a/capI1n2ysucaE/SmeRASRtSuxJ53aun5KtwHPi4upz+jEEUxImJDN7Mjpq
PRjNBn7qJbJURQXg0OP/j864M525C3ehxwhtbt1B/rfnxvXEm6hHNeACQIeXPbYEwoXIDrk2IFPZ
Xb1Lb7nOlAMHQyMmvDP/swfAaZc/gjy0YF7JQWDO7r/MNa/47nbyAEDhVxMmoHXp5Sz+M6NwRIeK
gTzTD+dO/8LFwkeHqycxZB5VHJWWf2qlQPSlo76Y3oTYF3o3wiWZh9i6zqg9k/tCTPcn5yxyzYza
8UkzOHskNocFuEJF16vIs+Sby5r67kQ6ZF08HB2kzraSBAuuzZwuFfq58aFZw0fERJTjdFSJAbq+
9Ra1t1GJg7xk/vTjMfGDzHoSdf9aCXsa6G1SfJOwgD63RpWHu6+v1ZH+70vDbAIS857j52MYDI2Q
7tdQQjRYu7G9BoFFYQ2hbkOg75rFfTKpW4Js7H0BNAhCgGnZhmj3Ut6mEEVkv5iFPsWHd3FrN1N5
IAuhONn6hqG0NtrOQ8qBB32Vumomw/57nR8E4C55FvVcdP14PLizleRfdKQ9rqhrGZDp7CZb7VW6
rPAXd7prVLDiEuFBKgHNT2Px0yxaOmczMZDgmKUZZWhy8s1ODalXy34/55B1BCHHHuR2LMcB1DQs
c/LtIXrbctGVNoiDXZGM/vMJmp00uTXLceFDAT3CWpCnIB8ySKF9Uor3ffW49bruN7R4FMtisknw
ehSHQ0vPo2ALvGRuhvhPawweVsvTYGfXiNcCvNS7EPIDEmIam3FHq+37RX0PiZDm5h+EXQgGsXGz
gazVPA+vLsongyo36dUUfgwHKx21/J3vMhx7JrHIzZR6Oz+/8iAULrsvq9mB0rGIgSabXWFcJc0N
5hmY4we1Jh9qyuCo9EWj8XXYZHF0w0SgK672gUxUsaSK5x+NwVRGlv63ieuttRBd/XrRPsltsgpK
UmlBeJ9p6gQxDqzX7+hkqB2QPMc0KQEChgDr/oEVQTF/V5ugi5pKLMHNbdafyL68sUJzsJg6t3+z
nmnqip3PIoCkqDKs5GCKVnyo17AZjH7axYCpAP9jEdjTJl9mDrVwhaKcOMh8LgDBpI0E0tIW4Dhr
VZIp2B+X39UkLy/Rm16VjJXCepu/IqKP4W//+cHE5TYdnix1XBTs+P9KNvsFdzwUQT3vM8SH29dw
o6fYke+JLKE0jSer/HEqkS53QLhIJztbw9l0FWfdaJYGv0uvCfTetN9ZYlGURGUUkj5sXhoRAW3q
MjCiSM82gj4kKqqXMcUju3GqIeNIBUddo3X/67xriJ1tky2VCipws7kMptMelQ9I8ImJHc4LjOAF
E1dMsPVhJgpvzvyOzkzEmqoh/dwJNs7FI16CLwape9G7qN8yLXGqK0YpOBDCWQhukNg9NPI8TUsr
vGT4jK7K7KeJXyofatT8Pezp3MK9q6beiYNnQSdDjRWljFyOdnQKdxdnABPtjCVwKX6GKiIJUbVT
gVIpV5IQr+0yi7UYsaZzxtzH3Iec5qGAJspfQ4aV37263AZHJeDEtboP/K2BytTePceAAxuzaSni
UdXtQlesto0OMw7ecoUVGzFrrRp3ZkMSY2dRR4fTu7bltNUDhFjmjIiu+qDsUbReCNWChXtC0CEq
GIww9xQmUKZ/MBEpsCDZPEDXVz8V8Xgky02AfdN6jUT5c4Pm/ZGpdXe2SI2v38Wiv0Ba96VZBhU+
2GBBhZC99ieY5EDtLuslasR1oVkbPPGj97SsWEwkbRd1Q1CgysOFh+qvA9oCmbRKkHZVzjt5eDX5
4aQPzTLd6B0DlAxf7XLRwbSmJwVV4t81kcIwOLTpYvHoCIbHzus6WTy2ndrYKX/cGRzhTqJgq1PM
JfV7/qxOzOwMDCLOuACvdw3WGVX+LvKFpcOu+G/izjTJb7dNNQByIVqgghBJ70xRoZCQOtPk8R6Y
CG7RuWa1zci5UcTIFgLxa1ZouV0Bi2wHLzZeWphus7twrj2l3rqcLNGWlQpa7vg59g64ZyKqmQlj
GvjyM/uiZp/VD2n17NQgkxpDiKTfKSfJ8MRd4KmEqwNNz3vBbrrKHSRTBNmrew8CQDl56+Mfcs2b
cO9nQOqgx4WBsclzYEKT2Vrj7d3ORfhZj7NJe0OP19CeM/vYxEdUpaRny03smVb0C3SoCgzO8jvz
K95vF65LlleLtaSF7y95X/x823zuzcCsEYLkpiXvRXueNr1rpVQvVIaJ+B+SzFiaI2HKnYMp2htg
zsEuxWKkKgF3EL4/dm40Jd3ztUpf2jMVCRgt6GEIR1S6VV8wre0+q9mlSWgpp5N5ZTC5PMigOYDG
aC4achnvjP2eaKD2h8sbbfdT+qw80yuThneynNCYW0JTJw73K1PyYTEimkArl36Z3fNIT+qy18sp
FegRsQFX/G4CKtEqb0SFN3LDV4R/AsHl3d6TsLqdcJhPSbul4H/B9SKtQSNEaEesWyOmnfVrqaj/
5epbH2xEK1BMCjvnR2QYTrIprS64wXdt9aklKbBd58N1Duch+aCYc3AqnnW0RE/cUlVEn9EBltgq
3/Q6hj4j2ARRXhm1NC5+RD26SdsQ19lGDwK2jSOs7L3GUprffdTWB+hEfSLE1lsdr6zWgw9DPBgJ
kCG7A+iZwCK7sK4d+Sg11Vde8YsXMF9t0n6Cd72soje+y93AWFWUWYwLx6EcYtG6dNTsUen6FiK3
Mys1q9zC+v60Mq1Nh0mXb5G2DbCogGwchssliiMXjjtzk9M4+5dW7SGj8rMd5owc783hY42WFwJu
Z0lBllkQ9W3gbIWn/3ISOapdvKCzzDknhVMphM0Kv7ev12dX21SulMp7iEmiQscnarMXA9oHj5Q8
mvVQdZ4nEuIsMudW97Mnymxz66CHEwmUzls9AQY/eVGeC0zQZ5Y/Ab4Fjm4AO+kW6bBJ+r+QMMW0
BQNhfPrOQOCDXxCD/QavNp7E5Ej90vBYabVFSp+mHoahigZfgFVpvS6edYa5KDkJuxLXb3Ajy35J
ljYP3dAi+FPFqajtowQKqFT3HQBJmV2jLkvAKp29k2/hh+MONHBhLuHAnWCcBnhiu5MwnPGJy9QR
t0lIpSbCpt4hqs5/RIPhOrIVu9ZlySb6HP+HQ77/0V9Q6WmyO8Gjvc5JBne0BVgsbVtkIKxktkNP
NT/6cthewDinyVyM280FsJEk8GolOPxj7hrU0vRUnpZmyrPaQhotE/82/U1Ls5Kt+r3Wpmor7VvG
nZJE9JHDwDl8zpty7enXqqKbNVXyu98an7VtAXiR+oxOIzegXUkx4bdZXrpJkVoege+/T0/7IBwi
JXzU+eHgFzHyf9+jonxTvI0KRpkD45L6wKX2Pa/v8bPYJskCPeiRyfe3tYzKW5YAIeVlMvQpwfCt
ZYqCKRtyZnJFfxRg8b9mkPitkkz46BQA9KkzcakRU/l5hU8fpo3RDcd7RrLTUAKjKaESrHyAQVuf
1k659WD94d6CeFMvEU+xLVdFyc5Z3AIDCqQiPFG5You7tKDs7sWRAh2bZcRpZxDyL0SspfL13BBK
PwTdRsdGg3Saa0ogpVm/ouzDBICRVEBccJfu+FbuHWTte6Eba5RvGIL//BgkSF268YB8XaWka1GT
JYmnbS0imEYDX1lpfuX/qR1utQxzsc40dN7FFDR4eGyI9yGNLa6PhpU5+yBFX51xuqs+u02QwllY
BwaKKeZ7fAHJ3pcFh+7QUgwLKBApNa1tXd96DQurAwgUeeVdY4xzb3xpo5+1op7mv3z/TNLpa1x7
smGEbcHkqAYEtrJdhq9QVFqr8gyE6FPGiCg2MSiMLuKFdMdsiRafyb1d3FuRH/4owfsP2fVFKPaN
FOocEV6QpmbaJuom5OiTD/uQmX57Cwyc/fPYOGqNRSkzu0QCWGeAMYgUmvwookx+XFVJv/bXlgKE
OCAMR9QfCWdgFX2582f8+ygl8oKYyNqHlyUM3QHxwF5lxzI+y58Pv0M5aA/wcGc4yqVIamJ/2NDU
kduFRvxK1PAM/u6JC8sNdcdGRcIc908rvH7ULP+OhISR81ch4YVgeNaKXspJSxCY3aNVuebHpaSB
2yeqBVPYmzZdfffBh8mLoMVlfbZm/m7SPM8qiQp7jFfn06H+ttapI2TgJMtS1M9LlFIbH708TlvJ
ljQCKZ+Rk+eUjA/A6tKGTJvxqGt1y8wUzLu+l4gy96xmPtp2vZ28xlO1LfYeNUI5WyZTntZuv5iY
Nf5W1SPoyGgAi088nAS7j87nCdnGjOedlc/GlZl8MxhhKeqe2KiCUfPYPM7ZJVuWw3drGVbuJxsw
Y9vTGIyTkFt1HDOJs2UymwkHMkP/9jOYDCQD7gUV1zEj8qhDN5jTMNO23+tuhZzqrnx6plupacr0
YMoxXWoj8MuOISy5YWBdHGHp6jrgJSuuOrSucnG2ofP2qtPF52mNGtsQfYBjAZTaPOtEP+hZ/QKM
CbYtSyVGosnbnrRmm2y0ay1ZhpIsjmY2bQgX3uJ4MI6WK4WiJg95Y5LSD/HKC47a8qsq2TtKgZN5
AEn+B+yfqaG4XrFObwE7nUm8xhgxCd0x/IoH0CMPCyapepLvdKfaUEIkSktH1yw8wANCfV2nRojK
3WCFw1TAues/dOcyZdtRqqIxYqS/N/VT9hihWwkZDdtuUhWpTZuN2Gy1QVm8uOJZywNVQkXOd5ik
Z7VtocqgESpdsvTwYrD9Bvefg5IAzGag/jbT0L5XVroBP6i/A8SOyuzRAlhP97LQ5RmpqLWy5UCn
GFBUKbx9F4fEW4tFRcNaVq5ZdHIL+efWuvHODtikMiPRuAeQHi3JEK9CrfFoyDwW1SPnIGMxEQEO
9qk0ci6CGB/vyj/RkedpznSLJmQ2yw9PXoVrUnr0V46jezp4xOQt65wZN5VOY93IRbBxyoLIm9pA
tvGiZlSQIwH8e69cGV/5Z5zw+Se1UswjKUsuxvGl0pwQA3/SKUeochieToKvWCMVbw0LR195INV9
hFEY/AmdIHcg/GftP490wzXA/mWAvl1vkW+XVFMVACUbavgnUmpdYDG2Teqj37BIv0iLaGirBLZJ
4Hy7hwsnxzdR23tOdGb5TuKw3C/c4/u25p4sswcXgoCjrsOmj21Ba0LPm3sMWID3RXrDq/xm0HWH
VmfcPNDN6543js2xHtESkvrG1mIuhUNuvyJttJARQEIfKg1qovCDX3mNXsW+U7lZRv39W6kQxQRl
Max8WxCBiTDJANoKg6rc7UQ08gUa8BNvnY+jO4AlHoJ4qNtY4uSTpmhB462eBYROkh6qbjhdsm+M
jZXrl6xAjJJjkDBGXplgRC66AziJryiGsNGmGqK3UkDmeulH6aC7BWJ1b+4TtDJXkA9A+EIAe2yD
DG47ynLSKn+EEOJkDqFkAyMWGCSFqin/ClMa9Cf34Ink+724wxoxBUG+2aX/kDr+hvYgnLvfQIAZ
Sk8XZvFaZY2S5Yq1J7U9ycGGjZ/y9M/iS0nVbXOQ4+4QdcliMSabDLySOB74ERO9C/j/L1dzszFD
OqPcVgCRWcozBENhl79tFtf9KK0jRcVBkvXq+nhwKwd0VNn7MX3FoPG0fmdyh0pr8qzoYELRWDla
reCI/jD+vuzg0pp+DOE8OhRDqoyzQZXXS5EQE+Dvi/6+iIGTaNjp6yqzYUWZgDy6KTL3IN7kbLy2
zmN7EsQNGm30UReN1c7/6ZEWLQvWfGP1ZEQRLemKxZpc1uGL9LBMJHPK3Xcagq5p3V2UkMgxHVYk
yG35Yx3N8OyNjYbbtO1FcCg9n7qyUJ9C1DFd2oB8hI6zsp/gqNXVGyhquNu8eHCJHUbIqOJSCkCC
EpmQTee98TGES6kSmbEZWb9YhslYfqmQcztFqUCbde+py67vTT6sSlozf4+lzqe03Tj55CIyvY7J
0VP/V4XZrV0ve50rXhWD44IF+S2igWLiuWOHa2uIKScD3BkuZpbeMonAFbl33VJ2JMwCnu29kBK9
KGulLC5kFlbshXxXa3YkDJJSVQi4kfn8rmqOfQSwwR1ohC6pIHuAO5oWIbqPeIImNL+pmsgP8n83
7wfDBBgO3Z7VNNKXXvcS4SHHomz7bY4e16SpTJ8hb+Jum1zXL4XcQQsPaQgsQZDkepsoQNXUViO0
2QU+ienYm3VLVKerdAlFqtmUkmSy8f9Rea8L/M+z0zvhwKhjKDjCkVaK3JveN81DifavpdcoKwuS
6Eeg/S2LU5ldKMM3lnpDVsWIgapDjFFwmBD657RnB6ih9bB5vkXQijpovS9USck1mInrhlDL5keS
CmZ98zSIsSfeFamKsscXQzB01t3MvjD54kSfl2wevM2mahTVCh5eRVOV9EYj4wZG3IPUgq0jjF6m
/ul4DHbuGA8bjF2J0d8se9sm9xSsesg+K843d2kTwoPCacewhqoekLCSmus+r7rqxEufciDLUuoJ
zrhoVm097v243bTQfJ2FauxTEa4Bn5dWY1QGd3HPhZBfbXFHXkHT8uU6lE/knRJqklNbqGkom6gS
S7etJokd4uW0z+fBTTZwZ27smqAlAdsac6W1WHxR7fhQzmvtj+6VNmoUHeQk7wcuwyhWlxxfTCS8
4uOXci0ZnBRqEQuPKRpa4iU1Xt3Trk1Fm2p8NFxzHfFu0SqB6nbpzFvn8NS+5F1IPLw93t5FZM0i
8MWl38+w0GahN48bYAXOYvBcgOecnecTuBG3a3hR91PdKMtm88u9hDEFzOfSGbEcf9vzJvVPFaK6
02pnFovBsAEoHUlp+mbvrFX1cQpwUsLqqNpeF7TAGtY6m/NIElpq2d0SftXFV75k+Xrj12mu71XE
kRx6HMk+ILdIlUikzzAcs/g5mztab61GBrAfzgbGRI7w7H1hznphq0Fi3lRN/Y2a1LZBfbXJ/SXY
dK9uxdBLwHt5+g8Qdj9Pizu4hdt/2+BwSLpHIl4DgcW4wMs0qOo83/5Vzdh83LSHFfm9fGa4wBRd
oOoZYV3AtVutXXNpNnCmFcIb8I1jtal2MK4BZuWcDAhTU2941HWans6w2PnvWpJfU3hsp9EMjrMu
l1rjlxCmPPuqI1m8sATye/SIzQnDOMhN8iMaNpFTwwzuZwUYjmgt1P+nmfUd7VaCUyL/AC7w90CU
Q3+oUHxXJ7NOpaN9MZ2Y4AUVPBnKyk61EdOAz/OZLau3I6QqFInRnc0sCdZiMyySlCSuGxVXFEwQ
xUtRdSzrmJP38NsbMf84Em2FfGaReILe1M4VXVfeDBT4H8lRfFizLnmovwqmnmMYEPOTbUMejHwr
12HO3ypTyDX73mKlDn/XUf/PoOxlSHFlzDXofv4n/Ek7XrhjPiACriATHEw7tTjL8DCAVHF5oFVF
Dhdy4JvQVE5/lXmUaWiB4HptMfOQXUPsQFCOA0SV5JOUfvljH06W0PrCmxAnSR6xlpYWvRv9fk5W
3YtfaB4aUKKpExqQfZWKl03rwjywUybjDT98jhgRuD8jUBfpn0u3Cm+pDFC2WE4TYcAYiTTNLDCT
1Riz1Ar61TPWIUCCWAm7geromftAPsLnYJ54FcNzvLDrKJ1zSNUpUI/c4u5kaebEFD8Z9TUQ+8RO
8udHbrxrJYrSUsMjt6+uujtOGNbvOU/koz7HCUxkJE9CWInKtBEKq5qw/tlEPZcwGWVn9A/EjeXQ
1cZjeJHle+tZBXfb0VMPIbyA2NJCe2Tvykmbpe6EiVbWwC/HwaGadsURUWQtuRTx+zVNwHTCSZSJ
rPOuoNbqKoQOl12vo+Vpqr5FjQZuZg6aQ6cBpjYJ6mXjG92v1Jb2nMIjiVcpkmlAVjA6X60HezB1
1dGlHFzIew/dJBU3giqPfGKldhm/AXqWDjZFhlMEzLkKyc1fhaNOeE2BqxRrDUtez40Pl8JKQzl0
6pMkx/eJOdYBWNyDBgk7aah3lVCA3jtm1Olg8miy0P7wSLnGUw+7j9kNsx/jm0jXZw4SFUrvol/U
m6Eahg1Qv6vKn1JsmMFfGnft0smTnFeYiBg6+OBnlcmruKRTBmT/U2Vmcg2mn17NZkeBYsI5799W
A92tTqJas+z8q8TGkavPwVB1uG0vARgMlokgqsKHqL2QGBqKaHUPzmWlYjhav0gMdaNt/ZCvsOoz
kamfa8xbyiuqQ5XwQuI9OjUZt50vyUl+svklCIpxJ/pGOm46wS4qta2PHxPWPnui6rGDggTQetck
NA1gn1r6+Bsap2ZldbMV6ePMN8XZTIsJqPRQHWZgY5l9PmSWwNr8IQ6yeEUWRUS17MeFftJJHzDq
mWYIPHARydnTvLmeUnQhIS5LlKvsctPLKRI2W3JfNkuvimyrzueNe+JDHwvrRiGFZx7eIxD2A4Ti
4QYDllycHHcGM0uOBrXk3CHSYf1+AWO7Ew+uKhPZjixMcWaQ1ZySedGICBSvGacyzd67hJ7VXKHK
qzun/GwfK19iSE1J0Em6ORCLgKOCY0291eBFEI2caLQEusQBnJsgTEntNQ1cKf5NR5PDQO3CFE4z
dSkAl2yjau8cJtSB3GcW52YifVXZcgAPDPOS7ZDk67XToZ/E5Nj/RBkbpL2GgP5AfiV5Ny2j9EZE
hPaldxJ1uk/qIdyyePWl9Qvi2VYtd4vD6rcg5dXjxr0Z92YTCmieJ8U7QBK34qYeTZsEPrDjGIsb
cuXaeemHHO0e3TPLFeYo4m75INmpeLpu6S7hKpmk2NNERpXnDOf8/qHe0k2zubd/yjnOg8XXYDvB
QoRGx5s8U02F7rQGn+BytZz2tB9Jii7p6fFxMSLhuOCtTmvaxVwFAI3htw1hADhlCTeAciZlNqg1
8gqKS3ujxjjlfVleB2WWulLjEDUsnYS4jQR4Yi3cXO+2McDOiJRn/cvqga/J/nDS4Hhb3TAZBwmL
OQDsTT8YTh20LGKNtuC+k9GlKIULSkWcFRJSWWAe9f366n+sO8s770RBVQ2n3CZ3u0hdR2oVIMvu
ugvjONCYi7YrM3PcUSzIFuRtOgatD8h2958/XL9iZugT0XyY0b+dgBswgo7ZCzSp9RM0hupgetDA
ILWQnot0UT24HCcb82j/ZEcnEXd/Yga6B5bgUuhyPlJHbIJkM30ZEqWQjL+djKrecV0jlwMd02cT
B1iGxP0ChkdV4ieNY6WWGXXkIO+nB73kY+7UJQ/WGnsPvFgOBWMmOUMsPKjk5xrNEzp9pCM6CbZW
SZQcVZLz1aJ/WVh5WS8b7Y3277q55V9mUyFk539uFgvafv7sf3qAt3Bc7UkMf293qkRijIgH+s6c
d61rAoYC//K1k0lPbxp0CnmcvfWmOtd05z6r1XL+MFB/aEU6WR0zcmvSXYpCvs0pgGkGIDYn0sF0
7a1fmERwypQztCJ4fLdZYf4NPNg1AHqxtJKX2gMk5rvIsowZfnQr5q5owfiyqUafiN5QtyzzuZ3r
0SiHCQMDACa49jTKm+RQbb5P4Q9H5xHH6gnJrOIB/1oEyb/t7MiBWf0LUD5t9BKtQZEZ3kbRI81R
oSxUnPKZGUwaC2R06BLhyOCitDH761dvG6hOXzju4LKpdFwthFG0mlHkT/YfYJeUlEjzv1pZQ3iw
FJNzaz9WTcMD7KsgKVyyH5Cp3YVaofQpyeRiW8cfaebLIqw58t74eqAXNcAUJjD/RAG7BS916z1+
1D2EraX035+bFlgfp24UQE/U9zJut64Qvo/qaNGsY8yCA2kio8II4hpc3IvEZ4VAF3jBicdYEOhN
iffLdJsxL9Oq2e8N60jtlZT/tD7gXsrLjJUIqMfegZqcD5XC4dV7CeXxRRtB4xaQMRomfGdZo3Dn
LHoqOYt6HLmnq1rU5+J5yNgUXv7DjnfTMsk5/fj/SAHDVIkNGBT8LGr8RhBO/YRKzXGWo7UOAAAi
9oqkwdmNablJQFplIx9rDxngg1I8EdlwC0Jwg/7nuj8Oo4Kt6LgXQh2vCg9F0XO4yvsDtJCj1uHL
Zz6XmZtkFaec7jJT/DPXtVDHOaVpPOPamjMs5C9MFPk7dAKkhl1HQkpVhNLZtzhxykg6FDNguEGu
80MSxEZrQbTHm9uOwdICbel1CyIUWZn9N9O4zCit2LQc/rO0soi7mdbfy3jjsOHBExCq+MKsRU1i
ciGJFG7UG0VF7H1yhtul6LsF7KnyZ2otudgK5yXNblaceQ5PNhOVnPusgKku+aN8Fpsh3GCHQYMT
bgx47X1GlcKk7jOOp/FAnYcttd0V9I8C3rRkjjy2GC7eEoZgYU/TcOkwdebVrdWVjway8hC26Qsh
mIIkyuc6V9qiLrXU9udd3SAoiJJkjGDar2A0WzuOKuxc9hGsb32yxQAfVg7lWnOzBxlsykV60nFR
9DEWhCIcO30akKpfJfWg3jE9XPciHjmKjmE6ec3BdFuGj/eQr0JfE8IRpIe5rl7PT8upBrM8XjJy
53E7kFufZakTynrCKGvJ5L/P6RKl9zzKeQgYHN79jbRJrht7UlQNg0Uv8CgBQBShBMKpRbzTmpn9
Y/Hieh5PGB76mLszOShPazYv1YdgbjPDPCOUKfRCrnBT7lz9XGp3w7ZB5o7rF9XgaaWB2fxxQEhS
CzR1TdmsR4EgQoPOTJRG2KDpUxJBCNocXz7/Cbyichcr4zBKtjLNxxRVsn64ZvTBsOOZ27JBz5PM
pS2JqV5+nkU1u8CnYO/ssD5me9kZNsbKowcaPUdfodj7Le3bzdnzOBsPRP9PVJgdxoQtqcQjW7sG
CrNfLKKXGlU6IcIv0/Er+tR4Q26WvUxsYo4oWLYzLK/DmPGTs3SPfyGKvo7Hj1kb6bTmfc6q7ptC
quyiKHTKPk2hWhaEsXg1swZb2PzNAGxwyI2xjo3RA9igdg0FDHSodCXdd0Ca6F+UKen+Uz/pmOTS
CBp6KDVs/Hn9c+6FAo1yBtJv0J9JcZdXkcZKgoRnXKGwCoIWzPbAnWXJg2jPaz7xTpPU0vxn2AWM
0LqrDGgOEIrBEe6YjrpOG3/uvYk+OtKjWfJeTQl4aXLjMDEA5jVehbmSaLW50ZdM555Zm1JIecoZ
9Ln1pKS0KB8DI1VDWbs3J/1O9J+GCR8mPyIK6qKEV9lXz/rGYY9ru9kGDoeaiQ/exjon8W/a4bN/
I9AFQt+ozEV4GtAuiT2u+0mbSLM0eebJ1LX95KY8wsvLjhrantOfBEa6r4sxRc5GrkbQkOlfen/h
+i69Ba9KqjdX8wyHUOs7f4gPhlVJpowWsWRW6cf24SynW0u6GAieLCP58CcPDs3ne2JeY9C2bMRA
BtGzAiu8MaZieG8SwqdQaN2odFasO4Ri3yx5gzpUPCieatl5GdtbhKFRAk779z/aAp8VXbyKraYv
W9qUwR21h+u4oiGUBDX+VXwSwGzWM0gSb02hRVV/ASANLznEamknoENe/nO6opF2c5KxlttItSTC
9wDU0rRNMf9LBtf5NvDv2X5WAKKjpG8iVF9kXt/cu2qQ+YIL2OxvTdykDkVjVVBu7u5d5cJtdSkH
4dUn2ctSTVJ7oI1hTycUq0oaaFyVSLR/vPwveC+tnmUwh9CscQSqYFq8+aATsIYA1JeQq7ERnLKv
qbFvnxCz1x7fVl5n7JN8T8TWI7Iv9oNnkxE+knUqF7Ou0/hblIDLwQUFbM2IerG4h3bUIFA/jgSa
VqpttSa7Tl+xCmrzx3jQY8G/PTyuel478dqn86BMb8np/9jPotiy+1G77oSGBl1fLTYkFIBRlS4M
DaWaGCSCw3yhHcHTLNc8uUWoDyIDcDFBwzwVlE5AMXF1bwmcgYxgVHuXjcnrBPW1beENiL+/7CKV
E8iDTYmQkjeBoEc7/LD6AYgC1l89YDdiLSyKqNS47uI02MB5Xk/GzWdadVouZs2ey/B3jLfDHk60
jQF+kbHAvFAfJLJKU+JuxyzIMoLHE9WZi3G471p4fGJnO2ulaxFbxedP4qoggrKvZstT2zYndV6a
Bpyl3YhocSSAQYMA+2LB44uuzFJyYZfyrKZ8OAoqv4HdnP+hQZ2/QJfFDy/kqCzOq0NdlO6woFbb
H2XOk3ipiccTOBX+OTk5jmNYeVVgK1lI7KBYroRN63VCMeyuWfTzSJyCQLbu9SX4wW2NVDd6HjNg
Uc3mhtRpn9C8yYkAPE3B3Oa3FnE0tmZIHaW1aT3qjcIAYnVNG/zsfVo96Z7VKJ8o880u7A8wzxCz
eFaqswdmemeuH3cuUMfuPs5JyumcL3tcaXfZ7RlcxBlqFD67CRi0DbFyu7GfP/nIbWl3MFM9h64G
m9+EqXeDkO1iKYJlWLw4p1idpi6mjxBiNWZqnBhgC7f6y3mZ/8fPx9jyAbbHtO2/p9ZH/8mQaKsP
LMB0oBn3SbLkYsDYs+ZQIM2e+b1Y2LFym6nZrz9aBKiso28KC+rIxTYVK8ikDL5Ses+15tL5EVu6
Ha/hIUpmmBG95zP9IIej0GXo9jonEcnPGkEp7Vd/NeONeHoA6EjLQva6rZKtpW6gkPQ9eLadetQS
YcaJg4dzecrDwJ3pQjYOtJftFUlV6kvcAmi46A6JNquCCUvmgkmG3qeW6hlBH2XYkogK0/JysDDr
nBIze5hTMD7bhCq1zksjMGgTvw22kmObXL3VmHKQjDNHsCeWJPGrpfe8m+MHQFep7kJq5FKFuAmq
lH5FITl1/trv+r5RRz12ceE6b2ogB17U2W0Nr+8HtjggI5hQVcj0YtP+bHSB9uUVum3fJVYOxFbZ
FDAQJ/xjrWJZWhIfEXL81pnPDE+XtheAfajd4N9Jd0O3nMNU45yAHg8rU9B+P92CPYFVrrDfGu7U
4iAIOw2a8oFW07cw96IzGI2ZbguTJV6cBqV8n6qY/q749THvjVa7COLjYTAIVIjdZRKkEL7FAA31
te0uV5Zj1jwNNn2vSvkakp88rbfYWjbIEEo/ZmM1q8UrnrJrVElYBqySlXJKFA5QVDvGkODYmrzn
IN7VJsVRibXH0gRLr1NvHkKPj6TYEu6q7IaERIesNgv/rYA8Y9XxF5BW1gdWUlW5HSzHPhH4abcA
wtHuJ/Mjen1S5uH33gPpxT8QsT0bklqru4OQcp1jKUSivxU2fVFFemPF+ibtmI5gMJ+AV9DkLvI/
MN+0SXudGZKYaZcEJti08aCUTzjxAUIB/8PQvHG+g925GBjtiyP2Kkf4eDKTYQo0Dy9E3kmyuBna
KKJNNnWxxeL41ccRvEPEE+9VKtEMqUOjks6riIFgiwxFmdroxJLLjSNo/hjd47G+jSTsnDg7MTae
tOt0klHZtN2Ye2y4qgfr6LXJq8JInsd6rT29dkyCnUXkixza0wRVUQ4fVFeg/B1KKhS+G5FnFtCD
qh7+IIlAIw9vCGbRGB0ZXr4YnQi9E8QqyT7prGY18Rk5MF82GInqdHZrIGsCKuCQAYQdK0HiRkmA
xrNmoN/Pqtt6PI73xsTm3sx/r4rx0bViFv8miTs6qLfXnGR/+727qIPQn2hpQfs49pmIZjPGopZ6
nS1/XihvDdKlE6+GLUDIsf/Tw/HDhNvyACsdf5hb7yymJHiv7xqCYMVRZm6u2P+9cIsA7lsUwlmP
jECHmBLLOrv+LjekSuqR64+dgTSome4ArnvwPtdux1ub/pDu6urLBZ9bB68Kx83Vbs2mmrcyzByN
J22jyi/mw1AFuG31CWRC8yzODBj4vnzFmFwfmhaIo5iOen7b3CEdm+t1+IZPnkeVuR5XJ8peCu2c
VUe+g6DpKKRXgq+sDpG1E8cFxgOUMNUWG9bQhx4y+VVZqlE8yqAJpSHhtuWcldMuNKozBgEA3l5R
UO1TK2L5DEUjXGlkBk94vfM5mTFEWmxnLOGW1HjKAuXAxcb0gjSFCYLhcZ81V0o6cW7wC65h6Hxy
pGtMxklu39KsyyehVoo/Dc3yueXCS6nL9cWR9f+HWiJTABgmEi16LYMfmBOgWUoaY3M/OXYvDSGT
YkoxrozkJTpqQT1boYw0ZU9XRFrPW+9r0S6lGByGkIYjz73HizDs9HhyBu1Ddo4K8aETSG+ADgRQ
ZXOv0gy9u2EfrSK8qr+Az5o4/gaAodv+hPdm/lPF9MdyV5W7jie3piY08LOisD2hy7JrN4/fZfvg
N00RmnDfiJhJW6kHFBSwl22sNseU6B5YgHCN9IsV4AiLMkUrz9DkzJAchM1IhaW9KkA9wrQdIwKp
YYdlNiYAPYtPYRdGAyml1riWNZdS7VXW0Ru+NjQbBTaoPu1L14lu4f0m9LK4i7TYt7CwTNBo6e/O
LcPte1ncUw23IWomjeidIBQ+EughrlXV7ufGxlhhpYLNiVnE2LngXoPmUQ/XuDIvl8fWlRwQ1W56
d7Vz74hwmyMOFwinQeEGnsf95U6a3mFMD+vpg1cdM6X7p/urWrXAZNzB401WmkUWEMFvPCbFIec8
ZaY/fuubhUo+vN5/kg8Q7E1TPWOyljjuWZKABDerO8xcjgnbMm7FLSb6jnzlxGYFZgnm/sF1WIaE
ciRcUtASOKQz8EonPHsGLRPVtIaKLYfHFM6LBV8dEPxNd913eu7TEmJaP78/AUMAQVnHL/H2sfTn
bDSGSkTQhwVLlDim/0RZHCLIubkNjSgaGy4K7dRWlfMLXt1K0WqiVkSrEnyGUrMjSR2E/XRmAstc
3Ukq/tMllum9vmTS0y6WPI1bFPVSHUb83kA81od359CRDykwwu/91GsClony4M1FCsqaSxzOiT1Z
CJqFpB+TUHylzlSWPJfL4mMsv+iP7Z1LPmt6TUa1Bf3UISwSoLeL9O32VI+5sdWITxqVK7Y2LVVO
5t3L2tLejKFm+QRTlZ+JFg14CQ8XdMZNwXoon5JGwD3tSOBI5xXIdkElq6fNHaOy+TlCgm1Gu9ly
7UBnT3f8dP2Sl4JirEGqydX4ZWlPHsQRRCQaXI0+gtO+XaEnPIeM/8P5DZaINEHlrhnVshL9PqZ+
Qg4B2jLJQDc0UgDZ46KAsJToknDiEUmn5g3xU91G9LgmpXwT/6IfUqVBNhRTGrFcKH5dLibkRHq/
PheTXkI/3Wfyv10S3+l0i6jcGr6Qnmaa1ibb9vIyAS2c4PjJB56YZiWt6fK94CxCDZZFfFnO1o72
c5BK+J5G+G3jyqnXcc0GVV4RRwr5BoJxdxB86M+8oY2qSCAo545oU6xnKU76NIa2BwU/HqSdpeG7
kv7L/Qz8h4Krk1aOShpdVbcyoLigbZcBKESvuACmg6ZzIkvlMhyceE9pybASV43SPKOQtviVzZDY
4fpNWYQt6PmGWst0nmIHFCjWAbS2lhxh2dMBqURWJhlZcL/gtgs/8m5zF21bVKPit4P3dUUYGfVV
XH/Lfa0j7F6Lb5eQqaE5+wdPPTvQZkM1YHvLhg5BrUHujc5+RXLFv+8Sdp+Lf7LbPiisYYtOxolv
v4pfWAch/DqMDkN1DofpSaaT0T/qeMifleaa6GwgjV5ziKANhJhfNWT9/Ax7ULmGtq/zwB6ARh30
xvVbbtqka2VTHymp/IGJQGUrOJmDZXKp7NC1FMR5IpZ1AHJIUfezhDiCuHc5OagkXYtQA93EeH/c
mb10pQgpN26CnCTBxFg6wAYdPkBVQH+57OIqw38R+9ItQ4m6mk9NDrpAZwbauYYQlES+MuTu38qn
n8y/n2KiIYdLpy4oDtyGN1PEv9qETrBIFaHfBkkctC3nD+8CRGpvovrDvswWz9xVgIT+Np/TKgGM
NYm/qO2Zaef7j/e7wMsy7CC9IYBQ8d3NsnOSwL6Wdtzs/eK0mdDdbIdz1swPigENRMz6ZE8/tkFS
EobzyjZCGle75FtXknwbxMDioyyEzGWNp1OQJsrZBgQq4S7Zfa4gJszs0lK62jpEooYe9sA1PXxI
hzhpG/WLnUuKFqWJWqQfJzoTfIadTn61pp+lVTN6TDrwrp6IrJqgbAsAzzZAwuuo+1V1NrpQAcDb
PFvldhNoXQH5NAO3M5BRkYfoCdT4ZNGIkfUM4qkNU7BBcDfdiNMgNqoqDt/z5n/MK/mq98qR5+2k
SvphMLRgMe1DbrH7QiKkw8ZniRZtfZEwAxq1LEPM8Vs9UbWMjqvrHkHFdi26UHHh6FPMRKw/w0hM
4TPBemZh2U/Mk8Q2Bu66Kez+qQ5gvfLDcQDForG4mgr2nJhtCJOWTliMeRpjr1O6egGIj0vRsIDh
cRWnxPoyb4qcqHNX9gu4QUAu6euA5SEYSkhonRRQDyq7PHQgmkgScEuIksUUL3IG2Yrf9Q24MAfV
rUpT9O+HmOT/J8pv5oGqoL/Lz0idqQKKmY1AK1c7OTJOiyAxpvwedyCyjBGQrFpIxCoWU/SDtS2t
uUNlXGxSYlH89kg5pk3KB2o231ZdqaP5RP9SUHJwMP/addIu8Y6EUV5YfNQO7vTwVAPdZs9rOM85
5A+Cgiz+iD6CxZg+LNpdc7jkXKB3ksrw+A3dRJnXahSk/Iqf73wcViC3KY4hRamExH4Ev+WPen9x
4JAIYGBV1kL15hP5OFK0x4k+mbKlneAn25VRCnCjNLTE51KvkTov+h4VLuF+e+pnrm57bibLcIvB
tMsj08LuihH4YTmnCdLzw53RRP7n30eSTgk7qyZ/7fmrEeSWZkKmnce2CYYc/l+ZdDgwSfaocxXA
At/1L7JVtDhEZ0Pe4bd5ueeIiWaRcW4x8KkR2nQs2OA3B+0CbTGffwEGSdWrdUzu0f0O92t4SQym
7jEEXtdF5yWUV/DoVqitwwB/0r4TYY69gIcU9uZaKkJvmt5KbJGUHyUZr8ShRFAi6MfmLnsZUorG
PPrTKOJi+lKtm2utXN8Xv0hrFgdcvSWWj6316FjDPaGriIMDvPlS9QXk+rAMo3WIAyOxaK/mEOVo
gu8OjOaoSlvghEGZKxvgZcetOX2Pqi5/24eEWiEUUDZYJo7wpr3N39h1Lh9JmOWb3x6BoKerO7O7
cgqqRwPiD1Xv1GSDxKeTopPlhdwKQcsX/UmcUbkO9pmxd/qQwPvwKA0JvdOi8EAPxRpkLpJyrgky
xgKtL2AlVQo5vwQ5zCpr1CUcY7DHWYS5C2QnFs4hqOX5RwT6SpxjA6eFRQqoHcboCbAYZIs3RE/b
vYvXoihk54O0xy6cbRtP8TWKKVWoF9drGui4Sd8gNnZ/VbH8AQIa8w+etujUIHA8RRvODbguoJMg
JnwYSgvJRPtU7VQxxxupeEcnlaQh7aZ1D4iY9PwxLhefiNDByeigq8StEuqviunhlVaRNVEdnEat
ZQ8gsnurHovuVQqC20rGrIJGDWsz83CeBRBA5U/UeGikMdVC9XkjYtsG08wcoPRrDzpIiXm7JW97
Ml9jMOPJsv/3mgXEIk8xMavynrWev24lvgqEkY3913lYejNzXbJZkmwGdQaUwD7rcHgCfE47SNFj
3ws50HjFs57k1/rUA5l3+YdcEc5dtNr/j2V998GnZvVGTtjEGjlnbpxIuOStB/Dzf1NHOFh4AO6o
km4QyVIWwo0eEpnB/Qjs4Dpi7qIE/rL3djQd8ptH2V69w+S+VK4lZxLMB6TsVAp0sF87rmI899eM
NAhKxhzC2isHvr+255KnpHF5YldKkHstvjjlmZcPjNCLm8gr+KYx61hDXclLD6UvCqQ029hAwg0u
6Nyb6ZKkAQZnQSKEdfutr/55OUae/p8JbhdrF6Ek8nM4qKRfAJwLBkn74Kskhj4HQRo7wiVzrskF
tLxFEHkKCcum9rUA9QgOeYU+ZQ27hf9Kwhiw3Xhm8+MdoGgZ1HPB7g6HmFjytKbznqEwDnSJ//uo
HtFui8EDYKegEcHv186KuKjDSbcQA6bdSs7iPXgGVR5sriuIRGXhNnw0ZwL0WUvDnHpi5RSUKvDI
dgolkYdAJSwu7hOr4okMNX0ufkPveZcrImfK87Ox/5t9jm6QlIvgSeEwuRZ5gx0+YCa76C+fzxb8
XqgeEJbKgEpGO5j4/VOPTOKmjC1mHRobKgFfrB77M4dq6KXv2mF03IvhWM0CgSpSr+5utUH/sroU
Nn+d6JScp/ZZf0l8yyHuIWLf8GMCpKiHPnvuU+1ICvxUDKvciiIeGydKmde34iPEKMgysYUOF75C
0+EBLACMNfUNE3mpBw0ABlwOPpMng4VqYxipGNEBjBieirgV+TUp7JSm0pbKoRGzC473n5D4wy8F
kLtPgd+bN6Bc4iZFCiuBvPD6q73mj3Q8NhMiYyO4nhzoMaaj3dUwAO7sGj4MmIMc7N0lcApdtf29
w6+wmzyfOd7W8lLaHM7tjbNfHF1BkHLgChigylGeZjnolpbc92UpthxBrqSRcX0iJzOBgCJEQrAR
q4KV/c98Zah4I7+yGYDAsw1K/3Akz+t+V7c7bad9R+KvMMtDUxLpxWGsZuZ23W+IToB7w+AVzUlR
EiiiC0877ayNuuZHjH5mDi7orZPKeCdF6TNeOXCodxCYZw74Zq58UvpQUHY18FW6kF59t0d5SQfJ
O7G2jM7dgSR3OpFALnGrnrPbIgcWG9zcEW5soGFclqG7TxoGP1rgWCQSYN3xmgVBcDUOoykICreD
6zxD6Dw3Wf01Uxio/qA/i6a/pY8fbPkXZmpdq6GxGym6EMGjCx9bybB6PMOf1GRsA8ocKEJVlnHj
8DKj7D2C0ptDIHnZ32+C51wsr4ECGU1pADe1NOzFCarC4/bJzntr8xnQHN2zUw6jIBIY2ijsqHai
xXm7MuQw8N9/Ey5NeLbpLg4NIimdww96l9w8j1AwPcU8Ig4jc307cLpmJkIIToBx1qU9AVtOiDYK
JA26sG3R3rTAEAeWclEOeHLrMymK0Fd7zCuFTCwoLOfkYRL04dovh8/1uK2Fy6bPr87yg2BA2T99
9mQfMfOsNPj1ZWCmWRoDiYHZmC/0ALYqtpsyXRxRquIEbb0Y+ab9gxcq+FVjXO7bfiHx0A+pQ7um
iCeKRgs/HOwi1rZXt2DpxFsIQQ7RNdQEO+kuezr7Iz/FoCbbwoZSKNeLwadJhxDTaONp5eB+ZbC/
7t+IsC5wJ7XHDn+J6J3yktxzykTQoNBYxWfyCjYhBodZTrkXEvWD2W/i+EueA+WPVEuHQjWChISz
rkDFaKOWMW6xkqp69p4TSFt36DpzN/7xK6sirc2Ekv1D2NRvo99LBa3I6C0Zir6QSUSIc4MtOj69
k7MF8b0z+S/KSr2ltl2uyjGWui3ZqzmGS/wIl43Ei33r+JB2b/blHdR5d7spHFjW35pkuxdGr6G9
RrDqCIjbjrWUKQJ77HBytOD4MFiHheQKyiHrAMvkJ7jk7P2tKeLQ8OxyTdEdYm47+1zi6UpBEK0j
sgGMd1apVqj6fwHwTomuf/4EA0BEmPJpmIQQQgAxoJp+dU5CKBcKZyZHcBOeQcm7+Pz1Brt8It65
aZbfPIH93Nu1GAEa7nZhJPny9wqH7zVpUu7fW2F+x29OCo0B3SX1lwxPBTs/iZ+pcEAqCnUcb5GK
UlGG+Yf9IA1cz//ertQR5Bu1TwtfXmQnx40T8XfZfdAaL3c5SFfK+o2s4267hCd4053D6s+Mfa92
Ww5vsYlufTWs8Ek2hAQm9YWvcgj0QsXiQUCK/5oM8Il7hYseuxsZN/gm1RAmWgj/CbeIf2kw/XNp
QLtaLx9pTz9MGzXW5O6zZTQFh8CiLQcJ8C6fC9trBV/W/7DItAAG1ydf3HqOBUVypwuckRUyF1ox
uifDlR4B9Ta6IC43iUAEnPzirc+tKRxIPj55mdmMyGt3Nvqj3NSkR7yFCOtcr/b9NVgSHsQhLJv3
27Pp/aHc77voYLCd/LqyU2/0VcpeavpQCOyYIcthyVi9gypFSo9tEK7jUud6yPTMaTaD/Dyg6iPT
LF1nTxPRB1Ml7pj0CfW+K/3914nNm+wpCrhqi9eOivB5cETbU4SMfvWWFQAyQ5c8x35gfW/IDujb
LSTpDyf6lt0TcIiea7uyjQF083pJc2JlXUFmo+Uqot5dSlEIvcbmTqdTbSrZ8iUaBA6xSxeQP9yQ
O3iUkBZfGR3K6wXXeBRKnzOk6ws0HhEcz/Bq4yDenOxVWg1AfmI2+GcIdYvnzhcjwGCNpdjA6q1W
0a4130MjwjgAjHmoVqwd8xhsdaxWj1eUwPclHb2pBKj6yRqYNs/OY6h7sSPpPWPLkTE46CkZiPMj
TW8nF0oQqfhfJk66evgPLrTLKvR8FrEp0N/TJyS8NRgE4UWaOpHzmnmDaQjXa3wlFGu+SfS9x6MA
dyLqQ+IZJQWhjDWEfuU5YKT+rOxxksiNKS8BZcTbBN7SoObxH0a/bEcL4StRQ6b+Aqy2IL5Cxin6
+UDC4O3YRYdyAHVI0IuFSx+15LuJ8A6Ie0+VniBvMvc/AIZklYWs63I7C2zbSn2ayZMRnFPzdKrT
mHdDu7bChLDqaawha0AIOrzEyMnO7jIWQk6PiQsqbKur35wYhNFiB9u2t175a3mr+Eoe1q5/vMwe
1Rqicz/2BxgqBYLCH5UnOyM7uyPdD2D2f10hStNe2dYtZywZmidI/ajRHatv0mZmFNZ2GU5YFrF1
fuh1Lu1cvoxiZbAVq6ZV6ZfkcDL1r3p6p9vpri+RaAoAzoPRh9nYo9B8ORMoWfsz7r4h5M/WWQlR
ajTeDZjjv3h1IEqhNn7SdaXsD7pHhBInoDwWJiBOk/6JwYCVSjf1Tt8PnyGxf/SlKcU9YCrRRCkE
ahciH9MmNa3Bx4VGIzP3tPM49eiVOqDboQDvYFJBi4+vBjxIXgrvkDN1U1bT3u5HXUeBQBQE3PCl
t+bjTJ+ZZlvd9kWwb8iSgoklofywwoSPnDdf+4+4tQe8iQz/mVGGbTu+Xe+jeXgKLQYlMqlQB0bh
xfNtvvJFMx8xMouBj0qF7oMQi6G6N29nPDD0Ed1736SPldGJi7JZGXE1UXa6rUhb8Felwv9HwLpi
LuGupdX9f1dm6i5KlKDiGxRSvf1MUDYAPbUShYPC8hQNsMSdgO9JjVWILWx5NYuc2KRk4gULBMXX
+AUjITEO8aE462DYMfZubWustxEK9gU5b8EJyeJNGGH/AhLPNVLwyFIZGrhK2UB6mlFanjvf1KdV
At1q8QQW45jEyhNIIRoFw/C4yWfehx+i2hLesKheC9HMt0DvchDJVEP16WmYMeDoHoYIVyj8Jq4C
c72DLEePU44UO8hTkLJbzhwCDo5MZzUsBbED/E4QuBkCWXwAQaBNWCLt992qGpl9Q9V7VdSnJQl2
TL6+pGvP8V0n7eQPbcBQ4VXBkrkvKeyexwBymBADkKeNSpJKAomZd3OSAekKGXfFsruImci5/3XO
EEJKpdxawmXibQE10+wd2q8/KCFIjaKPkgu+XQaoL3xLglB0dFTI8aelTfeafxpb61J38sHUhz21
4dkQIfHpmRM/sk6pDz6JxUJQQmKIr7EYDHOwBjP84OP05DSSjkl3vY/3hxqHjpM6mLAy0psJuole
Ewm2shi5T50/A2fTBaYuqLvJUkNDpUe93GJ+NUumFkJTR/WMFFtlQ6KsUz3LvLxbD5GHDKaDlFqe
VRvzxGBqjEOI/Bk4U3YrhT/DfbkY+/8H74KuAzkY/fTlfc0j9KtB3iYSTq+a47Yaq4R3ydjBvTvs
isHeB2qQv5aSligfGlE4TxR45RuQdZwbOV9Y6GY38maTAcgjtFGZOPLZvYEiqL28Za4ZKvPYclox
4M6uDykI0rpl3HUSxvf3KdKjFPLuV99Zl1dwBj/HhCSyuAum5ysJSeM/c9RfY7jncbTCOMgV0w44
kxHtsErdzuGXpCtCsCx5NqEMVq2MW11e9OcX1pEro1kwfNHk10hE7L/7uik/JoJfBqTxlVrJmZD9
95pukvPv8ZcdmzvZOgU/VKh+PO2QiVkRw8DABicWEknANl21icl8H5uTmfLtV2RjucbGtKi7ufmK
hRAB4vY6anLGl+TvqChk3kNcslC6hpzAFDkqyqBCBZ+gLnt+I9f8q5gqbDEib6o/mIVUTpZB10d3
V9RqFEiWvBiMETPcrZC4F7o9WLeVXEWfBFcT0PB1/qOQc4HwBGMAYISOAoULdmA27ZA1Qb6v7Jpt
9gFXCRo+EWzmt1YWqt2FMZwnj+j1PrcMUdiDub/YXeSW2gWlISUM08HibldxFozTmifU/HEXqbD+
XezFqRPJN8XQogUi3uFQ1XxPmYQHS8moDlvbMEXjismyZsFhJAu4IHCW70m4iY/cWzEXyxP2G5hs
5CUiX5F5wik6S2qxugrWavcUGgHb6oOCCLRF48VzunNO18nt+MPMC24+iA3+uF3JmpKvw1S1yD1Z
Om6schvefqmLLjcAIZ/bP5HLU8sySLNSWwPVMEhxPsrz25ZJrTtlam5aw+sbfd7JDVV/lRxprr2O
jlta8yELWUWcdeOWGPfLY+WWZ3uGVxTkCAyXx3nophnrHe9xkIgr8EMgDjMEBHyawUn4KkK1Cor1
mzliocexxALqngmKgVMHfmQFN+SdqX/1z9hQMJ8s/V/f+XXkkUXKCK5A2SIMrfK4JVb5oHchRTUY
lbmGUmEig8zXeXYfcvcKX6lG0Skdf4Tzrc8pzXAT4oKW+TdqWx0ZoIBPRxjPkjg4By8yAsmII+NG
4C3BtEo1v8RwzZ+LXfHWgzvhinZmox+zDQVAnOBb9qN87mev5FGQ5/7cn46e0uLyFY8LcHT2TUiV
qVtbQTgWjhNzHIbKEbDqDjhsLeNggn0h3FPKdBm14OSFKsJEa1UtKwuPY9zEtYi8c4HpNGXz0Iut
5aoT+4t0HHxJckPeB0n3VG3QDnR7ZVdhk+B92HlVIQJ7Xg+5thN/sFwXPOF6HCUNZHADRpgeVBMr
EHXV2FroBzXqobgSt9H2w4E65JliLhXYeQ5+wjCM07Dm+zC9eaWaCa+Ad93g9lPkAT5Xo6WCtbZB
rmngnnGjbbo09prrDdPFrSH7/J2G6HMNa6zpRglHV3/0uq9f2Q/YuxzH7MlTQWv2PGU0dyoiyDoR
+mVipYuC6mR4WNSxfgJDE4Z7ddZJzhfIRsdRFN+oI7cwXGTWXmH1uN8lOE45xA/eT1vnd/PVf4dE
upuaC4O/gST7KBP9RFcbevRZO7CfQI4F3OsAPbCCwerSve7jcKfaB5gU5lgvNXhfcdVsUyzRbv2o
/3A44AaD1VfwXotOTYE3f5fBtUQ5bzPhkSjiwqakn42j3x/7yZ/MAohCR99qEGCppHnsMPj1TJkG
716aqe6IltjgG+IUc7TjsG9WV4nhD0wM/HYfO2v5ZeoJlJfa18D5ABFotVfZmrg9kEGEDD3Zhp7n
L58idjseC2P2g9w2QOqPVmM7JlZ0+9U/+jiXZcU/cIzX7s1n98fkBTfnzwpXtfrJqJOtORnrmwbf
k8mo4mapiUMVkNFxHV9OEvE1Jpyq0zebnNXG56nu6bSVobGfgGaB6qG11SIVXzzNnG3O7xEecQdq
YVL2nVwPNKMJhiuj4CsQSRfdUbwEYxIAOEDrxO5OoZjVcwqE6gbI5y3AGDhCmJ/+JDHP9xc+lNo2
QyhYx+EcFc7y4/YaPEID0gWmwE5Knkkl2QlTEf16KTR0MEEV6qPYV8CR12YxHUjQE7EXoy8wTJUD
kQhSUAl5KdmTWpHbjZkYY4ypcGLyVCLmc53cC9n3o8AaEJONL27IiVv7V2azmAKQ1Nra6HGOBYts
CB10nX0MEyhsXwTtE9WlmcYeyhnqfP0bARuVO6jLa1W+f0lJgvq6Ad0M+anqbArNVTo0dRQtuNQU
DTrsEo1CEz53FXmFaaflr8EwfcZD/xvt9WrMfKf9+O4+JquuYnVUqys6qHadRK4JpNGDbLzRut4i
TNoCfEpPseTNBi2Cx4Ot92tCv297cQXiG1OWT5b3hocnGJveafOY7T2az0GSMvnRVzuz2uP39qPM
ai8/xtXq3oS519oDSHzPbIr9XTrBKR137Gw1zo218Fu54teD4JBPsVlMVE0RITTF/myakaI3KolZ
5dCfVKaTFVXI5i36Cz+zSeppfMUEeC8YQbPm9iUlP4eBGAU3SVZ+/npFAe4CCc0awRo+LIQeVqz+
FakmpGuSthzqQg1QVl/lFPw7tcOXgI7onX1OWoirT8TPKLFNjvFhI/tLhDLlQMLP6Kn+WNbE+cVL
fI41M0sOH9vKTnGIdgM6G1dSZmJEuInSfQmcujG57fVG3YQXgB9lWUMEg6OGesZVDaaX45S/uGo6
4YQbkcD7uUX2Aw1QafOPWfUDi2to6cdUlcXCSakWl7QEk0I7jwqb+FhS/OXComCgiaBq2biK5Hnb
UziBxzjdhGyxqoE20a/k1Ww85sHSL7z1rCcPRdr/vgCxz44MLcBfuO8WNXKcxf5xnJhgtCwLIl0b
cu9Mwn3iwjWxOzJS80+Jfioi5c3nAxx5QN1LirhPMwLBKJaMPfho1OAZROIewre0Z6NofXcrJyQ5
XHl/yPzFSby952dMHvsrXwNJfUltSQwqNk8fgh3sWr+LaoLPMMdNUc8LKAtkjCgu13gWZ8EVwMhq
c/LQmfPmGgZZK6IDWYdb9l2SK4jhn0Iz1ggiAgZ0DNaxfwkCPUh0vlLk6BV349XIzWfy6ZFtoVg5
F2jP7E1Ev3LwJW7Hc8vYCeqUtDui2PNVxgH1QhO/rEOOE7/DYdTypjn0fVLBwbfQkyB8R/rw/ep8
L515hA96JbCn64wANJCWPggmrrWja6ADPeffDcTOPFs7Z9eQY+GgXd3SLmxH1EhItoiJHDWD1gse
P6hBhJ3dtaRnYwXfXHnk71ykt62xYCJQrCxYa0Vnawe7M/R/gooe6eMgaA/5zS7L4NoCrvKeS070
d7Yj7HVxTcgYjFURxFrGicUExG7FSX9Nir52L0Ewta75lKZrCi/NtRRbmPC4TEL9eoctetDL+m/i
lR2X2xCevPt1KrRY/E35cRTPszQ30NiHS6uA125CQNdToj1P89dH4zaWpPuW3CRApSYlyvOkzZZh
WYT0lAgPtd8zcfrKW2KklsoR3llrqLEahvaKjVd9Q0oBlCCwx5ErrgYRRFa1ztAoVgZnWHqbytxr
QIE35TuC1KUgPXYMExlE2DaB30CCQec7O1BtUQ4AZT+90VRvLQtBC+3bFVN+WnH9r9w5jIvXsMi7
c3HuQAHYSRY3YZSANFtLalW+alNqK+KSNfM0YEkgyWKWmKcWKM2MEpA7QuCk0LdI8C1Mto8tfyFl
bmcups2ddX1i/bh3rSPjqgdkftAw8zUcvloRGxx5VdkiPJJP6zK2JM9+vc7wvbBw3/iuC1XTBHMY
dKDyODYX/uCu/TS4rPXyH5F26e8Lh+6jKILPisj8oo4cgeJufo8Z+ytXb6Dwl8ua2iXByewCfTeh
iiMZkxRzfPSJKbw0mBt6bVe4PcjKZ59+O4DbTEv1j3Nt8yFO+kB9Zxb7fxaWNhLNGU95CLiAnbaG
Qm21/VwLGM1EUFYNMyKwNwIGeRRCYM8swA7fnC8ySBWV0CQS57Gox/pufgaY7cDlajNUB9OO/G2T
uov+nruDBWL3fHgZy5soTMiG/ty5Ate6vUwbTsXYk01M6OYuXTkDElxO2atVSA5jCkMfnKKD3t29
B6EjF9elE24kkVMsXj41nzVl8Go5XwA+LX7LhHByZ8L56KetyfD5Y1FgoE6xuELC7rD8Eph6Odoj
xDSK529zcW1blJ3Q/cF7Iy9TH4ZYbFs4A7c14F4uqyz3CRhlzhKHcAMAwWesZAlqSXF5r0FdpF8c
PHJc3X+wZf6623MFNOWkVrc9Bij2ApBOC4od+7biQAHi23hw9y9dYWr0OCBlW97jhorpQpjhhfmp
2t+ybjbuvSH/FCJFL/gHfX5M0IfADMV3rewO30Z9FJI3PwHQ3Tpo7nT6aa1gmjQOLNBiXQlBzgYq
xVa2m5HansLTHH8AZ4Pu2P42kENbXdLaPfd4MOJjs6wjFuA+oS25JIUdo+AKFChiNBIs/QDEQ6XG
wtBkVlv1HA3r8pvC2pnoSdpdcnNc4icJ7g5vjINrYN3/UTn+hy6S+zQVlPW9gJOfYb7VnBr6z0H6
jOsJOs/I2+8x1G4vweh2SW7SEYJQ+XJNJbe/oLkjE0fykoqDiTcrEuAbT4DCQrGoyBbrJ6UJd6Hf
KjBtbDFjmOSSXZwlYzFcLJ1I3/RTQcIEsNELz9kdhK18oprqE+AKKLRbsNi+JlaLrjffE15d0Vfe
RzWpXahncbfRVwUOvWHNzmYiFjGlOcgGW3sGIBLrmO24+lshzMS3vKgRgvghbkVzaQ272GJWjCno
dQjLqxffT4vmhjynXXvxGEECrOONE5msUlqF14I3dI7fJ4nMPZJjWbp8F3rP2FuahFXfo4R4+hMv
TyeBtUSzWsJ727fYl6GskupZlaqnYzJE0GfOm7a0PB3I4mHYBvO1pdGSC+CFcu+vZ+wCxu33hkTX
FDVfqV45i+2YrKu7iGvZrZAGZIJxLBk9NIyaVTAxzRsm7Qh1C837bMyDsLC/h7PaI/G47j59Alh5
HrPykrECCl7Hq/mSfysJrvM79cwgaLl858BF13f6I3m33xNuJ4P6qByFzkS8ckZesqggS99vQTXg
8xgMLIAD7+nmZ1PXi1Lw/+oU7rBkJHn6QAbilGbC6vm4v27YeSV+IC270MrsyJDhTp0ykdZ/tvW6
p4iUiXfn6Me2v/+5Tj6CjQxUt28pHllNfl7RgMQuY9/2V56jAES7imkaFBlKMYl8YA3GK/GNDT2i
9zu8n4uAXzCiNg59PdPFaPXMvfuMhJ0Izg7yovXoewqcBEIS+0WeJ6YK2AvVQlMGXJTMjPKQx934
m9JqtgGdkm2M0ohmYMRXTjn/CenN8C1bSLdFMU3cOG6Jfryt0+7SEYsBXCZ9gJa8aGbNArevAYhS
jEUHXrma6INyv9xW+P375XSa6YAIh72HpmBtRnJH9beh9AgIZzaqQ3pQxHPbeIXvg26pEIdcee3g
iQVB7YQnOH+LKTdCVBijFmSOzCvXG0LWb46YN4EYssdl/CyTMnwmXl32OtCmttoMxjrt8f+DW8sO
QaPo7QJp4KuHHZVKLoeKfrthhxAAWGef4yl7OJgNTtLGM3hFj9R1+SWW6vVPty0syrzt6hgacxTZ
lrDQdxVrhIeFuFKCv3ilLrJSfmcsnxDurvu8Gywd3Mwjnm6NfvyB53HqQrPqGEGhsSeb0Nge7Pwh
uRSYKUQpBJLJTg1IRkEgnsNZz7/COLqGJjYiwCYLFaqXzhNfro7XEoO13iTMnNEdZPCbe50K0UCI
AWO5GAn5qRnikGcA+Ox4xEKzA05YtEFrCMGovRCXwFQO2RiNs2O31+qP6/8UkRrDI5BmTTBMd8IA
9Fsi1ODZ39Z6DrzCWZUn2UUUdupubE/nnYE+6QhfIBwfXR2cnl15SL/qC63+bdDpAQ1f7w4WZzoT
5BZO5ctT3yGBKNXCZkYXc/U0KBvYVoWmJGDeS+AvvR4n3D1n5PQ2X4npa60tgefwEFuehleIMHVG
+e9YhlWuboxtLB3wKgkr/XdWs/11rzDmc/PiCwWB/YeiqdE4EQbIivn+b6g0YTpeF/KPptTbAEX5
ED7H+2X2h4+iqapz1K7b15ytQg06nVx44L7dC57CvYpRvU8j0D9igDnbKswy80gIbYCbtsp3y1nK
NvcG9pM+EB6uJqMs8B332y9vuOyfpoTRhofFqYlYVx1zVi3KutFV1Nq8Yah6wR+M2ZuZtGiuWH04
e1DAIpwfQVWHkvRBo3BlxOBG1d3HcMcuf4jUvB5Oys2E93rZulkCdQmnx9JVYlj7AM/A8GmcZKl7
MPerEBaRo5DR9oA1EbyuFNmry8HCZTnfhzAQJB8pjId3z674J8NSVTlKclbeiukjJKbFb48Q5lCS
FTL5QmTlgxkmLu3Flf87iX1zScE76gu+FHm0ZEkxB7k2iX9f1jFro4zMjUb597qRyDyYCErCTVBH
ICTB6lx3S8T7HSf/8jlKeJlExz3yTKLS5LazIbDZ8pIo0HxQ5VTZbWZuw7qN4f/SgpGGszfTVtOk
6llCifWdsogyjvrq9F1ehCXIHIVETz6fDFQoARl2lRjhp8qmCFCaxslY+8hIf8WvbK4vwv3Jq5Lx
3NnTkDHozq7a5E7RC2/0SRqZGUQ7gLUaI6d4vFj164ztSZNwSFcOCaWReu8mMZrweN2fHN3NMkcb
XxfBZO32qUoNqS2yevC8veF2/AoUT1hP6i0cn3uEpQQiX5DCwJFvt/tH2Zh4TRii8ISRmOMnfFHb
7pMAIh67oaMXXOb1pvW1aUK+9VE/S7w8juaH/2Lm34OZwov9vFKjWlRJG/TaSAlYe3oXsxOX/7KN
Zot88n9vbgTStKjiOIHEUNdW2evAntqe4qbXvFRe70fH8a2SDgVakb7wOIeZVNLtafpHVudOl2Z7
U8mBCsI2CEK20gJ5aEZUfh0VIbATeZK9+BEd4yzmmdvLcV54krRJxiiq7aUADeHa++bR8dx1M2Z3
/FEtaoBVkv7/2u7phg3sjJwkqFSRPq1eqE/K32HgjEHE+fRG5j2d9+Nc3cm7O/WVQlDK1lRW3rn5
+x9uJPrPmBqWD8GM2++3yCKHY+T3jSWVywS8RyIr0cKgI/MGeFRu3AF/U9wXDx0tVympCidifwna
Phg15GV7Yzik/qs5+P6JGOwcoi0YkeEHs2cADCf0252c2SQHcSmAlgrB2kQDkU1tFGRMFDHTBn6v
ipiwrJkmRjyq+Jh/jChu9bJS4+nuxoGbt7nK6+3le+u7cpTrWQC9Jm3aQE3TyGP0rJUz8t+SzK5j
boW26lYHBIBzlcqsBg5xqPjZharOvZ7kJC6qLwjGDuuuB9O1LZWrlDqHiE6A+xhJ6nQ+AyluUgMV
/0cbB6QHT4cMc7HfnTbTWl0Oh4cIKTmePuQFQ5FZq2BKYfBKJPfKm8H9P3CpLKQYLDm1+ET8rchQ
y9bHgZH1KYaphwrat40lc/t7o0RSnwhxbBczvXRmIZvkReNIXsVTusRaJkczRYGKY4XPZaKfokHC
02Dc8faDFKKI572n4Mio95vfBAz0zUj+yBVFC+ojjd+OjQ2K5UYUcpzEvYwvhEYdW8A6CkSeqYxO
eyp4mmwZnwK6NhkYLibYf90gb/tcoQTwQyS5IKoyiEqprEtStcnBaKMI+Q76Xk5EACHtsf4rRmtj
a52PsGgpuct7frpQsBoMbwWZuf8KRKcO9vsPH6ftPYxVgQ/aAtJWhF36n+lIbrJtO5sDneJXfqV6
CpDzfohOruyd8j9Ox+AxFaiM8eq8gULG/TKqUmMf4kKIpF2od7BZT6eMc1Tq7iBO769Uqadi4B1i
IcRXLHKeuqUKhWJNN0xUjgAp+JZwmngmLh4snwl+ZdqOMieLuvoC43p+fmdkOzq1D7ggsabs2zhj
iMi8b1KsKoHKZ5trEK8wxId90KfGPuDH/TE4l2+qBFe/OlONOIIWuGuAHN3W6Fo/zFwkhMrSiXO1
LOcpIroI6lxm/5yPN3ZH2mau+4fKn8qx1Xiu8FkvUQLaYmJG2x8p2scbx+hwKmVY1VuUSvKCefjn
1IKZU1zV64EjzbftArFoW+aN4bt4Y+a0ZCfONxem5abi6RVv4TwJYAtlHHvljg3/nz6yOvKv50Ru
ZOz5M+Je6gUkHZ9Y2avltJdUAXPU79t0SDyQUSGF9EyKWuEHoJSjqHOZoXsx89uYM+jtOOvdp8Rj
jZAr7cAuHYoqVModCLvkXpnH5JnmH8zrwlSGsxwNDdfU4Xg2T+hYPdbFR0W4XhYe+wp6CYo8wqW6
dRhPaMLaA8lqpfG1MQpqRwrr8JaSRUvANlu97dXxsS28qXLy8F1/WLx4U/Id55pCO2ABhFeuT1uT
WhUUF0wYVK5hhdff6KxYQN9ATUYr/msDGq5a9enAd4xDjKUZieHPQssGz3ttRqGaunff/7AbeuDl
zGZniaZoknHgyYlu1YGY6R1cUN7Zf8xAK/sOFVkAWCinbnVyIPrDTQiTLjSBCVQF6ZbsAiM91DNX
Q6T6+o5KodzMspCgwK+k8jNBFiFZLqkCJQLBrxIOP0jkPKeElNjMwHVK8iNlKvIS0jh5I6UApkh4
8hn4faEeuUbDhbW+l9HQlPX8OHe6pZUIkZeisFKOZZl0YkcR1msVIVrTxq+nSsBC2iXhuBvUwkMB
sJaBIuleGwh246VsMEtXdZXo+GWzxvy+mU28bIDpZKIn37dis9iUfQk+xZjR9l14ZJUByJo3MqC+
uRVYuRu0WoLYbkSaLJ+H4gwFETl+QZD4chG5Pm8S/u9Xg7gUMrmKX1GPwwfiEuWOu5D6j0OvQD6Z
6+6Jrsp0xWSsMSpOJZwI9vr7WjtJuTmt3b1eJOv9HGoAKfiTVFpet4uylp4XVTWKjs3foMvmhBpS
gwRVzKsMGNmL7uU1YEzcuW+gSZaT49G0MIalfaZ3BQFeZ9KjsBZXOBt+Ithg5be9RUVfMb14tEoa
W4u1tbkMvdV6nYuPiTFOeXSfSg08zvlPBxb2ViN8swWeCxeO5Oa7uliddJisbDlRqu+hsUrOG21A
Yw9WauAaUr+KIgp3Xd3bQzeycS75rFSiwlIUBmP0InOLWLYCfYiozge6XJKoR1q6Rvo+nnFzQDEP
po90t6VvoTAV37f93C+FBHW3N03ZiksUA5n6e8a1xCdL5trmaEMk8JlhsuBuAy2mhz45YmZkU5l4
aZDqnQKpu1X1qRfg9Jj0eFrRXH3Xq+fsnk3MyB5aY0coI6OJWIGI6DHvVHbynHYrRr+6AAOSwK3L
Jmcg0Pmoc6TSZjHB2MogJrLKus8id2KOYWaKysxssTcK2xNGnqQcPuLRanTIqATOJpKv2NkbRW9f
n7pOXr6p5DdjVlbR7wm/SUNZQqJQR77b/5Cvf0g7NaZ/jCYPaP9wV+gN+ayOSQIFYGh/xZ8NJqqK
KD9/GIXguPijjjYasWR8hCxun7shaIDz6+CtP9NVj4qizI58BY49GgkPGkHdNcIt4MmXEtk8SSjC
lSjzR/SRuqoRF+heBVp/ZrHZlN/LKpPTi4lz6odKBXUTzXElVHR06EWqYB3RF0Zd1Ev087ivvHGs
6QriA72P/ZRBtHvjSRdIjqN0kwcLxutIuE06pmUVFvNdzJY2bLlNLF5u0W8zvky/xDw8eYa2LhB3
5aN3DZXKDMf11AQ1Uc/XaBYCJiB0vJOxcnzPdBC3Y+PDRHFD7JKwbZ4G78Naud9TgNG3hspxSsr7
TtiVAWC1qYbSgn6sV+t5qQ707YLXNwhfNIy0PRULWiKbsYEViKUpQD5qhQHuFACqHfCVb7WJP3hL
5nPSNvtw5FLW2k1zjlZl/OsQ6NpEVHx7jZguRigO1DWP9o5O/tQUesI5HBUF/aQp5g5y/KiZDYyo
vJ2PZuJxTILnMCdv1nx7Lrq/1Hk0guMEn1Hq8Nf73WoPWnMZhaanCg2WBSlWvx7h+kgH5PrWp1eA
iK76EYrHFHyGM38xOxwCUiyKpBnypeaHtdWycfR27BLaIg8p4CzPMblFYHNnqUpd79/UUjSpHMMZ
CNW8qFtLvwSbGw8plTcTuxJwhGVvQWuv5VT9B9iufLYs25u5M5XKbt8ed32ZjeUo1/rc2gi8Bluk
TgIxrBJYkfkJd4ZJppg+UUZnHJqOIueBvNyoPvsdn6m+9eF3mSZmdKuQn8XZ8P4NF2J08Y5uN827
0e9kN8CLfcKkVGjoS86m+Rgq8uY5E6blO6bsfg4yQqpuP1mT+aBNYsAIUg17cZ0YMqioVhVYHU0N
B/UdUtHMoZbD0+6v3SIDd1v9RuaXbMFOGkhIKZtxmWa8e4JApCnO9oxqDCo9ICRW8L2yperCt/1g
JmXqUFZJ1zNQAEiXvjVau47KOzgKl3GNCXpC9cUhRFOhnyt6yaFIIdVdutOo849jFIsqVENQc66g
m24y0pr3o54/s3+ZXFf2lQsPwDnhQubq+vn+UnBCd6JxUbSQ05to7v9s8jclS9613b3DC3yoUiyC
9LZffAdfSHTpZnExi11YHh3nAzEkT+tXvCXwvbzpM45lHa4AlENM3YiEzK6TsyMo5kaHdHmXlMMF
fzQwVDwwnm6fP2JHTxDOOA9fX7s3huCOCiKFczbUV3E0ZvAq6WKszLcdwj55+boo3mX239rZcWRn
9dEvGK57VAYTbKs0EOFD7vpvWh2OB04AIwwjIjlxpcINmGqLOgDdfB2bCB0ZjNMuiGo24wft7ogE
kkepKuXhAlFj4sXN8tn5cbu29XdmVtwo2P8k6Db3qiXarnCM2ZwQ0KqrxwPAZuiEwVioKXfm15we
mUlELPya5LL8oX3f9SQKPc9rUfddoOanhI7iSJZMpb78OAeVs6YHOYoaCrCu4wgrcBYL59dy6Tso
evfyh2Axa6eysKm5OM+q43Z0QAq+jkaY3qBEZVhBG2F9ip8NapnLVd6YXLYJqEGT6mnZZlsdHkNA
DbqIAnv8Xn8EyLjLkkGoPNGnCqNA4GiOu5oZu9J7XFJVVVRSzSPSlAR85u0PRX0SWNOwlo61HYy8
XeDUEniDpKQdSgBX9weklUSSVqIvWFwfABvMLIkwPwNkTwOuZMmo15WCCXUO4SlLzSsvqXkb+JrK
6Avu2LUsV1gkIo9JyQZX6xVDNPTwZj6CFiGo4A+rdFMmJRRSB+LzkixDBEOkdXHDlQ3lDpjPpvXM
b+U21+PiZqTaJUX0Aqtg+oDPi9CSPTnRB+f9vtpRv4Me1qsyB66ZUAPiJWQe/fbzkWNeo3gsWcUB
u8IDBXCTU4x6O3L8fGqp74nZhzuJLARaK0KEFK/dnQueBrqinEbzBctRwdcEUaIEVXa0tFZloaOK
atmk9BeB4i+MBSstWNdC9Do3y88NzsM1WKWz/ojsus0nyQ/CvEC8DprvBgWGkfpeOsXstwXrL1RF
V1qM8Fvv7C37h5+If87DhvK1Z9XqqdfKa645v93tZYFzY04bFMFBZvJfnbXQsqrE8P0/L66VKzAQ
BJKk0ChghdCT1iPUAOX7lXg38WCMKZ3SeIlr19ML73Q+xe8VSJ/nIPOkSj8PZ1Dn3B1Cp6DxIDtr
1G94WJPIgJbQRrGuSWv0EcazO6L2ESgPH17TwO9gpOboda0jK39rHom130EJ07Eci7EQvOtWu+8E
Vd5YQ40VgXKVFVkvt1SMTog0Nb9FJ8SAUhLV+SraZ6S358Bxn6RsqKwC1rRwnkpGNFIotZBuUZ8Y
bGQAe6X3wq7oAXwUS/qZTxwcCrOKdw253qW77VxBSTM4ymt+NRgQiVqqv/UMaI4BgVhA1GrE+WGT
b8QpqkyLz+PI8h6atEidPQwThwofg6vbHStgN/G0oCh96gxiSzRjT/xwUd5NRrS3D1IyDZ1YWgQc
imY/F5JYBdKvSGloepEdhJyqY/YYIZ8oFhnjkr5m7UkDnG0PMIbl9eNhNejfNKwcjDJqmHPwmMck
lXJOTxtk15NvszLyJcF9anezy9LTuSE8LVntRAPgRE7iK5348PdQO7UBongtNpoFqfVD8aF5b8dX
0Yfteux0NiAckdChegk5rxc52xxWJtOKRTMpBvNRHwCfGSPZWdf50q+JeH7icTTl1d8cO5fTMi8q
DFKA9BrBqhFfk7neISO+SyhiZDVShnDK6uG/Ijqz4Ty9PBIMTFXsn+SDXWB0T724sl3UE+dpj/XM
5QuNGzlkqEWqtEsY3MIvQ/IHM+H9PI9ueTwq5j8/pvxBt9UMRXbdG7ZONHiBfszT6TAEoHa/IEh2
+JgIVfliCIgqG8A8G6DYpHqc3OCGWWHcTU9HFV7c5HoZmAKEyLXJrgOTKZ/7yrBvTyonEUTWZ8m7
BadiF4Ttnq84pwuSgJIbol/ehOSKI4Ld3deDMXZJddfplklGacY/oQsjFkeVP108gFSTct9gTuVH
bWNmploB5Fy0gt0xMn1Hqv4VF49GVVvaWle0N9s/sH8qEq7Y+alQR62z+HWRfvlAHGRhjJRFBp4I
5IwQ3ADiI26GP+t6iZqZQNKHYPJcklv3TL9jdzr/sqtVNLVOCbtIXpSAY1j2ZzuTGglL3ab1oQYS
QLGbH6Dyc7KNkrphAXUGNLczwAIy/Gko0sB52mGCRsYZhr/tPL9Wv8rGXBZmOrie8Zw1KVrF5jMA
szMBDIA89dGKj8pa7reGlUnw94SdvVYSFxLTsPraGZqj35sWD4c7dDhJ6nHochObkFxpT9ZY5s2k
g3enJr9fYUq8AuGXwoAX3EDu7NSGn87BPFeE7n1Jv1woF5vyQ2ArDhRb0DXg7+FSYhZHrje+Jcms
Raz7TQcvmB8lM0Wg2c1/5otxLlUAKVIzSWne+hi1ykGozPfOWbUa1rxPoIB3XAtPDrdQqk6HEpgn
WuHZrVD8BEnGPWawUwOWxpcyzZuuyE6NZsMIt1hjtJnXYGAIa3viXx8McHCOky+ovnNAH5L0Vmy2
uW72Bu0lLGpIt5qF07jMZbnXwN6WhSbnxvr+xSCAW3Paw5f8e4XwRl40sBpoGRNenf7ozywL9DDs
6g4AAjEhhHEnYIhzOVH1soYkY8hXDvMS9aXahpT3XK2y0/pPQoWZ5XcMsnqOJTN90r78imxlRvOd
i3H5YMyw0CRuqfKMi52xWgS0x2xqCrTQVDXucwSh/pAYWtbAJ/6iueJHP5EbIibedCGUcGIpGrg4
jDqb70s/DfBHfQI9sWfQHEeHAi5JBTTyT53u9r7o1smnfAzERBWofzKenmaHcAZjUSNOk5UV11Rx
s6O/eT4byk3IlFyvPvnfILqgaJbY/xEvkEwZc3L/ecAwnmUlK0tEHiuN93x/8EpWBN7ttLOBie0K
Prfj6nffxPTpQQCbNS1zw54nu9sMJiURtTIlgW1rON1HfgTYxDoWOPgLpov8z6H2NuaMZ9VxTGGD
rWLJY2tAYM5UY9uRqkXQYfxGllSeeovXt2/pO+P8NtWAEzL1SHhnovZI6sefh/tqwfe/A4OGv79o
bzOCRC0FBBMrrDj0wAYtYGTQt8MCc/KWUHRiZ6xqVy8e78jVMNmm1FrB93mhY34WbPrUIBLrLxnM
R0Rs0ervJpbyyP9U9Z1lhTJdznl8sHtt3Rx+eDgvL036YK7FxTZ20991gMRYfMRfxlBZL5OhExvB
A+YoTIw5de0QB3plj+Rnl/PCy5DOjCjn0/m5IggyMdS4r+vutfo+vfrNf8yEFrEJsERswPOmqUID
43bGZ5RM2KjuKm84kZGHSZ5n//ohfiI01Io6snqObZUWsGR40Cn1Kl76jWj2SL7N+ApZrYKkK0yJ
6B1vUB+YblMTc3fuo513PaT25cD6Q1GBmcFgzThsQFZWL83lUVUXoAWokTzyds+cA7GD9HXgv1/1
u2fQbZz3JuZNSlaOBir7lYdes9uiMdGIoUA2G+vlBk3jg6kDsmQn+r+kjG3eqkCOdQFjEzG+8WVw
Ov/anqKV2NvUZqRxoMt0yRFHehKPDeJlfgMMEzhCyu3FJQnIOKR8cfHJSS9qV2wD9vGmwEbt3FRL
71jnWffnprToTmwBowRMNfr2C4TvTtfcgwhDHC+Da18DKEpNPqwGW8SYvz0fggyiZweJyLvQPsE/
mWq0HNW3dQk3sfQX8Y/n2nwEg6MgB4N9IbT5XFYy6MdODOJpLyLCDFKl0Ute89lbz467PgkwbPiO
lJbBj4FDaqhhQHTwfI0MsxAqvvyy+ve2Mw0NarThIPTwkHk4h1Al30EEPFq8YoznCcdzCg3l4m/h
F+Y6KmmZBUt4n2670mJLWB4dHFC7vhyMGNrmEHNY0OGMfJGP5uNbNmtWJSVi9vH0wBHNYfWNr84J
Jdzz3jrQrJv/cDNxIASAeRgSG/spsJtb3oxi2hm35X9yGIEoUSDfS8W5UMB3OClOVTileDwvrH88
Q0hgpMa/RHGGHQlDMGoj+VEefDahircXXfG+KtlxhVRzeHMZo1iqQkErFVL+FG4oA15yeUdh8Sr4
IgwD8A0r2TCjzlj3SoU73D76opRMJSOmIS9FYw7HSmsgKbknEej4PvEaAwNHRy7PBBzHmwATO/od
q0SW+lL3r4nwEeNhHq218F4RG/Gulk5WVR2JZQ1Qc1F8zBc9dHsWK1jpK717K/DKj67VrMGzbTbg
XgMFIYUbBfDLT5esDP/W1Iaqk1YL9qO/Wr5x6JXvSTq8AbgxupAfxKK63/73szr+OJ33rQjWzdWZ
xg00P2E3cbMZrmJ+P9YBQgzSN9f6DZ9qi5gIGm3Yqc5NHGL5HqoBDe7jrtPGr32ueuAF1S1Qii0p
XLr5f9I4qmTo/sDI5cnTENzkpOSV/1p2HE8wc+1p6b538P577pITvlVxaSjwtROy7dAkBoVuYtTg
oI1mnQQ4qI1ggCJFbUdV5RFN24HmhyMIiwICORc8XSxiQLWWqYVKIonCNp0ew4Y895NMOmauzqqY
03EYshKBRW9pOoANaXWopnk/ukHV1XbrPGumBNwQhiJwQ4I2c6QG/6gXmFKz8yPG3MEBXPXjZ7IB
vhcfKAL85bojxZEfQimDlNQ+HCslVO43vBgVZt9eXMbHAcAHuPEJyFyCHlv6xm+mPhpCd6PclIOi
OkV2A7cUweIW7C0QoswiRsc2iR4QYfNxs1S1131C3sil7jGOF4Qg03N4AqxOd9vtb9Si8yPm5zDS
qeVymW0SbuqsRrrAPxcVvlm0OSujVJDc5v8Mjdn3byc+Kxiz5EZYY4L2AQRrHECmsEsSdJXIRkTS
j0NLPY6N/ZgfLrtdoLpGdpBmA4l8G36wZWRsrnrzh3UW0joplpH13M72YGqhwGKCGEl2V2gGpNAE
pUD4EFTnWN+DvQnhE8ANoSGXQe4Y/1BWj5CpR0SB9FuN8RH0JE1qWphR3V+LgNamtv65mxjm4yfH
2zzCDVQ0fkM7z4zO2XCb1RQ03ImMGR7U30kVYQWpu3g0BjqoqiAoqXkU354HrvrFqMc2ev8RKcDk
nZb6eiU0395akpJZ71hgVRjOqtrjf9A72WA7M/N9l4HQteeeI+0Jv6vDkOWYxZugqmynVIYnno7g
MzBbkEPzlAZNMxDOndi8a/SKMilV3lJkepvU/vTY15oRgmDt5r9UZlsN6o69ri2R2PUaM7D10AWz
vs7Q/803BAgpUpUXboZmEc198eRU711tkqYbe3AiRrE2F4zTFkq3kQr7Uozhn1P8MHekUnDpcpE1
Z9wNU6RXv79lwcFNYp/qLPpd28e85uxx5XJfyqhag9kvFURd+IhVpw988hxl/31i8HTgxxn92no+
bJfIb4Jptqyeuo6nJSovI44WFUr7qZ+wJQ7W8myw0GHbr7DG/5OponnorDl7nwVmtMQZwGldHoCc
dn/W8FNvl/2r2R7H9bf1j7QaeXYXucdXXBLVhwHkeczt5dLTeTzfcG7fMGMwPburhsNc4WfGDyPw
fd6jC4XmD6esWWVEN72FcSp0eRtbFkvf9PhIrGFdrO3gEzc0ssXP0ZPt4WF+eeW2BUMaITpGSs5E
oTW6R8NLBxLe0dXMVS4uPTfCtKBMnAeskfdXHbi8xMSe7F6vK683jc3uJv1IGyt/RePRP2tKZqbF
j/V+iOZGaDKM2nSmOAa/lDzIs60ISvNjRvKDCM+1oU4NGfMOjjIMD2/lMXXRkCbTH/00LuPS3iBd
+8HoWeU9oAP6c7exZt/bwV0QVBNLDn6qBsmwgTR/See/NV178kRCPjIOTgYbo6aLC0FOSCSYmLU4
jBWqqL3mrBzD9Aoknid4//2cSfsuPtGwp7HyJYUtR2MCmDFnp2/wvq6I2Nyo5YfVMYVPVjkpJNEo
BC1a/luDO/cjrcQINvXJ9F3+f5JIRABLssQJskLuI/Oi4c7z2qrpBvAuhqk84FVp6CV+cAOXY6js
hVdIN4X/TeTTrzX4zAV2uDN9rnCBY59QaxSksTLiA8mNS+yCo8zbhKUZCM0sF48hFdhBDFAnmpz1
uRpQlTiH6g4nVMAM5OCoGv1QpUyMK0zjgmUNntHlAQkq8sLWzA62XOCx1PccgQb8QyJc+0XlXCS0
RjWCK+OulVQ77vRLJ1kxWybpQBB12kXJeK0aNc0qkb69PxAFREPl4IJ18ia1JA7D7WROxrR1vlqQ
DX3onU3UBg+k8LqPQps7Wf06+1MiNKpslFE4j0baHe9zAejCMTO8yjEyadRPBnCVoJUyy2/ypEPp
tKL9O0nXYPjzIr4pXLE3MqeauV5yPua1IE/HOKDEnZl/M7Rs9jM2eRnLePRsSsa1lRpMeFHQB3rD
mUNN9WsDa8bVvGsj86PdjOLD4qslQgc7KMKVz1eGdtMiDUOKu66ie4GGBE972NeTVO8iOT3Lj1jv
kU/yAz+U83t+uDgGs5YvJJdFajNmRiRlwNmiq71sB7at7qL4zW01ClrQUyDqffieNdSXhTVOffUh
3rXzCyCc1IrGaJ1XcFsENYczT9qnexyGgb2rNwswytTipRoBEBKiwuHAxmo3PHGZzgIi+pyNG+0d
ag3Ijd1s2yIsPiVI6W0B/8kHub85F1O5g7Kl93xEwhgmh3cvqSfSgTZ6UxvCkoI9N+h2otUGuBl/
AkeQvG4g+2purrze9zdSYoQL5JEUF7hNqgC76cFxrKaHnI1a5hTsjgL278g3yklL8ktTWe3TC8NJ
hAqef+gK4KF5i/qIj9sTICkIph+XIu46vpDL71XDz3KaOEH9bXwT98dQAdQvBlYjl9QH/hodaOHh
iWTZbyyof1KeGgMm5copNKwLQLsDvzdalLvFCu8rW+FA0GDqZN89LeuOslmbuuRhUYikyP7mCoKw
e0dLAASOACVy2o5KCGmj0K8HGQxxcyin60QA2WLGxfELGWWqKNdsuxQwMrKADzJ687wbGKO7AD7/
Mw48l6tys80szcsuw/k+B4LcnaZjgthg1Z6usIK9fayPT33EGQ7F4neEo1feHz9qROyEr/JkPgda
mWgnyR33WRHpn+BC+HS/s2xXKJ9cQ3ZQF/4gHy7TLMyGfuUkl8aVPTYK6i/Mg4D7gyt3MPqDIWoR
eRRU/4W05X78sKZV5Kn6TGVQg6yEnS/Agh08BH2M+Dt2l1syk25u+pKKMDi4vS24qofFgiCfXAHD
RN2hG20ML5Iee/M9daazD0gchdKq8+hdVXxrW4gx83MINKWzAPuZlZrTMwze//L8sXMTORibGYeo
FghHb8acq5+/fhdDunQ0qRUd8A8D/rH9ZIprEjY6mLyovuAFO7AQ28fOwaIJwYpeifK9oTzPauOw
JpNU5jIva+LLaqZqzAy85DMvRuqeIbVZwII2KyVSV53fAYjapuZqjkrLfV9GXqdF7huayvqI5fHd
CCPTdDcONl4JbRzT5T5l2ZSTurITwPKHBEVcQ9BiOaXyL7nZy8/OIG86Gbr7v+eVkcpb0hkUIhFX
f0FZ8VvipiW12iMh2HzarEXr702aGGP+0Ip8vpVLqNd5m8b0lR2WNRIgp2s479DCmSbvl/54aQoc
SKr+4BVX3iVdkLu6W9SVcGL62ZtvBubAeK0bdpwDdALX3+vEqsQ8xqXgdxI8wqXFIfn/8hgV2FI5
WAQRtDorCWmmS8sY9+JgLtWQ4M3dAKmGDBtk+6WqnZfbiDAv8NzGrGTSEhtr0t53phQVNajC8DzM
bxk8SazziEMTMe0xvcDXhaS5B7uZw2+NIaBdUQfaMKTBlHHhoPbVmtBH+NETjY8NAjzgrEauu/Fm
+2oa/YwDnCsMWXkYxzmJCDmDR8g/n5wwvuvWL2zB0rlTkPM5I5sKtJmrd8B1TpxMtH06i1YzjVvz
J0DV9vyFqL2Y9+wDXEKPwTV3tkJ4BMucFh+Ltqk0OZg4FWlT7MoEnFLULdadofBv0+xaGBWK04mQ
fCCAqfegTuLQAReXeSqBDRIb8+lLD6WItmZMqBlujmvY7C5s88E5kXdCtCORO77Qo2F0pFquZJfD
7QBTViOgbxNdqr89bhQ43SIzOp5Rn7GnwdkbUBU28m0FVXDX2LfbABOOR7MbyHw7nvDsj8g1+quz
3DIpwpoC259YAArI47KONNZ+ZOOGR1FPGrjO9C3e4HJCwqnIcVYGaafYCdUHRWok0NP53XWpVh/u
ouga8TQDCgYZq6cZWBP2WUTsWYeRBkhYFPmsr1TDhHrVeyfIfp0W2T5rq21LYvKYV0lkPnIEm0xm
nJIWNGO+TyWVDkMU3AGERQdgIhYcYk3Ji7ucoqWzkjVAdV7k4Cmfp3AsYonWSDLKoWdVMOdH5tr7
YzY29CX4Wc/u2ZMgm4vMw6Bb8CY1nOa/VcIapU+aBXawbvoYSIH+mMbkRzGq1eE4+9aAUxN9ZFTl
D5LgXWRO8MOXxbzKVSm4+fE7l7gnmI0qkNmxNnk1X/hozvBSN5vwiyzc1qiHUH+7ZnkWaU/Gw9go
SsF7gLy3qplmwFtDeA4g++z7YOaL+FJrfOq0j9gsiHpf3lOAmgack+r8PB8DDWZeCsiJg43tvPa+
wpiDbV71e04qNmlkIX//25lysBGyGl4+3M1mmCuXV4TZ30PnGtmWi+4qi5qvYoyP8Xmb9QGl8/V9
rl4JeP3j6b7Z/uV9KlFmlf77/+7kU+JxnDeEviiFiTugaGtkRU9fO9a1vWp8E1VK41lkUfr7VH/Y
6JSGnG/bgmzcQBDZ03HNZlSruSzwUSJ6z29U7WvrcKtSY1y8cBo4vFLx1dJznUAzj0AhBX0lTsYv
/WJDN/4b6yx29E/jsf1Zjf8uE8tMKO0A52vAu2rjQbj3lHPO0ggFeIZu9Ki407ucyM5al7Y2/kIz
jfiEaBxOgcjZcu+m5FPrVr/zG7USTPicl/4f6T1aUgQgr9RPeEiZMiXpsvlY6n02jgButaYa/gzQ
NTKrVUgJPzEOuYWhwCn9WQNdIXIoBM4Jci/Rx9K7rF5M96CeXhdggoU96eRCn9rq8R5ak75P9mii
x38DK4fFI0ASNkIpSo0xJ9dnCwjJdKpuCjH2pDT4ubIbYpU3uCZNn1Hnd3wMRAUvjcxeYN6OifFp
Aj1D1l9olFfHK3bvTOBP00NsWTOzjVPehDcxBSVrZeEuigDOGvd4QihXuH7H7TdFvnDJ5uF9TeBs
2CKO3bVHhi9wSaKytvihf/LrlrcusEICy9NTcGvwfNkyy4aLzcHFSuvBAIjVF+xndmnTEzHQY2Jd
f5TWkYeJkAMdGukEZpPMr+mfhHZcEozqb+yLGHFZ9lL/cVb+wY993yrtWErkPTbtHjerTYlKH6zM
9SdPU7xm57U4gWIbK8CEkY8sWPiYw/3s/Nn4mrWz01WuztnNr5qtua9p7kvO5XrzuGw8CYQ5go4F
R3o1JiAZWLuDqfaupGj2Z3xx7ZFvSl672W+da5Qjh3nsDyhzCzlO6hx5XGZuhVT5WyojcwC0aZds
JzxD/961iZXtdFQuHtIvFGavTV7GVt/AqtTv5X1lZawvYkor4DlCR9qIbFp1Gf43OXqrIB2nmUFw
YoB4+rQ+u97OkmBWIKFWY3kcDnaYkhRv+D8OXCc3Zn25oogjCGHzU+p04AbLQodit/Or7TdUf/oO
Hb/7e4erOksPl7Q79vI8cs9T10vq2lzP5cyrwx8nuG0Z/FMTxsJXqQ35aC4GRv2THaQdlTQ5EGYi
lkmXDU13Q4q46qKvP9hDEVUXMzBu+33s8ibcJ3g4YdUnmo1DzpnBf9X0rAsGwIHXNnOzO/Wxt+yV
rO6E1xUuIvppoBy6y5KHOZYRy22nfUpbwEstKGyHjjU31TE+n2ynMhYuzdiJIIxGJeNBAPOvZOHa
0nuhly8CuePXFcyLYSqAe5jq3mdTpeXfv2FzexGP8ZBPp3HyKj1ZEEJ1Nl8Vj7iovJpdHgSxwacW
RC9G5pB1Pt1ZJvU4V6z1UQorA6bBL/8a1KIGUKt2fbfeeZnZLJi8vOu5o7skPQ8RgN+aSnRZCXjM
XSaBy1mVO0hR5JdqlNjmURTrFyZ6/u2lwelpdsycBLctgiDQNJ5Jy5iaCRKyddS68m5qUwS9RUva
qcDahCICCHFThZJ0qoe+balf1wClI+e8whhfDX052zkHe1abL5sBHufIiu1iAdWKRyTd00aQTgXn
1LOcoliRFXU0Rz73a0Pl2AOvdlTY/0PK66zPWD5AsB/fyezv8HVOnO/6P+ccNdc9zOs5cUSpXUNl
KqxFl53g8EHUQklo8Zl48hkqKAbAcvud4y/9BvlYUlk/LKDb1pXWz8ytb2Dh/laajRll/EqYSlbM
M3CAyCcr4ljJQYRr/DmRbxvGcOgkKL1s4AmHuVSiHS9vZnseGWAEbj/OPTNnDwtvMetSKVzJ5foQ
fTbcR40q4sVaQh+PQIOyf4qLWl/mIqjD3HGocPoVqg9A6AuUotbpapDMy5elOOeFd9Ba7SiMIz50
fR5lPE6eg3tCKc5NC7K53qsqeqcym/AP2nqbXpLXEM5B4UU/944tJYF7p8V3rL0PAQz92BHASPrT
BkoDfpER0xfeEQSbujqRf1tUhLe+ZUdofocTHD33+F0ebsT4JqmtMuqR2OaP9LWE0gFV0LxjeVlP
GGUQni4BF4gJeRlkZ8SSPEma8ViI280JMYu/8Ju4SisTLsbAtoMIqbs+7WTOXUfEPI9OHVeiJ72d
PyzVRZbodXVqfmv8KXHCI9kZYeu9CP9GRF2NyKmicpQGsruASREg0SObdozB6rJ4vSawBoGx2xYO
kMr7ziIZQCtu11A/cTydGht/53r3TXFcYZUN4cDWR3jH/0C3Rw8BkYGJn4ZzVATzs24NrRBo7iO4
ZDWEKuuzzMk2AQBcR8/OQocbeQvaDnZ0fhIy5Sc0xOTtgPhEXOk42vAGkrhMBiXR/zfbFvJgAUAs
t69Ric054+EVCacvHfYZKxB5EybLnIj3KlQdPpCmL97uYuYkj79G+mq2JxFoUwUeiXqqtuCWeV8Z
R/K7IshX2HhCQvDj6riGiALah839VZpYLp8R0HtMTqDILH4fFB1x83Nc93XgJ5dgMBUgMdRlWdmT
Isq2yjmw+F8ToIsLY+1wEUngc7imXJW9ZR/1I5KsF8Atu+B+cv9RqQIja8DctbyurUyHnS/XDCJf
F7immnEhMQo2h9LqiylzH7mjSRI9GCN3Z/H6iH/6ljPhrrlh5WAdw++sH8wtFijJuHO1kZCncPWV
bNZod6oByxkvXT3DHX0TNzJa73u/3UXPcPXA3Bpq/TFzmsmoRFJxqjCWpbXDEafmimIDRdOQzUUJ
DZ0GnI4OGj4gYkl+VGHZYCmmtdiqP35FU+s1wzZXYkK2p2VmZx89/izaaLY4LXmIp6U9GJUsoHAe
JJl1Fiv9HwAZBwg3f+nY9gcEcqFxJOJZTEkO/JONKTHZBXZQnXuAM0MuQ2FI0dlkWL4m8szJcMMt
UnLzDw28fVhrnZGCcwLmEiVMD5G9J9WueJr5GJiFLXu/sZlOsPxHzsUXqpBV3wOX0DuSJJqdgST0
xCrLG7cgZrN+WvRtm1SN1qtaMVc2O27vcJVQ1gREO42Bh9MEUtLPcM+Mb4sEeTRHuZugE5xRUgpv
BcEzjLIaC1W2U7pHuZuFYfAvagWgiZ15C5tcaJjVgOH1eSW1pN8bWJFTaegTBexfNS/REIh5qn0R
IsMnDB6c5gFFhGMaVfsJov2RYDFgvoU1P1IFZmEM4kPEKF3cxy1Yx4XTmtz+rTpJ0bP8QXGAu7aS
X3yhw0iDYKG54RchX266gpWulWIV3eXFx5+nH9AqGSQTHVLZLkY5C0pJtEt0xFGKORaPhaP1rzmB
F6MociHxwGZ5PAri7qhRmQR+5z/0SaWhDpyivDb2TAiheTDFkNZP6t8ilA3/1xVh37QPkKZJ58BU
6jBKmI4BMYFdvhdkz8JOgo2v6p/jfBFGxuDSeHKMZJP4HFKaO1t4zMFaYW26xeuV64I944XOiTRg
IUh941Bz7UqRXIuKqQEcfddXak1eNAwhHxX8zvo3OoMoK7GdRxtWwRsER8lqXunzJeek6Qlsojf/
PuBn0sGErLUdSqdcYAE9Qdchp754gqM32KGTBN2vIxOfzeah98gxwvISvYexgWQ+8qs2pRgeJU+h
TVmEc1MFuJO5rzKboY9ujUw7uPFjY0335kIIUha0IgWO4Sr1XhT/ZurYeF5jR2tb32YCfqifAh4K
ZtclMSqCRsjlftfCbYKNY0RJurLYcNtfxF6dNGGnF25x0Vi/iGaLWBnuBI/TJ/aTwxdIp8wetnEl
Lg79CJY74iGneO0n8ZEYTzLfpRIMWy2O2nG92BA5Vrv8xj0Pki2dUsj3rvITzFGJB768xs7uTm5f
BZcFHOHeo/j2juR8447+TJ7r2oGtQ2ybGdTWIW1B4gJ65P6yvTangITLA7uoBACU+nO5zNBXHotc
AIUSCgSkk2YAB7TdTXKKp+9YU3BBOV83TTD1TsJR58c2VqCda4gJX7c1IlGeJIbPGf0Rvi64Gktm
QX8McLUYex0NDI7JZKVfuHLEJ9BX/13A6ycGEqAMV2YiIgCOP7XpbxMsMquSuOH48IyqfmGoYDmM
aSH8604FgYQIC8GFCDmCtZLmku8M8Oujnv0awtB7hDZjJ+gYJJ8fmWyuBiwgEy2d5BhjV+mNoASk
QuF1A9+ptMj+w8OAJg8DXvMDPyjIez7p+eB5Wtc82Kwk0cUMzE2eHupNo2DihLeUF21nTr/LgU19
ni8KSaKPbDEJRY53bOnT2YUxuHRVLSA8s+gu8cLz5QQYcVGCWnxYMSowpWuy2QOKJtTGsdFtQIqf
7i+FttlTgfi5kNnyT5JXNKtjy2yNGrbkOv2Waydi0pDKBpvYZQyEjbz1O0DEK9Tmq6VFq54n+fCQ
h2CbUa52CtKEo1TKN/+CIzobs6TBDGpl62hrAQAMfsEYxjtp3y15Bni6f1gsL4nB00wOtoJlQvDg
m0H4tzUoBmJ0fNknWBVpsl6cGDeGNgBwOQlmo/0rBLjjDkTX0Rw1ZXPOSvO2DSqEHMdBXQJU45Lk
LVS8uL6wHxKtzTPqK/wqsCTXgyeQ97+sAWbdU/C5Kq4Cv/QSMH0LqGaEiw97IXVyb63z2yNlW5wR
cKbNvJmxH2KcpicMebTQObHTJJG2sfqKNq17EnwNrHqOswix2DJFuyEl/7ShA0dgHtZxfzN8V2Rx
BWeVHJnyFqg2drN8Rl+TpUzdbHx0HbejX8KnvxCSHIuDryCI4rDDlZcjeBnLUCLL+vvhab2Fw/Jw
1KjG6ifwtcftailLmWA/iqESoV0ZQu2WXQcVsR0lEi+GxF4p2ZOP0Go+ooB2JbEHZkbotpJjldRM
8K5pDENbNEvnA714gj8HlgtRelOUeGEgkSq7wm01Ix74OSAfhqf44KG0DBg3bw3HftLftSIxvBgO
byDY/z9w7SrTpK/vV+cLIWUKzK4PS7/E0IMvUNCaP+FBlVd6pzu6cgNzWulGvrSfrLxEU1/3VWvN
6KOePh//OKbpLW+x9w0xoqiR5Q4MKUU33Sb0fAFdfd70SnaitIzi8nHyGWoiBQ3R68E8CJ+9GMz1
Nr9bhEbFpZpSMVPpxgSYGeHlYkXs3rGHk+EAnC9T0JB0t37wdDCZAwqoKbG+0xtGFBcwwIrXpp5q
S3CFYBSD2EckkQrVPUBCFJvGwuLsvgk1fTcBVJk2yIn5V3FHfiOXZzfnEo0UlYBTUFuH/VxHHWLc
yJhMuHV6i6ejYy5FOc4b1vGtlw4BcriOk+By9PxtmpKFSjYOwoj2FOpqHJ/m6KLvd0WayckeQMmu
/OHBL9mUHIZ3Lbm3KUNzKfpMz/r36h/hr0QrJj3t04qVAOq30HV0batZiXtsZXZySpNJPY6TYpKk
2C9NFRgTxAbi+0gQCDstr/dQEFGe/TiHFeWG214AOs0dBozUBbgM5wb0EQsSDPsG6Lyam34h2Jkg
unUu07XtFnetvUhlV+m9XzjD5WWFiWO1IkR1d800pt8IPz9We4588UZ6aFj1SkdzM1TTQoHX9LBX
tKPqoK9mHpRyM0mQnTPGoh/YDQcWfWe2yTPbe376MJ+thch1lkBPKc2Wtg0HpVAR54g4S9M2IZ8I
rvVYTFFngbnjVNy/zMfu6JLk3oJHfI86yGumgq/vWqug0vGjm3IV63KQKPC2QaehTplpQ/QiBaPY
uXQRVk7VvqmdhCgUB02VKsVub9YsfRaV2L1/2bjRkfkw0f5e1nGkc/1aXkVcyWE3IV6NUvBsjYfv
CTuqG8Q1SRS19Ha5yoPkn+SxFZ1IbttEKx4pEsRa/XfC0cQeWHRlrYFBMUOmStPg5wFhuefLMv7X
rYhPvT8iujLY+AjlaKbb0f9aZSQFXLIz9nGx9k9ERb/w5uZYoDRUHxRGdwiXE+k8u6TLqvz6iCPv
FG12bmNFoyikEAM9hTRPQszClOAmzMVyi7dReDWkGV29M+A5gN7xPY4+0rSNnQn70x9PzD1K91NI
qZv5MGdwof3EazOg2BJ7ahQk1kf7szhaIRmv5WvMZSu/SaA59ErKuBGdhP6W0UvSRscFGfgnnkZO
Ez3bdulUu4GFhrSV4toa/X5jlAKaiBITQOuLgPjSiabcZfgeqBKxxxSehFjl8AthFmabE6wbyf/L
tqoXe8akk3oMzNgGT2peq8pGYWLFM0GMSdcLufVelUQGKUr+S5mvaj3yLalO526qu0D7EujJntFz
SSGrKauNu6QQ5AM6lhmiWOv+Idu3oFOg2VqFcKcwU9T31um4pI6s/Wmr7DHR0mTfdYJhGNSsuOR1
t8icxdPx/KYjrwaptmAujbEPTtIYz9CJDNl3ocMaHrCXWxebMeuQjKJ09Zojb+IflPJqRPdvJJYR
Ia8fiyJAF+siuH5GVt5yXkYZD0Af0CwK7eQdT397spRwk0rXU0eC6noCF5YFe+0rji5RrjJ574im
LAQvg7Su/CvOHhCXJ1/Js2L1d8uarg2Ih1qN3RlEw3cARpEtdQBFHTX3Frh0K+TPrR+VON3CVEry
jtgh45mMj+jQjaoDZn9phUHFrC5bYBPCfQ7NMRXoROBoif9mfwashOYGlkjqJLbCuuU/9P2komx7
Cp8yoUiJll6144udVrDQxW47he1MBe6Za6uZ4meYWjJ4wGr/kT+32NkC3eK3e8yRWwsQuP5SgxSG
tIlYiGyL+TRfqeIsJhiww9S4gwbTuqJD2l70cwtYzATOZ7HlLAuBOGoMZcF/8oH0GQh6A3CwwtNg
FMmO0JprjuWVnxz3MmnbYxIRv91cVQEqXjFd+k51JuF63RpHv6kccIUD/HO8heMwxb1C/OgXLUMQ
vcc65h9hK27pPDhS8Ih4XOfRJrKsQXlv5b4ewc8v6mYVs9/CqdbNa6HITS7V6pj6lTI9pZG2Bks9
rhuwlrCrhwSjLaXYi/2R63TBn/p9aSeHvo9SDQFMbCZTnf8kyyOAB6Ng/u4r4+Z1lkZ8eVDtzmm0
sePmJYNXAUskj1PzLXsqQkPm53GniI6htOWukXpbs9630u7TVMEHku68FWdfHtntsQF6rxm6Z/Y2
vzCe678CQexqyUWWroy6QRdfX64W/I3kWMDG01FjwVtI+ZJVmn4QOOEFyFXXQUvY0TgZAvIe8/qW
pyeVnpFXd/dh9nj8GMX6GzX7hhcIQjruxB4IcFsFRpIUGTIzOPmCfFTFSVaJOlO9XjfJy0X3cqxD
WCibo16BB7j07nL2zaFCg1n0kaOwH2bzr+rH9a3l0uMEwa+ILZ5QcREQV3VqgDw5s82+CbgN3u3X
HwAIwV6Im3AG1JGpzTbr9GjghhfYdiJ3w+dOJLdW7f8g7Cls0YygRZB7rVS6xNhTKCM9X5+jjFgh
yH/Wq1luwUyUB86++2Lf1gCe4tGoMKbRUuwi3+NUuLYPDvHbzJ+yIQpBeJRqcYZqpwo68kyIHQKT
vkZiXdWAI3daf6yZpcwi2KexUVbb2fn38jgWQbLW/+4fYwdt55MvAbrl7qbxamyUR1rtBMocVdYF
19IZ8JCVqlI4G6pnuO5sF5Ahg1g5Yac8iU+qXxLbWOwezCw+fK+1nj1M7n7THYJ91oyBXYfRZ0q1
Un0u3+kvg3+oh/Yl1LPzIYdYgbbL/jNSVcZe1rmo86pFuOknXEMIcd6GS8nSK+X73EdXK1CXcHRI
YV45/5XxAQJ8TaYHrDm6SbdwzKGL2avDmS4NJ50S9tpVRFiQZ1xcXGLzqY32jZxYJuKYhkAxXuuP
LoDoE7qDgxcG/uc5yy1Ucx5wvbvj5m8o1QH4SQrpuPj9sNT1MgPOvlzTF/gZ4g+p01+R2UpV78Gn
iAvMhwmziZgc24YJR8ISWKH8Y/Jn61cTjWLVbF6h+T+h9cSN82sKqXkGVXCFxwXc1TJo4s4upLT1
Z60X87JijKqEKbdJG/M8FzqSPlUcFuJyH3pJzMh0k4oUKoQQRSCYCL/4lYbikvRbadrgSz/yxJ+A
xD2Xt4+3JUMk7H20MpULUFMfGPZuIIRDjYykiry3bcF08xZf0FYu7+vXbdQS8gTZF/8JmWKFP6Gf
N31TaiPhKcnP2JqhDcEiDhnMp8RoTp8slDdfpRmposWFYlwsUcPiKBENFoXguWClGXkv3XJ/PNeU
NwUV/QQx4+/eGtx59Adz5yXiO9MvpdgWQbTx2nlyHHHQ9iXfBZFvCOzq6dW04YbsJyJWI4BHGyGb
nsnpyg/VtQJHMwqHT/BdLJsoOk4UT74TyId2qesLWQypvRU6f+oe1Gi1r6nimiYIvO71a219Xyni
sVrmv8uy2dNeVWH8WUq7eqaU0mVXrdUMEzt8ybE3q6V0HOis13XIUIdEU0JSs2qIPUT9YbwBwU2d
JuJ0/w790zASf+UwIA2mhTalKyp1ATVohYmih7FGDWNf7//wuBX5M1rc7Mx68RgilvZ3HyxqyjWS
Uhfx6calOY9wuG4vDw/Nnb98+NM+qJAnWWIVUa/W6PP5PaCyxXG6lDopoRQcp+DcXUV8MUcrpDgq
+mLxBmKkSbe5WpxPzNLlIM/9MQDoeeK/36kUvtHLMF4MoK1r8x+BlzGJB7xMhJ8LxfG+2fcbkP9R
6kQ20ZjCvs06BxAeAfCria5PtfKXhHR+EMGhNSwE+aEDKOKuMCbrg4yWahddohD5zIqdsqTe48Ro
J2Bga79iWXGCOFeAcQ3sYkCV6d6iD6AIxHWYJfqGXBHkePwT8CbgNjHewbZ65VjlNk7icnjxrJ1K
QIj78MKQ+wP5I3vzD8zPlO9a8jdJ2JUfvxmf2S5y/7xtm6WtXgf4V+esVBLvpIAmV4jnrEWyDK/m
cMIil07NVrvF90FMVN/1rTj9f5h7JQfMRrYj3gyVGFaOWHzSC5VyZvCPIC5m64+hQARUSPoG6R+D
E0fLPjwJdnFxCdAV7MzsTDYGpBReg1XmUoNp0YZtLNjfigyqT/ROH4tjC/T2AE76k8TacG1NHPDN
dfPBJIVe5vrWQCzm9yyKyxLamEwfdmSVpMs7+7zsD9ttHCtTIOjQ5eVGjV/KhHqYqTn1p0oOACtI
snaFyJ2a/rQ3dFaxSriQ4nN/eZJQPzyjE5zILl+19H/nWto1qxLiwgp6AXI/0VnW1KzAGhq5G4iG
r13KffrvhQ9b1jf8lwhc2slVEZwGNQRHtfwpuwO+j1BaqWtzCFF/fTbL3sLT2hWHrl7H5PWQ7UH4
QfxeiqkREIuBg2FgqJeytTO/AsTVBTrvi4/7Y1TXxxYSOXy4YTnyDZOB7Ontsw+q1aOj2Hr4Oph7
a/hrnTzq48kM9ZkVbZBzr1dF2mSuYvgcse45UMkKYqZpCwcrgF6zwkrWG9R9dwCquYdbRHUglR3l
7g1o2E0VT0i3gfOmmUIHgbsXH2aOzRDUcuq6QKysDScKV8Axi2CjM5DnPYACzgyXnzPOwlUKM2hU
Gd+o8hHl+ShHiridkYz8UBT/jQ5X9FDBhpDHsCKAB6aXzUSJgEm5ATrDItfS8e9q+DMcIaQqUbDp
gN/jxMfcQK1OzbF+qPIcpMSfpoG8BdyMpzxg1vb5da/sYo8b6nFwlZHe2l11ofGdN1+hJsNjTMZH
7TCeLqQClStT0Yl6I/uuCPvO1d8xmP1iLfHJeiLbj2Uc4PLPmOlQ4daYqKofHQsaDKOhi5UpcA5X
LZvRKzM5P6epeBaqnB0iD+B/smg87EbNNmgPduTg1+iNRYzH/AvAXgU5R9SBDZqLX8an3FIHhFlP
e6Iev+N07r8Rt5NdeUrLQn4PR4rN6D5aYiRmVxxF3agJGWw59TcumLqL/Y7MD1RsaNKm3HDLVkwo
FwgLXZDBuwOx4qb9wFq4tE1fro7AIbPW4BYSYiB1GshtZXo0d8/fG3JenaUPNc/TAIWwULBxdm1X
JGojdAJKXvT0wmgKdvaUKeOLGSpkbVbk/aJvtAs9mVKy8TSSANZ5L6v7eUnhlLc/P+caFiDVb30J
H2ctgjZ2negloA8re93hDnQ0YKr0t4MjOJLlC7Klqoodfudcpd9YLp4Qs/aNejrzRYH4BFF4U/Hd
4Ytu9gVhFsvcdX4Uf16nzOp2b15x9ST2XkVEKK5bPLSgzRMNaYWjKTeHJVge0BT7pmnh4BvUz00B
dbbTMNIdKSXq83dToQpEc4FR5QVOhgcGBqlp5BozFDw/JpJYzd7PbrKLFt/MeJ+Y/v/U/v+q+kki
tb3UH1440y5RC/+G0kUzlrt5qRHYeswXOOkYnoacnqbbHnIbOm/7c7IpQX1eLdAfi+ZMoqNJlM8p
3LGKpvf5YNHnMQTp8Nel8xTYwP+aySVht7E3LdmAVy+asRe2FKYo2rwRw1OnKkzof3c+DW3rZmdH
TQM1gD+4DXWBz64MhiURAoQTy7qJyP5XwklDXkcRNR2tYaR+zvG7cWelfYnESnccCWXWSi6k/AK1
EF0Rf7dIfNPicmVx29UDNcf+Lomz3acq9oKTj6RS6PXEJgP5txDn8SNrGQfI8170ZyJSKUUkNUYt
FzqQ0F/Q9C4Ggth0MTDCUVTO6OGN07ns2K9UV6BHvrYt6ELKeVQK3k8iJnDnhEONdqzwpCCb5yG5
/jDgQLaFVoRUQ+alCo1sSpzk/AhO/fB061LEnS0zcRONybm8zyc29AQksMpwSEzcxltNqdeErp7a
P+l3jBKHh9Tbb7X+q6IudAWCB+ghQPXqWK8niG4UWsJJOV8AT1E0sH3H9RDtF7qc9lFPEHvTt2Y2
GwNcAvFRJU/bcWbsIXwNVTCsOUtgbxy/aL7YaTw5JAa0sCJBfrjn1mUzoThxG7RieKLM0AmInrjX
3nPO3dPd3i5zEbHzs7+WkRDcjQC4bFCvk/55tLUv6thez7/cZbdHoaZ1jljJCp9sDMBznnFHuegw
uqoPbJvhYsliXNjp9WF/XTc3dEhWz/P7kPSkjBQ+eSAGT9DUv5/PRYH4iJcdO7PBW4I5ATB4cKTl
21TGFFfL+zcdSraUsmSyTR7/7wdvG+ctoNw48WTl5Fl28T4Q31zZvpj12zjQbXqngjw93k7gO3Nc
fKM3G6VIK7qIx/YRMqMgAKSZnkH+q+0BCL8xhn2QguWmC7vQvk5NOtdsRCrSymkb+vWKWg2b+UPo
Mv1qWD5NxSeR4nM4v+DTe+XLUuP2+7SCDvNgAVGknCM4kR8doSU6OVXsnxrTVY6gkfV0gxJmFszd
6BehxuUbwBSQpFcp2hfAtSUEh0k4os2MhTqTX33aRuyLmWfpM07RaAD9+QB7fByv7ZRUwqTM7QJI
8Hyaaz7QPZ947AI6DMAsCFxIxD57XHeRuUupHFlgdmZ7zOd42GxU++Vebb6CDuljCHg1/10vF1Nk
boJP0fVi8WFcbjZM0U0bJTavX+/OdnnNleBlmoxHyBv2NZ3lcHIn6AsjTxW/Vl/jYRrSxp4GSLd3
sKmW1QqP4kUPbU5bjg6uaa0WfqESWGHKR0Tcm8EC5zQr6CU5VSTv2Ar2ArEL0OcZVECjMn7BBPH/
57YDD+5Zo6bF7qa3A3bujOhW5KAMbckB7DW6rqdb3oZsYbdXS1IU2TUYyU/UWgfsPgcFkCUPDNf4
SK5kaquXcc/d8WQXyIKrbyuAAidJ+O2/tnarpC+6Qx3A0Y6EvjOA4FpgTdNXLFrFlvyVBCVSppga
iXlU5aTo9C5o/8PLFeo0j/xpv155uq7d0gAWWWjeB9PvpsdWsVldgfaynIDJi+s/Cyvb19RpuOdG
SC1u+h7EZUMKXOjLB9yNg3T4D0r1IPLnZVzRWuI8i3nWfC9V37k1ZSqAD+akpb4bRXveFMhVrzg1
fxdNTgIhKJxPdliVysWlgFMK9utXIWqC0jwA7pJgDagz0ggHA79RWwyX0zDAuza9t6rEpbugx72c
ShOEBtvRMiooW0dUXB5H+r3G9fillsh4wmxPA8zot2N1e4gfCxjPqdm1W2GNXiWjd7rRfjlKoosk
y7NZhgugBcnbYGkaZ+TZ2rV8aBzybMa0mG62fiJfWw7oqr7ZIHvOkmWqw+GCuM2JZuMhaE3IJyF/
vFaUy+8CP6/HiUNSueeSgkv5tH9o7JNUHAbxgegSZ+usPAqQzJKVeuCKHCqYKFz7LpaqoS7fCP5g
BSp9fQ41GGin5smGfAghKHzHu9hCXCZIOerLYHtQP6UlT7Ve7kkr5r6/Y36twQ8yvW/T9HcFgLcs
4UEZ7P5GTMhm8ItZttubYrAY277ER0kLoI6jC49at3yNwtoC+UkIes3GfvZUAsKBn8t40Dh35+gW
x9dD1xiObuChoewvpeCJKMefyr1dgoKxedJfJqDy+Lat3fceCKu0e2oScNZwow3MO54Q0wJ9COg3
LCZ+Ky2cj7nTdVZaKxOHLZl3NnJH8LXMVp1wFPbkll2/UBFkHDDuwBrQ73c+dHJQsrhOyg9Erf2P
jG+tGYMTWqMUpMcnoxjGu3u8PCD5MSQoAN2cqthfp9Zy4QX/kjzE/6qp69p2R/ZvG5LCM9byQtgT
j6oJrLV0F9wvPrV8oXcaWx0gt5yMTTWvpRgrXv7F5IWvnztc/Oi4OB/HDTENK76y9GqGABpBx5Gf
ZYntw1s3Cy21oS/U/xhB/RMxXu8vCFBBvlJHdJUmg0NflrdMkx2aPmb7TSHC1dvsbCexou3kqK0H
y/8BLsPS+6COc713rd6mCQ3CYKqNSw7IJSykYIqSpHBDjKkddo4nBpvyG+aMruHkjIUoJyulTaUr
RAk81rqCw4WW22idK3oWRGmdsWGsib2oeOBZ+kqhDT0JdMzZI/eUD25v+UPN+URNnMrMevWp7lZv
iGfp4+8yh1Q5d9yGx9ynwxDMBv4X4X3koq05YD7iTa/UTM5tYgMXtUlR6QQaaaNlYLLSBvLPFh1b
SR6WhRsA0HvnQ6pnufns5PWdJO3yEBMTznmq7B0pit7PWnMO7ryAXc6yPFWkxCC/I1gbCG5E2iaU
iakXIq+qlkD0reXSFY6/CIpHPVSKJZ52Tt/gIN7aoAqOV35rTdDZYRzy7ecEVNPiZNt4gGZPNdFW
dxFQAYp2vZ9TtNF+J7Y17U3vE5/JCkcdnKwOui2ltJ6NzXvchBAYtef9ILtQt92i9VBSOyUfA12b
m9OShATQDyXdQTieYczK+NLf5fbpJTzDUggZIcbzI43UAPNbcR9EeQ61UANjUXuCtxNnpNFy1d9o
iwO3xaB2Xn5CXe3dNlo6j6ThIETjSCaiXHRwZmLNoEjLmlSHKMSL4NqQ68MRsEyS/s0Yl7KDGRO3
CHFQmv0OvBpROfckSWldijXn77Se2Kz1iuDpT9lNKYS3HOKte9LpRANWrgEtdOvxFRViNTSlvMFK
ujkPw0mSl3jUmjQbXbsDbA2okzuQdgGYIkIjgIVqQ38B/gJk1mFjguZ2461iTKWa8FAS/BJPaYrO
3pecIZMVKjCby/tabnan1QF00uMFLHSoGI41vmBbPZTDjYHRwZGNEUHFrpHikHR6k715oevbGOG3
bwpbmUYfWkIsP3M/qTU5ABgVPvlJEdYncFeGJDGqMwRRDj/MOcNURSVlkRxQNP8vip4vhE3x4LiP
c+FkDHfcwzAQB5nclM2kf+pgm07xB6DAqHCoXt3Pjjgu7Mshuy0LIcDlbZDo6FO4VIW55UHO4qQC
rlYUEBD9utQkQeXQkC/lrSxces/FjJLZG6y1QUW1JUaYz13DknSIoUvVW+oXUkw+Id9+UuO9dCkd
sthItI4lyPfrxiUoK2SNCuoLDuX7CUquJELfxUdgXnw6FMRtc6ZQh1ZKtwvZVP+UNO62Nw9UTslZ
s8VsMqL1ZFIgCke8juFv6v5TDXgqDW+pNNfbDtGbEDNsZ1zPEubya7nmSO7udU7Qh39iF3DGwO/C
vLuZyoRhPfmmEKZaDtrKkSXA2CLmAsrgwv2iXdz8Vih1X/U7dMb/ytR2FaQnWJBt15VUIlX7bC/l
Bwa0L72ddt1/YfD+vXabJcjq6G3DD7IThmOh4iJM96uX+AkUutCdCaKQXD7xyb3+VpODTHy3eoXU
ZLHqU6hXewSvi2KiYaqI/O6MULjfl7QIQ9YjQm49bXOSVdil1ygqSeeJrnoxD9hX1lC6WcqxXpu8
7F6MYUim+l6b+8tNFo/vdop0rxvQoD2hcirURlslKBhlApY7wlyNvYF59lXjUXMostB4PF21jDj4
urmC8TmCNXvWQWvti44Sv8xGYJjsG0Vv+9i7rldBZutuqqD20KqKF08D8iHDjWiVbSuJSSfXvQpI
hWizBEjflyrcKMVQsbGosXlqaGsHcKlvpLXPIrEo8LVOFagtMob484BFpZd09MkSlXzKwueQU3V5
kM7zNKoUsxNN7aRd2OEizRZpu92J28hi34XbHETF+G1s4jkOTGVaZDG8LF4K+kCB8AOmurSQGvko
9BVYv0zGq39xYiZZUEyOiof8sJiJL31Jr4c6TG+Yy1kXv87+5Lfh8/vCkGktZ1Rpra97878327Li
Co5E8Qk2gvNz3n1kSXpqe1N++bao/ZW1TYPx6m41jhWrddMJ31Xd8VFbxV2pZob0SiqVB4KMPVxO
GAfcrM9jQOhfy6G/hCk21IDGHEtBvef9k1+AAvBNEriUo/6hLZo4leXws0QLt1f91AaiYeCMNCT4
Od7TTQqqhZqq+m7WTKpgPTrmt9LnRn22pTizf0e1/T80bX7D0VvX7aAc75KArdLxD3gPtcoekHEm
4AmQKg/zlNSoEQjST3DqluKhO2VjNdMz7LHACbwfNNiC4re6OwC2aO6KsdOLHM2kbjCvQOfq10C0
HG+A5aYWTYLNFwIhB4DM1uNZM49iNDBtXCPrY+voCFAPTslWi4ckhC+Jv1PMCf3k/JsEOfk6hBXx
YASuKB09PzN7/u82OzPj6v6dq3nctyqMqxNweVtB/BcrAC24pFw2Eiz/ukmLhgphtNF2HIYc+XmO
7IbCynUlxVG3kLzExIt3xJc96Fn/gokrLJi1h2Wgxa4bbuvIXDYhXtWAHBg0rDh6Z6Qia95m2DT9
KaBmvLIpkmHN+CPoMu+6GEtVKFzmG8Lx1TTjgRS1aY3VW4DOl0PhS7+23NgZ0Lz6J+KPO9JophOK
Fxc4aq+MUikHEbFQI5wl/3ii/eC9TRQNqAz3vk+zuImMZehbEbIP7YSM/OJ9HNLIMI/CwR318fj3
/7YAjF+PLyIx/ut0CzeGPsFRKgPffmQL2iMg3Nhtccboj5W6mVYczNA2UfkdFdbN/MXk0T6Kfir6
9hHuDCkbK3/2pBN+Soy8i8SBmmKgrbYEy0NESct2rljZ6P8dEO/p3PhDiWsbzW8Wvpv6NxcfwzVy
HEtDeCCDZupQVhwd1dfpuc8djFvPMOvaS0vj5qZWNYuhs81AGrIaqsGWC98rSBUOygvoJ4x1qKoh
IG+g5DKhA2JHwN6mVN7VqWisOFKZFkbstnGdJr/uJwxndIcvphBRpl+PT6sdn+ADxABqTsok6DBE
b12aQ2tnn9FtuwnWegBXTTKQi4HWdVGRptOm2wl5n5sm9r1DUrnBKTqgN4oqnwW0LQkuBd/pZcl9
ASDibClqPVhA5DhLEWkQnwXTJ19UN66NBxrFfkWIZJCNcQuwdXrmcM7vNEYXSteuzXa6uykyn4oO
7FcihVwxeSvqDFlkdhptR0wzStWJDIeiPFYIgumhS4vxsxfNaxYhoh7O9otLZJ2TgnLqWGQyS7qN
EZgMzVR0hcyzYqh8NpUqqPTHYP3cm8dNnQB6JecxmqwogbsxPZzjj3ccfTKSDOJScxvSzTg/VwfX
NGAWgX/Fqj7AR9CNwFBhjfckqE89z8DYB5eQSYOFL/hggPYMafcTeTt8jqmMUbiM7EF5Qr7336An
Bfc2/KxN6azM2jwWTWi+TP1YzVs3MDVUSpc5zG1OK8mcXUJB93FBl8Z10aIH09qWexG7hy4fFGEW
aToijW8IIsfQ6MQYkFFkKB7fVCVUEU5y6UYbTz55FwXqvFFpPUJ39YvuX3YvlYEjHLDgOdB33r9k
2DqTk2eog3XEt3v6ojNNDJ8Ua9lnDobM9gr3JdjWeIVCNzR2wt6YwuDd6CgTz/TviyNC/vWI/iQX
DYQjF+kSHS2acZEdoh58FeATBzsJ+sF5IRC2SWErPmXkHU8Vo+DRo5Wm+o4/A3FS8Zgt8LzGW0El
oRgqq3tEYoKANwT27QkJ9rRF8fqVIiBe8VBHNGGAzF8XoNt3n/ZXwxaUpnT2QOss15jv7SoD0igR
4j1oRMy4JL/IrDyVlBfLLzukVBrL1lLyCYaC5NtZ5QIiMGf+YScY+FbIJcSCD/WhBd3seC9WdBqb
YZm5YL4hB1CNtv0g7O4ItGgLu751srd/NKGLWnGWgfdma+gEooZGqVKiShn/IkcVXC4VMFldxYln
TMWF/qiG/5siDvw2D6OW6ySvjcyM8GMwjcRWrIvXohu1yfZ5CcPwHOqdt0IihHNbVyXDeQf8i7At
cyr97DTdiiq22SvuffeW7AXJWhkZyr9lB04vtkkLz0O1dgz710TM4IS/TMYtGun5GPinCrwRDrnT
07DKNZGdP69p4y2H70A1Zii4k3b4S1pkAcQDcyv98ZBhMA0Z/MBGm3vo409BzqbzH4TB49Dvx6Jc
6SMiHSc++SRO5t7eDMzfh1l5thU5gJCcXlOzREE3GKW4TGB4QXjn1BO66ApIazeJnJ1ZD5JNJpfi
6z9MpxppQ7NSbckz3eW+BvxfKeszXzFfIn5HmLWanMg1//DIapYdcNa6jdiO3VZLwz9NlhCVQgsg
2BSxgXrVb5Fc6m82Yap01M1U9R9lxtDCSKwH/NOrESaqUYbSNSIOdNu8uwIThGK++bogsj91ToWW
lnXe8WJofkFwk5DVpUVI42Sf5mR9dST5KzvK8NWvXhSs7YUVPtsqBtxiprdr+I5xK+JoI/BKxGkg
icWeRv1ON7HnIqmQlk+Dll5MYM6pxoFRrDrxveEtNSwdDtc4flRmY3zZUq0U+fIkEhZAyz/Sf5yZ
JbeMklmVTkZ/Le5wJ4os/r116Wg+IVIozB8kO0Z6bPyUWzxLnauVDG6bltq03+iQ9GThudSncvw9
gWBU6y74s0aGDkSvaa/n5u6XXBIJ3P7Py/fXP/Ijfs6x5L2rbagC99l4KaXIJvwsTYh80Ee9M5xr
CX3a+8heCFv1K3h4HZ1TD/LC/ztBQjkFMuyDlrbvURpECYoLNsjARZ225SQseJrMgIIicKTYBu0G
bMIfM4N6IvyMI2SKDLWTXrstThnP2XCFs1XTasL0j7lhN0uai97zB1BZqBRqR28q3q+boMb0QFmR
aDz0MCNnMQmRqqHcejOcyH4BTv/+RWoEV+OH0ci/ft2prFMJsudVWeLu6ZVGqtUDUe+IeugbV3iq
tye7hS8apHdy9INoEgFXC7FIkdAgyVgaX6dHysZamvB9xd9sRSGIpUkZxca/WoA5oeqBJz7ewpu+
IgWkoHuixzDSGNzFfmBTyJdzUlUkp3Hp/6XmdsL1p7jcN/I7Fm/HaVug4WUkkWmT18ITp5jZXASO
NgroN1Cw2vPICHo+F+Dp3ZaRspcNy4o+SxdFroRCOXauksmCLmAPl3tieFCKclw7Qn6idmryRwc0
+6hRUP1ITEhtnxC443AiPkn6cWHwOgaZf3S39f6HvDo70H1sbSFPNIwPCSkPk2UYUHCGj+f8Nkz0
cw2JlBDkxo1dH6ZniBi4GVMe8FN2XnpaUVMy+8Wq3V8EVi2EkptlWPJh+6uv20aa1rLYMBZ3wFcE
kuduMQRqmX1iEE1nUUJhQnL0cnn1HI8inasu9u034Ta6cfRv+w7/OQxvDYmE3YNBqsJGacOTmH3i
Gx/4oPedZLPwXM8k/lxN8/j/CCR5cuCxKJMzO7/rGk1Bhqmu5gUgsyya5QaPrlo+HTD2UmCXav5Y
tx5jA4sAaIp8QPOFX2MK+1YQ5XMBuJ+pa3F6FRogMebCdVSIWT6EU0f4qbRand39yPjpgwvBsdP3
ALt2DjWTYCyeKbWBCPuv6l+LgYLzFVNNnuYgbeYlnfQBc+nyKOYc59JbWfkRe0KzDYk6nz+AJa0m
wpLGJ9Ut7n/4ErwSaSxMeEuTTGbqaEHxG4khStdBOqRyekE0TO4WZUvwESUalsnXuaveEUcg33Le
G7pi1xy7IrduQ96LCSva6Uk8By1peT0iAvQBoT/fpBWbhXpsken3Rmb3L9rmWVWCO6cUugyI04bm
W6Zup1NW4lsoISuqOb1/KLzm18LK8oSwHrox8SZBI1yEBcYLI7xHQYDXkkwVafuKIOgNolJwyfs1
VAe8sIE4XSuGmM5jms4gbN8bhiSXC/n1kL0WMuY2fnegnjOe5UritrTOZ7gNhHdfPZLe6rjXELTE
oZJosggxPptYep72TMYm+2KbyEfVTWka03LJGHIvlVjwngzSrV9wq12HAQy3vinm31hG33o3Uy1v
wlL9tLKbbPDPZbtjGw3+LxyEcWFtqHqylBWSb1sKK1N8EhHfZcw5CNlNwEfYxfEFSGfs7CPO6nCT
K6ZMKq4TTHj6bdt7lwXAWgh5qJx+bheS76plvLr8vYYLulT11FZQsLk2afbBQ1U+bNaE8HswLg7o
OMusKg4GgOzgmaXWQJqllOjy9RRwl/CtSuNdSFmyZSvwbOWOCaXiQBVVvrPAKWdaekLfNAij+NYL
9LtTVf39/OqCpxV5GCg1ekaJARAszRouaZ9RtuOSpaLRPOIeDTH6sqAIXi8hKjnuG4hq2G1l18NZ
Q3f7+5HfA3amDun+GgXqtI3X5sF7HTB24sGdHEkgshTW5Ra/t+byRa329gql4swykNXhCHO88Ct/
mSKUCE45DDWsDC78FAjuTVU6fA8/TMlcmt+yALkvwHY+bvgeaaIjt1L2TPwRJ6hnTsLdjpT+DgQe
ykaeCAJpCJAcnMAt29WxMnAPnSwna8IBHCRXclbXgxK3Z0cHiDNc666ycyQ54nCXbUQy043K1aEM
5LjIFnELNDmMQcbW9yZtXS+PWE0wjoGTDumhuj8BP4nSVN1etXcuCy0zm6x5E/botnxk7vfGGH4i
riCIoTURJYZUqeZt6xKxbG1Tq9PX0jI+yEWIZVhMyBt3rrw6JL8Gtq4SWJm1M3GtoZ0L/K47+y/G
65K//h7G6N0jJuwO8ziG1ci3m2I1DFBFCw7ZiRGm+ZpmVF1UwIplWGoqPvQrLAo/x5mLGV6zGEtB
Sq3fudVbtXrOEtFFcW5Qazbje/lAX7LUL66cf8oWaBQuyhp56oHV+c5buJy9pNNqBjMDB6yR39Gs
yVe/4TP22qEMiVKF8XWs9+7Zg5etLu4m69hwbvypCEznPyxKFEPYV8j4UpeWtUCkoG6IUtjfFpwH
C6yPDAezvS+m2ENPUjQlOoMz0mY83YBmmTqYEITAvx0+xTsh+ZdmOXqzWVROszLCYN/CxWo8XCCt
Y15eKiDT2n/zxmWLLOwcCOeqoRKADgIzHuDfkNHzY/z2+d5cYn4R7/3qXPthAIpwjpbQFJlBEhXZ
k766oyjZoSRe60FysD6yl/HY37nEtc6QVr61nOLD5hqhZqeoNxa5EnE0jrAFp4sUDl4R9MoYiQFW
s9b52bt9pTaBR4zsxfpGnRXse5VS5E5GmDHF0OziRzOT/7ZAz/szZGqNqbZpCzWx90q+y71dZtHG
sxUWjOySruEZcgh9HxdvGg24TMzd7hhzNS7QcfVvtzCRITfYxu3KJEtDpaYDfZrz2Mh4inCivJFk
u327WycnWiXIgb5pHqrPpUjLUjp/Ebng8JLKsUv63qKAU/r3mcYHo9sbjWaw+kFyMiITPePnm5No
EM7gctnxbB93EYzi0HYXcZ9e+2XkeRPHn71ei0MLe3IDEOdpLymsmV0DIfK7NANlMgA1eYgCVaiu
QmRLV0CYs2NwR1uU+GJnoyCe1CvRa3qgNlA3+BgSe0YrSIL4yhrw0rJNx5015UhSmOwgiIgpALaG
G8ozOQSM/sfuVR/9/U62UU3V4ZFfc5yF3c+R3y5KO+H2qZrxWhMwEVSMaDtfiHIAoaSKotJL4WZS
94Oi4Eo7AAL4IMqSQPtHg7VkVt1B7ztZp8UYHC95poVn0PrvqCeOLyAsBBysMd4IG8CNXVoWeYUj
RBYaFw7ANb2SNR9xMBjgGtnLJYi/FJIIlVMffG6H241quvipyLSf3xXFTIfMM7kJbH52uvxgTjjL
Yj92Du3LGLcSqwEnjJ+7xKNTmBjfXjWhLzDXbzNXq4Z1y/2Z5tfHGadJWpoTftcSzNswDNTU3NjM
HO9RLaagESoGUDVlTLAFwurYKqIY9r2BSunt7gRcUzRuvPfZZq+AY8A6iBHrM6iQ/rlZlD3krznI
m/y+YlrsrNxyV0U5wdNjf1gaL0o+3SzABiBZmZjbBvjoQhITZDDSInfXPpmsTGCEBdrozUFWjOGI
pA9PHcJ7Kr4+68OveKN45j/+g2JbkUist1a9AwPoBt/5V/LMFgfhpRq/etjKk7c+QC6c52eoFhOt
/RQtmqJa8lOb6jWlHow0f2AP+YzGZPtwPGhQb5NDAdJtu6Mj2xIhevxMwUSWm3OvjgTcCz5KE5MV
NdQGKxB3t0/29oYFT5F1+36xH1jHQ86oAKwmOnFVyDztTJ78BdwFHO8stzgH+e8HaKSPwdVD6u6Y
fegELL143jbATLE0Sd1Q5qzAvhPwQz7vVb40Q1oE7JXSuUm9TUBJ1s+/9eMbyUGJKJaLOKgKCTtv
DIXToCbofDJFKRXyhrlSm5prlERIr9job0MzV6DKfFKjJ44ppCVbdNBgnaPN9KZE13VhE0Rb5Chc
oHa6LGd2YYuOljY652rHEDoKz9c/jVgAPEltCtMTEV+8Zbvx/pkN8NmdS6aD+QJ89QWOpSY02mdR
L1cZF97o+Cs113GZ8OS88fe3r2cSYeuffGiMMIh9fO9FVaLhwQY0CSAJ1a1g5b9aXvBBjx3AHVDt
u44RWMN3GQXP0VT6I7oOe7FSd5VDAqFzkWrmdBC6OybXl5awLnUsptEJ2M4FUuLxGYboon8kGiO5
+nXV+8NKUamddrh0YQm4IPgT5pXjbmvQ1nL+5fDDb4SUwDYTTbS2m6kIqPs1T1Eapic0ZoxcAhVF
px622Ylqh7NsjwH4zBYb8FSdfyCovB5itb5bE+Fp0ZroifVDA0B9+6ANb29P0ojvNiA6vyPw1976
+LaXCpg/zr3SDLiYrJmJlkN2YI6N1go/q9ScGNU1cQrT6yoARSMF/RiRGrsjh57AyNPmfFnHrE3y
9/vNRU9XRVlket4c5doOfQNAjIQ8gMWK5Z/XbbSSfm1oFxiVZWyyMNKczkKnGoDbEmr5yV3QnJAg
3pRrJBq2sSnGln7g8TIGglku83Wmd6S719I4p2YnW31hSQKN7UEypo8jrVy5Conb6AkqyKB/3p+P
O2dMMrJaTE7eWzoxVJZG/y3tkG+edAD4VXHfr9NoWnFwFLDEEV6ImcYJczVFSQ5XHPG8zDZ1nSHi
BDKX5cQIM7tJR/JPiqONjrXdirzX+KNPrDD0g25/mXGNAyFhvcB4pVv8gXQyQMW0Sy0kTr7RnzfX
+zKfAI2TgraSEdOM8FHxEwE2nvFgeTK4OT04uVq57Lzy3wzE9T1ZI6YogjKHPyr1OxpEJ42rNUth
TYkYhpFKkFM3NNMA9DCnN3oCCvl/yVF5XBZu6kYSPdRkTGrfmIF59JUNJ6p2Gp7FgYT46j02KaHA
86xoJHd9PuRjVKcfAi8syXMVaCFZBqlH1712/Hu7hI0GWNkHGbaibVyp9yA4G9EF3kLdmoOjhQ2D
vYzuyy/UVKtSOUJRGvhyRgopVNy/CFL/ybFWrN374+KyC29T4XmILj40QnnMKlkHd9ekyCNz3L6e
R7RDv8wERdkS6E1pTtZ5oW529USMrYP34jyecfMekRxkpbkW/KwJyq3igOikpRiFJFuG+G4M5X4g
iTqlRNPMkkVsjU1cGGkpQgvGhTnSxTUn9kfmwUcj6b4MvBodRiK8iBE1osKAwTZpoVhcRV7HhP1O
stFKONCPqH5VfY8Ncw0W+sFRPaQmMhbnM9xic+oP6978iSbVmRGrVVML9ruPHMDHi3UZhRvvp67c
7fNZMXVxMK/6W1HwTTFLBMT2w2sR8C0fzcdzlSrlXhxf8A+1d+uyhUNQU/ZVH2CBnwfb2b2HUPLd
ffTgUO7GnQtDn1kUNPWkyCDUWcVGG7u8DOdYLFBs6Y63XSAM20A8jxNphilSoAA2r+PSnimAfN9O
BwCwPr1dGLh274zXGr5sUnOal7G+2BYYqQrwVnrd6wwRwUN4Sv9MNrVERng+PO/33K77oJ8KaSF4
jMf4ZFwlpjVfRsq4CmsPgCB3Sr+JZQGwrPh9HUtZ+7VpL6RkyZFQIZ40QWe2Gjuq+xh72otZPxKm
AWhxGmVNjGFtxxdaXijtYcz4dxL36KHY/jycg1q7eSNEFzwDAbUFGWDdOj9884qe7A9gA3s6F3Ew
63QAqX3VkwReL1AU3R7sgJrJ6Utwx/Aa87JvGsw+zSBVlaz1Xzr3sA6neemg9DgtotsZxFShaPTJ
SP01U0dIuZi3RSybTbZIea+g+Qm91ZlpVHhPq9/xdFaQgGsNAPlP2vHendlhN9PzAa2Vjpl0G6Ko
nIMmQCLgYBO7l8QDVYqWMAHDewGPOEp7hm74bCTJK9tvcofgRhKrip12UOdY5N0BPBkrFRsZ/3W6
MgeecJNdCB+BVHZz+8/Y0AWrtMjVYE7ifKMBQ5UCH2/p9AgbW80iwdUqFch2+8f2sxcjN0/DkQj8
ObI0a4YQ5viKWGo9VJqNGmzRQ7kUoeOy4cyaq/yKkKliA2WX9JbIkiy83Vlyi+7yd6qLOL8pbWxx
BDZBq1sKYPl0SBujZ3Bf8kpybzEF5v/kT0aQmQM/5X9ypb+enn5actJ8BMtX4l1+T3KUhBMeljKT
s+kF/v8vP8gYq41v0dX/lmoH3unBcBT6+AQHhWHCAZY99hFlee8FQUFU3v+vY2kNjPi6B1Gdp23s
fnK/U7Umt7IfiHro7/sjBGTvOdZDR036P4TqPIcXNAKa/Kq0PRN1WxbPHmvj8mmd8gjP31eLMQwY
Y4KhNPz1DNnO6XGkEwkMTIyigZkIC/wcC3ZddQ7SWqn/c9hNCx6W51ED3BScrupCIMetmz6lgJD3
JxTLj022SkdoWxPIqOhjghbvUXVHL5mHMU3QW4yIJGu2VPfMe9LRLBr/PW2Vt+Xv6wi5bfetuAm1
Nk7fBSANkIgxdJlCiMvcqNpeTpsF4ARt89+3Gm4Q7MIxBIVwvtphC0Jp1gOcAgbKlLtpdZQfX8Fw
3KMlJW0/j9ybzbgnyxGrk48+iB84OdwoPK3v8jdzRHpqgIbHdBJYthinNxPAL704XL4Se9AufGRG
lsZvKPNmVoHCTkVJsK4vDJ76iW2XzJcsZqkCxYifC+AJsD79iTY850W/tNipcnj1wenznIVvYeIW
MGNDEu7GKqZjQiJ95hySwCjEaN9xA8kw4Bz+KWPBNYbthDrK3y1F8yajHeAVnQFhJWMiHbGVEcsV
vVr5TX1SDGR/GhMdLgUGYqVWmQwKv4jt3SrvE77GLkKFrwM3ZHI1g5JtGbx42o6hNGDfuIihq+oK
8C/Kuh9kllLysynI1Mu+hKO9NFyGuWecfDckHZjy9BZYQuL+PbIOlJBWityB8Rl9IPZG+Xl1fznd
/lxGDIRYvUxtGan2r7vi3XUXboamVppak7xOO+Uvy+IdtsSkezUwkHCTMTLaW0aCSOws852rfhoR
ncyt2NMMAvx+1iZtTbD2d7D8YcrsbyEDmkT+ssyxcwSzNIHZ8zJU1+PFeW6Ab3mSLGj1QJ5Z9yhv
rCgFBmrXO7WYbYB5PeGRXkyh24HjbCPQS+T1LjukTE2/NAiMOIotzPEqX35WlNv6zrhckjBxPLI8
exGzxw/Q8atO3Ztqv5ziSwF0YmStbegzETcsED59VGc32XsGl6YB186Z7RZOdbt2ouxA5I8pAR85
Nx6pXvqVjmK8mrmI9DQI4XZwhG1eM9aRvAMNDm/G9Ijjz2P6mcU8Dnv6pFtB4Xi+1gFt3Ve5Ljvf
RceWfI/5orm5XjivcdElbaBqHsxjgwcC5p4EVhmJB7nduQJIwlMOJnzbRTMIv5Hfk+y4K46fVJiT
+8YSC1WibodkGqUGvKfVyjU1dmCWY5eed9cHxcSZGmgTWZOm7omCR8GQxXKsx2XsNpvL+JQwJ9ys
5Q1pImciduiPt5WHC+2wB8c/ZqN2k2AkpvAecB0QH7x0+DRA7j66zsUBAOPv8iJxd0FpW8XJEuPQ
TfriGGvgo8nO3AezuMpRKA+YH+LLMIDjHBRQYtLBq2zyFpkeDyZFUalDP4ljqOCqrZ8zNUlk7a4y
e9CxebDd/JQaZ/m7ya0SHSmhU9lNHo8u2a08YjA2wm0Jin8aFKhZQtarhod+cZ4Ats2v0VEldB/U
DJXv/pmn/Vrtb3OOKr+9rAObn/OI+4EV5zMvR+eE6wvrv2klqakEUByOT57uM8BJwBJ58cu4XgcG
CtjcCgBiV0wRMslNfAJ1FZKM15ExhqCg/6dumbdLqdzD7UnYSzsaaHvh8SJaffnD57WawqkExpZp
0s3yPrdZdnIk1PRz3HDUVPtF/uj5Z+4el79AI6iaPIixDz3bzq6Fte437Ibugjk9NfEgqb7BM1t9
5MGWkyKcJBGiFAd11+XyREFuJmC5s4XDTvM+lRr+JB89ExexFnWcD/mIdIeXCIRR2nVtfMPeERZQ
D7doilOX2ypkFhwXciDDYZurHwewIhBmVv1FBKOKOEEvYlv7nhVeBacHdJDAy0LIT4aQQhBkq41Z
8hWca5x+DhaHIj2gjzpQ5mr2giMobmQLcRnQ6IH5ePc80zgHzC5qpr6aOhojqNAUVtQKt58FYZFT
Zum44QuwZI5XzVIuopIvlIRlPH7snyMF8jvWHN3XAPL2jGqbIMNsWfSksqCaPtdzjKgXgRyodUFB
6v05wvunZ3o2tPyN2PcASpvbRlIefdfZ/UD8RSqsMiaSFUl/kFmBMD0N95DfjcZWZBoBQWmfMfuY
R6CAk+9E6VZC0eRQ6K+BCzzKDrr2fveY6cyg9UH6VmeIuOeBfU06+NljTMkSlHAGIJD86gugxDbD
M6cP/6fpQquctXeizH5MrNf5PUZs/Ipl3RHfrZz2PCGjr+lr6bBlVMqBYqhA4noKdKdknD56Ed/x
G4dWWyzPFgesFSv7Nn5b7LxJCKqTovH7QoB+5K4/PKdcZuJz9uBfy38ZKgV/hyws8UkEkgUyajLp
SlwQspJpAJnrStqVrM8rsCAynAWQ1FPpFxLXDWFF+QizFshcnTqtvZ93x6NrVdCU8YwtTOMWGXaN
jxr98L6L6gdpsIVJGYw2U3HvOxFxzId37Jn+1eDnD1y84udftcbhzI8QpM10Asz+AB7v7mJOx8NE
1mDOa/IdYcF+iBrtB9igZ/CWjO2pc0N6i4J9EzgvmcwFBy7+/DDjvNA47DI4k/tr3qk33G1svq2E
GH+HuUr/Lmv2/rhDJJplLEWlGZVtFZqJTiPibb7YaFF3DuI+MGAE9Zc1l/sTwJrGOZTdztMg9qqz
w7FCqiKFqYt15zOozLI85jRdxhED25AH+75YOrcJpN3t9HOA2lOxW6h7b7QZd8h1FHSFiWNKOw0a
/o6A8KVu84p/ctRuTV0YLLNxRRtPmwRCwTEX5uodeSTz9dioYKnpqPfxrynPbC5TmxKcGjx8FKP2
rtQmf1SQqMG/DFkHlnmtpyPEiReHYv0M4Lz8lX4RHSgiQClJeXzC0VfOOXZvrKIPC0UiaWZ7tCB6
jPzmX6VJZ+Kk4RnH+aFy1xyEHzRIOx6rEzAeiR1YL5YWNnP66eGK4eJ4UBoiLR5I2SfBo92zTQZ+
Hr6RYtBl/QdRXZnIqTMp7i0YrXtrrU62e1vFSNk5PxxeVjIpvwmbicPKYAaHZsrVnSXvHHg6G8GH
+8hk08zLtcPuBrBuQ5hsApq2i1HfHIJIkUeIx/XgEQJDtyIML6+4jmzyBhM4xs1YHa65GyK0xiHA
cad76Z75550NU2OXleR9aKtG60T9z52VLgSYoTU0OvZxwj2Pzn1BNwG1R+RDAF5yPC2qDvQ9gA0m
v6uLdbhwR474mwt6gEKAxSr1rN1/GBxdh7EXB5W7M2KyZ3eABt7OYWdw7oBcW5D1IDBpzQivatWU
ReheO/m3TwqLmfYwJQQVYIUIB7VQW0VWtZ0KFySu1ZRWcOtLqzmytJYt76ea+ps+V/UGcp1dg+1s
EP/1Ovc/lO65eYEXmQkxHnLXjD01rXzVrroffLm7bQnJrjAKnBr2CZLrseHTFjK2QQPuGECOKF86
F2tE7yGL/2zCkN9JXt/6hnmD/PDddQmYRiOW6Uu3Yx7tvz/QXJJdWD4xgHVwym6SjhMCNKVMZOwD
GdCg+1DtNI1cMv6268vBV/xbJMKLYoVX/+1BwtQwJ+LtcPwdICH7azYH6ymu23+9nmoPczlnO/8b
VKHrPqx4T+E8DdVQDVPYugp/6A6Z/Qh/h5VO+yLf0WpjLMMG07OOOnYXW/TUO3YCsIBNn7WbmW9x
L3FAdCL+c127UF0kiEiptQgMshigyUB9NzrK6RxIrszs2hqubMykjIxdK8zIFxEFFbqkvqhe1a0g
9WwUXeEqWrxajdUaJm4QTuBhd0jO0U1RJWCrxfg2bUDvC2MgY/l3SluySIxf5w0E5ROPQPllXKjG
t3ceZf45RPFqiWbevgUn3vryo6n/8MdcyGMJjXmNE+QNFmHBLWlDlehsdXC040j6MfFBpk3306ET
wCEXjT0Fe3vfMVFRvPEp0JKDAfU/7j7aPzO9zcAIwGCngTWHSFgSDYEgmbZ5eopimv0dEdlthxqy
GF33fAzM7FiKxglm7S7Uml4ttLSLMcFsfoSXaATuESOoO8x8rdOLp2z6JvjaZqUaltHnV2WqElpo
nYmgeK/HMFRQpglYhWHCqmsDHnt61U8ZF31WiB3EQ4A8xTnREkFLf+jsryAQV0bO7hfI0ILcFVSb
WnboQvPLTa9g8pa13lWsWCuHsODFHYWrNhBHgxOHlbL7h4FLZCfCN87KWQETX3Hxaw70RhxuZzDl
Mzzkcbo8o434miH5ANp/zEFVGmZ/vrkHZeY0a7xumW0QB36oSwd+yotbQm/XsjQ99utyA0lUeofI
o+rs8+o3ELg0iYYlCrE44/3gDRDvSABO9ZC0GdyZ42ykkA0J8jf2p3TUGK1MxDE5Pc0VzF2fXXQ+
nKif8/OP4mUWnNdHkuSo6RghCoa7F1MvNuXSfAAjpQ5Asj/rTlz+yjaQ2wlJALHXp/2ArxPMYsoH
DqfY+IZ47XhSaZMvq43ZH+Sc4Bk3eApCzONgEoA2Gg+F8KfJfhtPjDIaDiBRS7z/LfHu8pLl3uR6
vrR6YH+KDbzw6eBqCWx1y/hmXgyM+5OgnzcAL7kN8Vg/WHo6ZDRrCy3Pox5ajITEnLoaUlFO9PKN
UVOw+YBHFnl3PVN8x84Vq8YI6kt0Pbo/Oah/rHkYp8ySnr73VFepj5SrEX2PJD3w8YS5hkBqXFtQ
F6WdCBlKwIpfNUqnC/O6MyO48PvXjb2WT7Nxo++nmHF0+N6lLDwnYaytgYHBDFi6aCKBoqC1t/VX
sYvLJO09+pNXHwE2hzHdrt4ID1npH6+8Y1Q7zEixDRyrRBL/Q/dL9tLNVS996rnucoJQyrUuSf9x
nGL2zCoutRxmqPE8OweNZg+3JK7ohjZPRZJTde51BQEdy0V1HW9XsMxTwpTBmGdq452rgqbxGSYT
7dwuNkpywBS20w+3Uq//hJIfhRf/VHfNZ3xPBsB247MD22/n203JoFzVaPWbdIIVWucz+WIm8jSB
Rv8Vbj9maxocnQnU3ikXsCJzvy4kEoNVBaTOuEQfhBZCjXP/ZlSumXbzJ6yXvl4LGuka8S2AyFAg
0B56ah6NmqxfGHG6Z5Xs45yzz2BrqVXYUBIbmRYBi9GVZoWZO3hzM9OkdD/zVX6LfbSRCM0YzzWw
zkUzl4pOEwfdDPABkHJhNjPXiDrOr+/+lSGO+3VPOtE1ILs117dXxHQ/4RH3z2cJs9BRL2Uqm2k9
JwkbaLn3vGvTvcPux5rJF5gBJ+vJ3hXzkmA6L/rWW2A89hSWxjz7lkEhSJ0gVhsiWr+te58Wf4R0
BZs4swbjKg+QneN3V8BYo2LueBvuhr5WPFfpKmv0yjRQvystkk3b7dVPjnF+qKYVuPhvHngLfgj7
u90zGYfF6bk4IAtt2u9ZqQxoc3HeFtrNh5GbIb1rlEWTB9sGCRLnXPxPI1u4YN4mo5Bcs7iwYGQs
4lPfUMrm9l1VNP0tVH5mz0dzrtM+z08HazNMB5y7QYuPQYNJR4ommGUR+ZZ9pYHlKGnfX4EYZS/D
No+wTWbbC+LrgaX9Od4o0UlOU8zx0h4Vz3uxUlV7PTpSf4kY0lnkj/9then5RxYcoeW4QvcRiRAt
JrSikDFNZcoR0mmPWChq9qVn0X4PJ0DpoSeTi9JG2/TbW5HMBhUp9SaAprQCWusrzoQaPRvZTEMa
aQwKMcmw9NtDi2lXTIsn+nTFS10BzaXoihNoYIVDJHbLS3tCSGfxcbGZmPtGVMsxyn0kA8Jk4T9P
ob0ZYlWWnRyGEmQnBVvzv8PabQ1cd3/qbTdrEiMZDbyo3kFr0SVUuElDHZv7x9tTIiEkRkizh+Km
dlbZWpbFTgNhO9jNzG8lWw/jUtR0c241Tk6ls1cmZJK7gpAEcs2fAXQkZe9EnEyde+K9xJ+GkPnL
b8hFrENf2kQPEBzuay39KFIlfvfa9/4LYINtY2cEAjveXgiTiwurPO4zqI6BfAll0THsISTROXmq
QxW7vpWDXkGScQRMmEPuybHi+rY/MwP6eOEVwy9E2UOFYZdZEDMU7L334qaAKGKU5g9s2/OB5uES
UQWjO8PGeUSKlZ2laUGCPpHhiof7GmMfnGybej5GNqp/ynHl+uVWQoIQhiRtAoyE2VPKnV7iPSXU
czhKU0+CI4ERZE0EQUUQ70NZS6T7cap/ZUcW1yiIJpAJ92psPWSc/zNx4bg6me0Puhkpjufb8Em5
YApMY031gVS8MZUWfuLhFpWCcs7uQhqk2qzc71eNkkOUA27yXUvopkmUV/X+FasUmi0mP92A33Ty
7n45GHp+Zs4CTv7Ien9RFhj4gEZQAqkYzPwRAR3Qf6tgeRtTJsT82X4botnQ+XYMgXRQLjTIKlII
SFobyNwhVgxhVsnPjlMcc2T6xQo7AdnZe+2LfDt/eXIHLhHQIDzq0acDEj2W6aENYtLWnJZlNKmC
UVT8n5zOLFb3Dgo6uytSEnVeI5oo38MpQGYR8c5Fkxe2YZS7qDd6gvWjBVAcmbr6tXWv2CwvM4zM
CmJ46ZWCXzSnWa3yiVEdum2+v5XQJjIMXCO+7o33ub25kNJx8iA+2odkeBUEcq3lIDXQBJFCaAOT
MkgcxcLicG2/mR/5tMGHzvBpAz6FClK6nsEEhjVIJ5+/Hq/5/zOYvPRc8C7pz3NTCOoOeL1MsyPj
tRfCCUEnQmFf/hvuocSmoLRtFDZZyfk7ZrSthr/Cye0HX0uatjsbX4ohyzG0f2XTML9W6EvV+/Bb
NFw7IYjTX70PNNakao6UBNZNiT7VK01FtTBs+jtJ2i/avkLg2IbuNKoPl2e1n5oSrYwuHADoqshW
TjBi18R3S7X2HMv2ZiLgNL6qnMHqC3xAyIK8HqfL642BsSoFR3U1PWiwlJBUiDZFwozGM1c5jBNg
YCJvZCzNYo7tqf24S6ZU3c1sPI9upf9RIg4lsmLum+kLnFtYr+yi04hlkYbAkHYueF08QLOdnJzt
Z0PZoU+JCE6GZ1jIJAB6aA2b3SNHMd2ZIqxW7osbhaKgni127VQRug3QIbFAVqoqnQIbpRf2kUNI
hR3SmhchjkfPsHvgcZ3dVp87WHsO9ntDYv2ChHcNUYxRy0/g5gdDNFy1XEYtCRtW6xDJ8STxV2An
Bj4kd9wvYZLiLY914e1roEJBs8TeJu8qbDEoHVl5mi1mBpODM6EqXhRVGQ4IA5paZVGRHdfgAd06
KGbwWbhLIH2NLvtS148U8WcCuGLSW5nKzCfuryr53XoBywxPxs+837DJz1ZAm6FE8j4l1Y/f96km
pmAA9AJuWdrFqah876kREPIAx55qGacrRIU+eRQ7U/uTzK+b1fh15IBWMGDLYF9KvhIAhwjzUUUQ
Fnpzu/NBTZLoH+MzsAJ/lwRM/DYDd+ItdCRYFSJJXzL01ugJOmY1t64fxPJr8/c+0mF2Q6tXDwqr
UviLkdi7aBuzJoe+I0nbFwhdi2Dg2E/bIG+LMl8kwN80Hrygv5qPsAxBLyflerCyf6VNcyyr/Xbk
ImybYopP54Reaxg8X8gOB+t1yAM4MrZrVXw2JuFqc3WHBllJ3Y+ZFGzkY1H6fK6WBrkAHjHug0h+
IoXXa0YVKBgvRA8XZOjoHeQu3N/+J7mHx0Js7c3kZgM7cghLTyImbkKGKh5XwRM4HpmN/ghhdEGJ
Q55KK9G2jAuj98+5UAl90dI8zBn5jw/x1uDQA6MG/4y0wWEbVVgB3HjNiskW2KX0WQkh+d2rhDTz
5m3eW/T0DuVH+K4Dpo/p7fHhlIPUuhqWTLDP2pHmy8VilSpYPdO1f8h4s64lQhEJHOLK+DjnJjLE
h0RH4E/lvxjENXOr7Podt3NStQmKS7rUs0zHafrvGkBcP3OqqN7PeJgoA6R5dSSpwXMZ3k2lILUO
qKZNa6IA9h4Nios3sv/syH3kzxpcaYsTvolvwH6aL0BFm71jlwoOFGU5osvncKjK81uzsRytsPBf
47IHC2Tzgws6wRvPYhw18cVqNmbdAW7sDSjsZFkectzBWD5Wd/8TZ/lZWMU6uhqMDT0MA1lRHF88
OMGewJN4I3A0tKanUdVF8vlLf1mi/ZzpeCDCS27nuqpbhXktEyKn3UQdMeZ3qrxj5lGv3+A4X/4f
jwBbJDAXQpVbaBCANXjsWPCX3tfkMRrn2hFR1qZP7fpTge5NyVP177gcBVYKT104cVcGLk70zAgF
LurHfbGjc4wOkuyv79CMJmHVguID2/TEGLwH58+go56/Pss5F+5+FTWV61CRSqwKEvDpDXQ+i5FA
czN7CYDitf4A/pmvXlhsAlXhgGHxjW0JQARPVqt3dfXC4A6r5vLv2n0A09W87at/6b/GprKY/yqe
2PGvHjnNihhHK7IpZsxgbWVSB1jyGplTlQZcMpYeSFu+QRj1pO0Qt3Jey1KbArBTkHTWxRzizH2H
C/WiGI0jEwuSQVzZ4d07C1CXR9JMu9gYHs/DEI02yuKrRkG79MEb4I50oVe3WMo86dqt2UMvoApz
B7JPvBv8veupA9MOvD9MAJg3+9pG4dMZPunjCqC7unepgdRmnQSBtol5ZJ/khsK9zW/iZoszZc1L
AOvaF9xXVBzLc2UCnODYW7zk62m834A+NmIwSqjeWsqT3Gcjc4jANFJFUTbkf9EBbh8DAZM/u3Vj
jQoyRtrpTcF/D2x1YGCYo6/ud2J0mg1gJO2IasC9QDa8PgH44GDeap/MaEtI0wgHiymHvNTalYxs
aiHehS4gY9QFkmOBmhWsjZYHZ5NbucI0hnJ+04WbszT0/zDjMkhehCzBCYo/FPe1DEAqvKWOkBqc
pyIWjAreUOs6Sx0sl5SKsJP2OeoCRLz+hsOb7nPGKG4L8Sa+foKyOU+kIyU+tBQgJQ6/QN3hE2yt
l2fL57SuCJol1D96yMnB8awgnEfgSAGEYmaypegb2J3jcKWaVCZiBxkSPtPsIxJhDlzfHBAqoluQ
irvEmCIKgWbgSIcdtCRKLPciAiBma6DB4rGWXVMoArhs/iOfIK7vNmi8768cRDAd4syOsIAaZv5H
7+tElDLjzdFF7pysoRJZ3Gh8lHMg+MsMJXVsnN/R4guMiSBA4dCuctKx+hejjCMUIlOB7F93wjIs
wLKePKXCPaLxqWFYux+TFOWR6QHi7M2NHD0wAV+khti0AZzMSVs7xMOglYkPXLT2Kkw22PymgpEP
ypNX0PId7CkhlQeGPGoUAqIdRuqlCrgrU9TwfaMr9onLY02+z520ML6PqW8+ftuUxMGuLG/Z6ZdD
8LsewZIqxolRQkj6xj0CSuIL+jB8/XE7XnrlZ+asbKi/xJPcM1ZrV80Q3FxYySpUibNBqMkTejGI
AJeLTk8TV3KGUsIK6C6IBnUjZm61VkyNQN5xCEyzGsHCR6Oib2rh8TRVSHufWJF9xMGcxGVgz1Yb
GyqRMxSpiWBEAp+Z0mf1fyxeby89VcX3ZOd7dn3krQFP6vW5JblEfqOfHng5FGE04lmzehOTcNme
RESIpmdf42F7r13g/RQmcgaKD41dJSLJE9rIGq4lyxqmJgKqmQmd0c2AHivC8hPcdlrla+PG6XJl
Ep9jlaTFWb8tGn2oRNrpVPiNmB4kof4fAGLeQQrAgw0YDoy9ePh/ss3kJqOoR5asyyvrLBj8uy8/
MdrntxnZF4Ee4yvbIj+4UAo5y23AI0TtBgUFAln3h8o4QFeI0LU4tpjoYO64lvt1fMiEJaDsqFDC
bsUaprPGRFby7JnutzoC39BQzLadEkspkCow0KPQ/VH8VWYMGsGskZ4S4WlBENKOT3l6znQ3uIjy
XcdTiPQaygv9Ri4YrpAkhph0zAgVc4ipjccGysJoTvP/WETjAPF8VRI0zC13EwLGFekl1LwPpIWZ
2qp/ewFWSczfQqYH62xDrop1JN7N5ior2Xc0fdKBeYr6uCeVRA+KcwjiyLGnrzEVbcqUCnRxJhUd
V/Kjvh1fQuAN7KtvuP5RoYFZ1l9adR1ujuCLFUl2gUmcTJw0W6kDCqFdd4p2p+w8GimNfhk+QAWM
gWvx+iqrv91e30bETIQUHP3tFaWCp7EY6b9t0vqaMQ6XVGVamTGfgpVNibWc8VbYMEr/tj/Ffrvw
+Fa7PPWQA1jO6HOUo/xnX8vPVIFiTuFuONCq6OIr4Tyzw8l7pAleMaJBnUkMqAGcvaAbKAKMbnaj
CY2xA7twwECTFFbna+BcU1Du3kLSqljrmbvL1AHokAxXnFWRE/nN7nBfEPqyRtwVLnIi3Re2xsRO
wBqhC+luuuzDK+9BWb+F/Mc5ci0/YdegQ6blT4pVcfZLxRXUaJTUGQ8qZxZ38qwjHHfBewkM3DSW
rJyrPL+yaZGKZL6jFUB0K5jxEIHCYiD+QBts52iKgaLms8rVufNh+l1HQtgtr5A38GAmhzi3N7gT
Oi1In4gqvCDQ8ES6dkWXNjWnpqOa1B/tWvXIFa8z2gRhtz2csZcyEaHdGskEl01sWFTutUDBGnM+
ehGgXZCZUjfyEGk6hLqJ1CzyM3VRG84OvmkBeucYnga6z7gUYsN6bF+28LIJfRBq7VyZQAPiFkE4
wAyj7m5qbPY/47oxCdRDStTjdnlWg2Pt8CBcztKoKLygXw6cVlnCBE2MeI/z8hssjfckxT9WC43m
zr3oJ/szKVga8oa4XI/5tQBpAEQIg+1JWfK8Y63YRS5TaHs+/+6O/2u49oci9DkOMTt5dDFt22B1
rYDSOy1caCllUidIKihkN6GwnB2g354LAmqum4C1fqs6y6awGgDgdn65svodUX9P+JarXudHzBlx
buvK+Dryze2gYhc/h4M/ZbCrQpETFVhwbzZy28I70bUziiEjnHk4BnKPuWV7sdF8rgTETjwYYAtI
Er17iMXBvgoVdrjFWkj0HgNMw/RBOWkvn9cs2ifUMCtLoUbgAcLolqzXjNX565KTtF0qsVw1oYu6
Lf9SoEruKun0+isZinWLMQ4BDktNSGb72c1hdlXgXrO22bws7idmI5YQ4yF1G3vMZxCHkzamszPt
BGywNdQeF8val74se0EuTh9iBGos02k/wEzW1/kCmGAqwspJAWMIqngecnhdk7UEhNAUjBJ/hor4
DVqQzJt3Uq4MQtyw3fqCprJI+ynfmJX43jX/Od/ktjYe1uthU/TbK6hsaBsN0to5BGkYqPNlwhkY
V4r+hzjBMEwFiiEidYraxrCcjMI55LQphNVDcvdq3+qP/wPls0EUM30clqFACg3uCPITjIczUmYK
LSvwcVwzTsOGNE/DXPliIxbj4G/oLObGbRlLOY2/nQ7m2lSgfeL1TRidDD/UDjDArooupLA1b9Eh
gY+0kxXN0hktgq0BZfEBy20qWBs+CKZ9oRMh2+IaasrJ19L/93/UO2GvOwVOErsLsw8AES6adkGz
HrTnKHt7mpk/MR2eleRt6H4fnSqT86e0xRMNqN0AuHg0WQ5yMu7XaMdPLJi9J75YQUE9MwUCZgNe
pPG1NUuclPCCJdEj/gEhL9dLHRGsJkT+sHxjmiLrHo7ecASnHBFQjogAc2jDA0S1HQOR+FKoPSd8
cDqMKgiAYOutYceLwrDGtB6SpCFBRm2CB4Wo4X7yXMvBkZ9ZstHlMYtXPa8krLp3QQvk0st9e9/k
x/gzg6QIj9YIsK/aADVPcBbzaduQCutcN73U6bgGIT90eNPC8JmvZkr946Guy1AQC8Bj9+8DtaAw
Us4eEtJk2uFCU+TUeyby/pcL1wuIaGvNxZRBK+JoSQa+jraDeqcFntaoY343goZx2IGOjm6mi0QZ
i7mYUsCxucvbjo2TtFjUEzNBXteOEjj44QKatMAaJRAo/wFKzdhLDr+WkhZ1IixDWyYLL8f/uCRd
RwU4SQlyEvpfT02e+D2O1gD/ANHM/XcpsIGnrpaG2mHzZh1W2Gs2QKkw8Jm8RX4/VK9FHU6jzVuv
pMCeoHhJQ1dJ3+1iV9xgepB8GMOu6beZzBtkv24aNuoYP7Cnx4AdpPCOgGqadH3eBtNQvX1kkude
Vpj/X1i3+9DvDWmMwIhVPbAxarccE1NdYupdyHs93mAllGif9kObgbfiXrX2izKbsqs5bblfanjh
bYToQZlOCUlQcsHmITaLORn0hCDuzC6AA1SXM89K1kNz/5cOMVZe8rB8s1z9Yw0NQs7XcLnJBPNA
hA12ZBYIQFDEbhWBl8ozI5wSdXlIjdxMasTzo8/AEfZTP2syUQtF2qGeDrqZ2ABTmjiEk70k+k+g
BfNwr+FMqQ80YrqdCKv9lEVXANaqn009sJsZbdtQRccPJ6uDqmy/poZsQ8XKDKaUn0y4FxpM83F8
pYXrDoAIJ+nFIQMIhFSaT+ws15GKf41Zg4Gp7e5Nm4FwYtb1FXZl0cD0RGZwW5wXZjoNFrhHt/E9
xoHtA+ZzRBe6aTKzYu90e9wExLkZqvLWu3EJsUt60rpCgL/Zjr/eBztJ8Y1t5BFWygZCTNesCYLw
AnWtYXEiIFo3CIOLCGQPefqghjcb80ICBkgKiHPVUYUQ2TvOZWAA77FN/bt+KzUZNICG+MsSTICJ
4A4k7TP7NwoC9q3/NS+BAcFVD5uDVrVqXZD1ejZTGpom2prdZvji8UwhklPxyhcd5vjfCaoIuvNK
CSgQluP3GHFrjR374T+az8LEB7vHGR9v+DbVGt9yNA2JikjoAp4SvmDIwmeFvwjz8GRIInTE6n9F
auHlk1wcoTj5Fa9+aqvgqXzJUofUfzkClPZKBDTLqsFT6UsR01Bj9zrkXV/Kj/p1m/sf8yikU/3N
ruU4NNBH7kYcHDLZJObXwuFR92pkjUZGfv0OECfUj5FVEWPXz0MVSyqDyZSKt6K4g9rK4rkDuNs2
fl1Qbks15ERcCHqSiuvocPoNVI3TdGoCsc/KfAgwWXT0hS/Ve/FT4Si9+zuP1qWqaf5IZ27gR5gT
wzDJ3vLB9r8ZLEFbPxDJL2WdUrRUAD9CdEMQDmAFukcQXjLNQZi1p4bO/W8pqKw6KPebWewf9d36
mIWtERFR5jFhTPkdWXxWkgPZGPhI5OjISK0OFGqNmbitrltDK3D9PZLJJCuOaG07kN2zeV5fRPd5
FAJguL9hMa8i6TPpnDaPc+urdhmv5UneDom5NVvbQgKuPy9k/wdGOzujSE3/eNqknp2MHJgfwLR3
Whu46TVPvGy97T1/M8moHm+8ACLMurQ7YNpHuaM5fvNTcQGRKY7O6yC3eYtO+5+FDoc4ohBHd09B
uISvVELwj8U+jrlhOES1Yx2s5yFPcmpAQCjp/ZCl12hnDvEnnm7EOGZXXX5Qu+tB+sBt9MV/1HBR
rgNGlsntgJuN8GBxJj1J3GsQrk2quKBciptoK9bgfVPbKqrxcER70YhfIIg+cSZHrNTKIrPGD7Tw
PK29xqtB+FM50WMF+k3joUblSy3L8YsfP65zFLZk5mUHqgA1W0eWhhY0lXwdDG2ly2vdmI6/hkO8
L/gg7baaYKaX+1YV/ZlxxwOmEvNFAY55rM+dehe7wGJJtenxMqcq3tiIlswNRZc8jKgYsqW6APJK
n1XbV/Gb0plutquYXmY8q3bAO2ZxE81hRqOYZDAV3wz7BCxqZzSYWUJaJj5wzVmrSplfUyh7chLt
HpfvMS6cqPqnAUF56yFIjR1F1JoDlbHu4N1mxGOIpfi4FaLs8Tam6Ylg5KPjN888/5keLS4T98Bl
w7xiIecvNBENfTXH4ydFSY9HJiSnwo6KiDvchO30+cQqBSIP8yu/jaCaRtkxXfCz7GSvZzye0cvZ
NKCBOu1tYpwxhIAQs9yprOsE+PEHthpZzU8hagYA3gJYuNvd8VyNmVAAYI6grNuA9k5KlTFTtqS3
t/2Wd6lAOpgd3gtIlTuDhNlC+AJ37boYe0r8Bm3jt40orPnockyS/xiYWnEWEqKoMyEieaQHkV2Q
/HJGJrb9cUJnXRGykTXFFnn78xU0QxnESh4+vTSOQsLwiqPERX7734g+Cje19+SELhr0QeQPPkGU
IvJgyIDui+r3kcbse+EdiOpbUv0D0g5VtTaBfS/thRDeUCavSDOO0HhWuY3aihI5HO3aJTrhmck9
R3AK9DGKC+aFCTnhQj989KH7ZkixiQxZ2X/TQl9TTLiK/QuAB6FJ+8dRy9cnT4ICN6E+lzAfLCrY
aYSfyxa4H2JD1Fb9+A3yVhzkRgm5+tfrIenwvejc/pbza6tgewri5appbTVU6HSwaFyqgJ0g1rGx
UTEeTiPtil6cboErH7ftBIHqBQHoxfmCIMwflfGglJrjyk4wlo5IXhjNGx/7mIBpRg45HvXI6ACx
/FVwUf2nz8KGp++7E+lnPFwsAEmpVfC+tnRiKzHr6pKQP27Vvm1TxV9IjVrLFMxt5JjF2wPANFzW
w2A2V1suJj7JeGWUPnVkFkfJ4j0cZIHOjbSN6Sx5KArDUBBpl1FFx/AnoigvjaDkbsWH9KwNHYHt
1TtEGgpV5XXjEr+2KgCAGK5RR7CmEg9+uwr8aKdStR6mCeT/qWUgmfhTZUm9emRkhLzajrPEt3IV
Vckv5+9JpPPam7Orm2EHyHNDG4CXCp2mIaco/Q4cV24lDs3+Df2ODPL64bxSKMQ9eQlCrFgnqrIB
qTNje43f+EJJN8JnadHdLepd/XNgVhNFa8gky+2+rJtA4pmslTQ1FdySG/VTXQdceJd6nang9clI
/mMiXHQDmdabrHbw7rQtpTKjZ8K2aPcKrmceBZuFt1E0v80RCbxRQuqPAsWh/MqxxHyHbeJwXUHP
GQTBIEFkRQgZXtGhvRXymIcO4v8Jc4A4HtI0py1ct7Sk/fvbyMs6aug/qUkzg/+J5610bh6z02wF
86kadSmPpDhnCOmzAcsJUXtjQmTCxjYY7pFniHGFA9E6DJW2vUtaZ4PcXUz6AOXDA5z8pOcRNZef
7wjex2yg44NUpBwotlZAmO3GSqHglM+luXSwu0ha92ekamaUCimTfHWh1BQwWeBgaS2VejFDJkGn
XgSJoZEFbsePGsQFry7D9dP3Eg6lpGyIO3wZhZxuGwIQBcaw9rJ0869pFdvJSJRu/dbJ2c2HEeGz
VbUGYIip10VVvyOqDH42gIT3HHg1uQDvrV0sQaxsf1HlQCaAAvdBLHUviWRIFMr6vFMRgDEe27gs
URxOZoiwvjKpy3qe9ae8hjfZ+aJXy2ZRZaBsKrg2QdPediPjTEvwBvd6xI+kLyQJCyvPUjAAcSYT
H42PKp6RTf8OSFHzucl7vh5ocBNb6+roPkGqZ1Kh+twoccVLzX5jvLbaxldqOpOkA/LH0/vF7nH3
rSgNUzMoKayUEdGb18amXRO+sEf9vhN39KaSDDrY4pT72Q/x76WA7Q5kBS0deKL7OHZ/E/wCgY1z
4NS9223JAWnAR5omMcf5OmeH0M1Z9551xeHLMWjs3eWC7hXz4/+/goYr5S/CoJRjTNuRFq8APlo7
rrq0dbeMWLm1vqi3MRenZPokdAzvZzk1sZDXL2KFvZR3cwKQHLIvcgbVnx9hf+LYn+V9XgVttHYs
i7Izf6+3+Zu2n4o+4fzXjDUIIYke0kgqmJM1FB4+wqGbZ5Svx8q6aFDImysLYQeWMLIxA8HT9MMY
NhkhVopbTLypPLhizynpCUQYQMB0V3Qx7ADh/NO6rucmYikD6U1FzR6vbyal2WsHXbamm3xX6kFs
GFPDHxd4ioZhwe2k/FRi5CerKsL8M0OSg3aH8yu4EM7OZhgklSs3AYyFjNGvJwJBfsqb5UIVp84m
faUMF5b4SY+EbKdXhgCjh1pTCOnrPw/Afe32WwjYiRiP8+hp0pN/Kd/NJV5xSJUZXluTakQ/xuXx
VFmuHYQkGyj4cbDPAQAMKlOaQsp4749vTMBeaEnCV/EFWKLBHe4dBIFggV8ZPrHWTlJZVgxwXmyW
6xdzBSADpsXytbcAyOgMN9c7pqVCDFDtvTMEJUsgU3vQLyIGXdmOfgDswnqo9OLq4juK1PZJ8D4/
Ebv0eBTUn5Ae9NDr7Ps/s7qFTsN3e4R54Q5eyESQUQcLnrk4XcqI9gS8F3qEcERLC/jrTnKlc/x7
xmOf6QidiaOtagTihVfd66ALARE+qzMTDnmzVFWNYehuFe4GHB86ygGFnQINVoi85gBYptZLuxeQ
7ziBa542Y2M/s7lltcT0rBAyFPEomWHxLaxVw7qHLY8Xg7U5T/iGtqoBpw8MkjCbl0RcXhzg4Bi5
lL+1GTZBBjmXrkJ00V16xFlVHxA2jPmdau7HvIe9mtBYesBZAzMxWTd9OUAcCt9oaT/e5g6jWpQF
19FR+C7pu71mDXJ+ZVlN9ibKSO5idMHKrNwVEqm24NTGrYSAaxAylifZ2X/ROjiIFIhSDq2LyFa7
8LC2D3N42fnCD/O2zlvdcaofgDnFjVK1tjffJZ7+HvYVphFYmbSmTvDND9ccxK/OApCTd39smNxs
WQ/FYqACYjFiWq1f7/r9n+ccEXOYF0p+7FNdOFjgeLexv7H+25xkPqVJnMmiXH8HClfz0mjFA2bY
3bvvvNhsykru9G7qM4pkY1uM10zGwk3KoHWfXc5BXAHBmmhsJPM2ZxcEnF9kL1WqiMp3zEbRK0v0
mg76R75bWsHxXhgBIph2ML7U8MI6MbOMBejRlrXVQ+DgpblL46xV/lGMLuOpu9QLcYUbyhwXrRe6
gH0IDXwlepxqHXF9CpJ6v9wajQFMERlZ8gkE2TGPX4ErklguUcnjoc+8HR6AFPN5+qjdsk92n4/3
ddZ3Y7fxaF2/7A6Y3L8v98e7434iMmlGvSQPJ1lyfDBN+tY3ngkPCkCaDNiqQn2eX1sIPG0FeeQX
j+PtNUaMh0DuF8nF3Beu5bse8NGK/HRTB400YIO47OGU7c/V7G2awIQnY5J1wAcCNpMV8MdnJfWq
WLKHunRCqq8vVI/lIhQvvDeXVrKb6ogIrE3jKpDprxWP43V7CGq2OXv0oCLNdmpOu4r/hW+BXJl1
1L9rEMugMjlONoNpdkvwgVIh+gQTIMP2s7/4OZBsjjD03ZCGnIyMe/gjxUU3qc64kzsIy6JtrE1x
B+B+AWfuaM2r4Tj0prZ4RuUZzk+kL4IBIOGcRtqeUUd5oQasUtECeZBSZwZsIAVD27UzHFjqJTRb
jd7mE5uHXEwzn2bPN7btUD+9AjAtx+sqm6g2SN+xRVPlYyB0qKzBOsFIm9CZh3lvZ6sgrTzhAk31
amOKx8tzVq7f4vzATzfgWmGUmDj1ycorPdtgFhvsqyrBvh+7SvMplzP/o53KXjXAB6rU6r+BBuww
yqs4vvmIno9MV6HgSRY1QojkFkIr/A/vAELLWisd7O/P59Xvs9EQeRisHhup3SZ/rGzctVfa8EqG
Hd1ec8gLynXxLuPre5haQU5EXNxZg2zxFKWjTImLOWMRLYnmovAkiQg5Zalga3ZcGlKY+UiPDntq
NGFUtDI3EtOgfpTj0c+QWwybidTfU+TkcvV10kyQCkn8hChdysnuURrVP2kzA5twl6SwA2kpuTMe
by3gHoh4Qu36X+h4+kkkGURthpo4H+CCzIBFF3C6UrQTulC3ysTluBHtGu5G7Uc5bGVpjBWgzBI2
h3AaOxU6aEfBv3wspxGExQr5j0NFtW84AzNjtef9UAThQyWByglurP6VTBuXfTBjUPkgP8FXpFTz
pt4jtMojPN7qz0hfMQ1Q7WEK+f8DCxkUiauigTTKpBiS4/MgELJXk8O3604dlVclpXNuM59liiOi
HqPeYOTdXztyuruSs9RWL8ArwY4uYEy/PJetyi3AMfJB8SsJgD06Vrb8pv5b9/q3Bdf3wdaua471
1uh3hNEUg2HyfBPZh36RpC1twjsUTZabzL5kbY/vtzUt5o/BP/eV3WKC9f0/IC23ScrQj77Plbcg
zgHMcleg5QhaapZ0VYCfuucmLADwBbOC6LAkxSnqCho/sflNdPJaQt6+K7bJk1omnwpz0vRLXx0e
AtCoRKPBiMY1CYMUA8nsKdCUe4OvJ1VtFNBOM8Uq1OtBOni6oFLUTyVIB50CbDq0MWtfGUhxbqPX
PJgVmAIV/AKSyvoaNIfnzSbFQ3ciWutS9amk9Pp73W8a6HR+bB/p0Bw6OtSl6pv5yWpJ+sVQzcLN
mJGi9NJLh2rU+Zse1e/64KQPw6CaMyATI9tS0fw3bDExF3SPDXdkKhmcN0oM8+fWs0emwV/R5JH+
Cwu05X88IwbcQ2+mJTG1w+YQ5CJWayOEJJlPCuCYwlk9J5lYHD8td+3Dx8Nb+zGK03PEm6woTeqM
re1L5kdrQQW/U7xqjeAlOAZq/kQlET93xUiazFHM229J85KlKLSxL3R9ywER/xES/kcUtnQC63jd
HC95Bft7SKdoUPck6iwmDiny5Ao1lhaxNwJ+Keag+OYc8SNlcERG80QsHv3yCMjEf4ZtO7CnN+vN
StyfhEFJpCzG4DC+XBjP1WdlZAYX1GD7Okhgw12+QISW/OHEkAzN+H834GXgbDvmlOpPvIKFHoXP
ZcVzWXIOvNFtGmHHFG8LxPzuqSRqBzP0xE6CTo0/0+FSLcYReL8PIkaoUFpe6NyTkAN1UBTIpBVu
5plj6ffKtK5dzNwhHA6MFkKQimZ3QNFmOICTtm31yXIuN617KMBgzjhK30+bnPwKsM/Ry7w2c7Bi
ZIUriTFb5z2EqUgJ/HpKt7JNdjxzAtuh0UR/A/Vz+WcK+mIWJXDq6gBuUaiCMutXWU9n48bNiSpk
u8gnoKiUG0TMSgeJYQvphS9YJwRfj/3RPg5p9esgvz2TPQgjJ6OailcDPI9yJYiwTdTSkmk2SdJK
QWQvEQslRkU1YVY5HcExy/qCanlutQTtGyKI2++qdaQchYLl6BwSDIeWlnJXfAb58F4L47cNflUz
Y2JB6GKB9FEv09YlhbhqFZYCU/5BiEyxJrt0dT6cxpTQiIaOnXge/Vt2Ihf7ObhzhBBqcmAIqyGO
1hSdnlNxAqGvsy/wYNf0Mz5ZLFGdpv9lKM3IvmqPnbyd39g93xZhg+wjQyBzSQRYy/UOwwpXht/C
8UdLmvaeQS6SJFm2FpAzlkBO5D/P5Q1LIiZHLOhCYVeF3DSITPjpyHQdUxf91CukjgNurg9nZrSD
waoHMDMvqQD86ixmZGshU2VzsmMINWYRa/S/ta55LMzigQDlcMEojVoGVYO4+GSk4l8DxkqFsPr2
7ThKs3OSf89oepKOro4F9W41pu70k8sok01KylUxr2fIGsBK7n9+HaB8dBvcz9OYVnRE38gWSigT
5B3iS9a7HnbvSruyjqjHUgPyt20Urk/FUE1Tf2C+ORpuHKPRqoPRuysxGSEOmB2hFjDDpC5A3RuL
diUd/neQPwFwIqj7MSKtlVa/MDiCaeAxwBrdTbRPh1YjOZ1GFTyglmK0QNUyBybbD9x4ZLKi2QHq
SQtOmXmX6GgwDqS/Iv5LGQiDCSsZJJvv8Yatyb8Z8fI973s/MksgHaIdz2MVQc/+5zCHxYOi5cA8
dwAIoo905w+brV1izD5pBGjdLJ6uJkhlayPzoUkmJ89cbNHzWNH56QSUyetlacyQx+DfnCux+fFw
eYFOOQiU2uv7vAXvcZGcMRGBEZ+aka0ojK08Fbo3vBVlWa5f6O64173CL4VFyXgVs+uzSa6mbX5l
51lrpzPL13/hPIp2B9BoURkXkE4R7RlfYbHEd4Kz6ArngY/8OZmQPZpD5GjBjvjTWvXnhnf3lfsk
V5lYZUdJwYdrdQEwegrwzfNJRHJY+68nHSVoLqdjzf4+BCzXRFCEBE2cF3OpNZ5XBqWeRgDz1WJa
C/PYJYhLC1UUBviSvH9k5/AhfbjToedXQVw5Kq3m65/k14SE1eL4A5tk/LEfa9JOGSA7T5XuOsrM
H5R+mk6cXzHtZEtWTa9tFQLzx5v4rXT4EDGmRJMKmJoM5ObLp9LRm4P9VO9Yw6QaBoiPZjKTka7y
JwU4VrXMnsPqbuKYYT8ioE29ypHfDBoFQTx8td08cl8plq09kuwyzSKHIy+ShwaPbvnHFZuTulWu
vEa9FaQTWIkxpemFuVHJPAzuUKyy+CTWNIKEvxhDltP42XaY0KtR7olNyURiN5YTgHckEA90S1gR
mplQYWHX17pmiMS8KxjWE2H8X5IGKgxROYjqcARlCzp+r4qpCCAJ6dvZaVU0obtynYHBF0nRRPLI
xcECN+v8e2OIOZ/r+G78t9gGEQGAPT+y8A6fi7O0Oq7hesla2rBBleaVD4a/neKsptiK+EJ5L+P+
jOdg+dDEaZ4cR0Ve+Z8K9cKFXaVmvJGHT8yOhvUYQIOODov6bqZSOhaCX2ynVfwZ1t/vB2aUcbxv
ms/HhhKZIhEF5iZy4M0LqbAMXsiHGpuznY1Fq5d0FTIeTK0wZdTpZ2EsTiJJCoLnoV43TdBmpJX5
ka+cS/OpXdM/gNiEhRSxhQ9uz+olXlOEFgUvAta5jarHZTtobkTuUrVxHxgx6Ce7kQCQDQJhhe7g
XmuGDhu1/zx1jtVsCreI86oaaIchmw68RkxJYpOQAPkEkDYAo3Lw97l9aOOeaafmTNga2PGwqjDZ
zcIORio4nA4tpLfC/HGdcImWsMtHYeSCeCg5ftHtlylKTtWJO8kaSkpYYR9qO98zqpPxoP2ByuRb
Grr4iGEWk7mYdKYIznk/NPzJvVR8W77MOjWi8IXSQsCh3NClBc9suanJWRBFsPkDhqFLr6lt4L5g
dltGd5tZU6QimFLyzoBCM4zEzC0wA+hX3Quz+4U9GmyHtTdhG0VS0G9eJl4qJ21Ap5bc3xzhaX1j
rqivcykAtZbMkqf6Eopln3gVhQXF0NDncGikMcx+1CuQa8U7cC8ojdKbX+UIUjie79bATOJGz7PP
v7avAGAsT8rixSWLhgOEWPqNvqPPca+7pJLsGnXIBAHCfG86RrLnsXECXt077vTrlCTuLD+MDgTJ
GUaipm1WP+GNUiDfd80u1pGCdbJuPtvExUOiS8PPTANI/QHVwPS9JlykOWdUQ4yH4FbCwNy2kjGF
mpB9aAJIsGopkOc5bQcvJSuYmeWg802hy2n4qFC9SWX9tAFjWrV2EAg/S3+A/yZ7jfoTlJd9XUNK
LBLgy6q4aNicfxSIw1hGLfm/WmX9lNSGZ401ybqCrU8UIaoT+SrKLzoLDX5+0rhsYjbO5lNAzoFT
n0DQY0qn8+BH+UAtUnanBTDrVuq96UMQXkj4jDfk6166muBB4BefVsSV3bLIzhYrj3ez/PNiX9hQ
B4E4Km74yE2bmuTT5bv3rEiA7559M8f9H2oppWxeYC7x1MjCNdFIWHIrX77M3z8vmOPvJ9w/ySzB
iRTs7ZtF53SaoeDCsoaTeOQwVrtrr1xgoAGix2lnji7hyBRwEAIsREq3sgSUal3rozXWU4eRHLSV
XazWJxmDcYSvjCCL5afA4WuGE3OSXAjNL0HekRkRzWhsx63OYtfL/BI3Hx/pKnUX5hpMAODZGTRI
kHQ2P9pEU/v+jwfy4nfoJDtowetc5wj+Mw347LI8KGd1K5kR2K/f2dm1a2NpKFNNCsDQsRCL1X4/
+HLzpD0p0jURs4lcSBtZ/qSWodogUJYs9zfkpbQMX+xlYWyxp96atPnpTNi/iR/MzJeue43cuQeZ
WB2PKkp3hzafJFijXKwGmCuxwbk3JvuqKVnzwuKX5JpNv01sSPhNKct85PN2pnBFE3KVnYRzX3Tl
jHZdNq45pucvjuxotMChecUNw3gErlTWLERVEXQxdTulUt4VTBy2d46Yn3kDOdEwsFy+mLuld7Zo
qq6nBpRIIt98PubxXFDoetLFFSaeeKqwhEmwAZJX4lpIk1epNc34Mjodt5HC7Kbp54NkZCY7rTre
gH/1oai3PoMi97U90ia3IKe4+buX3HbB8OjaImXcu0huVZL6eMTJfIV8E2/QPisqMbA2OKwZe2Q3
ot/AwHYejWjwR+w0rYc0U0Ajx1ncHnPTiFds5H5JOpdmO5jp6XXUypTOAvNVomU1U/P3IkztOap0
6FI6f8ZHLHMsvqaYbwTgWjdBV8i555Ghkphswtsqg/4W9STnDc3HlYQKB2SxI7v+Xr5tOh/2Fc8J
/zx/jt14W1hB7PAIAs1NVvEkwdPXH3GoptEglOSznro3uk6o9DuCv1OA4kgCqY9IHqVMgTxKos8S
1b2cE5H/0wrqKwx27ptnXTo68zAzs/X3qX/lWcZzlg3P5oPkjDwC/5botLr4JdILmiBRGaUi7vlm
JQsl58IOnlbm/VHIucoK0C78JEgaghoVnWb9y5wRzlsNRkyN/YvbVcFiJlkMThEUePr6L5uD9rKz
G8Hj8drpSP1jMfobsGnczmbyt1CmZ0tjtI1+ZS2N7kZ6ypOOhUm2yMnFp/VG8lYLXHl+DMeT0dsi
BxSKBmuJs/YrQ6lVr8OT9g2FNZvzAh0cTE/lWc4kz8jj7yqgDLP62nd4QJInQy3KX+dsO2EJQNUI
jvYbXtz9180kdO3ZqRCLvO9kglqcDJ1YiFWyl2Wa6ndzvgFQZmYL7xr41rjarB4O/GldgJUbncAo
TaAanBWj/qnbDRdPt0P//NHBWGmWBO6lTRAmGp/dnUi6SwygwDet8PlDa2CtfxBCUCyfshZwh8uo
iNetkJ/z1qDXyl9I4e+nZ/LRBMoVi9P3zvYaJyDJHqGxRQeK8NQ7D9+xGeQT8//HEDcdgHFDZs4O
tB77+igsqTRsLWlEmDdkTBago0L6y+rIuRLa5YhyTkxcQXkoXogx6JuyaQcvXW2fHMb+9bFKN39s
sQ2uagHDFUmmc20Ih0bB/iLOCB6SvbQVii4wgSRPWfCEETNtmNwrx+1l2DcsvojlWIWElt8PEsS+
+5mpThYNlAgY9XEDC2OJNCmt7apJ0hm5ZSHajlXLp7DJRLCW6XIyDjONNL0cZjEdneI97n9Iv1Hf
rlETJ7YTEgkz46qXHRiR1XkegMhCh7WXZFGZiUUI/a9TUmYQ4u7dADxltC8YFa8RBFfBkMYDPqFc
fPeB1fG9p6wy40sMG86btmTeFFT0e5SQUwXbIfYOwD5fhs6HN4Lql3y8/YYX3Kw4xGlAYBrWUO2o
tI/uNV6WgS3L2cL2pkVSETre2VITnINHys6OrYA5gWu/MZKYRLzO4vhVAxbXmx5MOdxzCXJJZpSA
2q8+qWWOaMBDGRFOx2m+FEUGDO9WI2mvA1k5arQdZfXPQxIJo7z6X6hkaI43Vxg0s+aExH0ftDwl
ZPkFFyhf+hibrv5tgsGBi6IHJhWG0+pzQB3GuLXfAH/wy3rmJEByKmfpn3CTgAclJ+Qk6O5wt6Pz
z8NDIxaejqfZdNImdDlIvdVmKUA3YDlmK8tdiOZJFNSY+s1eJRQvyd9jkf8U9OXpzgScsXvOV6zj
8MmMLhuvH1VqpNO+5+//cKa2bUfEcmy1GntOC1YF3DZfXjgIFCl9GAqlQtRZ0JopwgRZiB/L4Pq+
TkIgUTwCdtv8yaAkzH96n5vmLn0d+/HkCmisKzf0PpZZTxcf+IqNHIyPe935B+eo5EkEjg+yjeEV
PYKVBcQE+gz07luWnj/i0QZegijstmayDDayrW6Wd4r+928t5kwA5lE1JYrI/NQNCUYQC8QWMFwV
vBuCtGI7SGz9l/jst4/MJo7lsFh223OoquXy+b0fipvngAhiRP3/IsHDDTsmM6aRg3mWNqbWairl
y03hqTgss4ddZsVvfq2DAl2//XW62cWXRfRmsjp3aAbnzZLHc4cNIFYgmaTmvfedqvEzG0YcCZaJ
XmZCzgPdAx0UmZg0fRS7YcmveJWac7dzVmAAaC4obkhZbG5yarRDw5ioSIs3TMRSUJBOBd+s0Yyc
iU5o6QsXE0beEOldjGdF5bmjnYwPbvG3UaBEiYyjP8kiAy44KU91Gjylu2ehmYwINoB6KIZb1TnS
NAb33xsesB2THAXmww1GjEHlRZB/hmZfgg4ovP1hOM3R0QYe19eu359EBc940WsO4zwLG1ZFhQlA
EmFq1JjkBeTvx+6jrKBmFaFPwMVnDzHDBYXgDAkjJhtuhT0qVfTWa+NnTDuC4KUi3emF4GVMO4y0
y5sQ6m6UyETy/bTNj7nyn1e9662Q0UkS4BFFY1IcwneMMUS0pKEZuIN+R2w4teJjGzfou9SKqxZr
3jwAbQotKw76CTXZoS88JRge5BgDgYg2kR5mwiLNcDIvIgXDcPYVDgNoZkrVSg193GfU8mb5kuQk
m1nF+VSjHs9rnXglr13QmeHV6gTeG1OEfmf871/UD1lsjxSExkRL2968Ob7If4IWT4aR2KSLrFYl
acOdNqFGltQNMuGBFVm1o3qiXbuqPVIcfk2WGvK6PhPiXOwCMkewhnt55YhjErU0B1VqvWLP+dA+
wewDB1iFfpfp1PPahPYeyxAdRAI2ktkX0EmV40MA1QvpF5TW1sM4+DSpS7ZfmtzjLYPnyfUp7AVi
sJJlnbSVyhtm0t6PPbnjtibNqZEBTR5r+RRaLj6bBSJXRUK3GGTOInu8uSNh2DVw9bQ1T9+qzaVT
KAFoqdmrNI4bu9RcoTU01qG9fIEDALmL0JpqKBb+V3GvtnXAPARPBgc0XjIRF6oyeP5Cw7l2s5pm
LCZce4m7fXDY02KykQXhjRKiu9P5eoHt8oP9tIXCiTocAN8dT1f6FuS76NBBD0nB+LwzWttofBxt
J4ja2HlJa058pD4BrsfZzCkCLW4zbNp9s03ehNZN7xP5AXgMgnMTASc+oRKs5X0WeAS6BzTq5J3I
3TZaCGeFVujhDN7pZMC0kvE/CVzhWk5BQ9oObdDOx6cu0cHZIRRG0YtCEPDi5XuNBs8dkjvjw63D
cglNPVYY0/aSM7kQkxlC+3esjSXOX6XsqJ8SId4wAbyS9TkweVxp9vtvALm/OtKCZOrexEJ/WhOW
Thd/tddhXVxRSRfGu6/jYkgSzLHiSzozyfnd1kR3twmXn4li1NL7TdWsTK7NXsZbu79aJy86EJcb
ERutvHC2S6YamTjMT/vDfRVdhvt5Wrk544x8fOf6dN0pcgtzB9C/gPROT3ImNCe+vI9ZCHOApB05
TLHdHcwmL3fQBIuCSAD5Y44XfDZXidsgWP2XzseXhy8oeSZlCl5F2JiVjO2HlqlbGqLqZCJfDedl
BpoINfE3sQN6LSZviVZRZK3u9ouP/NeIPw0Y9rg3aKVKvpku3QlrpteX/zxVzH4LxDBPFlIdaIxb
Y9cXDBeOz2zdt2LG5Io/zznUEMGxBBMLa7q/9WW+JwShteglQBADAQl1gdl/SihybG92Ua6Snl5I
HV/wIm02b1liJopz/YgO4+QBquzjpubDjkVUmHXtWqvd4fTPz2kCBrTDAZbuq/8mp79dKqcdi0t1
QhFv3oBWRVoGb9WRKvYKna/MfagE+bsq+PjBaMcCupSLpjZNOjl1IMr5kvDOBJ2/+Yc94aJs4aC3
Qzbg9O7ziVVReZoQDVDc4fqeUvju+Y4s7ThRQ27RTQieiy7zoRjov33cwaFYi+LHGdSfW6gbm2OE
fzGP0z7rGhiBQc3bW9T3KJZ7FzL1MGoLp7SBmtKPyjwjUREirCkcOv+eoHm51KGEhrmorYeLLIpQ
h24ynC0wgHpAlgINbSK3wU6H4ZfO2INj8DE52P2rJkz+xCrHCJAxIcMvps1M4u4SSGJT3Eac6eJ1
baKs3Q0u+CL2XXRtPshB82y3cGCn58bPn+WCZFbySdAVbWNH4xr0H12mr7nroCaqadblV9Zbe0HG
yEUG8hplItbcKXcm75N5y4F/Ec3aHYJJFyIQDRI4T0tMWzxtoe0dK9rviwv4mdktGaSHl2pQDc6b
dDO2F9P3DJu19upRRsSyVdJVlzqI7Kh9+1kv6QOufSD7qYG8lAE2DaVg7ObcZA56klzpGqurJvBl
F6qk/7VM6G3ho7U/UOm9y0VSlH0bnw21E6OvveVf6npu0P24yR0B0KQkprFIfGZ5eJ+H+ZkhvIVY
15uhGH7A8lYB0mP0lPfBb0uG/5izW/7uk7k99VmFvklL/eMjUIlAE8/PKs8jXRsp+NEvWghCNQcR
Y8CsrqyOWNwletDjqI1iTwV66mcml1Xsx9Pl+wmoE0TOTgdEKh5kHs3CxXSvvH88E2zEHyeyWBW2
cCmLhEa7iABoZWKW8qBWGwyLOrt97AunvgmHmjKuaJQvHweTGSj+152e6Zot8XEIuDlW6d3ewC/x
Fy4ZruCICC8bV3aymrRUDpX6QtwQmH7VkDjrTQpVibx1oCIXWdr1/wwyeawqKNjJUvbUfCEGB3EM
qcKxCbCTTadS/Z/uVDLDT69xThkywJxWrmGvrhNS7ER2w2BFqkDKUuGQbI/1H33tj6W2XtTHpUiZ
sPKIr0xtv5IELPvrmViUYZn6K9VA7XH8+8RKUMH1kuczLEFV8gry8wffooUnUh1xzrc1tvjEeuvr
/47cS3/GmDYxQ8WaMxTBnRcCMtHKWaR1xdrAZDHZSMlI3BPRzY90b5LksW1wiM+lGgN8+qxgCJSk
o8Oj76D8Y6R+aivQsq/0+/7qIfa7waVJX6a3ztk5dHaovhJ5lLa4rRvq+5pz8+47mXAUpob/Y5yq
NmLVpuEEgPB7Y81MXPBYFevaOIyyQjf6IPHhbXwRVBJvNx/UOEE4pcOUTj9byEw8hfBLItRRB73N
vWxdPDcUPLBYbjxikZAvXo2UDUHQvgC8o6FZBdj1NebXs+1a2QDYfvleus+q6f9DDsP+togHy5Ac
uzzKO7X6EG4aTCtwVx9S4CGRVAtTf7EZjtByunT4uwK7i4YWdUZk33AhO3p73CAAfrRSrTBbyPxT
58rMaQFFw2AnKb2gsVVHAr7IkFVKgPcELo0enqaJ3nk9uxs/cYmSrWjBt0R2VB5t4WQQo6gfKeJi
mg2znK2CuvKPKv0UVxqM2WEjRW444ccmJO47+tNfVwlBjWuIbLP5h3ciSP2aPCPpqoXMgAfpumEB
Cg3RN3jR8/YzIQeRlG7tNJFtA4dOVEmNNJxxHt85opzHgVlyeLAhdfnzb6JUiw5SyrYZGM5eR0md
EmXdzKvnSaqV7/fYRI4prHnMcmB5pTzasATIgnbNT+omP1w+VlKfFY2wix7N+WP7ZbeCSY9FP8hJ
w2jMmPC1dO3acdMgY5baI01gb66bjUTprUfyogJc6PvAMpJ9k9TFZvRR6q6+2sVCq+OvYzJD4A4o
NPZ0UlkggFU+0gBhI7M7JmWJ4moZasSM5Bv//M01aC3v97dIZ7+4m04aPEpXFvdeGDzfBY11Vn8Z
nsJ/eBUZpNPf0ccEe9e+pVLhrtnVb4AhylXxozsFI80JzlTKSDMQbWjQgFphlCCPvxbm7gm5rR16
gTr+BZLKRFiqn2oFtMD5stSpv1tYIwo58lY86e8iG0JIM51SUq8IYsgk4IAgSjJrg7n1PNd0tFGT
aIKh7QLOgb6NVxJHxeB5FsGWB1dwAispJ9Oeg3bJLWWprERsu9lRkhmWD+ZtfWaHEhP01dDV/7QS
++Uie+t1q6DnPnkR4sgwmnNNtjZOGbns0W9Usm7VB30hZqJdIqmXTgvEKmhkBiDMbAlkFCS1pP1Y
c0Miv1NkvX2/7+YNF6unaIBB8chUVIMuvoD1cUO4OsPWv1GPv3RK/AqsXgw8Mh3pKRy22LTpd/eQ
e2+PJ6Qqy/MipZkrdCmArFzzeRNyJX7yCBXMhBBHfVa0iyiuxPna3YnyfsiZ15fSH14w5Kgp0EOo
pZKdFtIFJQzY8vnuj84rW/qBsKiZWspqBYPCmCgob5TE8KcCQJvDuSZmU1ZOFQSWuJA5Zcw0GhJJ
pzqgjoGduheTLqOFHnxu6FkWYloy7wr5I1w/K9+e+I2Ys4gGih5Z6CUK1zI5uqcLkYEvuR8RrdMm
dAwzEmIUFMN2/MXkxLqTB3qsIOWgPKGtGE9xucpoIVmTCFdSRE+KOtUdBAd5uNbKCNlB+dcB6oOu
PonYobRKfTWOyKDiLCdg5sGwlj2U5g1QxxjSe0SDfhbTPM2YETyrUTK+oz641tn2qtW+G8Bp0NDu
rtDNsMV+CpX9IJ9xzjYWa3S2t0tPzrx1t+7IDhRZbDyO/bXQPsA3X0wwVaLLqhHmb4plgHheBv6s
kGPtW+r4v5KqhlOKRFz6v1Yk2bTS1d6KwTTgLbThzwPjtdeO2INcLJ7ooUmV6lucuE8K4ev8Rve+
dFwA+lJBdLF+LzyCWoOKg42HrIhANM2I3R6t642gjSkwgKTEnuUhEJHM+eqPwtLbEO4ZAtyInwVT
YRW+WRRffYyVnqIkG/J80ACPJy3mD10BpLPf64L1HAPtHSPaYI6XtxLI3LMm8sRoJdmOjDkiNyCZ
Nvel0KgLJ2TGt/d/vGLDu+W2O1PFBSwtBvgPyDdJHJ6/pEsTQGig7pho+3BDNMo6mIDaQq1nnkBc
IzS22coTz2rKcIEu7wzOeaO/3oqAPzmh04OOR/0CgPwz7SZgCNFxNuUFW+3av5TN04z7xz8sxeeu
UO4vxO7BoRqzgUcwy3sXj/q/b9hO+trTW9Z5qgGk9wJqusbzvxXeKriQfrC2TPL9z3YGSuYyxtKV
C1KAOcdupFq5corKH9AxbTphmVdTxx/Pc5ha2JiyV9qezEvKNqKCILFTntynzRtxw/KfkU4szL9K
h9Ilakf3zVIgNgtBDWkUs71bbzZFdYZTlv+o8PyFrku5TFnGWYI1+wP4Hg6jWVgey8aMXz1XhgSB
dyTop9G/jpS4AluwMnMnGKmfmjn0fFm2Yke1vO8f+1/cnuyEPlsGekTIDYlO14NXdcu82qum89AL
gP2MSCzGV6UtVaHMi1pwyBvGwaXhiC/fxgcvQh+txKrOo+xEGyDO3d3VCpi5ctV8Zq+AtQNhSbKX
vAIP3IVYYQ9ZBcsh0c8SXKPwUSRbOnLF2ka0lpS4GdvHEqjpGRtI+S/5PL1kyifIOWuEl4PZoCEa
m2u4bmHXadEu60t6y4aOzlkMvtG/+j4NXWrOvslJDdAp9fmgAIH1pHLP3fq296BXP0FBWDXGHuKn
kr2PkYWrIXDAN5hqpT1YlFrGmENuBymDbgO3ctKTpuoTc95j7V4ZNzKH0IJAYZNBXqr4/vLy1ot/
9RdgXj2mSxyKsAv58OEZF73t4vEU2itxgWkOa7kdPkk+yAIyHtf5pjvpTT71zTSv3wGJTkMMgSNN
swrCNnwsgR9Nf9duFz4bbpKOrcgoUWlWhk5mVaS010v3dyCCu/1/ht9PROcEjZ0D0ITCAy/Ks7ep
4MOW8Tvzldglcbbd8w9e0zudTlG0s++BWgO1yQgu3n+TY5Uv48CLX5LD9cPMfML0jTvL13f01unF
yv4SHFYTRWGRekQJy1kxlIyNsXyF5JvmPk89RpxoUQzLo8lRuom6zqNMxGjXlYTtrjcVtwEzohMh
552KW8pswk7iC1CuAiavJkevr/AVCVFnlQRY3C1mz1GX/u1IkWeWErLmDEL7RxZmLn37YH7YCqZ+
EJNayhfZrLF+M8Py36tEkSpOciqlttU28Nft/j3lxb6oMrna9r7Vzl0IwCWrlPxFFEHMPLK344/n
0NXpvyvfoCvTB/flraljor+lo60kL9fsrSk9iLBKV/moWQxHg1BzPZhA6JoaaXaGegFc6V+FVhzy
lppjqV6RKXACgDHVy8YbgdMA4CPMUXwcwOkBN6JvcGxC2nUPoo6Hqo1YqWKu1hOzEV6EXbj6sjRT
TztIKXtOHJA7HhWqbTCpa6F+ldfE6ZF+UnUwxru1VGTKlb+uhZd04kSn9ewPvtUoF4BLcV3q8JPz
lRHZ9ZY9pzMyY7nq0ITtcb2GIKnR65FE4Jz5mWKljgRLGpvriJEHFF4AxIbYj7RgQxNAcNQsVSi+
qp+9sJiIorWxH7u2SAuFKHywvNSClTlk+f9hvPql3t+5AdrjAx9yXXwGen2O/xg35DRK5krVk2cL
zZsSEQZZAERhL3EHPB72umXswzVoyRolceZo7i+9BMnXHx7dDibQxEcaVQSzITuXqRq4w3kMJzaC
BSyjPTq37ZfpTzsQz4A0CQzPmbjsvMdnyXFvsPhchck9p4g175XQapRs19X7N6PEWiMdo3jwzfqv
D06YyCH9qoV7khXTVAd15bpcTstX/vowQEBLbopF4nb6+v6W67/kafM08TeSgEx0IJD8YGeDFrdQ
UfwxrArKir2tWWfZ5uoBQMSbhZfd7TPqqt1bnW6lyMpXBBASAF4z/wt5PgDorkn/gzzZYLpdwbUT
NLAnDvNpxRBOd9XDOHBtPTOczpUgORhz7yG+l/byPNkkc9TIyNAJDHpqwUHIV5awpmb4xoAdZmX7
aZfPBk6s8D5MB9il8LucJy/N4YZNl8xz/IOpK/PgjnH/9+w2s8mTeGfY+SN5jqoN6ht5I605SSuG
mQ73E01rZAv8ZjNLVDETRx+ABJpq58mOBTv27+BxQuu+EDVnyxaAOag790/E1bXvIvdwYhe5/aVP
78HbWbcS31K/BbPxrwuFMErGo+IHrX1oiQUit+3aCB96F4uMnVkq5Mpb57pYqEL3FofAT5E4OtbL
X48YA3wBWtbjBsp62o25DU+uipoXonp7kYc1VaT3daApcDEdCSKA9mQ/+V9DHjSMYyUfLHQEaw9S
RK77vXC/m9y/MVWj3gHBOrejl6KIqWmRJwC44HeYKCLaxDi/Iy/Dwv7S0jVxw5j1SUf/jH1nTS7V
4yu3wq5FuwAOHDBWfEctOyTE6ddqAC9ckpu1XWEUL62Zke9IUdNc+M1BQ75O5lGYndSMEUoAHJjg
4nGFeNNPIIqtn2qWsSXzIoUP2PtIeadhXukQyxHlvSh844iQ2uRHqLmR5rIBHsqj78OgwhoMGufD
Ru/Evn1tEF3H+uo8wtMEEHvPHcw/NJGqw9lSY28+Ja/lRiPfxP41XxmETt+zWii6zj+hKToupg2e
igdDnjiCtO7gSukvYptpXylrOVWwTF7rJK3FT4CZMo67MkVS6rKNMOE5Hgl7htlx6x2zAmQdsxp3
WCS0slvLbeZM9cGGDIOm6PjaitX4vapHq6RKy++jrnQjiPiqu7szKk7Hck8pf6AkyX++W05Cx6cr
mPcVJt3/Jg8nbXxjobfjmd40WbcKCZqWkq5wuRDmLtWsSYmab2e63SkKX04DDtvGVzzppF960D/o
7Bu4P+lyBCWo9lu1EEKciiETXxzooCcUcMScsPf6c62RgC4AO21ps3CMMDC5tKYMmhithPo0NnyK
jqoSpkzn7Esjx6kMO39Ap+FP+uc8HDhJiLWA7NPSJTlgx2TGn/TeeKfoXn4ebDHJMzcjbxIzHAw3
mfr0M4lh1KBfrlAdjGW17wHpRHmwK2Z10fFiGzbHahMA3pkGyD0nMgZBUOmtglKR0unUaajparyI
gkg8fynHKGr/PXc+P7aSrBHN7sQD89hzh5sB86+ZxUkDZqgO/dMAUFvpR4Ixokh6gp1SGs6JBlF6
NQnQ5vTLC8va2I4ZAyWduyRRFa/Gy2qWU4JlvVnocJecmzDH+JRfpj7YxbkLjSOyLaQAvuFz1Nm1
srwHZGfaEZbcOYgHMm+Ti7E4Fa9o+uanV4t3NzvtddTzj4j8BLfcQAninACEBBuPl8rscKE9S7ii
9seLhd9M8UUL2GNSTKgn51ay7Pp1Gcl+xDss/pwZFd5f3tNHohh0qubuLlIM7wXefr0NcDIcVESa
vR64fSXYyWfZ+T6wr1NRbdPA52wTf7AGtzy1gQbLDHUjK8qHnLCDYBn9ocKfgx93b1k5Aaar7N3Q
HuoR+uIoobQkfkacBBERB19B9nF1s3yizxutGVhXfov7Q3EueFcpKDn1dyrYBiP2/Blf9NMudRLn
lPx4W1ja5PNopu2pxYvpR+Ne7ZO54gooMeo2xOVSSgzpmd/x6QfO9ODF39uy5Mh60LPK1ZC9qaAz
nyVmNtJ+/dN5h8dlRYaxAk+IjARxma4Nz08xF1mC7ETsOJ17TotQ5tI7GONdNdVp15RashBWyRVj
Oy5pEwgVmzbBlC3g7Ah2Hrox9TIFYS5k5QJf2u8jHAlgrFT4vIpo63CekUoeYNiiLu52ELO1zOMT
tHkZoX/1Ay0mt35ZZswFdm9ngDx1HDaq+bphPGEV2pX8e65qp1GKjd1xwzifAvaHZDL3pzbJRbKF
F0RltYXez8phxuqolV1eqEHm5NqD4jYdspFIOJkYIeB4pisOx9YCJsqNBMH4R45XOruccDJy0jcp
bO648DykH12u7ssYhtzQZ4d/+h774KTBcy7tDzKGJzWGuKmoRur+jM+OgzEucMRDyk3dS5sIBmHY
zDuarH2SKzkwP4biSnecbr0SqzJTnGWkgXzRV6rb+AGfB2kZsnySstIrile/CP/LtoBddKTfKErL
9jWWBheniiqysc22sjSkSdDl1KHWwUlwQ6Ic+Utorw5KdfFjbOZeTW+46z0TRhvYFFzTDMLcRwuN
c9e9DBxpnw5/WDkZFZ1ACfSykon6I0mIKiHb366XsaKGuRryiL/ut/pFi/ppX9q4/4dDwv+vWJZV
nU8yguCai6TJNR2SaRUEOJ77X2kZzhy28BWUeFpcNWbXT8KCRTNoohSVBDZqtlVNOwRq2gZELWPj
dbNrYwezG7/SMaNXnuxW8PGTbQRUKqGK5RPPJ1mXj2bAlGd/XZOFsebR/ANYTrN4E2XHhn34yYFa
OkjIM1NVvQeGDaJdRYzK/+9TLWAJG/BSwru7s/TH7s1t4NBXRzgBZ0yy7612IzGeolD3qaI2tuch
QRO7Qq5TN9GMtRl2l2MYhKove0MsxrEae5joCeLaKtr2RV8w9HSZe3f3hLLZb5lOcXFBMrScg9xB
QJrAtniDjmUtOFWxpSmi2CPoyLIFF0kkNd5myavGsrMUa/DmHlrfoWfe/qOo9GmoR+t59PUIu5hG
Y4a9JpAFNbA7hRj34rWtArmdaDdVjzPPS+8GAi4oCChyfFhRyaRyhsh2LGBAvYRUn8q/9nF6zQG1
DZ6h6r0PbqPMJTl+s3+Zr+kmco3YwUH9wsugbmGQWVCdukplw5l+/Yp7wxp+aNRoKq9lHQj3/0Ms
iGAUPG04Ly46iHYJUS/J9VDXp/veMT++IH6K9uy3bb625y8eQbT/Cve/lxdgZHfs5TaWyTVmIF60
MPmGQKSfZpESW5fGwrQCBGQlmuKbeV/1jwZq/RgMIusNjBkqg1cEHnaUgUq4SHjuFBR/f8RWt4Y4
wVDDLpwi8rPOjrBlhF/jiDkBHSgv/4Ud/JW9hi99XtPDkCVNHZIhvE3sFVrFr5kqsGCsT2UbjaIL
nf219QEjx6sfm73sHP2GogPo8fDfn90c2ASdgnL7ZiedigAq5uQoI/fgx4hI0xCrC/Mr5LYjpTuI
FnXe2Gi0mtJKBrA4T8TEBTGE1F/uGUWpDfO6rJNCjAnSNJK+Ke8K0FOdQdhi85vkFUh8RJgqyFGQ
oVnufq6wRVYZTT/gyfAIxh38EcflO0qyH/98v39qGZ5tbZD3qHkYAW5mf4yUS+bjorKHeI12bg7C
Uv3c6ZTvBlS9SpuAD3JPQ9KmGtbdw/ouup5eNJbfeKcPWMpRvteo5nRfjzWZQaMmB6d8C5FwaOzc
A0xqOuMc9Xj13Pg+yESpGGDlMIHj3xUdlakUbLaafV6KuBCstva3RCmjPtgbka9VZlFnqHmAodJD
LxDDckTQx7VIVCFXRzjhcgmtQoT9ncjUEkY3WipYfOjgjsiUf3bnu9Ftje79HvzujBgpN3gpqKVf
zbQSfa2sZCkAclKZhmJ1RZCfOM5+b3E+6kDR8aspJqSyiyNluqYMagyavqWZVy7q4NoSnkBHqN98
Nna9+D6aZSjcnhMjykdtY/eIB6/u0zyqQGa80cCPKuehR5G4tuHofus06p7GaoKMMNL9KBN7RCfQ
0JVkdIPyLmAl8YrCCaq7pJ6XEIHA6qOBYzDLO7jqR25ehdMm0thfONUtkKvs8Vv71wO3uMJwiKRP
1fLrCNHJtUAOSy0SjfJ+e1LyXNPkFcwOer0278wumXK5mb5OQ2aDGKwwddhmJu/cB7j4jdeQeoCR
LyUPxRD30zEv7hwH1Udz0Lcxe90oX/22WcPSNVHkpRkxaexr6O2b12kWeoiA95t+Xghdr7nQ4Zdq
RKYbjR2svif2wggMFiSUw7gA4wUxEQqCEwH2rRPaBUMpd7WHcoG7huUrwUSG69ma42bcmsMkxOD/
2z3h4Xf4f47INfOvPdel9D7MtYvCZx2cbOOi8e7SB+E79EsqQ1UWkt9lggZIUXyNwH4/drdwGH8g
8o8usQMEBW8wFjXGwv0D51wzkh39Sq7P+X4Lix9CKDfTYW3dxO6vMTynv720/4F/HpiBHMFL/rLV
X/5r1LLYL7E9gDI4/Lwq8J72SRn/q1gxE4RX6M4pJKSwyNZySTf4azXJT2hx3RCovVvc/wZMT1Iw
fzoYT4ir9AQEtd8g3vtm6ZMUM8hQVN23uUnYUQhCAKxglP8qix8r7TWTmTIjv7mfHk56wkJrrOBG
mKoRaLA4X7yCRe+gtmSLZ0jSaPcCLMzsL4EolVbcmzsRlqPLQEgEnp/6tD64IbbVn01R80Hlxnv/
9lW7RfVyun4/8fMVa3eQJpKCaO2oFJangl5SIKMCCXmORqQU5uK52cKALJAMboqj7eYxsQLkiB41
n2uVACmOMuFGhw9ZrAkluLuouyvL34lkCUPE/bFkTiebf9+ugc9JYcUmuKbT97TtcKFcwJXffbYa
EOddTKEfj3tPGh6iu5REuufkQAshPLWD1mxbfPnmDqPcVsgnocq6i8KXAjkCOfjpY4VfnQNrqVrg
LVyQ7VfpRBo87UvZIO8FSnwFoJwYtsepFm0WRo9hiLUMvHcvyqzPOHUim9bxzCmvwLj1vc2zgTOs
emf3kyjQkFsuk96fJwstN2BopXIGVVX8sJRgmSWhwbXj3JzeF/OjFolghzWYCHVSN1VcTF0td+aD
WeVDmwdhk+ctUGGkPyszotSrFs/AojB7usJYIOtigd5gSFEoBIvVsK6aZU6gZCqez3I1sPWi2jQG
olcE22TRQ+Ddhc9ko8Y1DYvOX8og+sDfo1n4kDaKM09pIzfAP0S88irQU2T6he8fxlc3yW20ZLhK
f/vXwxo6O/d3tNJOasgM5zbM+Go+oZr/wj8lIrWMuQ/uuJut3KsIHqqTw73Zp0xEfufoeAOefANi
y60fid0GSnbGPrWKxrstKogxUPvVUrB4iWxCtgl3NP2Qz3QQJ6CjbZyu2LKCR2f6Y3JM3t0Bj/J0
tT6BILjE/yF35Lxx5QF8NcHPRYRtwbMxrWxzI5IltbZ8mhHHvC9lllFnHS7jW4oiwh8khpLLtTby
95bIBk6LaZbkWJCijXjE4BzLtWNUEB6sWQ7vhN8dyNf/thGY4hxzFvU4og/Ti9KzdnVsbdlamyzt
/UEk4OrrGuG+HjYhLBU8jTPu+lDyO0Dw1R2iRpDVzFuykAftPCldwkYnTlHfMSMB7YExusDz2v9R
GilpwHYJBuy/AxcIwwoydeZYjRHarwWMT5kvlu3tiC/ln89+iqWQsZ8UzhkNc6GoZHtdAJI15rbN
8dVnU+yR12Q75V2SG+cWGb2iFjFXE9s9ITjbulwS7toRWplfHMH7X6cO/dGCYAE9wQ0lR/kWCCwY
Mi/PCltARhvup/Y1Ia7zEfiwrrwUqyJazVIkzGPzd/vsJ8UsAtdcLsxRaQCZsKzjyurm0CfeiXBZ
NXI1RhWM9LCMnZPAVz84KzrP4ha45L9aMHAPf5unUWwpgyhV071o/ft/IlEq+tL4zs+QuYqlMgq5
X9KilMkrizliubTCKxQDMiaPjgMDuMS/z02JxeWLBsIgZgi2Td63l4EEMnUKcuK3Ey1iUukXcIXC
frmSrnavjPTTzdk6ekic1GG2JUtC4zXIP6rW6YR+EK1Zq7qQ23bLnVB0PkmjyzOpbGSCSXJiTw+B
nHFnvld9ttyPmj+XrQ22qBRDyAwiw+2dizzbmuX1hod/EBUT5kVbOYJdC8JXtsQb8O8OQR9vwIZq
FpHIJTn5vOhCZeHrvFZUSBgbJwn9Tq2Sg0n85A/GISJ3KIuIk2/S9bujq3tDGWczG5DJsyrX5Lbx
o8z8kndfxpsbvzUwJZxEoFfurf5C5SFzunf573N3FkWt3rAnGMDY0IETgzz3dmGdKqKZUGM6461V
ICauMwC6uMq3kpdyiWcSM2EyD0JeiEwK3HyVv/YEDUtD2cEZxMN3lLA3tMbLto0CrWVFOzI6HEQW
lmuHyJkM3jWHpIqlvDl7hRjsH2q/aXg0DNOxhgSDKr/epvMVKQIvSWU6yB4BGpM5WVWOpWm3yNIy
iTZ8J3n9e3FRhK/AZGiFdzLivJXbqqSaQQ24DLlzpNfVZ7zAjujK0U0LB7As5Pp70aY6m/rLAr1s
omKSZdva7NKmZc8IfnsfkGtR+71/EgHtZ/n8lYHcVvzCa9W8XJbNvE+s75KojrF6NclLWM3F/xcO
X7WWHDS5u9bDqIVChBLGBUjq8upyT+KT4ir4h8YOzzRdL/o3UmKg4fOD2302inWzJJcD0IraeV13
99ObItHgldG1l4zSrh/7Eu+bjTayEzWlkGlGb3vVDHO46aYkgpkVR1PejfC0aw1ED8fGn62S1/zr
mpS9epV8jchsqo4N4mbiPKtL0oMFaqnvCBFnTzAZuC/9d8C8XSqY+JTwUgM+yP/a+DYWfLDSuGFV
ItPk24gyyrRjg3ItTW0l8xI1l+E4oEFya6lvtuU12kYKcRisBnLFZQonOUbGV3ZPR3Jv61gQwoia
kzT4qPX2WLBdkxZ7c3wGQQ0+LYU8yjJ/eT0EFfNcXlFMyKjIhm3XmIgfldLHrZs4XqqlW4vHBfPW
i5CsIzE5I3V2NkIsL6mTzC4IKpvTP5ZcBaxfufmBBEDcoQlCWGOmc8bb/b38lJ13noO5ogfBurFf
t/UxFg/f2wE94oSZUaIdHRoI3OTiECRL57x6KONUncvGk8/J+OWLaa5pimzXzeDzvTsWhwwEnsAq
NHyABQrkrLjLuuYPJAw6FeRSgwBvhuzFvUddVyEZCfOVZa3M9hHC02bVgxUYIz5w02J0Yr2uaPvv
pFkcCcZeJIdtMu8bJjpLKvz7556DgxUEt8Kfkr6gFnet+eH+J1YV/4+IszV3TiiNIJzjPfkroXwQ
l9+XQ7MKTBK1AIM50KyAH/kH7iFurL/Mv9atfb2yrcGAWL1+ScL8XVm1Uen5v1y1sIIQnw76lrUN
V4Tgk4xJHgHsL8PW8lMr6OdTwAnZcCQgklyM//awJ8WA1hM0UBEPx7BENjTw0VoUnIfvPTDhb+7b
ItK1PKpkDaJgSTHbWwzyvBCtUGWP4hHWlOzR9Vqtrqk63X5e9aFHsmITWTfbpRE3cCUTh9kMqaF0
cs+hRrdIavTyykQg+KbqULw0xUU60EL2kkkQkHTKDwkx0/O2QsHh8/SMl5SA5gmCcHhMUGpPahxf
dLpaGhjisJeN4DmgYhB5/ogUK5N8nDw7tJtEsFkQJU6oDTfvkzYAg551cM0EXY256RQ3gZ1seiXE
i0Tm3amTVWdoR2U4t9KmQgRss3aGEt5wn8ZSREK2jjcd16nb4xbuifcHXBXRACPhaGtdmedt6ekc
j2u+DpyftQZdzBraFPYSj4OuQ7DcR1OF1UAI92IrKk2SFoI+y9q77UygNa9s1ee7G4MhjPH+2SVH
AROw5pdqQWpA1P7zw1dqtgN/fKbhNZ2kVGmyAED/mSDl69zymhE34ppn0mGBQjjLB/sFAqeyHDve
+uLrt0MMUQEiPp21sEoAvtmJgURr9rAeXfLBAS5xV8xFhnDcTAWzdp9+nq/lE4xQsk9swztW/4cr
xtG6AmL7gIBTSPl/urq5KbTeSoXVfMiu8cTjrrKWscQcHBPLyXSX0aUFwpfLv58zVrF1c3Nklmec
dWmOQOpTny+2MNQQOCkTx6XYZe4ipTuZtIPCbQbE/addHELY5/e7giTzalZuCGxMTvENprbBku0d
E9g5jnOxKWm3ank0F0d++j4c1q7e4/Yeg55oZRh36xxLfeVZCax4dbbmSXuDAaozp51OnE9rAgNE
O0diQrirOiheaWaTnY9Sf69ESbTOf6DrxH3jaqHUUigH+HHw0mfvv7kuXJb+ovtk+Mt3l0SfLijz
6DNvte0EEHP+Lnv196RLi4BB3V3x2WZWisXjxComvD7yTKPxbTFmbZDekiAkJC5mcpN5omGlpht4
VTchNDVJ0FGaK53AZ/Y0wNAaYpzhNSLHVcNha/dRal4P1WCzy7qPewe3m/nY3jsO4lMv2NMSQfMk
GTyw2tqMW03D7N/RZYzYIlXi18Ty+os70xQD0uD05nrL7fXItGYZe1ACN7QczbSUZAv9FMQPJxQd
Q+ktrKNpG+rVmrG9wy+RpIhZfmR9tWqhvgtVuUsPbul+rJgnFtkSyAz6/D1WY+7hM47aqcL3p7ob
nODuQlu+QJGpCWSf2TOrUksXWiHcV08NMBuLL8Yl/xWy8mmCEulHUnaxceX3V523VjL6LaJZZVb2
3bnG0IV5AzDb58kzpsfGIdJob9N5opG/hHp68UtJJQYOmDvqfF0cjbHJ2SdTphUldCY3tyZw3kJy
ez5gJCmRhshIsGHzRLsN9dIQGXMvbKjmxRWwmzQv/OuvhTLuS8joYyxFzUIFNBGwOik+oFMDRNMi
N+57rYpHW5vp60wOjTfGKBlCk97NACsgiTiQ9m/XS+KkZGF3C37IJwaay2nml5Xt8vK0rzQR9hOH
Mev4DCylompObYIspUlBRhP44Amoelz43XQ+PbM7ejKJpGoTVPJjGsUzyO0gr6jvssVKj0Omy1Jk
qLfH3sQKqirk0EdJJJE22UcgufSuM7eDdvtxqfQnf3qfmnb7mZkRpplZa4h2J0+gHfWorV7Q0Rqw
siJsXCs1eUkH1kVuxcDBXhzQyf+B7764RTdVgqS0FUiLxr7TiBgsq+kwDaYuBqrIoWcNRaxGqSoL
nuLKy/yA3VfNIgOfMwTaZcFMYOoAO+j0psTrst50680p+izlOHz9Bhnn+LH5WlpBiw5ghcyMj2qu
+Tt0q+b1+mkFsehnkwtXdzGOoFy/hRIuV6Szz+/+5/2Al95KLLp8TvnSCh24nOgeEC6EDyPPHcgD
w1te7Mq5rJhrnt+IkwAiFeAHXulm35/Cl9KktCGr3fqKk8BfI5pn19/EmHjT67FT2D+pRKQcRXlb
Qnl8of492o9nN8f2IKKMESOcnVAb5v+dRUBW+RQ9j/M+2ca5eJO4SUigZ4/rB62HD8BEXn4i04YT
0ZE5OY1hmWPIhPaIsXgRlShCEQF5u8Urfy+Ht2WMIKA6I7MH0URr2RaXEb3Xq2Lzmfg7iyf2a2ry
9uZsNALib6F2TTUIKKXecKcWQ6AahiUX8jKdHgOPmbvNtHVIMj1XTb0DNHYWOZIJwI7RoReN4fkl
jI+LMGegomtNC5OD2gSOB++I2V2vSKQdIRPKGtm6UFiPWNm8xyrCEL3IgMMRpPJfv4ReFlcieWN7
z89CVUh/XJKx3wAjbGHGqn5Ex0xmUMW0K8NMPbJZ7Ih63z3WrSfLW1r3XyyRqwh7BNtFBNmhqC0M
REd6xOv5LtDH8QU8GlG/9SxHwzi8NLWt4W3pJhtamCIT3pbUjVzbrTOxJyvndtCGBPEraYeH8Kbs
glqLrPiLagctziXu6xNnQDtKUmYH1pP14Jux5y3fr9gRZTRijWjeiIyn/zI7YhgOhCgW9LsAcbXn
b1FWOb2+LJzNiQ3T/2Z6EDNDKljjRujqf3zgW2DOoa99N8lPdDO4qww1EhXtMW+fn3V2p5brrADY
6yNj+vIJ1ZfYJe0nOcZWrPFIb5cqUR3VGRmJwOCeuFLT2wiJ1cF8paEd9uRwWQfcPGiQQrXo42By
zWTrrTNIDTOaoa/9MBiXvTg7Ev0suJdtcHcT52tVCtHFUPFS5KyVbeE82Lku5vvvzP2c1pVMCa3W
ajXNWkKRx78j/RuvsOrqx0bbAinoO2o0G0Zhn5Qw2L4dnbq9mQ/Qnfi8APlIx/ymQZeTC+9ZNUoK
l1mvdgj228ByXf3yw5wIpLqKSKNK0xc1E5t/CDX/HUy0a2a4sGTkU/sjrJxw3CoG6wdgB9ch47zC
ElUul5vSGYMa4ZaFPMpAx5KYtThSWrLclwsRvJZZ1+MVPY4yOvlT4E6d8GTObTMGp8bJzoKbes9X
V0Dcy1WXjdEQabh5Wi+X1yH1PAIeZ5UvEw42wdWxBjt7n+j10mHdUPBhgD8sHUigds2bHf1KqLuN
GBbtP1dof8kj8OheIrFFr1jOsEfrjeWdt4ElpOtXf6/6jgHeJFA4V/OiGzB4hsu63idjcMQJLYiF
edg/LdPv+VXI5Y0/j3yfXr6OXin4iigd4fEm3D2VrIFIJ58rhd2s+SwWYwIBxm5Spla/t+nVe+/s
ru4i2qTWsIj2+Q9Rwl7G3xkez3QTb8yG8+TUsm8BFeJiwL/u6U6R/H8nggs9we+8vvfKfMOfsPsH
aV1me7S2WzxTKAJJhzkBgQsUMbPz3UVWkva1ETWHtt9XuabAFlzD6NrKlNdUC8qHg+ATPxEnqy8f
0payoxEmaGTZaa9d47t24LtuxwpEib6cqVZM3qG7P9Vsn+1VwQC+5ck0FvuoP0Uj4amKy7+YQkhN
FH2n7yXvzoFLNsPbGc6nCib1ohe9UAc4n93yOfPlccceARg+ct9t6ojBSQbe+XBnVOpDKlThkg0e
9dOGjWootHEMCq92XRiACUSuOgfJmpqlTRJvbynGbuQ3H75X9hXt3R6T8ab5YD+5lNGh7j7Y+3gR
iglsUVZsSgsgtSrqM1iF4lZgcNOrAtJSuryzEBpwrVGVpsEhSXwOTvmP50II/EhdZjRZmL7cPMwN
y/OWBCJsaeN37UrPztvOaavHfGdIEbBHr1cli2ajJoZ/lNu4ZS0pLckbRs+wBrRj2an+5wWBUINC
GT965i2+P+IhKw/TFCBUwfRkIIvHud6lDpdW3x4SiAgPXVUcA/ksE76iBDYJkH0Npd+pg24mSzci
gLb+7J0iCJKKn7gBmG90gKDBdw3QcLJ92CMG6QDbKCiUc5NA0jQpMsWW5wztx+4+oTQeMk8Q9M8i
n4wtNMsFz0K9IVhHc8e/+XV1b8s6k+iG9vephCqsSfhvp6W2gEG5my5PfJY1DGOBCI/b9l8sohar
q94YA2MmwhdcYbJRkUvQuQ+0dMlecfdZupM+qGvCSxMLxVe3e8L12sa4+QLoFfwuxXuiSwR231LL
EyuTPkrA8nrK6dwT8ICrmLlv2Oxo5l+wt17CO2wEl91nsdXats66GbladqGF+gBTGy0Ciw95vNQi
VN0Fs9nR9W3QlIIEX1yn295aZKNIg4Z44e2sI6SsxORaJ84HuWakAnVjA1zI3cnfoldFSxRtmoEf
4LnZGeZpjkjpPTUYbv2vyV1zFktmtuf2ii2VMx+Lbh23/2tk+3m/Q5w7z8xh+Z2qPWzoICFOx+D1
5QT4/YHjMpKYiy7gJSoJI4HTM3WVTMX3OytRpme53HkMYNhETyEoWDMVFjogiGfuBa/XFLklqhst
JJxYDGa17yBx4kCtcpbAsGr+LV7nj/jjMWURcLH4YKriYA02Os0NJhylAeXStx3JcwWBF5cHN4gY
Y6eTsHHjflngA8uC9okLw+lKC1f17nYmKa26QXeWWa3jBOM4SXLmn3YB3erGvn/XyQEoYWMwgCMy
iihOMQKL/1fe5Epum8QpEg6Tbmjr52OuxUnqHDzV0xOfmXpsjf+ZP7cGK0GEEG8l3fKzeINn9YMb
NQohK6mGpMz0I6khDv0J37HDH34Svdip3itgHTX3FTai2RZBXl53M7Nme2bOqI58mGtKQ8xXfLba
Y5UezTnXaXMTM0Fgj/QaAoICUwbMnTopS7Yh7YdpLCdLNZlVLrLTg10Z3KK+J4kWgLQwPr0k11uW
V3mUCgUJMcHmyjbOEIubC1qdSpYN+a3WouPybUgKEuVo8XSSJGl5yKKKhCBWf7xbmII2nTHoRYjS
4dUZ0Ys7FA4OFzCqiyWq0fE3M9+CUOWyPrcefDG8wa8uMISexhmFeiQe60+TIuFbMX7ffOvPXIL4
J9vldfJ5cA3JDzZfXybAFoDnoLSxSKiEvRzIbnLLkZvaaqWIbmgb0l58g0nfOoniowDtuTsqAjfU
xVkaFKLjY66AB9OZAL7H0kZ1yaAdzoW2xVe7sJ7Etkv/3AmeO6cr92+7aotQN2vvNlZquhm21PKM
OoPAg/xDu2+GCBKCkHxVGznwPjIkDWJHA4CtjXXuWAPId3LUJA9hDFDgxunO7N/9OcOWYMaaNS/l
fHkBWsL5HayLB8y67O+V7r94RZ9DM2wYjQM6rrvBUZz07co/M4WAHS0FqSxC/aVq/hCbKauF48kJ
kjprQ2kw+JLS4mralDH4mmuBpK3Zk/Ev8eB+0f7G1M7tCM2ur5UCrlDEdlvVsjLEkR5/MDUdGhEU
gKYINLHsttRWIXY5OTLERf1U7HiSbJ7j1sohscPkTntgacoafdLcSduQRWX4Br+N/H3cXGImddRl
xgMdTIffJ8vg9aOyThA3ouzuBJAiTFlQ8SZc9fBIiBqS3BFiGQSXFUxGsuuJw9hknJE2fSqhBMNa
H/7M+CT7XUcGAaRX6Sj2RdxaSDqe8/4ZCKRoRzda79RLV7FzjG00CYctolaeiOuCixowZ0oRq0P8
ahDIadU8qTVp6BU3rYC1nyzpbtV9i6J0U1DCRxvCVLO7gtf88hjyJMx4sl0oY8d7D2pTyUl4A/qR
RPLNKqOAMVmL0eRyDp79G9BPrgboDjeDGYt95Ruj4EyW+o3UcGD9gcVgYbDHPgTX2z179/k0AhYQ
XEOrTo9aoy4xEVh65rSN0YN29po+ojR3Istikae7c9khpkLpfMekW6iadmI4R4A5D7Z26gWqgSj+
0iyBdkAydC6ckH0I4hy0HhPwrIOzYaLyWFukT/BTxpdJmFeoYsmIOTqPWCjF5kAYctYEldTvSLMu
pSKIH0T5UaD+/6QdAWaZBWUKJOYtDnlehL7iGJHlwqla/3/AuGCMX7AOOeNECLdGOwcvEI1JwwWH
7+xA9Fl386Xq4RT2Puz3WQWOfgiQ0GIKoQueQO5Eide+TAC+4sBpVOC2gCVI7rxtLDH6RqLRH9CC
k5QRrp5VKQTM+kQu1qt+wDaShB9Y+nLh2uhw7bBzQ0qMPKsSLFx32JNly03eHsCgIvqr4301jUkg
G+LqQbWUzTUpRN1Tt0L2ZCHODhYv89ZGlI7sxgHiVVsBPrJ3nFb6w5Kdm/a1Jn6SOEnrN55yRbC5
+fkbA81Wu4rhmjZWOMTmEz6ZQKTHz7oTgAA5i7L519rt1XCjM6j1QCF4iEd5TcP6rpQz7VtEjRLA
xoWP2P/T8KlJSJQmTN5weFHhus0PAhQHIebFMmQvfhpjXFJqtlYHkVqm7W41UqrBdkqo84xYVFR/
3J1zGaFRHtcKupkpPAM6DU15IUKw1U6UjeFt/s1emyyr/y082ITDkzCZDrEV+TMtRHe/PIDwrEOP
yWiB1GiBQOAzsRCAp7YHVbiFX1Mqt6NHXZcDkfufNrm5p48zyDZVBxaF4V+HFJbEI9hdfL3ltpKd
QCOBavFhz5DTGYyW/Aegjzq7s0oSx7mCeUgbyoXbECdt162lGHcb+C0/+l5LoiX7kPGxTAAGaXX5
fkv4UsZVW2Vwk6ExLkfra81QEi+lubbIjEqdYZMS7rPREvhH1FU6JppHX2kNT7ZUj34h1MhMqBoN
SKdCKQIhkfWm9jT1/B/qtmamXr6ZxAmzN3PyWBxUkPAFP854iiH08E2G2oMJyUfRSqMsZqIiauaF
/ilb8yi8d1S9bA4d9k3TkugdsR8YHBVB0Nne2q1f14X2D/npPZ8Z14aYfnRsPTTNj7ESgHsj8TBH
SURbYyNfikbu/tD0T8sRJsxZX+60+0TVqeBc2RfF0ONmbgtU4e8LUqFn/ltnA1cNkumIzUiQN+LW
QyIuilbGWlfivR847ZQOiijq5lsWC2jUncs+1zxmEn6dUqwm00lLfbjuakIPvT1sPLacAL3lszSR
WOZB+Dse4Xgq/kMl+8PAuLmcdcasKwUthUgeJRSDLLzbycaEgJwqO3O3GZUB/6atPoJg/zmQmnCT
2jmj9DS28CNi3qv9uA54GPi4MMrLlCY+D7qLvMv6AV0y4f0xcl661UNKHHL3Gvl3VZwGctf2qsZp
T9i83mj2kjpGhV8UCusun80tOYpHn2nubc1pPKe9Evd1+vY8OjqXn6OQQsfP0KCOMHL5pW8LJarE
zZR4Ysgdd4NVY75wKrzEyy3z0rYWQeW3VdeRXFPVpa7IzgsTCxMiU/b7WmjbKYCEeQrURP+RJ8gG
eg01HMul+c3N/0om8BThXju4ysiHhf2jmLijQU6q2R3dtrOc+wRPSXSq9qv02zcPcLlx1bDZ/Fpl
B1eN7ImNX/AkT9QSvbfcBDucq0YqslMOXdsv6oGa4TcVpHe00F/QRC//d/L6480VqjeyH2xVP6X9
sX5kTvw+KRGiKOEjeaMLj9C5t/X2c/n/ML/WQsDt7CL6Y17gEhWhvBt+cNvk7dRYyEbpGC6myHCP
is4/lQhEQSGW5tgSkLc8/AVGfEiCTsUhVupM+wk/RsFJ8XzesCX0xm/Zkan6ltQuMR8tHanGrXXD
tAYdNR7sF5guNslniY53Fy2ZG3+Z8QKm5T8t3h6ElomXFS0Zfu9Ys4a/5RumNzMMSUnGqTUINQSW
VsPf15MmGvAvcNHuwhURHM7LTSL7MLaUP8MnYjcrxPfDPWrufvEzAdROyJEzjAm2f6jMBpoJuJle
4f5PAi1EXgpaDlCt8rbKmivOxJf5AHPLbrax4IB+m6o8+JwCI3inALNlJ2njh2d0i1HLQ8ukmDRJ
sM7xCD30FTqzof8IBoMZZ0X14IL5hjczq8ClEM60S5JC3RgODYe4tTCacHO/PO4vlfOuzRvSbjom
0Oo81EvyGHj4QGi5AZ6D3HiAuw224Yp7f3nWQTILdJRjxQkRc1QiLJQf5RfHHPCdmie+Ir+kmLr5
LMI4P+ti8Jl2Qe+4xdnUglIEq/qKNAwRpbay3xZGf4Nph7N75S/gRKTgSKnBMHffU98sgyS927S8
7VxzgLVWE16/3hwqfB4xOVuLafXmB6VSxjGnURBEAZBuJQ0B2LENoLu5rmB+Df9JFq4mN+vrFyMv
VqK9wGOObGTmNyKFQZY4P+aC95Uj5jRBKPOr2fFNPo6NM6daH0cwwnWxIJKT6x5kbc/oRgEZBbSA
Hz7yRiNXyikYg1xmf5zXHAB3nez+gelX73SiyP1HeY7D2nNGzZQLvpd8E2ljJQfMEKYqDC/f+5dY
yLDf26d3AhweReSDLlzQ/NK5/KksYXjCnWuS7ECe2/pvDcgA9qYlVQO3S/9hjq5bSXp+cV8W+Ud0
7m1zxYR4ZsjT7AmfZWspTrv6NSKlLyiCDPTcCH+uVPPn/P2JADEN1NWWZd39TzOeD4D8e1uvmZhE
qhTAEdTttWh/IbO4Zmlv+M/rB8rJT3xtM7EtGAAQYaBnzqdZ3n0KFm3ST4bHa8yKF+xRtb1Szzc9
YU3PcFuOZOQNtutp7m4vjbE62Fpfi45iN0CgrYyOcDK32DJi9OceJUjWX+DT9r+pJafls9lZW6Pj
6Mxcy80YuOOF8/4PAR0rR+3Pi5XVfl6OxFUb3vKLBpTSdpo5z42Fo8ZOn4J2bnyXMt94GAl79nJr
/+uEZL7AsMdu4VjQS6uPNIAqzqM8xapzTig/2VqoGlq8OztoLfpHXevXZ5WgxJK2qiQmRcHW0FID
lsTYHcrAWOCOqwDBg63U5rBiRyGDFYWmBdw7rCOoiSKqKeaVtjO2snfh6rEupIJjTqNFe78VT3Mz
zuhuqt5drX5YYoEahF1B4wT7kw4oRqGCxTYKFyaYt4mSCN5V9/fYCJxU8eVolXm+KLzh+dM/I1HE
3WXKBFkELBJI/n/t7lsTT0HKp1hwwE8shhjx6m9TO6NaJzb1dY+A4FyphSzvfv5V9XfO8R7IatgG
Qft/Hm+asComjtdw8yRR3Xi/fuC7YGhuK6jkypGzJ3scXm/n4rl2SEtOZ6nm+s1NHr0HePj/nvRT
b4ooexGE8k8KBs5yB+h5GY38J1c7TKdsWrtHwj4RoYVzHHGmjiBPqzsacTAutd6kzbPxg/xZ2yEM
HpRDRC3rhyTpBLIudx/4/QUxqaEgBWYtb3FNwNhMOb78fAdLhbWTSvz07WTSsffY56TVAksGX/uK
JzeGsRPtsVxOzqpOOuNJhRtMRuvUu5jXm32zOYwBN7jAgD3eS9qhz7X3ruhF/iK+COLfIuU4PePo
5Y3xc7LbRuaytGOUfI/yRWaqrVwo62MnB1P5Qkzf88rUEUSOG5DWxQ50hEr5Bh+kfJdWgxDPjsdh
L6U/WeDSBEoL/J1tuXvxqvcw25oeSGS4WnPHS2V1LjGVu8XX+FYMRblMMEbmuaz7Zn9SeqQaTaA0
pVkTzdx0Wda/cRryiV9EulDMQU6vnib3suqXKLldhSTANQwpWNKW7cKmbVhmSC4kRCmDPfi2pFGR
R74voyDipS351EFKoRI/9oDEwCzYBA6p8RVZuBJV0vzqvDvqPA2nEIHxj9SHzVzC0yWdHdVjvJD+
wLwnZ7Wgi5i3dD+h6705yfyjizacoY7d6vOokfXbow3asofraaG9YOChhQV4TxVDXkYp19YEiWeD
z/VsGnraL8cFjKtbaurFFk3BiW3uTIR7x0Mu8Ed58YecSx7hdgxN8Yo12mWcu9eXoQYCJe3PYwFG
IQUzH3uowudIAs5eO69AP38aYTwO++mBVpKpaSbxm4RKz2PtiTU35ahLPiCHn6vQ5COdOzvXLint
gsIbKVt1wh831uH7NdOVzxeGMKpuCVfwOFhwFgJiQLHNUZrgE34iBxBFHAU4sPy67nO+vxJuapvb
9+ddpOlS5gFFBdu+xAubZHsUMNwCyKjufSQtbxvOSrm4stbjgSV3iaG8BOygwOeNmnFlLtnROKl7
cX+/V79Em/lRek0VZOyAuQv3sPJ2K0FKndfyEOQBsho9pUQZCUS4n6FCBFoyr4EHaDNsjDva2bBX
jpHTw2ZpwFiCub+mmAIKBGeyf/tkvOWwJeg4UfUdLbyN8zHi83wr49riNAeb3caHMOQadzc3VpXj
qNT9CT/K53sXhZcfuoxBFlPoUSRrFXL10TPaPSgKleUISU5dhZpbVYNIpgMrQQEw5maoIqmrOIOd
jrgONslArXWU9aXpjHKqPSWVHGTjuCfT2iecyxmu0Jqysy7S0/+PDhzloSytPeiS18xWMWZmtSGD
dF2SWK19S40i8rHa8DxMRO0aEzfKnVXkX5K/wMgrl9lca8N7id989JArqVeXbiv2SAV6tjshkBw7
69k9nfxKB7aefAzy3i23dlpb9DeU65ApDelbg+r+iJVy3soQRuEYidB0IYsXjKvtP+PSy9cO+mLr
cIOEXKNg438mZp77vHNXJWB4E3bQBMPzan4bpiRc2td3i5+3LlzXy8nIFM+rqB9dxDvm2oQX/d3L
X6Z+TZc8IOODldmun1ZJQmlTjRwpUhIqegXS30bR438OZhBavHUFX7VRaXY4ZIZhihujHYf6bELO
ice9WRFnP9oai7fJAYqBhePrqSOFN8CC+0QGjzJqocR5TEh2R+rvVwq4IFyGWESV6LOABN576fQW
Yu1qwgOCF0GlGEEAcKW4XPumbHU7vf8G9gXtfYb+IzAqmwxOVrIJxxNf8YQkKDvncAb0EgVOGuFT
vDcdMNHCvlFk3fofuQVc/iaw5X2jdjV2dadCO/anNxzU72ofvOXOFtzAFhE3044GRiTQ17+Zp2oz
ruIOhr9q9fgIfoKUqa9G8j7/gteOy76iNsw1ctVsmLq8bdYkUjOfBIrGTK0GSYNod+vj8AMX5qfy
h23KRndX8K8ZnuLLjrs2UhNee1JbegrNdkJJFtiW1Xw8CznrmxsPwWFwIaNO73fGl36/ipsq82lE
gP1Y6iloDTUX0aGWUbAz9c4xAutu3yixK+k5DNctf2O58+RzlXZe5h974OuPSxVIFDttHEYHy5Xn
y2Lvr0Rqek0uKWyhwlLzML+C6D1ZtkUfaL6lKYaTWyCrrGGeRa2clX5az23ceVRzLsh6s8z4lPRJ
nJKuHGMU2uKgYeryQgG4Umt1Z+5l6z3ih7OMUKRz8uQGurV9+CoQ4CQClqhUBGPrxk60lGWkE6jJ
74CdCNobsMbzSzA8Vgoo0uLoSswLu9rDx5DypQG5wWTOcrAPhvhMEtEVCfMfJi2ui1OX5jovW+uN
LXVlNKWM6KI/8Ed/TQFIBXfNk1zk9FkEXQ9xfcdsC3CuBPSBAUxuZySc1+pNSyzU6L8E9wXaEAj2
KjNm6GeK4BUc5cTDHiz5LzhW28SdneHyrNl4IfM5c/q4wS625f6MiD/jEq4khSF/UUOIiJ6n7ynz
DRIFVskcIi5GOQV2CQvaqlxkw91zyfvTiXkC1tYSsW7oT6LimN6m9cDCURnczmkclloLttqETUpC
tFSRxS43UEv3knC4OOvHs0CLHpx0/gpwXbgXxi5v3I2bySapJl0BlHpq8tqha09q+ljxitSQIn+T
t3+JjSpNhdIR/bUYL8URq06s9jSLEfND2TsyR4ycWVnfd/GgOPVzXEtgcFES4kFhnKOSi9S+FQtb
3uhSkboZLuCJMn2vXpDCQ1Bz+jewQTsT2oS+51VcdrlAjU6G2x8YnCva+xM+8+ruH0SsZRoHPYW0
EZ9imtyKSM5axfqD7URzfIJCMz24YAAqDsKXnWSztYsejZoU6v6fa3RZrT/6JzVx7ocuiny9aIgr
3gOZNX+JJ7Orv4y4GEhGFXDxPaI9wk6OuwkfYi+Rg2w6vvlnCTSaMsVE2yVvUtEginv1Imlw9nij
PBSdNDxE1ZOpFUgRu51PxMAd2tjDS247I0Ob1b3bdXCWWCkZvGXGcQsH5jHYmYB04aBvjGrJSJxq
U5umcw+CPTSGMa6c6eEt/Fu+dOdsAwaZ7Q6u2rKog3mAQX2wL2PI1b5XGpplMeumbbPlSeMuR9zK
zUUe550ayHte/SufhnWkgI//1NN1CSi8eIPi2E976ymIam6Mk9/rq/bET/1ntgLmOxkWlqI24omg
SRrWDug6SgVeQjTw3ncenFZSUJYm2EzpnxweS5pOEmaT/fuzI61G9aUnVz1YF+qcVO4lp0+h4r+K
NRnMR8+eEVY3NCWIyoqrF3G+1DgpKnknUQUCjUTcKotUdGesfa+oxaTFNBTopURIHb8ifmKn6dyY
LI5B9hMGEOLPibxrWakCNNOXqVJzK4bYTcDYaKxh3TWesZoQ74n9yL+/63h+bJgI5kqHxGunBTgw
FTJNLUVum5iGbShMyQbVn4CODzBVTn7eT6DN1JlAnGFi/Sbb2SjPTb3m3uQNMjLQugyptR9vmWmE
ddx1sHBkboGdhIav46LSSfvrHuawFWt2XCu377g7XeIgO9KTs2HOBxAgYuElIl7jEzwaAA1+y6lO
hLlSM3Sb/G3tmV+8/7+3/t4kvQJHKe84mVYjVQQRSZlU2zNbKu5I/RjweJpMhsCwdu573Nrogmly
CLAD0fAGy/CYHaJchig+aBAqh2EVVdMA8i+fiDZExA2s3b+lZC5u9TlXOR9yZfzeaZK4FK4kGLs+
4jHfc7nMLBV0CsnEezCryc+/RgDNv0UEw+CqhXm1tpkz3sWGzRQWR9uhSm4F7QMXv6UbRhD1kIUN
6m9jl+EOVA2dCAKyeIHyqly2TbFkVgRI9RNEyyj1F9oUdIL2vuHnr0RR5Pvvq+sAGwPbDaiAgUIi
2z6cNzCVMAhWOICvWxabHrRsuVsmMZ+c/m4dSiXCyiSb9XCetEhsv+myXjodSyAmPiFZan0LtbEP
h6o1ZumqDdzxrYN7RkReSsXVX7iAXt/0X6f4nV5YMkahuuuScLEsmoQzS6r94VGhbZjmI1PmLYZr
P/CkVPYwIF0Vannn3rn9bpn8EG6r2YAVdBWSKdUOuUEbzEFMiQNNIY7hSxL658x+ahRxlU9DzM/B
Bjok63udkMc296/vOGgCfT2Rw+Ojf1NiZQdqVcN4tHyMdGghc8HvmC9T2ZBHHO0+zukD07kBDxut
zFlg6I1HEDKW4fOABey7Uv1IXjCnlBXgX33/5QChMKdEZpRTGJvZv6bddz4Mzr4w6ZBLl4MYQE1G
xV6A00RRWjSMVNVvOLU7kp+fE97JiXlATwvl8ovXT93kG714LcLawBMhSBNxxU1DVJSdebQJ59E2
G9sEYjgZJekSYJD6/NPBTueDgyKC72mKqKJIw32eJ4KjICdZH/JLyl6slNbv4ZAwWTETqAkHz0Pe
AKFGiQ4Dkhtgdhq9x8DZlvR5PAT93TfAfLdJqpsFM56zgM6VmgJDJ6zxSxFAkzEQeq5noRcw8EvS
VY6hGHgFW3smgRNJFeu7vjdLd9aMqQwBj8vBNeVL8oHUHo4wwJdD5XGF+gAb/t/1dtpB6kttw4Vt
aUnAGP4jN2jke4jXTbjg1ytHmv9tMbi/1tk7QXyL9HgAZQ4m5S0g1X4hUBGvjV1wJBY4h/vfL3IR
/CUC8Znd82Yy1Cu6Wzv2YaxNrwNy6/UnwZhznOgXw4x4028FgCKC52wJmMTBvd2qVa7qA3j5tzz4
gvtIXDvEV4CoFNrnA7/XY55QWrwvH8H8AlYc7ejVInMfH+68Rz+mnzNQwXZM6a46hlO9rf3GMUSi
28ahqYnYZFzNIJJAXvg635gC9vRF0YxuAPUaGmxiMaL53IY+qnhvQotLrMtPrVef4e4Kk7+9rES4
vRPUUOa2Hzbsi0/9btstNr/Kj7rynMyAWRh74jjMSgxjzlgPFCo6y/Gi7aIpki1hcHlkUOimWyT7
rp2HoZnwFKcAzbZ3wi7Z5rX0G5pQgGtYBnpXIYXIe8GFs7eLqHT4es4/mnKqT751gaXSn9jScISm
h80N274PqeFVX4xbA0Y8mZLupQdH3eRTz4EKdgDBs9Zs3tENwTdYzJwB4EwUBryspi3LhOJcwSgG
/L3iBBJMBPA0Pqn5m7w4X70Ay16xwFGSv5OkJVmNLti40gfACtztqDcr+HzhzJrt0YnUCVg5ahta
Cp1oYgpf16Rm2hh0hzdztSffG6wGMRo7Iyps41iN+vm/FJLfkSMJGDMeQzi1P3a6WEUp3/xgtI8n
o2dkgrarRNnN1Kc4n8JnkUt+JbHgM9eR4efouK8XQHk66Kx49jPKUILdbYnAFklf0T2g2Fnlql+m
56Ar9cfgLMbD6ilTncjH6dx3W5VSf9Q+zQw5OnatycLWqzVwSJYF4gRyouKO+0SMGwgcMJu0nHut
WcegvxqaCxKIh6MsRoxkFDfgXSioQc03vSIefBsM/oZf64g9Ym/paWNN9QYZpse2SX0pxknD2UBP
4kLUvdNSMBloP0nKc/Soi2sYpThPFHctymhlnpAJbRTuSIfCD1owl9+jbbh02dm2Myn9Z5YK7oP6
rteEyWvv58sN7D98DvSCWQ+1miqvSGqOYJzK5v0w19KphXBIFPG9bU9w1u+ozA/5QWdT+M0BJevd
b7dB6DcIok92/IjiPA/vJbIgb7JpnFOSzjp4xl9ytBnh/pXCruiJ6224gd4tEpgY8W8O2qXP1xy1
6WT0OBZBOXpelsdid9nbR/unjUKa91epCVnAWFg+k70ooJvOIj3D271GAyawnPAJBASZjNNvWaSi
wa42seTyWneuaD8yvA6U6aOhVNnsR+BqkMs+pQ1HeGmPSFuAFm63yl90J9dZ9BeZ50CDo88nOxUy
yDm0zSART5vb1IrjJzNACAmyxmzcZdNFXkw2NNChsQy09/jWRQzMEMp27lsj95FerZHZzw/PZsnl
l8iLmQxvPqftqpbbvrO5tdGUnbOzSuceFyZi27cDvl+CGv5M7s7e2ZnGtY4nD+PSoGreDcuYbhZb
jtvAruUBum6M9aDhC+G+uVJz0R3Hn2YojalBWg9lebbw7Fxx9lZKS8eJ+fvL3+Wu9M7NLUblRI1V
rgVYl17jMtV4YGEH7poBSGDFkoLqIpBkreJyXaw+6aKXiMjphXs8H7HPUk5oYczhrcdA8M4U6ZVc
FiTIO8lPz9g3YIE9ZIt/umdd1JCohJOgLirYwuZhVvhORM30ZIx9mkJBIePO52WtGap67ekD5464
ibeS0q7SesQvxofTUMQGVqJ3usLvjbh5Kkl8qIrgUWv86CoiiNd4Iv5+C5nrkU9u8CoP3VuNkMMl
rDCtBB+MGeFR45nb0JD4dFBpCOu8kEe5RUB5UjNU/u2g+JOKJRcPAGBePUf/zyWOBYBdUdvE/iLO
0Vz8d60mGGjVrjvzzz6Hwx8dA6zuLXZMP3AcVzhUCyw1czSnZp2CLyGt3KfGkvyylx5vIAB0PRaH
bJvXA12/Zy4btx0e6tcgdTy1UIYBkLXtkwIIt3VzvFz15hJvr5qqvnbnVgeQTbzefTjumdB8s2el
6aBWshTYJ98fwuydLS6xWh3Q7YbMQiNJ7zqZMuDjmnyvKgC608ukVrF9O0yjH3F67+GlgKSKA3zE
n82lwF5dk62Ih14agP5xTJ3tOHwZ0aiJc/e5NnrJDmd8MYKSshUZGyjzr2iTOjuizyznKDROM4RO
DxZlVoLJ1zJqCecNsLCBmbCHusL6zB1QbuBFNYqMbNxDg2apACa/dFbm9aq6mwmXhqRiAx4sUOdP
3CKU7scKf3gxsjD+1KGTRiuf8HHGhxZbvzhU7CjyrAI3RKZtbGDBMv7aYwUxXJTDE1aLKPxL6lj4
RY1J9JVeXSQM5xU0j5icppGjBpq23SesYUJuJAHyMZUnq5w/bFrUX8/mI1vSNzyXwUnW8NVr9LTv
EffCHRXX0APQ59FqwEB8ONzRJ5fnqg1o6GSwzvPYzj9/FLIythIlf9xVEEZqlbN4NTNYMFraFNe+
Nj8FdAWigYp1jydaECB6Xy2Pzl7gCeP5yYlbB9DncVQ6Nji/uDcxRk2Bbwp+SdqJr7awbxljSBZg
bry2OvT0FT0jBaCUul/jmU//P1r3674spAxJlQ1nYSDOZsGFNuirfWyCm0u394RQDKJ94qbaXjLs
taXhaiU7C0LqBxEHRLkcN7kGLh43MomM07Au39vNt3agRcbk/eyrPb8LBakBTso+6aHVcSyGWa9T
Y2airFKeca+cC0Id7+Uk+FWHMnm3gmUQVAzqlAfDABV1H8D2x4L560GwJzaAJVRQqeai1shcd4yr
YroieGb4N9Htd4SvCzZtORS378SNezF9rG+die8rCqjwjIdG1dN7bX07um4CfsTMS1xPcm3xV4BJ
/oA0UX+2erYj845enSn337DqP6tGzgthfPicH/EtS9oKeNSINdO0qE0t7ZO1arVab7iKH7EHX2I/
RNhX3rdfuIsv7CyOLO9qLOFWY1enYtXBR1GqNW4IRWmoS8wifYZjmdag7baqSSPqs9n2AYN5OYTG
7szw4dM7hx2+LhSBwdw1WsGOrOMwnIR2b0SoH3CFjRZTBVcy6gPEQUVRzDMSwsK2u+Mq60eAxyX4
wYvd0Wr6aA/2RWFEkmPiEVsmLi/eY4f6f8LF8RXfvb7RUQnLSKetY0MmTzuR5u1/KpSeepN6GR6o
Zs3QUVxMHkU4qhuFJ7tZHdUA081kaGBmtDaj87FVhkQJcfBM39DP1XOT9stClBVDnrnOhsz4Hsof
TAeZxrr2oD8Drt4ftnvk1QvkgIIwXpMXJfsPsOOLaL6rxBhdtwYuNk1awZC1fnmAdkWHEGIj3387
scElBQgcVvW7cZl03XDxCEPPzufgUNSd33592lqJ6IzhwO7/vQLNXLoTnhvwFekbS5PWFsLi+8Mq
O1dL6hjgKjvB5Q9U+YvWhY7lseC5yI/PjLEM/gMxcYvsClO2xpKD41qwH5r7R10r4bZmCzMkEHPV
xHytJ0jG1IZYvIHYtp3Vf3U2R7HGEW4S5rkjiUI7IxDpU9x+R9M0h0FxUTiDb8syzU7gUOXu2Vvh
HO6LhhhurUco+55TtR5bPr1mVrVUMkNzM0DdHkmHNI2CgL2kia8QNZJHhMTNfQx65/I5bPp23PDD
ZUfKXv4wdldzbNtPdw2vg1SSjShK3I4L4hXyZPMGdosGFSbXmVHE1OfriHO5jYDZyM6DMs+ztQ1H
hSPGRfgyc8JATZsDBP2PEqn0ltV+MRvgNKaeUdPZ9h0cIwtgRQdh5f5nRiwsuQyqdyq325ynQH38
hd5FxgksvPwx9YDHxhItuUvDKIVrNWlnnEirB4b9Tc8xoxBCZcImmgQmSKOe2/podjX6/JjB5bh9
3hvtfyuoM34Ffy/z4B6QJf5JI9YAircOj11jfdQctcimU56eGLU/1f+3Cgmv+5zFlyxyLQDWKTKy
bhsF1mUlLFTb9gj4PE1/dRIvPQ7XyGATyR0tOqjQ7Z8QQB6lRN6uCNcPKq//PX1+OGOpsQYGDahY
i1y6GrsgeC0Pv/QUYkttEma3i+9Ht6lbxk2ydmNNQPNxIoTrGKMBsTi6xSQwVLQgfBUhXu0DmPw6
YRB4hXoRfDbXPjOzXpD/6HZL/LW2REgEbwwEa6V89+mUVhCUKgChYOkh1GCIQ6t2BpZLa7cOCG0L
v9xdKR4ZoZyT3sVJfksHtahNJJQhUYKzI5YripsxZwIVmS92dVxDgCGG04nNrnGMu4TJnyK5wL1M
dUpkfDkY3GMY7ZZo7f7TZW9VbbSdvk85Pu2NuxOGPhBjW4PTi1NG80tQdYpprqrDkIpwPhydBgMf
JabR6IJ5moO93sqrvExqHkxNqbf/te0BH234Sas3HznXYhfkpXwNd0iUQR4VR4KU0eI0p76E9TRc
+fYQNIJN2UT8JJGRpYiIkJRUA+GqrxJXVeNtpOydV6tjZgOr25XoULkDIoLMsT+dbF3rTwy4huBf
LzeDwkcICqjplCujFuZPopdYKvbxHI3DZuQ74/QCYiwUUlPC79zdZMl49nhHJc3zIVuKJhf977u9
aEcxdTw30GTEkaSFxY0zT9/+7gKu+c6NJ0hddbhKzrkwzpP19/J7yc3glTFxhlUxN2VIEX5+UX/7
wqAPohwvUH2fcMjeSH53EFhRfVwU3jzFNR8b4ZBwOF0jH6oJN5fRzPjMnwqpGQDpR7sG5SRVBftZ
2VGQQRovA/K/8ho0Nbi1PKHWfyUtGXepLP+Zfl1bE+ooytMK/zNUuHkezEsGgmtUZhD2ppPmtPp8
YXlqktwhwUCdP3UPJbWo63Zs+V1smGVe/mBO/JkOPsANhdXznkRbArkPxwxs3DJO3Ph8N6NGy27Q
WK+k1d6Ous6YzU7oocmK4yu9Iah9jqPbuIbzfZ1jutg5pD5+PyiR/cBeFf9n70N18zxYkmyPd5Kc
IJI+5oESU0Cg/2lFuavBGAyC4hpKg4qJv2tnmK9K+yPo+kMPhCFCCmmKwzJvRrdSJtYGg0K5VP15
yiTOWQPm5/zplzh25Bh++uR0Nezg12oKhIJWbdiUqD/icZBTwiNGVcXPsRLukKXrVO1ByP10AibQ
sEuLaZtsnOUyPAZ3WEOqwFQdJykXIIgXMwA1XJMsMUgbFcTIozzctTQPl7sdZ8f6TLtUDFGXsZMW
Rnvh8vXp96/U5CARu3PGwCSIlXA0OyG0gJfZ2Co8U7+xzyJFV5IdjbUZNaKTxtEyhU79rdZgj4Cl
LZu/7ayXddZdfXKuZRkrvMB2fp2RXmHUhA15EyOkTpi1JA0kdCZtKYE3jp4G4Cou8PCXxDqsI1O4
/yMgZs1ULls2ieky2dmJmQCKa6oTpSsA6ZumIbszFitwhyKuJhMin9B7OdrTMcr4jh9jlbYqWQ6k
otnbeFTz9zgzJjvbNb9CvcOA7xsOxqTN/sMQO3t3QC+ig2QX2cCJ7GHeSs3FXuFCdfUnO7etJ4YK
4MoN/eRQ8ZSbIEJI8yf9r3nhTuei4PbNi1pBhd0RgT8n5W/aKdbe/35/s26ZvEwfMJ0SIoMeCd93
l3NenASykBkNIa7D8FROQsHBo4NQfuZUKR9mmGRbYkT1MPVlHsW31yyOYmHVQm4TlPzrMCQ5Yagf
3+rGKsNHk+75lqbv+5Z+d1f9FlZV7Oyj2ivduNpwzkJ9iyZoak88tj2/zXm/iD4gg0m59Fk8t434
z5Uq0ArXDm8RynM07+vbjVGe3ktuX2S7qpagSK+oYm4Jy2fI0wibB/Mk6ZuBhDgp8KQjB7i+VtTA
WKbVKjj0YGRsaYa/4HsTn7FGXk+knp9B3xwFfllNg3Tlo40mEtEaQwHY7Yc5SJ7qYsAtaJocqbBz
TGgq+2f5u3axuMog7Y5wBI0MnYKLPJ7ehjNmfi0nydR8a0IVTAMMpXrsFbrwoE5PgWEhwZUIOEeY
xjXd3jaYwOyuHJhNuHrPDO/PK3T//3BVnfua/2ELBYs+h1wGJtDg6gTj2SkEOfGRbsDv12sj6isE
esWL6wDrlQY/tHLH9XWThyIqpyP2tmHvfj0/nCEtDE9/Ax2UrinhPYt3cNYw5EoMV0eC7GEaVcKY
FGBgMc3za0Tjr2l3HpbZNvHQvC0MWCtWtt3dil5MxPlSTWdw3NnwqjGIMdsSZSGxZt0JM6R/BSd0
lOW0zVMW0u/9XjFQX7IYJ2XQMrV5Pj2OyPtt8UH8uUdDPCtJvg/MYmpFcayGPmXUNs6Z23bMhwKO
bsV+78HjdhJJpiYC0yyGf8/CP1S9M8SWLiiL2aSC7Jj8+tUo4ADKNBGzbcLW63rQ+mbdSvczmCfY
wJFgrDbiiLHWpTCfXmRTM24zYahIp/muSKxYVVBQINEax1q1kp4Z3T7X7e0MPs/tSWxeKDgQSQak
bAl062dj2Uo7qUOeHHvrbXpGEMcVI31uUGZPQLwqGBjQzG/i16gsh0UrvBSh9pvhMV14fcLmtc6J
vO1sxvEVTWjkCewcKFLVHWwu1XF5AG3qCW7UjMqwvaJVXlt+bNLjBdbVS8dIktykNYhC5bqMED7q
keg3WRzaP/0HdsxAauKbDydp9zWOivcSthnl0J9oGbuTJeJ7CZxPXFxzakN9fl9oIaw7fT3WaEcK
PTTvkl/L3Y2dsJDUFysAJLqdEm6ZrXFK4QzMoo2hQPAgtmheRh4AtMk9V3RwopnU/XgkzkDB+WJg
yyBeFvG2nnL7vjkaStTnnErhonS0kg/QulAEGpjkIpp/hI5goQ/Ujc5hcF/2lw688mvJyao6TvX6
ZOIkUXL98t3P4mZJxlV4IUp1odVKfZkrSzdWXEz7Nud9okt5E72BBw06H9EE7HCcBvo7AinufnSA
JPGRwcjPjadR11wnOkv5Z8FC8Vj4rghFlQsx4jXqSjbVWLLNfSY4i33TR0wbIeqllcJ5tIUyLQXo
ioSIBO8SZ89Yut+UO5FtbkHfzeNlP9HLIuS5xAyiHiyxUbPDSiRxdZIW/tODzJONqjMyp8KFAnQF
NB0+2908hqmtAvPMIgaRerTyblSgi8zFnPebCfDp8rvIZ764+EaqDtZCJ/ouaMJKq8K56FAjk8c9
TDRZwQWFvMbrpjV43VbDIdlZUGmU6f9FtP+Pz7YabXVfJjFuJAU4W2R6TbFnrcfRxOG371JSKKjY
RqzDedclzDotQsx5B+RRCbWS0mgDrixL8BKMvxRyKsTFR2CGgn92B0v9mBufs0R+O1lIFoRxmGkE
c+HG4awqZys1X+2snzCW8WVsLNv5LV0kYMcI091t3y3qWQ7DHAeRMzxBRSOGqJX7zJRvz4v63Tkc
bxtucsGd22wN6llbxtnO6YlbJW1lI1EwdKErUvDBhS9m4uNFF/MFfn6Ax4LS4pgxXZqmaEOh+xXP
EIWuM5toDjDDBNqp7fgbrd23o0N6m7zCaFln8Zue0qzfHwdxH354Jzz5FY6Goorh7+TUSglYa/Sd
dmQY0yC+KBm7n5UWTdiMJse4skJuDwfqD8uBT3g5S4sWdbaVlV20zPk6xFGPDQ6Oi829BALl4oXC
JBjklx241JrDVBXpYIlQTeAPjqvw45s6wP9CwluXBAlRp/CCKHtxH97JDr+5JrqtrUTsJxtYQsK6
w4FxMs/jwa5GCsAGdrhC1x9NHMB0l7oFUqkHzuzKkBLoVNapcThdwgzTNvB4/r44VVAxv9tspjlT
G21oRfKzTd5NkWj/TZz8fcQrJdUAO7+JcEJXC2o/T22JT51YPY1zmIvc0pCQY9QIXJGjyn4D1VKB
Bv317JofsrZKvnakSzObDxq8l5HY0WPDxWyyN2R+CU4zKFqVOc7LWEeHzneKOiczPUR7WxDTMP3t
yP+XlvfHVwGtnFOvZLxI9zCHcT2ibuwatiOzUtXAaPEKq4I05OqKkYeis+TbBcGaapUH7mReeUNK
knX7o6Gj6kV2Ab8q6ZBmesTriSowCYz9hIPGh8/H6qq74Id2V0pgAX5X49O3yV2cW0kHzECqxKlX
ZwQt0524M1YQn662RUB7MEq+tPmuuAAiuObT3kbLIOkH4s+BX4eaziyfiyzg90Glo/iWii6jldS4
PBQleAxwx9TmxAWl6wUXAG9PY1ip5ozbBYU8mnpVDiSWjgjG1A4iSGit4ZrYm2AHBHKrKNKPD5jJ
2zw6p21YyAoRLykYNuF+KZTjZoFIe/mvptt6sXxiz55FNopqxhTCaPb7ppL9tjxPFj48ohYO+4bB
tWasZ7ijf4lc3w3mcy6742Lv860v5Og66zecgrNRmnOyhahu6qIk0J18pfi+rrQOl7CZBXaD2PYz
GcebWe67O14ZqFJBZnAVhjKOFFCMCEJBaIi2p9a95XVQ+aTDduLImnN6JUFkQf+xBDAfcqVzqZls
AQ2bsJ1EzTDgCZhuYAyn+ZwE3LdSsdVtl/fitxhjC4yPiAx8zVDJpgoliHMntnbc88CFJ4kyk4ub
9XKR82i4mIPHUHmFJ/rhk9hnHlkcteYAfQ+6CE86mMFegbgfugIThiopExF/Q09hrISkpcMr0lKj
Mna/rWVP10FNP4MxpbXPT65Kf0sOiA92jOGAd4ajWo74WNv92THPpXpznwx23dQhvvPgA7iezR+c
hSpgfwIec1I9/SpZXb7xS0UfIfB5uxtYLAnMkSezArnl9pAqqJZlr3PyK4SE79THJ/+lSPD+zWqg
+OBkWmUKLx4SVHe78JGfKqK9S+0vucNGeg9AeFvla+sWZm+HfL8yShpxNrLQ5Nmb1yB1DYr8UEAY
2HqIKed9/vta3SKGhtDOqs4Xcow20EJn1U0lbrepfgXy7MCoWFk0GFpwxkNqK3V1eXe8g0NN4VX2
8sNMR51aynFc2Agolzoz5O38KdosQwcyfc1vYsZpDBYNxq4iI83rMqhwlSWwAg2yAOTWGh4UvTv8
VPUcN244dR3o0amAOtFsmx2nKJ6lMeai5O16Q80KlyBtU7D7E/m05N9COjsUifHho1cH0/fiYQ//
NuMdn7Pjy9HW+b6IIO8RorB/BJJYvNqgdE6zCB6TQOQ6KkJ1aoahPxVwHkyipXv3N8Db+s3DLEfG
N/8jPSgKY7cBJE7e9ViXHAyxHztPzbn6v7jtXIP+OwkB+Y/6h8kDrv8GrV91/p4Dmo8uCL3yHIzh
qxpyXKUgwcatGu9xYEOxULnTGCUzmRcqw/zorAaDmdpogD/f7AOQ2XSbZNIpuyEQ+z777L5g5mBN
pH9NgqZi+neoG6ar+qYw9KAIkkw9+Xu8ujQZJYI9ki5tZsRBsMGuPyX+TBwvjO2neh+GjSOQ5yio
EJ62QgrhbkaZQMIeoApclhUaXBAjBKMvthJYjIrweZU8U1JyQuEllw6Lxx7TFCpwGriHGNJnS9XI
/XKGRt/LBflRdbw2rQl/vqRh5a+PRwsFa1ZLS3o6lvA9KanQ2RRRk2s/XNFvkJMYL+cJaeqUyz+A
nylPmRVpU4u0tF8TOKQm4wkvseCA+3iN/yjMCJE5+v4VDR1HxEVqcWon2H87BSUuBLHx/AqRn6/Y
i+92MzkcE3XpNUBZelYtPLA90aDQjH25MFWjbBlEO9QhnEydpTaijOwtx9iuQ+Z9kF4guI4MDM5O
r+eTArOxK1lObaamfAuN/pu6DgXVjtCq3iTzUPjtG19kQycQAs4s46PcpXR/zfLYPYfFhAvske3/
CFTigi5/KDH8RY308SgtrX0a95RdiiesKBis39ZzNgmaSLhNbyyE1ouDi48mdHFSuW02MLOTft7f
lV98mD2xeX0bVvhabnVtyoSVBgDPkW6Ubhq/6TMacggaY1wvb3v1PQ5SLvJdQggM5pmAEEr4lsnr
qv7cIG26zyUGbEJNyOX+h7Oswa4K0845y0wGPn2PpSGNFmb5MBkmAJmEEPQfxWoPUSqx6Z+l1skD
/YEb1pRviSoHNaTsNg0K/UPHZ1FOjjPsN1mMjPFlkyZheWMaNDkWYd1SRtg+8y2PGHNge9IGBpj2
oIRhOZkRXwhyj5G0QugUMjd+vfizfEqvmzTIWmXcozvNZXudH/HO6Z8lDc7Az4hrYA2iFH10ykYJ
ZwaQNo9WmCiZ3raooxgNw2LJtq1My8YkPM2FNxytPlbOJwwoAhFUsIhUOPgQXRl+/Q6MbM7nK9D8
nDgxwxG9KNb3SpRoAlVfVz+ZGUJVFyEn7TyhGvABAZxeX7W/k8fnMAgbSALTME71sSPIBOg73yfB
LmWjBg4otmVMUywCDkhhLPfEJ0BzWbO1R6ldHbfoEvHWeau40289GEU7N6ccBETn8dzsVrfzmHfk
2RCYX78C7h23dlgMVnTijFdkQPBOz++fjKL3JhO3APcjrGUuePUwyNLiFEfTDE8eV6vE7du1FBCE
lvSNL4ebXW6lwpuALTiSjA8KrT0kewUNDI3cP/UElgqbUCeGJRBOU/hguf9ca5nyvI4eHeVp45ES
2TtYbyn4C/p/K95J44m/xNSDGli1cme2P5sb1BBrut77g/D9TaB9nmg4CujxU+RGmr8v+e+VOKev
CJEib+SdaWTC2oDFuVB6uzzWdoBSHCpus2gtkIVYruupkBTWkeZXbgnCM+liPbmxTMrtTmH6kzjl
ckJ42tl4QjuR9mKG4Di3D2LX8u3bVDcOpBXwEMGXfr/i0zoMcoStLg8Eh8CUmarGdymz6n8a5kkK
T8dvDTGd7OFHkcIFHYvlaHyuP5VFrb9ZLOWULZN795PCwv1Am1Vujsxsbk6ySnUH9bGr9I+lLlG2
g2SAVqvcoCFmyn4Ok8aQYKEobcaWI8I8DrEh+pksY/3xB6hAwX40MqDYI4nziFX4QRrwYsUqVbmR
U6xjWDFOEBqXh97+ZTXrxBZVxVlO0HcHswk6MAiDJyNDi/agVfDvv8rS+OP032O2oVptGzHpG52s
62ladKtVz94QnjVyN6qTSN17o16FKp++VNAS4Dmj9c3D2pJ2NOwgCNIn1/SDLjaVv7cZsVjlNNaC
jYXQ03+1G9sgujcN6AK2fwUAPFuQXeJ0cUih8l4j5pvkMLEG791aQMIPIq/3rfqnF299k4PO4zP7
5EjkJmkqVVOQl3mYiPLpTDg0JxboY3/oeO7Q549bzzUG0FlVe+oq79Ww/NyyP36DMGqmHW6cDQHI
C3aVkNYlhkXajah+9HatiTrdZNcl7D0HlRJ+ZbhfKG6QiFvqfgLTiXbmN4Rg3EB+f5Bipr1QvElD
ZC/i3yqT1SHkEyT7S4dkMasixncmjegVfz9nBgPiBPhMHZgJxFyq9LgCwaAsAtSAeZWLvKhrMjjN
klrwNF68Zz7T5BOu5gTp8XjSQqKYT0BI/iMhFlCMSIvPNCyCmGprPR6zp8EY9ELnN5EgFgjpPDlJ
KWDyh5DYQxv5Uud/Pz6e6qDeucUvK7AhV4r+/9JKkkq2XEAdCS4R33PW8xB15wO4XP3H76tNwwdi
hfFISIzry5zv0iaykcRwwMMKDV0NmGKFsMrJ6gp1xWMg6g1mz/6wrJuqhXy7Xw12ePoiB+BZfAVK
NK82+gt4PNbPU8jFNrrwmgoLKFxZf/5UIlMfeG2gxduM1B9F/pV8+kwB4zgcGCfvjglu5yFoiwpA
kQXnz75zpSjHvhZv+kQZbp1llGHgIwHssXOBJWI278DWKTmv/M7b5DmsOXYAYzqngOxMExvMbpcc
WoM0DiQwjca1hyVCI+hnZxEA3HDw2HWfKLs8CAkthIPcpm7Gn6SA5Vhvuukmpma0xVhjC5SopNi4
ygXmKIrKuCSP1BQ3TAuGS9vOXCsae+45tw08qq/LROqkmWsxssvKOOA/CbYWx69DsU6mQMUb5u7G
Rcy+CAOcgB6xO8FkW5y7os0SzHCoZWMzuOx3gDMihq9bW8N7LbwuhQBqLpvfnHc91i28qQL/SR6l
U2PocsrarRu+3iIQbu+uU9NwI7+ttdYkkgRmA17o+rmpA/UeqD0aT3H/iTHYqgA+l/N/iXC+2N/l
E8UEReCB0d2LuIBYMJrsetISM3ZK9tvcSPDosoHDzlpP/My0kVpDOLhWBrxnJQz4jBmPME6CkidZ
Dh7RVgO2huV18dy3q+7jrGYek3VzDfXeBcpwo8LqzpPEvQ4cOYTOXe3aOzEGyAIReC2jSah52wL6
HfHjpVXhNm+Mz8Ha+WAfjEKD44hsQvGiUUcOWd3fVOq/J98dRJNb1AEXF2SGucYfbUbEtkWEL/xO
NLAEZLwyMSLpRJLmJ3kBTUNnKnWzdtuLeFNZdyONGUrvB0vKKZENWImV4LvPTMmLr2WRFNQV2qpd
t+NdaSoI8nPxfnYtw1FXxjmYUgI+iGNxz6Yyc0JqvYT8zXaWXzU41+TXwyd1sP4PXl9HatMxG+Em
DDE1FkD9IT2pcFEPuW/qUZxqRku6AkAaK51XSfleflMW06oHXLzts2Ed+O/3uZCyxD2B+R+F3SSZ
oT+H40tnMCmzLd0hkYsPrYZWC5eDduJwf5cELU31ndXbTmcfKW37W+Kpvh1TLK84/4C3gqtiF69P
z05WJOmVWd3Xn25f4zwud/HgLoWTbUAv6QzxQvroSD7Xjrk4sPDRQHnTYpPOSHaatlGtLuja4PR8
/LqZ0qL6k+JgF3YXgyXyUR8Ht0VfOPNt3yAo1IqyaIID/nRcmuriwfVSFYfm+/n5aXXABowk6gbR
0JdcBMFtx8+ZhU1XXn1LvcCr3mz3ejM56C/GJwGucUKlGrErcxiA2rb6B+uTPANa6xE5P8Nv+Dni
B2ZQ4j9gU7yi/eW6N8bgjr7Dx9plvCnfRgy3bjiglFqkAcJ0cGmwxtiRCUM8MxecoJWjMup5xo+e
Ge5EP/c7loVKYMp38lVPOC6smwMqz3FEFJsBMS0885+Gx+Db2mbv/Z7au8BSTfiPIdwDOwJDW3UX
hpmamjyn0DKDfHeQbAzSBXpVSjtffdE+45WGwdwTh1tdB5xaUhFx6fdBhK+WdA0Imylo/fnlC1Du
jdIoQHUaxCwffbk9SaJcZT2+wbDCbWoerWsOa/Q2a4sS9ax2mDyjzJahQEtzhKL4z0I1TXHPUu4X
YqnJsEQFBAEo8MoBnB5B/yvUHyRJYm3lmGx6KWytN3HVOlW+sXjo6Ph233MO+Sznu1MKjQUK4WPm
XHIR+hgWZ5BkqzRIN6QO6CVurmyzr30KIEBuowUdLiaOVPCfSSJq4kSHdlhDWMseG+78ccbETMOV
dhqpOE/PEcQMN0Q2/Fc+6mwKJWWOCIcVxwN6ZBtY80l03Ws0Kkg7VhgleW0/CrRdl10RylpqBnzj
OCIj3p9wTD44RT/I1T0FvnxRE6NHtIdhIKsSVGcxpGmY2Dt+KgztyWSIsb5mHjvN3+l57p8gkm19
jCa/6C1zZoAUhAEY/wTFbgn7s93OnNozUwGyWs+3f+/HmWC6LL0Gxux9CII7cV/FxRaxlvr65mmF
X/wTrOiJKndDe35MHGtDbJRD0Zotu0nMTllI++7pXCr8kIzQ73KGv2EW201pzYkCWNIB8eXhHJj6
ygpOOAWZV44EgLtZKoXJg3lq+nTZm9iw43ZuwZqYjkOmM1yur4WZlspXhtK53wdDDCsJFCTyTEA4
st8QkOaRzguabl5HgVSvZWyYV/iqPnCnMrsdrDqQ7vrSgv1WIN8KqdgplpnsC5lg/XbCzdnaATI4
tCjZ22tMyPlcBc3JRLoSZ3mqCAUtqho0Dzz2r8aR7HT7fNEbVeQv6F5u5h8U20RFErjEiboMhiAg
BhDf1gSQIpssoDqRKy0LZX2vFVZre+LL3gvWnJg3uo8B8KIWb34Fj/c+X13SRC9a3pSoNao62LID
7GcC9mqNNmCcujHTeqqMGJCinS4maTBqIspNycjSQjRfX+rThemeAWrcH7cqXpJjiigzLvWsYUEL
PiW5HloU3hpOygDYXxe9Ey2zkArkJd/vyuDyTbo5Tur0Ip7xNCO/1aCi7TJIcweZ/mJFqjoqH6ov
eosVcuYvioD+y2WWPPB6N7qPWzH+xPEi4my3HcthdlHE7sSvqWWpbeSBH69biq/81bI3QnjkoUvY
P485SESIXg6td7UoAtaFUOTEcOh+DI55oTlWNdt2MtaZUvSrCGcvjiHzDJ5/Rn9CndyXm94KnM8o
PRaCWG6TzNd46AJlPs+kFaaqCMCBD3B8nceI4isib4RT+CFPnzvXAYQlsnPOEc1XDyX7j/lL07H8
+xGXoULPwaqcvjSqXjd759Qci/pelt8fCBojmLZbp8ZFfsnSK1T75ZANQvk9uG81yK4iRJlIFegZ
VuKf2M9oFh31ErGmsErN5Mub8BGRw5ysX+DD1AoSt+XIcslXcFfZsT/P5/rvHuBZZ9rW7EsjcZrO
4lZxOTGQIcc5kKuIkrf4gZKbrE4BHPZURoGkUOFvDNDk57t7siL2KaGu4N8l887fpMSyukUFvl3c
hfwu6n2a7IdRdUbz6+6Wm77KaeErdQE295rsLrkLLap9rCdFzAtNBimDMgPyuo3Ef6IR8HXdMGPI
gPT45R3zOeHUoKQXtvNE0+Rs9W+9Vu2Bcx7PQMhkezS9M096pwAKE8Yz7Pdkq0HObqpU6xiuOl2x
E5RvlMr/zYqjOSXX4TejGHu+sixuiUXITLvPI+wBt57is4GWKBD+V4haY7+xyiwRpGn9WmoU161j
VZb1rfG/Go3IyoYyUJjtQRpEVJp4IspgguH2l9IqSg8i7trfGqoIuShUm2EjRL91u/q1GGTwCtGI
1Y3A3ImhlVcjrUs6y/qA2peMjbWMxpmLOaN6UrZbyb05i6juKbyoLNYBVgxaXyWIGVQKCQ9ipRK+
nCVupYLSWlZwclXA34i8uDvXC7NvyCj1eySNfaSJMpXNfhH3AqHsMh4qnnJN8kkd0V8LTzO21h2T
SHJ6+aA49B7/oRKYstcOUVPUoLxAGwnaSzT4km8lEtDOKosv7hsSTmv3CDMrPHHb6IDFTmSu7t6e
6VYJlp/A/DUq7OWu97m+S0kWCrS4gLIEutoKnuBmsL+f5Rw0aHoHPjS9km2kLZgZ7fokqas+znFO
tNrEieRa6efTMRLyIw500GPKs+Z8iIDykMAFspW/C2MFhbHFt5wd9/0Ms1tI+AbKIuBr+Hw8/Ncw
jTKB8+iXgs8wmnv7H9FvGdd8VJhbepEPR5ZEMEfhl0TpujLhi0eGLsrnhm/d8PBb5Gop2IejgnGn
FkMNanJRfbaKgAPfijE1P7gJl9s3aQ0+TBVJq+2ZOJlNVCK89/mZW1cPlfXN5BwovJ/dXjG08vfk
8W2pVG5TSuhLvaWWwElLLVPur/+KSbmYjPvoMqojmHLrHRoTBTxzeyI7CnHkuXTF/597cHAqFXaN
mP3iFGWgaAyY4ANaYIFhr9FGP9ZNO3i8dwPZYG6BigbdKDessBGnhdFbB6N2Ow0ft8xAiz3E9/cs
NRQtpSn+Lz2kl2aZ6DjgfcABjvLg05vNc2slEMB5+Yth715tyKDGEKJS5hQrPKyKIRJESsj0V7Q1
T/mX4XTZOWCju9fqQ9WznEeZWjYOLG7C4qa31Ug2ZSnBHE5NHPvfzdmuxtmVrito1wRiMSzkdVYR
efSIDunP74UBi5fXXsD2EneyaCCBg96tUm4gBHu9sYy0fsDmZeiHqU7TniAaJ4YqYw6Ed3sXI3lO
hQzMUlW5+0MN/Pl7EwP2kdXA8YaGlzTOXm4FVTlOn6hAVd43cB8jankWeRnIhU95Ig8QTDipNNMp
+0NM2seQl5y3sKvPaO0vLMZ2aJhnlTJ8LOHJSOUQe4LUi1JbB/Y/9QU9AeqcqcvZQH1pJExtlgjq
08bqx0v4lA1DSUWWcCERfkirgLtG+/K7gz6MV/ZsKMwheTEVTCN3Y0cRPAaY7yeNFpsYiN21QX6B
B+ZYLwORAvzepVvwWUFx52kHYOg7I6XGJJ5SkXSDCw80C3XrzCruPPgdNfAfTe9b0vbPVrwCaiM1
IGpRZWZZ9AERv0bggx9t7FL2mUpXqC8ZlxhO1aincjKqGNHiRdrdYj/92tkj0dPC2VaB2wbvReDP
xKBUe2l3rwadQyMRXqYld070HN266OYJ1Foi4etyfFt81MPikb46/xUOMHwDcmO41tBXUH86CcvV
aGI1k0TQQp3htXipKCTskGlrlcAiZ8YBZ6w8clAJHqEkOwzJlEMSja3daKs9l9Rvb9LpNgTXnmIf
K/gKky5Ftp5JI+4eoEOEjked9Y7AoxFGsmzBMZWpXwbmGfbtRQKXCg51x9Knb1LdBYPQtqEFF36P
fxuDPNMp5YuURX2CYzBTikYqmBq8xusrIj69vVcUpi/1NHa4ej40lt6fLzJM2g5/lNrhGca+09fP
ARJ/XWIK76tSPpJ2IT/2gRu3lsW3rpdos91ACW+vmw0a1XOKinvsSSzgpKxn6h1ov1OPujAyGiPA
H74cG3ZRtCEcH26J/JfWD5cLCZfkPd32CjLgnFAP1r4JN5XqOz3nwLIz9PDSPnX3kFZ47yMTxrFX
GYDjaa8SyTmCcqP/MSAgDTK2aGbycekBjEL9zYOjBYPanwY1tIICsFlXo7UxdLJBDMjkLA9JgFLH
o7ml+agoMs5mYAiKDKsPDN95YJS9b8LoP9lG8YZSJrJF04Yp7w4IZJDJpFfB3g7CikRAZTgjGczu
X57AyXbN2S8MVg8XvMeikw0BmyQe6MLqqpD0sYik8BDq/RWe/h6mwPwhg9y8eg8xfibB0WDCNiIi
/t3fek1PG5WIhkTfshxFATeJp4ZAsbbfgU3l19/+fdztQ8QYkEV6cUGj8sLsKv2RvpXS+whljBnE
/47l0e8E3EuxYQfdmcC91wtM42WmlSAyQz6AQE0o8W86IOUPWTaOkBjEU0+YmLXPLJidFNxSr7mw
WGFP6jL+1TN+otbU+56x3d39st8l3CVsPo6bOAcninoOV8Aq4fjNYrytSY8JrJCuMcA6SXTLp3KD
o5zX/2d0pEave9beCLMCzqw7y9jXLhcWCuwIaOsR4P5iBs8c2YpBSnatbE7c3fKDHyvvxkqdDX3y
hjq1wYa0pMexawSVFB8dpBu5aIg5RwPM+vRuaYr0swdH7YVU4ads8t3LrjZ51g1GlbryFW/YDIBq
4OlvdWWv8o1Fv1R8uHUWwV84UKNVZbZoNkXJ+bqPPn7VZVjGWLIRt6CJDyrH9FCCYlkZEVHr9PsN
djbNdKq5lk1EaQaYzEhsHQdrG0QlCteUfkHycjAOMU4YIgmVsUb1MM2q9SgDgQ9iKP1+sPq8x04l
VctIo9wkQ7v+nlRCKYsROTE5676FkN+5HLksF25DrEk6sk8ox1UJ52z8RWO+96oHjaWQB09IBmEl
v1pAgcuSqqGdstl5x6h29Svd5x+4kfsjSl1ULuqNr3f1/Vj6zKDPbPYsEEtWmBAxmX1F9X4o7Pd0
/rXozhFGaqza5Irn97lrIDNP3UThxCW0PgIoC06ZqNt92TxTEXWpl+ghDyBBRxoe5Fr7DwZHHiXU
agXOsz6OFRD9E4D45z+DRkstQljNHz5XOnOLhom4S/8zlWeQmige8ul1RNOn05qDgfo3KDagUb2A
9MAlU4j/NUM5F0/ucj48Ld7W6+ozHBmHOHvAF3LsIENGT9uz4fs/joEz+BeQpuj1d6VhFdD86496
sILxQHlgEHtLiyI/ejYQ+kThJ3UZzrB3p/N4HDBI3pwOkfpBqNy8t++ifUuoDWlPPLI8JiFZGVy2
qzPrxXlmyoBvMxPPrwf9zT/sSexsGrQFAblbrMSr5sWrAfziVxBGCEPqomSAtmft7UmzOtIV5eO5
pzYs264r7LVhOL+ZgpLChKJuKgkBjBopmRAUiMs4/+EMIjf3nEafYuAU/2T1kKrkY7Ue9ehIQmCX
Ti84gDgDgbP2upyiOI8Zcjtryuk4WUNcFdweqerg9LTn5EPt3m3vPEtvSbPtOumrBb25uX/ME3RN
Bfl+lnXclwa6WT1SPGTyxwM7oc3eZyzRMvDCEUXSlDwfoeLGUkIDTfS1xuXe4UXm9OlFIFn2snqr
NJMr6TmKxeeyroyJqo+VBG0vmIohrgccsxuExZLDMWsKBD7TAKaBknyo4Lvje2twTffROEiwJRuK
yJWeBIMHQU3VtSxrPY+CJ3ldKF3t0qlDKW79WV8ACWrQH/o39ZCfZjcCyQDxIBiKhOTxwbI0vXMC
bKePq70KAfLTNLeESzOscjr9Sg8BRnItMN3U3bakUdbwvjDJDM8Wbf4dvPOAjKF4MDl52i3b6noz
YZECM0qgwfdNBkrVkoTAIci/RpJ/qzEk2Iiwg++a3ZMEUsVP8LyANmBRZ11q7SD/aHhyrYnKLrMD
KQjigdb4pY4YhiDoHWS5BTjF3yrXbPZ1Y5zGlhFyFaya4zYW0C7rz/8sgamjOw4rNuRLpOlV7TND
LiMKx9OAmuvjA3gST3WGnndVfKccDqh5+4ag/tlh5fiKF8q+E+I/JMCaXItBoSESBYvMGo0zzvAG
GkTQy9laSeDEELz9nfnPSakjfzQAWqrHfHbRinDLur7diJI3fjMB47zJIBI8TIQDaouni+CYIqzm
qIkHcMUcqN+iFmGTN2tDFlGsVWOFzq2diW246XmcxASoizs4D7qYvzxdLOqmC3HyV9X1ROXUXQRA
5vXeQpsg50DqZKQ6Io67MkfZd6IgexvQZZSFQxllj35xfl/PRL8WkCUPakWKzIQO6MJpYdMcn4Sz
Ha8h5J5rnNEd8CvMTe5eqba/YShHRqb/YtqU1HD1iWcn6JwOrkAeaXrIppV4D/l8sZTpm/djSb44
0dXDKH//9N/XmkRLj+cJNcMS9zvNhWRQaNnvR7y74/ry/63quLpyxVHqC8QDSgu9f48OCo6RKRr+
P21zzpq2ZZjCYCmz04T4QLP945oy4iS99Az7pRDgstit0+XoOzgB9xJp4HQDDQb7wj45fUQ4yU/7
oYRUWFv/sXyjisFdKy+gaAfTlSNo4S++Xvrg0Fi9/5O2D9J+xH9NDqQle3kKmu6elBzVHhTP09v8
crAHm7wwPmRY3eMdxsyeQ8/U1jfmS0mbH1w/BQIh2LPShAtb0iDtnI7g9cQqDOExpj5fwKSJBoAx
4xeca3+zGqUM6ew0eVG7qdiBjw9Darrp50w5J0xjp5c9r/kF3C1jL8wm9IMj4t7jsBAHfWEcT0Cs
Cr3Op5LgGOrhUT43+cZYYye5Bxd/4ZGNYtAIKdLW0mQzX9YB1rINvkSK59ySRCNimoXGVdgrvWXW
cDOhqxNz2oZcnN691+yfusCdmsHFaIsIKxd+uvbXkdS06HKFJs2qFikARDZb4qY8LkApdGTzLpfb
F856oy5AxHbAobTFjbMitEgeWBsruRaWSnWabB3qwD4nwF5tCiPK59yVi0XJDOG5n/sUFDs+0cUw
AX6Jq3+oCxTUP1EFXMJl0HxpBwV06AkJXaWouaIYhtBs7bQntycCUuAnqyHW59Ux/G1MP443gYEd
pNmX+I/cLFzIicRpmfb4YOZI3lWk0eo179YjIb8+990CW6cB19XK9Sp3TL/MQbbQQ9BqbgoTl5Al
XC8ZpocmlDdHaOsiN+d6Qwy94FBSDIZOPPxmE4yUvHYlnkGOP7+QTnPUslo9C5C4uS0CrD+To4J1
a31yuVOZ6k7ff6uu/mtE0N4ZPDT0Bje1+EH7RalhzWNQOdDxyiqcceftRvaY6ANstAw5+I2YgvSj
8AOyCQ5OuMvmXgg9yvXtzsyRSxlwkH6tz6pOJiuxtgxi6Ipnrx0rOdjeXHQDEsze8itxAGyZbKAY
ZlOjRegQ0sV5stayIXiUFx+xEHFQXlHx5O3VDsZAJJwKdArrRlCX9FHGxVWGEuPRnkEvo3bSTimq
AtqxlvrsUFb8i1ypXz02TRvEqJFTVqbjvrir8RX3m5goGLWAyta9zB7wkngYaNyQKaSOZZ0iXA2W
mJtH9UoScDTGZr2jNOkwBzTnYygzCZZAIXQBSW58BvEb93wAacvxrr7IE1SgK1iApEG2ZXfH3i1N
YBCLFmnN+iJW0fIzPQO9iAXKCts4bW8a+qbrowY6GB1QOnwjjVmgRRX6Jo1wEqjBgYvSXl3L7WU1
APYPhD6FUa/Wa3SerKrS+BFB8Djp/lWiLIAUGx89nWQqaS6rncAZdP4lDRiyQW1/sYxPpOhjX+yN
DF1rJhprpMioBoMwrp3xAN0oIBaSb3OeOUAl8/GvQ/NA6+G8/8IVG1q/pXXTTwm4g0vr4XAk7SPb
TY6/SWB9R6EAB2Uo9zJhBEBPFELK/FpVfiBL03J5Qsem7oz3abILJTlJSkjDmoKpJlrFRopSsGLZ
c6OZ+l0yceDdBZVEuSu6zKg0rQrgoT+dBquvU7/FxC/EKSlxYm2tCJgNqVjZwQajIYckSa4DfzYI
1HzUjBD5LGC7EqYHqAZjy/kht+2A3t8RzDB1YSIraMD8AJTb33XWH2lH/TrrSQK7yA1qD+beL4Fb
ZSONACG/9JFqF2S1+WkyI8RWc9IeeRHkYRuA7RB5HAejPZIv2e4wFKs2nZ8T7ZOXnGsD9Krxr+HP
06u37HRFc3Tl4Lx9canBIeh/iC0tvn38O/nJxpfkIfathh2uuUMqdMDvzGOmReQfK49lEoUD7C2p
i1cXRIFTCrOuCc5eHOiTYtGqk/W0ToClbbPW5dHbkjlD2QJXkC40xQo1a3CTNwFK/mYG4VB1eSqx
ZkLXJU1ZrREr9cNELhxbXm8kj2lpug5n7IiEwD03H+qMtt+YeR93LESDxaPAVGpO7ymbidsrA0yA
msm7NPPcE3b5g1Oc9M6HWDcJUJAQv+Y3vORHe9/i9cRQgq8/I08dVxwETo0BWIkXOxZJQDCA436k
i//JdLTt675JZCML8iLpVpf1U3Kt8wsuWdccqz1Y6YK/IT+oIEVa/xDleGhs5If5kdTZcyfsNl7Q
/IhLTOK3wS67GRx/JyAOMq+QvGHlfDZ61R/4kRrO+vZBFByAdMxgBODvN67zvo5a+gGn9jVKPRvc
pHvhPkzvn34oy4p3claoJfBEQBItCTDWoXcaMdRybk6ZM7vEDfaopp/irw/Va3sEiYj5bPQ5Vz6B
xlM+tI8J+VgEEHhwF1xhjV0LbxyS/sG4011widkCVISXTdzS3R9sCw8ec5eleJq5SIY45vuoBw9c
e7AGyR/Z7oUS3wrk3artC5SiSXWNEVCqffxSH+TBFiekcfbdrMEwtLk5QX2O2qZv2VS85uqRpaHK
BmJJ/eV3yhAps7ZL7LF2tKnZ4dw/UgcyGoN3sLxEwwi27LTLeHrwy7rZ+YtCqUAZbSpL7tOusx3f
W9zSaxADwBozRNGFhZt0zCSRn0JTCL+WLSdmXuAmjWmLLoaSAUx2D0pEXztxbFb+058AOIeHI57N
p2LmQePO0N080QwG3F/zx1NXNsl+tHX0nFnwyYibI4voQFu8CWhXMpiJtm90uSnnHuqXF+yqFjXf
jR3ch0ipqYv6qaF4h4KKo0gAMBbYYddJIsK0elNnx28mJoKdYLAR2iqTbjKINrK1165nbQlY7YI7
Oigm15IlgMFMsin6DVuaw4VG9M0QZ2o2hBkUCIDpcaeCM8FFb3S6WyYGCfNVbbDoVChbWIhLGKl5
npK7QWtIYTC+MSW/p1RptbRYlgf+dwxORF/htAVMXZYaZ7dMJ7+oTUhL79sG6NRYS6ebSpccYXmP
YuZp4s1KNVp6whUSYUDPWGi8+m5rFMvJHJV/r71A5bntJEWUCFUnycGnLJivOXHmhqznuY9tCK/U
CWYmvWyq9BkN9xT8IzIINhXqnyz7DJNyLVfgy+TWAqmBdqlnlrwhF2yXptqEGn6Ppz3jnJR+rTlE
zMIQFSfm48/cq6VTjoHVfWtf08wy0URmAz9cEMFSy6Ng+98g8KCGtKWzhsiLpVflD5+7MYCutVFy
MWTCzzJS7SBfNLVZLgS6X6Az0IZQeDRmBpU4vPzoZ/i4B5hSAp76rR33FAEekHHZjuXlfHSbhiDm
biwV02d/yo6mH8WwdB+SomCmd3ZbXtkC90fvctOAfyJ7fwsN0tr5ND7FRsN0ovi4kI7fyBm9dLRt
iqqnYNUenf9Am1pDZpu/MZC4hlrTKw/xKIBWAIpN6cMr+5EekcaGAVPeueiN14dfIz6GB3auO+c0
t9ruwD3tsJFKb3Rz2HtW5mZ317vm1q9O1Ztt3oIWdtaYkS9ll7PuPaV1Oc8wQS2Cgh4fJVyfTxJa
+J4gvFa+Pi3HaJN704mR7QGQAViVUKnkU8bzHc/+5jkkhy4L8kphyRcnCO/l60Lk6Zp2XQfxZWvT
3330UKiKUVMVWeq7BF/ImX62JYWGnqGouwb+L6QmfK8Rq+lSTtEca9gy0Dqp5/6qjox/JkVKwV6f
s1tGP4vgQg1h1WPESYFVcBpvUHmKP05qkYbeXjFJF7DGef1sv85txl3Fi0XXZvV/ZN358054czs1
WjSzEqL5XM9cZ6kkNP8OVmw+RIhxbRUPy5ZsWo01Shbtl7oNQrltTksYaLuV023cQbOM8NBkcRlK
CmIUReU/JO2nzjEKSY4b9BYaQYkFuVigja5AYGHq5yQ8Gnh3AKybSe/KTfsm6awYLnfqna5EH3B9
0taDfcqQeBMxKUeO4imaW8Yv1UQmVSIvUcEWTYP4VgxduBMkvbXdoaEyGVotF10El5xKapDU7Iha
FOy75kxOy3nDbpPKbQvWgzXjbgJRDMhmNXkhxECLN981nFZ+Ct4ROhlrg87lO62QrUBIaqhOtloM
16D0OOTXnMbfsmxGXPrM5KJG7bFL71DEYjBm1duAyQ3EX2dgYQ+LDKZA8yXj/KFIaGqwQMiemRKa
Ff8oI/sVyK74XnwLMAByVc44g1XFNQMr0qH/u3UDWeGXlFH6XWja+5LYewS+LFX8p2jSeMuGcogX
uHXASJuZaKf/+JAna3HFAYHErj6qpgyJRXYudILVw2zDX1TgZz8trEI1w23IHumP5a21k3llyGBL
iMN/gw8HAsHeuqTXUHAkFUpPtZGsRwv5WvAmq0W8ZTVUsOnh341h/8yBntRiRoOtZybyWbFnh+Tu
a8LwmNmUqoqxla42v9vFR8eYaIiV6WG9xSIdKOtS6kvOV56b6xu0bYvFpK1pMQUX6fapJASE7Onb
9hHr35JRPn20luwQtM4RBm5LaWFeVZIXQk3L2Z0a2NKuoJtS7tvieSS3dH1IUGN6HsUvfIhLaJnx
kVrsfDBLyuqQq6DR6OXq1Tg8uDA908H0WQaOOM+22Hn2ekw30k809o1d4PjYa/NO9TSkJ+xoxOeA
D94rwJkxndxidTxqZAEWlen7C16LFso0p0BrLIrSsvhXCTJoP4Z/wi3XGjXt/zqqgdeewJWuhTXz
/v8oCNQr1IYASpwnb9Y9oSwtUYz36LmHrjPj90xLZstz6br/dQML+q3YBS37hupDlNqfojk1aXPY
ZOxPDEAkdwSyaBsc0eGqvzw49VE2vbakDkGf4miX9aCeioH7hO6dWTz2eGHfEW26r0vvu5nzCT/r
je1SdreJ54MHFpmL7gqImdLUbH4qM1lJxL9JFmOXfsX+6atHnxeOuFo9W3YhZAdxKAxiUufWI2uB
ai5s3RWGn3DOzwDuUzTIr8w5GWhiK3wNSjW0gQUow+kRce4atzx7CqwPQPkBuNGlIJ38zCN22qd3
VNXSGh/9kcDsFdlikMUqlXTNcYRxefe/rr5FR1eG9HY8gAxZKWHj9nDCQQaGziNB7IM7mtze3WXV
nUORPRBQcGTA018wYKoF8xToZWt2bYRszvnMTAsL56l/hzDOYnAdqug7sJTh+RZuvqyTlcfZakka
0Bsy8BXVf/9sYkcCKWcf6ctugTQ53fx2J4UR0MJvo1AP7SYjq9kJ8SSne27NpbCniGTho5UbL0de
oa568SelVIqDZWNS27ZCMSwi+OouNWmy/htKykyYKHR/GqIhEqQO3eKQFiwuWdnrGqeScA48PmC+
VTgr1SzRJhqGQckCcHYV8tSunAPcYm5Q1YNOAIh2Yd95Eybz0EAs0sKjk6qq7HGNFwTelOTcHptJ
TDkOqkv+1Xu6XX9WAHQ1VHGYORf5a5ndx3Fs55GTDLHusTXLWxpJ2SXTrIBObvBEuN1bdQx9GVTx
riC7JO0eKvq6Qkiwqdw4SChK0RdF45evgFRvws6MSaGwSlVoxLaOAVHFoFd0SMA8XZqt9nEeUwJb
Oe5Xk2Jg4y05eFm4+smmp5V3FEb432yLOjCTKrADhn/r//QNAtjMuf5B3oKjfIAqL5nl97oct2CB
bvWWPXvC4Wgr+/HwCj9n954UaLgwzkWZDpKxNkY/iEe1o2KejlDTS8NX7e1mbxy8/Ad/4gTGWma0
6XjPeYEDqGxgmMi/dczM+YnKznpCwOqUakU0LqqiljzpG2KQmnyIEV/eAvqbTSEPPg8/UirCeoqn
PjsYYnznQDzMLf57qSxB6cNICBhpzBNJREGwhR3kCttSavC8K8n4ZRY/cjWJy0DKKjV6EM4Dw2w4
eKzckpzP4kojnKey1lsKamgnP4KtGYZHl+0d9np7ZCmuq772xhRc6Hjsz21nJl5yaBq7i58THoUe
PVdtpW2rMeM6x0DEO3ykjKJSdR/tpovb5qU1KywByK2Y7ZiNCzsMGrMyRgdwRaQfhWxcaA338YKj
SkOqqLiAAbbYL+e16M9duYPxHDsY26/xct1fEePmi6HXKW54zghFykGRmWoBNwe8WULDG9VBL/pz
s9Zysw86d1ZyLsyHON6slmd3LjN9i+9UWjUrLEf8JzfDico14EWcxHMJt9y4LydBtzkDJcO08Jod
R05VKYZ6uSnmeFvqaIa0o4yf5Jrn14mD/hvd0QJUkQOgcc55jxh92FOK46rdvVQuIrJqgrV4Kfgb
GOpaDb9z2at5Vz/qqcJ5PKGqcgPT64nIm6rvjASn+pcUcJT4qBVcXdx2v9BWh49oDOibxOZ42YRu
LsqpaRjEXK+eT97zMG9L3KSUzS9O3A2Lvikw2QAJ9R9PK4qhJvfjjU3NgoiVx9BkFoB7fjiGJ66O
DQtp2bCz0ciuDLnQaiAo/clmIv4LWyzpkprXzBt/m26qyrVAfDqOPPHf8CISpQ50GSATPwlT5Ohu
5VuAezh9RJRgSJufNvbZBdKH5yX8trgVWABCm+1VsQeru9bgZRrRuqn5eIdLc2wSfJXI3dfZQZqd
oIixonkvRrmB2u/srIk++Mp9ttwPXLkfNF15glWZ2GfPPSqfktYzVNJTI9zNQdmf2W8CMHvO+iNK
Q5xyekPMvvuRiEoEOvkFRAsJ7jTPQQIRN6ZR0exmoWlj+I6f5iFPb6bspFZ6zLsldXvHVh9xD9Nr
CMjbhvrjfMueBCBHzpZceY784Kxy3v+1xxnFVHJRHSmGZYWv9gbOR7rOk7bSt2L6EHF8r7EdKtO+
0Kh+6V+ag409eGP+KgflDqOcmf2WkDNlu6eGKkwIiLtYHAQqxTByh96ln91Q4F06FHWjBIJfIrQP
n5OadcFgwETRBMUc+wjEmPi5ff/nji4GKRPRw66Kjgyi4SLV1LmnoIWgJEC0PlbG2nCcPu414M2J
0UNvnkfZZ4sVT6BnNAEpHtU6gPGO/XwdIDUXQYyxrT1WV2KwRhjCx/YSh0XN/F/tnHxAFW2F5g3h
SX+11Msp8WoT3So4GJP6nfqw1SkBeVhHMXDB2Yu/ghm2QmW8OP01jSDWJnVfa8CiyuWNDDxbYE0Q
umE1hLXGEcCdcP0rRn2eDzzMYtlJsKAUJBj25w2yCd5iGjjnGrntPbGDQPdBcrcEIPufEOUf8cvM
/VGEEBJKPjY0eNzBpynOIf/ikYfboYu9lV5SKxOJM1ZWE4oJS4s9I3/Gb/v/D6tMqS9chM9OkMKN
HY8V0IAhNE60GQKMFedtl5Ks982U0BuJZh91CO2fL8am20X2TtXmHzO+0OVLBToPLUwBb8oLdnLr
9BzKI5SstaIYBFfMEdC49BxKJ7DQuWr/XjgphEf/Rci61msy2aGM56rEK5j5JiZwq4mNWsiVcVEb
W/VjvFhQbE3mpY/C+SEh4fMmN7nx2+tBOejjZPjOdic5YVIY5RWVyXFyk7hQLSUpWTogAjLI/NhB
GchTXFh6RFEqB9JFZASC8PppYktdjfXRuIZJ7/MMWn7BCf9+LUr7coahVWsthbnbPc1sBQSbGwBe
234WtCvgWsd+uFmNxXUq7RzlSb4WVmhzwjaWzglGBw0sHmY2+wuj/79w6eOtiZqvaZjuTPIBebdD
5uDNTUu/llazZ7QYqBUKZlriouTNOcgPhp5GFC4lrifTlhvXyj16RC9jwH8DCSrmQ/wyZrSyPVqV
EXb3n4hAo6O7R4NbHmPe4ucXeBTtKRE1XFyZTcrwu6oWPu7OsLDCNyHS8HDipwHNm1bIzKHspZUZ
L1Hs6L196knT2OL80djKKN00nE5cXlgFB6oHnSXca8zzeBxvI8kraX3bXHblV3FNh/7vlRQbtu0p
JRbiEWZ1rVteSG4JMu+MDk/dMh7mwPnR2GcEKkCkBmjOwQX6HctFhV4iXVEPxrr1CE3DDPN0D7fJ
MiHmTIUNfRYNTTPnkmCDYp8czQ4g8hwph9Exhnog3o0FTH0IV5Rb1A9xCsLsfI3/OxYgzmLrMvgz
H16brUW4PaFZSMhb6DzcZ2lb02BncbQJGVpDfzu604HlYb7rQz2Y3lay68226SUIjmwcM0oHPU3R
kcy2cMU1c+1vuuF5rv/tcTUrp/Bplz/I6asrLoj9HNK2/kmg6nFw9rTcI0F/P7/H/RklYBdlmn86
u2FsPHeUk5uWV+6I4Wp7VIRo/hipizCFS8GFL4pWOvjbZ/zZ4YlN4g1cH+lp6gW+lLi/xsaBY10C
/c/Add9GPrNvafi/BPqm8nXJQB2YgDqgvy73wv9hUTXzw9jxTTecyPzQMCMVtCdswI1d7gFab/FX
VUQ2gwJYE4IenGo8/foTWp2koCGQrvtPPEJFWXG3FgKX1PF1ty0SPG0Ka6daI+pPNvAtpbs4rlyj
mM8n0fxvYAy+dLe0RkD+URFiOrDQ67AMI8cJN82pRAykD5cREbDj5ETbXeu1eEsgK7ebO8UOXoTZ
Fx3gKsKiN6THLOvxARmQMXuCgEJ+GhZhoOAyvgCy1/DebngayYSsyjWfGQX6WFMMjJI/sTYAMXjQ
uAo3prbsIf3OTXFlJTMsQSI7g8P2iqKd+HRGLyqHXvstBCy96lNKeXD5Gf4v44Ps37ChNkk0kR6H
5gZuji4Q1nMZKSGBZZ7nNwy3N6i7epC61eDKiRNL87r2p08GjCP/59GkHVHs3MlvpWu3HSPjRAFO
0HwkMZWlW/ghlUD0ulcHRa886+sIqPve51bU2QaoVRnJLNOkRwdZ/MzwkXn0O3ptPsvXYco6R1Ja
yIYupJuNO9V9ZOOaNzY8BH5Yf289zsCyxqbVWyuUdex9dqXPIqjeJ4oTrdx+xhK1bS/YcbIUk7sa
pzwNKm/wtgPjQ3xa/2BMliXyqmOjStyHITD4wgkV0RRJG4wK6YRQiA523+4NFCxDBs8SkcHISb3y
kSO4aEdMM8OBFv9r+xeMa3VEOGZ6YWt5JVd0rnP/gjdXKl1xX84npYlCMjU3723LcuXPWoiiMAmR
y96pUrJV64xO/bkGwfsC374v/Q4zI0550VA0woGkdFSg9XHjafByzpaI2F9Iv66xnLeFAFxhxFxK
gI7G0rFD1A771/jdl0f4eux/lY7PAJ0grZftEB8Bxde+nULls8b5cX6UIZNOYJz8rROEybWSY1mz
PhTtnPxCiQsfhfnF4ygYevzcPcI7p6/L6ALal9frpe9t1zZRWVn7dtCels/xeQmvQldycIGHlV+M
N43fUL6OEgVnNyAVuMOKnSMIZJAenHWWdqnLixa1q6J4YLDkDhuFDhWFuanI8+JIt+JHz48w+e86
w4jpK1Fc57FKkbTQCByFraqZ7oy2hBw6m68QD9ZEVtAgBF8JCcg6+JTTsYjV975HsWUbWg6Y+Zb8
fB93JlXHO9w9eGEnwa4TZdA7iwK2pQH7IriCzM0ntv03df2lkB4p4JhZDDKW9kjOjqD8DdK2D6br
shdQFW3RtLzmufaDEKKdFXAOV5qEeaiSxbtQCNhwo0ObHW7Xysq/3dCS1Ovkz/3XpZS8J6SibA6Q
Ig6RVSj/XDyiRPkDUivJkFsPBkc7J+z1QSESqBCjw19O04i7cm2viR/umgvh3OHqKfKZATsssvo+
NqmebGmsD4BzVHkl6wYEQmcPMV22p0dAx9Z3K8Xqj1po5s0+NIZadhSDgHwIJPjzjW3YJeRGT1YX
Y1WkH/dqEtiDVQGPptB3W6jt7PUuWNcJmt7yDcV0yEXAcfGq7icn9Em4hCkuINh+/CvnfqQXMi5I
KWP+dASErQ1DrYJ2OadxVam+5y7Iq3bBLpAbRlOKlAliYuPSudadkS+gODfadtBjHDsyD2pTx358
E2ASU5PZMYNWd6jqffQO+LrFkLoM0Koj+DQAsGMYIN1Ntx1TNtzg0pNWOXvIuCFf16MYNaFais6E
pcXsgTm6gf13w2PVMNScvCeLOtOYxO3ndNjdOGQwLj5pPeDpu90o3Ea836uucwohnbs2OVH5Nt1O
VDe6OUvrztSN3l4WlvC+hNnxpKZ8PYoCVRdIF1cy0EFUyhjgYNDvmCR8F3UUr7wBGtZchejaLueE
TNvxHpOWVJ/SIApl3knhAA7tOEavKWixz1xCrNDlmtPqsp6vigwmv+TE8X5lcuaTUEY57d+kSchT
fY98XwQN5c6mnuG3yiuMp7msQrXIAsHzsNkhZwAbUk2iPKmeRSLvtgAbXllUAS20+3HPxOt7Lwn7
e9W4Jz2sV1xHK31qW2EUvG4OeCD/H8zIBj2Kqug44IFhk3JpuMZFlljNNuogIvTDuuxBrwbPInBT
1ijZtj5VO1lL5urAao7lqSqBgqxa4BtqRiHnyALuiiMJZ+ezfELA38PUx/IHgheccgk7PwaDiH67
i6466rhB+/a9sBPkRfj6Az1xhGQ96LycR8FSlt+U1RNaOPqX1MGaxRl0ijeH167zNG9w43GA8AKM
CPRtnKbBDtZBNtFGpjmPCZN80IYcH8YLByDQ5QYWsNFvAvkSo8vmsyqgCw4tmfIDp7Awx90h1z/X
avemRqoxu/MpdKYEYj1QW9ZWGC06iVZgbIAIqcY0Eyf/mxw4tYU4TKFPH3XCrcdexQTwk79ZkcIn
e7NjYg4Ut2P3+DwHQ2+Yas/gwxrA5WpHdGHOaMNs6Mm6I7jkD9JuKxlZvKGVWqfp1/MJIoqWBLDc
pWPQUiBrwx5pjBYBXsFpa/mqFXLewkoWIan+Uw/m/EI+NyFpMChTEirYHtiG3SIeEQ0y0XxDNbLK
rIXrOKWOtZUXjJqheIT3cfcvy7F3b/4xLRl+oiPj0FXeF0SZON7VznT7k+216cYzv5S7zl+2lwwf
MMFyV94SoB+8kamu7ycMr2+k0HleyVZnMxkwAGH/OZZZbe2p6qmcp0ZandjqP8JlEKHfY5xAqz+R
tBUkl7ekF1Szi+GlbXRiS8JwVQmfJHIkgaLJTXNGZ5Wg9m/s798XjprzrK5MiNM5h/VkjbIvKNSj
xl4JIMxYbNMpo5Jx/VVmKh5R9c4UW2l6I7I8xSUx34EgKcAJDXN1KXXMEFo3wojCPT4aBUR7cEEW
Bmqop11H3c+qP5C7lRDDEcuygPYFh/artBXH8SqoHlsNowHoKjbkLC4u1PCNsPXv80mKuXHXeHEM
ypFaf1GiEU+fJtlof2cRbQyMxzy13MWjI0IWJCbroBr897VwuZ/p6q6PVf/fkmSAIW/a1geisC1r
thXfFzlQztX7UqWnlG1LgHkQHyyHEwi0HN65kKg9o43SWl+qoW2ZbFzhEzhUOkz5FNTXyhh7fYz8
Kd81ASuIjSxLuWbQg3vFC16+HZ/s2yg62XQ+A489f3CLUWV4erYZZOPsZFOkaJ8nAxZ89tlGu9p6
KLWf3xTgDbdP2NKjfHu7FYWNA6Hmh7ZnVh1gK3Na9vGU4kp5p8glKW9A32eHm8f3W8Tz3AbRQsS8
IPlM3n+Cb/fxBSAfaly+XwRioD99OIuThMUtwRUn53qTZBlIgN+FnvKX++ldQJ8K/SUNXMH21D85
c7HmmZJz7FAN5D1H8kmVji3n7Cp4TMw9Se2GlA/7dwzsHEVweK2/CDLlSSQKPwSOSeKcVGKWUX65
jzDAF939M+fv+p0FAWbofo4q1w2uE9vtPZRKP0lbk6maaIXVCXWtrHkePN2ckmxJht+lJTKhP0xm
9Zy07tYScR4vcGnej83S+sEQ5ey4UU4/wrnHTRVSYKetxJgYMyj9jkYaEGT6ZL+N978XO5UTbAgZ
6ZI87ArzbqeKmGTpbM/dj1+p+YbVHIOmID8NvkQOPC660Oggf8HQqjg+IXmFDXpKOb7vuUBxvuYE
yLg/C64lv+vgaw3/URaedJnM7UmvGPs84hJd2QUilVQaxRqmnQm2XfZhDv9/gBiRQ2bSPqeVqJzb
T2Cxd2i1JblATAzkBMu6+mPvEO/aaa0yubE4uLyctg5LXIjq2FH2aKX/Flr3ctu/faoJilo2GtGl
h/PWMxm9DEtrMqfSR6Fmpf3y/663FVfEWRT0hNd7AKoqRM5NLyYukp/rFvoRvXoDofwXzSEQ0SlO
YNVsu7zxYmJbryEX2prV1BnJ3cU0+tnlfKUx1ovXiH/XuMK3Pnsx5f+qrJy1LHdfGKlNvJno6bsf
QMdQqfxQc61kUGrjWguOnauzG4D2lYnvDIOUn6Fu9P+g/YC7vqBqm4JDeEPFB85+fKVic5/gvzrL
MZ2mlkm84NHetY+kZCsZYtLfYXqgT4Jsag/OBEKzqvVrUdJcFBNGJTCYaNYNTPdU8UUjAgEwSoce
HW9K+aU5Wd62fKBgjBS2d/1ddnI4jUVzh0wdvrw4LfalZtlPj9/OPcrJBVauwldjb9TadCI8SFPa
YXEnkGyhzZkrtsPd1B33b0Z2xywU9xn/BWKnCl/WPRMPkgbXDwPIXukY1PyE1R0wMDnWAimoJ/P2
976gsZ/k8UCAiI1CvOXTMDLV32UBfe0o/kvrLsorLX4vpQSPC3fLkdrGwLPiTmao0tSTUsfQ06FJ
PDe9jeDAkkMsmUdSX5T8HA5x8FdUOlBj4C2OmONBiPujmYJ8vKcEm06pRZ7zynkA09089wxSf0kl
QztrWy21V61ROzsxgYPuJ14VQ1yzl8i3K//4KBllcPw+dLyyoqSxZ6TjlHjgnWnoOHr8KU4eq/PR
3tR7RJxMA/nsTLy8r0Zr9w+Mb0aG9rikJfH/XKu8oXJbqyXSdAY6BzmNmxeTeyshna2nzEdkQvs+
hMJWdeuQ5pAqWJUXJC/EzB9AzBljmypzvLW73hhWbZeWcKqb3EQxrPhrEHVCuE+PxDeLJ12fL5oG
ONMpmXyFtxlqVOxCqQbosHwoZqekKeYDozLAW1TkeoGzFEcEbdVJUZW4LZSrPaWYo+1ijEcbKnrd
WEDCfku2J42hg87niA0hvx8oEot4FnKYgJWOL8U5GkSzQIzYMR2LovGPqioFSCo4oNcwAaeR3USn
wQpRJCMx5FH83zkh3NdRMHxT5AUkDGqb8Qht6Vg3IwzPcNuda/tlEEefJauZdbr79uGt0DbSH+8u
+FN5lLPa/oc7OVSn1i9savCtKx2xMVVd2pLoa+6nKyREepgYMfV1wqOHd0XCFBEQHWMzHj1wnsMC
9iFVpHBUmrbN+EUokLchrpCDS/7ogfgpQp/lA0qwaRM4D9CcyrKsdrUWYNIbR/j97UaO5u0MUhW5
JF8M/3jglq9swP5Ik8oPSe18k/PebVNoA64mvKk/USrITBSYsALRe0KUhyJ6zW9cVJNktQfB7yLU
/WGzpeTQy+Gk7knBBHGA52hjrN/9OThGZnHXuLhnR2a+rhEeR+rF9ZrastjPBEf92v42MdPlibwS
+nSs/YC+0y1E4XmtTKuuPHGEw+Rp46fMuevJju09yWVjLNsdMHBFIcg3DIdy2J1c77mNDG8BcHPD
OONcD6UzlOVZX/sbQWjiEdzeaWzxsud0CxgtpJ9m2HusMsyuizraYNP/Ooi36dn9HSDNHcx1W5H3
Eq80ZADTfgeRAUil6oWA0N2dTZ/TmYSH6fX2ldHV/mJFOkiqaciXPU2uvrvMPbcofqelBO9e+AIm
4P+YNQR2xfCNVnNG9D+3udjRw5+ByYJI/8zzDaA9SqLrM6TfLohW8RbGCKRj8ktTvtf4x0NRGiWE
Wr8uN1LLoXStRInyaW6bzae/9rD++RQHLBVFlgKvM/T+ZxCPw+ko7dThoLOI/0pGas3HSSAOlrVL
s2QKiaA3YOnJITYZGSVlZ9Wfb4brTYZ3d+PuW3oWMav3AQUcqtsgofX9yRQZFzbwnXRK0JFhVmqg
xNz1l2PAdc94pmLGkk13MnN8zN+v+RNvfaq98gSs15sfXGR+SPnawPEomaURxcZMSju/Y+pNKxYx
0v7RDw8By+qWcc7QF2jYzZunkvNuvWoAaIklu/zW8eHewRMuC0fYgRaj/1mD+aWuA9I4IcQjoAHX
DtxBMMaS2kUvrGvp2EflpDbyUI5kSDk8VoNmeympTb4mBTz59sMRzbE/dxPj441+MnSiHFtrV+VH
Q1P8RGY+Yc/W35jURMTQ4AVbmIo+mfDxN/pfT9ytLLRUlcjyqbBj04xFqVXYQMi+iGCVHQ6gDl+d
72I+IrVShbTNtdta3iYJzfBvPjqMPNE/v3aa4YKtAcGBsLwkTLTsd5txmxBDmo3etfi+ymxcveNC
IW5zTgEzWx46PKlchS8hX+rrCwbnb35IlcN9SHeQFKrkiWL1hgW+LZDm0+g61YVBU4Tea5H2yPLe
ejDGkAfU7586LhoJaZTKgAxWm4sGYYL/9TZPBieLRLIEhXT1sav63HO9Rpsl/yzzJoQ7hiMsdvpR
6DzyeCYJiv8vFdEvMM/7aJfsv3pkcTtXsnu/fLc9lK+/hEtm2ybcPZbBY4AZ+qh47eHD4CeVAteW
F7PrK4d1eoglK/uuCMNZHQRHagR/KH+s77unjRtkCV7WOy1Y0JzvmnE7cVlcQm2pq7eXqAq5R0kz
Skw6C5GifbwULSUwnTLjU8F6apWViHBTwz4cHSLPo79/VR+F8b63xQgEYxxqGv8iTdOWv/LBofc7
oo0lHieccZ+JVMu7Zq1b/Aj7V9Pn0UKyWNA9RF2xr/Y/ewePbUfszQzER7Bv33ZXqiXWjNXWrOaK
SC0TcuwryK5FyzN+9ZxS3YUjPmd1jHS+mb/EOglzbvGup9MxanaxcwCnGNZtQM+9YgekAHe54AAJ
zPW8NHNbEH2OMO0o+U7IXPVgbHk7Y+ebgbsSKBmKWVeZ6na6LH9ikpsRGKeS+cLhHkM/HgPbX+BO
+maiNI9Lb2LlZdGc+6PHZVjMZMwe0LiW/xMSoUimiPmYXm1IBsdWINQwK7Zs29XCkeGi5dOv2A5C
fSF6D6CAogUX/eA0TluGa/yULd7EBGWkU6DmX1XzneDO6blzMa1ZqKQ9dEv9Tz2gxHLG+g1DfjD6
9QobCekwTh1lnmp7omyJ9Fh/+0s7AcXI3YS7e0yOFTzXt7oiFn0tAKO8Y6SGOLVF+o0/MCPuXTSb
064RZvBhhhykYqYcRYjgI2WT+e44LimcvWj9jV7lHXJ6eMGxYDdbJKn0en23Z+Fe/q1EW879CQGl
RsxxNoPPrQC5s38QMINZja2eTdUaEhiX4Dc7soFu9deLlLjbfOBIn3z3jSqh4MjvLPLogU369QBJ
mdqHWP9sgXZdlwbyFUZ+U0z30lv6H7z5yZK1NC86XCJHLSRL/XRGDBzO/VO5ll63DhbgMG1F3MK+
4rM8dA3W72k3+31R7ZzbMsSJGOEL9opq7XNEWQ1A/8tMuLDHsXB5oTpa0XuvI8GSab87AexnO4dU
gr7RjLjNhBfoQEwjGE+f/+5f3eLo3SNNufU2PsAX75dyxjY2k7KY/Ps4AVi/hiGFaX9dhHmjphao
R3cMKRud7qOC2lD9zTv81zPz6kLibp8vIhDR0rzRzMeNoQSiYyC0esKQDx0+51Rwf4rJNIS4dx9K
zVJmVAZLK9VMoe+t2OSkZ3KxZySbT4PlCg5mu5BIWAfbk4uRs/Pirk6GsNVw+3PDIYEL7gfTLwHa
uPAIRGmjOmTSSHOBFoj5/P4ffNY0SReEZXVD/qwiekIjamCFQH8XDi3hS+FScDHypwP2IFW/vE6t
pYrE9gvQ/JCY37qi65ZkcE9MN462Kv5ofzikSizoems9Pga6T7UkZu2N3Fd6cYQVAdKoo09s6/ka
gJml+3nn/SAyi43+f+LH0Pjq1SsivOHqSKLRWw8p5hLceYmMtnnN6hkyo5OICkw0f2DmfAnJXT9R
vTEf+clLaxC+ToJccgP8icKvH7sH3k9NIdnA6cv5ZTSJo2oQmT2F4Ozd4SRzpQcuXWRUteITm9Ih
T2hCvwlpzbzeTFl2XIeHR0Whiuh8DYuNlttGtKFhnA8+4RCXePkcCt2QeX7fuIrmdZ5SYe9jGgHe
jkmFfIQx6nsLr0v67rinwBgRtl9M+o+LbPUSgyyUXyDLjdQAMFVykKU2NiHC/dcKCuc1SuPF2Aq9
4RmmZcxODVOT39jTn4eSupLgvNLEq8mb+ypshEwk/iprYE41eKBUNR/0SruNzvWW5lWPhUnOOu+s
rTfbBMZHsmomVXFo3umAZuWnBz1f4ITXcyiuCm5m/zIBV1JQxqepQ3jWwVY8IdRJSJ03pvxbX44X
mvz82Ga9Xw5DmMH+fOV8V9mOMLKiIkv4LLIrENZEA23hpTW9lvZvDrB/ag7UDjWsQLbsjPwrpMNI
W8VmU2ZBVHsW4g9Be2l3RcgOf7MJyHxMot6lh6g/E4OglTnQI1q49CPIX82NhJbQQG3qjYGFesv2
S7YnwM4ZpfblrOVTZ7PiazwvknXp9CA69Lb7r3ziwBGwvYXVmZgzjMugMCtPDKOC+EXkuNWbE2g7
KEeH4qgBxLo7LG0dCyhmrRcwe66MUMLjvVdrwFWyyD+t3Uh0OZbBLLcMIENcLTU+B+CPuAXPa5Yu
7v/3pNwCcGW/uSBEeM4kysOR+VgX5gBieYGecJ9SQnLeoNa9Sdow7jME0Tb2gPPSCkAOfLGOjf1W
F55iNge42Sz1LGz3T6Qn/We61LKsrHOFWu1jkoyMIX50uw3wAHxxQA3iGkO+YCMKESlXdixX62eB
IEvSYQYSx086szduU8/oJh2vq1TqFtUMRSAT9RiEanvUxDMdwDoEld3sFgIkLviKX/Qry85OeaYU
qwF8+brmPt0BEl8QpFePToNNCzhLleXrf44pGOGETtQbtxrq0e2XIGQN23MRPTHkaXGVTwZB7bR0
QM8Dy2E9TyHBdfZXvCsvSVFWbqB+pu6xN2vmFt6/1VqrSW6q9H9FszJP69OH4jOL454ITewC5F++
yyzHDQSRh7aK7LDbdXeq9W9g5yxHlC+DzdhcJ0NFlyI1zoszDxQQQ4xA3SBD7+POQ3QWfYbYaEk/
XQnXfA5JUjHJxT938M32kfnbHiQxaKhESy4gEbrBcv80/+muUmMjxEnwsO+QEx5yQgpURpQqSEjt
dtBRA8h79G0uX6epBDmgYGeKoLyjXz2JUhktmJPt9I/cqGbF+h+Tkow8VXkaet33xFlqkzSId65/
D2g8LwPdoiJq+0NmaZtKAP4uQt959wRAmgXmxqsvZq425dRGNvZMnPaYohfxVLCV0Y1CEe+2naC0
sMO6jgDTYNxGvzDD3GI16fWepT4zGEjth2INT/Lk/Ovt9SuGwLTbfzivjSSMrzN4oBHcCNAhyxOy
uduQXOHU8kc7z5mAH458P4z/aS5EyWeHDEXqibjbycCx28/M7sZcBRgWXaAGJZmSL6SFy0S8gfbj
CHf7BVa2Wd5m4QMIoe2cZ0UHJEgW9Tork2TJDDqskqhGCceeNnmNOBZ2k/v6OVsHD7JTJmCjz40w
zxziiCjfmXLl7ucrcT5eMgdMVkIReunGXa+TeGXRTwT4vLfbnkkX6wNAOZdNvgJfdooHRoZfgCgu
fXM7wf1oO8FR/cGvT0t2K0AgFKO2v6b3+VFdgJtGl7KVvKLh4bhekMr5KGwaFYJ7fHrB5lHbXla8
N77+xjpEMM6QH8aErFbPArzpBlYQogTzqJPrrwWax9XwIYlRD6tiqjmYhijso0k+kLj7mRkCtFVL
UovU5m0eUVcaOq+Ez3++4t6/kjHZOPASl31koepXeLWAAe8YKvzAMaRdbV+Uaji7FlA6hdIMhKLw
Q4YgyPFPPOJSpTHNWIad/L54GD24ZqWAJ+dfUnVxPA0V59lFL1rpbRUGC4QFU/GiKiYjHhEvguth
0gOMmFOthLZ3yqu30FxfLBlx46HbR+6RPbhN7mCETYPSfWaMNssul3BCUNwP2ZqMEN3HnVwb+F4y
BLY386ogT6MSDPHr5iarwznZmtuFJMfCNofmjmvpTmgb05qRI0/h8Mf4FKYO+F7xwwffMWws3AFf
2gzYvwamHHFYCsxELErtE4RvGUwyOkL+PQJeXe3/uOA5Sc6dd63H68sAOOp9F7/9tjbpYk23AVJ2
RoHz15HlG4+oAKWje5zRcTtiv0mC0JEsYodXrioivKbMlWpOYxMyTE/vkBbtp63Vy5SCbyWPu/BS
k6vo1YUx/wEtVeJOTTisL4i+EyqGBBiOwF6UhvWGeDmpXn2goU2sc5ZfIRK2CodAaUic3d4C26bQ
Vj7YDNiag9rcjdbr6ShjkGDDQS8fj3/1tkKbRd/f3z2N28M5RmgJRG+hGeFy/OYb6IECXGAcdCVx
kCB5DakWsnqyYEZXpvqYWF9NH8yT2eAWFUzKWEfCy7GRfEiXe9NzqRpQgb6FGOySPTxRGJPji1KI
xnGwvjVdCvhWpqPocPa6APolQbuNdeUxLSNx62eV4T4m2t9WD+yx1NrxLs1cE+MU2Cz/mEITLeW3
UjBgkzgcuae93na1YCfUN7DTvXax38cPOU4ptbLVj/QbyITrIhAg1RMLuNYbUu0vNc7yOh04qZjv
9NdXIs0pFRtw2wABD2DNa+OZ96ZxSGrWlOTiz/WFqR1EyozEfrF147IdkZSVlEqS7TlySsC6vunJ
MLwAzx2qNR8iv/DBIQ9dPkr3cOH7/mdp33zuDfUCQm7ocXKWKrMEPJecDfizfzzLLPSltb5W8l5/
2KNP8dt6AHnugHzn8Flehmo2bO22dwie6dbyjPDUU6tGKhXdvkUTbbj7GL3NkVMkqiT88uXiiBME
f9UTGf3MDEP2ZRfEzObFkrGNGFygUMEoKmP6z7Exyh06/vRSL/YKxXSRThwRcF+Qiic/hd9KWO+z
d37mciUsOfNVFTHptScYCn/53BkH1lHTXbVUeHFQHtm3bPBUqPh0yyLIfb7u3aB8fnZIMeOXpslH
KDpr5naeMX+4BJB5VAQ8QoWKm+sLy+v3oiG0F7iYs5Qn5LnsRUoqDUxGMY5o/CF4MHDXlRx/H3Z5
CaHvWLWWiJO+bLG5Kget3+Ee6DbkGqzUzB89jKw3jY0rH1zbJlikW+CRWrUATlK2Q/2hcZ9WqUt2
L7R89KQzl5s4ej0XZC0dfkaOVAg9wf1/XZIR0LpXpoCDr+Q9KHU7fkDAXfE2Hd/+Z2efG/d54SvU
y9qixF/mEdurD7VNpdXrmYM/FCYFiFU/qRByDHEe0afKKUlsVyvMyCXZlWO1UmPa+VtQN3wocw75
GuOpU9dbbjt1Rl7M8XxRylF+tsqf91O37QQHHJf6QZrh18pqlLgHAcGIXuEiYHS4FjUQg59RRJL4
P+mMgEEN2AK1YH8bslzhNxiM8gZkduSGGzbwkToJsmYEuVDtLrsvCKaA2YMmH/XDM6droUjXVkb0
ob1uny/vUPUGSTfk81r5h+317ODrdH9uQjHoiwwVfC0olAzWN0GjZfc/eUq9+5bAhWLHe80AIDId
HVYD5mF/cJWXCActokVp09PAhS0AgjJSgNk+tAwh1sCygPIregRAuFwe+BFTSngDFi6SSpx0LIiD
oob3iQz6PyqwnNJmpN1egellqnOpR0VtrJ15V2q+z6igd7IfuY8lXqDNkIEKikbwi7vlJhiTMMPu
Tl07gxUNXMWE5T+Wb1zI2N5HQUA+y8PLhFOeNaeP6tsXdfA0lYOIr72OptSSFMJpg/8Ddf5a9jiq
u0Xr00YqTappCtxRx5oa3XntbRWiYMP+NxPZHhl4Lq5+MoejztLW4n7jc4em9i/zBtB4rCQPDrK6
F4WqD1hoReoWIY5FvSq/H6yx1mdTs06YmKOM2kUCGsa2Mkr0OQfEqwPX12vEITKdEl0e3xQ3dcgX
MQqBLTlrKSyR083g94wki5EUH35lgPv1nsgTpK5k/I0leWpnDpZrcILwlB6OeWi3T0HZnNgpKA9Z
E7u4/G+j9Dv6aDdW2/x7cFBMWR8l1s2WG4tevmBMY72EU+A6LiAiaUUY9gUb2nXaVbPtZvm3ZVkC
Evt1xnG3lxTh4eaMFL+B+YxQbj/ukm3hLpd9PSwTppwUskwnpVt6135Al1R4G2Vnu95xfWEHeMnW
2zkCC2DcxQdoOBrvnRnjojQSdBeZsihEH3I7S+F4ZcfMgMrYXZFpIuOx4O77b3a4wNBUHlCugXAC
ChBsoLNCOtUZ8icku042utKGgO42fcBbuKVHU7YHYOClkZw6boVhofluKJ3x+YtXOAc5tHrd/wu2
FGnlG3RxRXmZCHQJL91Dy19KzLCkOmvKEIaK9sTohKDpQk6M5spl2hkJK0kgIQXBq573IVH0Gh+w
BXg7mle79uVcD8qSUm6RqAg4b8JgUA4zKsbt61TNA6AXyPTDPtmv7WTZ/5E9Y5/Z8Rvt3BmEHr3x
39qj+GEmYB6a4sZJpEnZHiSy9ZsQ5eKMef4P/b17Oerpx1+6svR3H2Vm4Vn4cPu+lbihq2jjKXca
iI5dFpcuQfw9tjSm3DLR9jF+udUcymc6LOj7WIdqje1NOvID+9sFtKag2v85jYFsJ6jPBrvqPfRd
Mu7HLD+DyHNW2UAThNKj8/AuJxyHiTHAi1zuaW5zr1kX58sAcBxDrdh3javyFAtzwRPitUUht1OQ
JyaneRiOP8hoCaAbj6bDN2qV/2VNpKLeu/JmSY7k+U1BVVR+jQElmgYMfKdKkNBrj2m1IY7IYY06
rZkDbIxX+ClTdm3y4KJ/6FHrmEzMnHSqnV9NDGs90R7tyeG57Xa7VkkobcksxeszaaQxp7Km6TJC
SPmWn161FeI+lKOtho2cCUQtaF6YnbN/fjZ47LRCBWHF6BX8EfT7FO+LF+G4n6Z4/rGNw41dbxmD
lQm6ZFeKTsh7KDVGEHCoKu2qOjmjMDiRLfxHzzmyzTM4PFnbkBO86l6oSnOrC01jgT10xi33Wmxn
DnST2hRqq4NX/zBvgFHn529NU+hhOEmNRUqpW52i5PXUgEzvFr0vJ412+rV+53brKsa3z/DIUxuz
WTCzsXYVBuckFwyx1roxQZTNcAPfPpR66dPFdYTKtTfowjICpMGB0uqMfnR7Jihd44ycM6M0Do6/
HHeQ2atF1/Ow4hlKz9WAokftqzOz2Jc7pnUqBvn1wgNi8X1L5376hOjFAC7WSf4rS6ljgOG/YuT+
MaQN8GSwKwBXY9VTb1bTFwqnP1ONSb0hpQMTPXusoeBaQKibQ5dp0fSy/NqmnDVRbykmDOUDfKxD
+/X0yVapxok4KBK6djdILC05HAoop+w0rAtsnBRTnqMBtpLxISAhpoU61QQXqteHmLxKBG1q/rC9
K/nE9w4od62cP7jV9Y2bRvV4yDHdm+23crQwaGvEMYUAQsid4ADgCDjwq1IEWbWvDPSSXQKw4S8r
njxdHz79aoNfZUsMsW/535QGb+vBF23eS0DCmDwgx5z4I7ug89G+f73SlAQi2QGfkFETu2BuA9fS
YB1Xs8Gr7aG/dcFJk5792GfXFYwRwvQNyWxMiBaYR6eGjYb+IuY990JU2k3zxToOqgr4yyYbEcTj
1oTd5OTcR83dV2gYfYqawP4qGz2kCixf/z1P27pWROVH9QiFfY/HDHJ72Zrhw0AwVazb1dkRNJGa
jLz0H4lhZZh2U9P+rZEW53+wM9NuVp+uT9qMCMo+p3YfZ5fiDXncXHPcA1mkhvpsRjL+kRV2gnQA
7nCIc4MCyFPjGh9sH5GTtE+MigqNCVc6M1c7WO7jEKuKYfWVdeQYZy137EGR6T1oLyx8KQnSh8jf
wwkkp7yV0+kMC5srp7aFjE2xQqSO7DDK1n8EJ4l5r7yLrjxhQ017snv7/874KjVGPIYz6MWjXaVl
LckWNONxoayubVEYW5h7yJDq4lo/MWOR0Xj0ewdAl12NzSIJO8NIOeuJ3+8nr2tyMaK34uedixgw
jvs4vSVAHGXpEk63KKGgCjriCgP/dQkYRNbsxLzTRsCi/4IffK3d37zsVjFFzNMdVhqN27hw48Av
tG9uCtYScFDqdGlY2JFIqMG+d1r/RE8XHIxVWeH+j9njJ0XH+Eab/1/QyJl0UL9ffwtY6TngcBEV
0cUxahwwiZCAahHIoPb0vzAyXoVR98fTQsWbmujzhHatg0e/F/oQsvCNVXAEdsVViTLTHaVVZyuU
Ddzq0lBixTeo/LRifNjKJADAi6ohkA3rSMMDofY+jBs5vK8li11I1rrMiaYVMFeH0ym3R3/kRNA9
shFM8ezd4fS95m3ZwLwfh8nbnF1cNQlfO3sS4u4U1V6BNR6minO4w/hRxlUlAO39XUMyA6/khTDz
dtBqfNvtUGv3iR32CUGQ/aXkJhO54t3uKEOxUENOjwDX4G/OQFwmDepelT89662gNsAtKXLjNhcy
EMOGKYgymVJQJYcHadr0l5ou4MYK7UOfnaKazHWivD49ZS5p602FQ9vEMiUvAfDf4yD9w0aT/omk
V+szRc+5dw6v3pBSrlsK95aywy6ul6Smb70MBGhZrG6gib98NNsPFCx5Tg1Mjbk55yndNj/kBJ+P
UI4rlZYkmMQkHHc6QZa2o7+PbL/E6DO7CfM2nQcUBc8dwlj1h3ejXdSSmVZgHRBcRykRqGytXXeY
1EbL2Gqz/k8e8GLu7L+h2OrM+LpvGtducFLIshFMzFHH48mWnmho1plW10yRmD7CMjzn2fYDxXXQ
/OKbnfC31xNLyznGbWdrPnicmA3egdROzMzHR2p6l1jHGK6s/vFSWnSrVi0AYOALG5Bo5TmMyFVj
Y9ZrcCVWwXOEHX47yjRbu7tZUsLowdfMG1t810rZGytryy5ZMVBnWVIFcpG6bPfJq9WWhJj4RLf8
cV8Nq3N56cUVu6fuQADLgfO9PI5u7rOSMjSEOCVCioaEJI4OmwuO4bBl4l8VmDa5v2W3DcVvyq2S
3POW/seMCUCwIOHia5TK3CQFl7mKdM5wZE6TB5d76NPwSe15sPoB4e3CrzRSH2zeJBc9D5oKaZZ0
skJdoritPSmK4WrRO/Zdnn4BS3IQPIsolxnpwtSCTUkkTnhvwEubEBVuTxgSnNivLLeGePYZh+SP
76/GAqly+xC8jU9MDJmcqDZH+Ovd8cqrQQluY6f3IlBpxGPqDFPnC6lXq+QAv9dvbR3QltIVL9/1
g6nEG5v13ZklkpxSfldWswJOay5OLh7c7TT4DpautbRBMK1XpoX2vaZzB5r/QOhKbS/r9s3odXfS
//BrD4U2/gFdOgSC8N0QfdZsqFLCVISc9xfxUQq75D4/349UUPZ6HBXBoAqk+8cgtv6WrHC9Asqv
VN9Ys6s2Lf6KqXQ3iQqiBdFmD4T4Jz4Wn5NTkpZrIVkvCthg7Y3EmqKibUlYgWYg6WY7vBnlXN7Z
tX67NS7CjJWhaufe+scpfDEAS4GArTGo5Pb3xj4crsweh0/Xg7qkA4zvCCraCUemjOfnZizS0qD7
MBVsa8CBR0cvLiqbTob8c3SX1rAdpvueINW6tow0jVbaiHwojYsUBUd7pW2SjtV/KxZs3EFqCTwF
jccjMJceLkiFTBWb+0SXCFqHN+fTeWbuFudYYIfygPp9GSWpzbG0ziiPl6GuaNo/jBU17AsOj73Z
AsCeIk8B9SYJNpAOsxIAgcezYfBkGWeRpESoMrwPuPxe0jDNcdrF95eSRyWUMmlhExhAJ7SDilTm
Iso6XeFeRb/VUk7W7aUZEDtyMIQVs9BXvtwQy+elD0gNkmcEKaB1LIsqzUSEHmf/VcX2ssOio0jC
aIrF0kcIEmdS8WuXy3PZy1X5H2zosWS7VSljI13bMKKaMAp2ZuMEP/Lczkdbrpi35G3lD86tPx1F
l/QwRcAdp+oZUT/eTotfg6Ggjyi4bi01TYmg86xQbOaI5I3ZIMhLRzblg3A379p6INOGb0jdcTbU
n3NqZ0QTLcmOq8MsPwA+Bt3fEwqH48BOZAFmEhvkUmyvYbft/vUyFU3xidB+6n9b/rKrauMwbPBF
3us0F2wGv08fwzOBUh9S2l8PwENuMaMGspiMqhFpY3JGblKHbbF5EJHJ8xBRvCvS/87vGuCFMbpR
oO3RjHnP+7egIXy+2NUyraKZUMxYsqzPYIFKLAUM3xDS0jxRTtTqZp8qPr2eTr2Mo57ArgWZdaMS
n0EjsuqypXA86zlu5bmSJQml6zILPa16V+5yIDu/fEKsZPG+Jfvdi8KnZm4h+Ck9fJh5ObGtx4fJ
b+QmV5ES0b9o/Uk/tq5MM6ZuulnJhH2jBmSev+6wOBNWaCrN9JAfbiDpHbzUydIn/NWyCb1wnIJ0
nVCqCIGYoX3RnmjFooErsLPfSj3KlKqhE8eQLF1v/DwlZ5P2HDnuCBJ8jYTJXZ8JTA4XIXcj+ZLn
J/tBACpFWRombby/7MnG0/IeqNEpFsaA5ypFYwQ8+xQjLh+wcA0ZTEAJF3iri4mQzPOaQzX/2Jk3
dQ0/GU38t6LgFpIPAg0qxejWF8bdvQzzMjKpxYgNQJqPW+S+4gftgJglrmUB+RWw9oUwoUIZRAxa
CfXnUEww6LZRjVN1+CAUwZav5z4zIpn9vTjXK+TSXg4xVnmez+Hw4Yend+DGs5sRJtkxbMbYrcjY
+vq0qrqZc0ueUK3I78GKVrTTj+2v7L9ACaAq5D4z2dS4DGyuqmk8lilW+Mz4x4NbPTWQB71Lrwwf
xExzeFOh2AgVhKCWyM1AmllkPq/j7/RhR9IHcvredS1qgLlVR4iC4cJAn0bfUWsMDfsVdR9zXt+z
nJBcbu4dXbfrYHOcmNSpAoj3U9IoV7A5HBAVJYhwUDdYKBivwwsMUYBztEwSzDYXeHJwZXMHVAZu
R+T8PQx4N2N2M5vZBsPeHSDp8rGd7Up58YVt7+QBEknSpMau7pEi4Q1aJTT0m0M/zX/0pzmSdW+o
2nJZizCDgAl9MGt8SVwwvW8SGkLp/Mi8A4MLRUEc1XzOTSdWiLhk7fBAOp8zKesPhHYxEa4t7g0r
CiNEA7h+8KlbNm+7yCz9W5CqeheGRQ2mXTprCMQDZUESBOYMlBJXFBaq7+NeWZzSeHjT/3CXpns5
oF3ymDRB/djO26jnyAD8u7SmP68dc6G6GWhWZxdfbGh/lzWAQJR3ZU8B+WvY5NcA7gdzPmmB1YTF
B77+BrTei8jDaizyUKlnf9pwGDeXgsVcDJi6ikDcy9pJrnD9tvNLOwPLpt9S7Victuagxjgba17+
lvNeH4Rtq/PFmEcM4Lvi2bmJXIBTVSOUAWpOELMcOjKj7xRWHHtjZgc+rDnfAjO65AzWahgUbKdt
deE/nVypkXuU15GIsgXcG9qmrW+jaPFBemiVML0XmWpH44Ht7iXYhemmwda81gVQrJ0R1yB5687Y
t40LsWxWeh2nWUe8MtKRC+qFDCUJEqYXn4EPjPEaHZGr2UDCv1rNbJWxFF7UUTmbWrG+Shhb/kEn
V6+TzX0OVc8tI4hwWhP5aatShd5MNf+GI9Ihfa7b35ZCuBdgpn43kCGPC5fOFk4TQ9DqxAJQYGh+
IyZS/j8X/1QSKDTigCDq9kVzCinM2HXI6old7XkO3tdqN0zg6snAfhDvv1aYOL+zR+eEaDFeX76C
BiOTIU2WUUpqkroQ/bCixcnyNUIZu+nKM2LuPX+qS91u98/FjsXSkFr6BjM6f5U4RJ+Jz1Patgv0
r3QkqoSZWuAV+E9PVJaOiEmFJqonnyFk8br93Ri+HvJ47h8CdpwjkmNquOU2llovhWqkWOJrAPBn
uc98J4fGVns9rChOiSvBtmiizaACF5i2w1XAJM0j+jDCAusbMOyylstAIZqdz+jNCI41qwhiooOJ
qeb1sO1/+67vdKO4KrJT0mklYyoFNtjGNJxGF3lNKfvBJxM3PBOo9NSBcSIEqTabFgMqqs4XdykO
7ZIXpqUEXp+0N1WSJHpYoMVTnW23ixfRYvRlYI1xsY1eo4nf6VHsxKIHTqF9pPIlFah+YQ8kykNZ
NkDIj/igLNvFuYZN5dJuRGZAjOGw9e8742VbZNewPWo8ouBpWEPF9kgiSXDXYM5vzqm0kYScubJ1
QeSC1SteWIwbyAwF9LVTcxe5ZxYHd7dzPJhNOc+2TOCkPnQrxcBSp/7oZqqRvBrqBYMqDXrWGY/+
53pqlBTjRkPKrRE3udM5M6gLTY+wD6rBSrwy/qbT+DR0SS/Lu9oDmclhmJaxyT7bVxsgdNiMi12h
cIJyDcfXhw+UbjTUNFc2TWsU15YHOI5zX/x85A3PGrAZ0fWMIkuw/aqtXArYDANtxenYdEaqFf+D
wYg050QuYN0TFpFw2DbE6NMEypUtLDSLKSUhHkd1pqkreG8OeEE8X+HBCOVV6oJIsPg9s9NElBs+
fKpTpXma1ZvY8SU1undjErTIkp4GdluvqyuxP8m/jFCUn7/1bzkQoduvToCMSUXaCY2K9nLRR9gS
bdP8lfMk98YY/ygmTor03f/8mGHxoOIMvbewAjUVEUbvcaR5qXjH7ZW28ojsq7NF8oNsML6bXxWD
sy0trRvdfuwKP3PhqVNifxfHcPoOLoLGYHB7clnqa/9iNBB18aKPldO5q6TDqgGazNk8e1b6e6Yj
MuW2R0L1ebK95HnkAnPpxMCzYmuvTo2vt3sxkELi9iKJNqub+jPGxB/2Q+893ThFnsPzLgVRkZP/
D8WMROhraA9HgZMch6WGWQLc+EhixNoy8KvU+BBt5PUrwOv0x9iEulyKnBMw4vQAjTgqlMpUaZch
Wyxs1peNK5iKKlrz6+CVnmWu6O1ThN1NsHDBuEW1aSFaXQDyY7aeGap1I76TRjv6fHiJTUo2VacU
We/mWWwpdl6r5tdk7MYkFIcK9R4mXbSmLKfA5vYtAVfXwKFWlKVmWg1e6sednz0MUlqTeNFwBqnR
XycIr9RH4LleRqlgh9p94Y1oN96wYljs7HYqu5riAifDbmfdiJI6iRcuLJANdMdVDiAPb9fQ4JdU
cwJEkai16a5BWCA6hcUeAr1qVLaKDLOyPu0TeRssA10xaFz1KGQ6w33ywfsC30fnPCZlUW79rQUj
LEQU/99tamkk8MiQM4+KPw+LppfRA2F6Sl0LrnuZBdNRxssISCcyEZ8yNPR3XfiR1sVBogdN03xQ
kaJJ3sb2i61jieQjgwW25aAlyhtBjijJ0MYia2Bz1uFJUYZKBpBNMwvfF75Kkchyy3VSTqz+akje
/2CezImALCoOLzz7hJpFTeZ3kDjhlSm9H8Pt/cQHl2ThcN7kpGil9XOYEctOQEmryKrf+oLwknyo
tY8kdWorgZ6k6MacVxgS9g0OInVjZn3HFXrp8AVXCiFymSTPuieYxlDDB8QkkdfEo1ZLugAqjpP5
s1tARqX/PQhSSWO3Lh5taMsrsdZeOHiYudLq/7E15j0lYDjTl9uCkGh6GK59BofM7sv1sjhitaQh
lI9qVkopyHcoil7qy7+y0kYx/w870ehY+CmqNI0Jr4lHy1oyAMEGP9f5+uLupr9IygXqZEUWsukT
x3v/IJ5TLcr66Gozi6fiZeV1ZmEqHEbXu6yCQZtiVhusfEURt+U6TkO+et+ldXosJBc6o2vJQNkg
1ewM8QgNSOvHbEwkQJ+P7BTcNyYg9a4801g5lW8fZ8Lc2G1OU/glZ/aa/0djOonYGuJCVdPmUmRv
AM7fpxorsT0QIfJ4R2MKMWSH+184WBcm+QnjTYlJxY+QK82XkJo34O7zlg8ZJtIsh9gmGISyvLyy
ymPdDAD5AEJiOZAufCo+s+wPFZ+ADLdPC4aEHAaMTCmYr5Ny04cr3pqkkLz0J1RFElmdK+/923Re
nuUJ2neUdoc7PT5J0Omegj9Zrfmtykt6dP5Uzve/dRbtBl5Pp5ESU7vTlQR7MHXznQBfEC4zBH1c
NGF9VhOlDgLcHqUyzN/2l/b+Gd9Te5m/GsOEQbxjrUBDK+IqMHKwCZegLMb1p/XQ1yCDGQLHzvD5
dIPRyvc2FWDNJM+lUdj29SbBZ9KeHyFtKzkgsGwv20knEt+Pg+S0v/s3Ra86WUzA1bNW50B+Ofz+
cbFmUMwahQSQ6S34FRpsaAsIuaotc2AJT3syz/W8q84pA/RaZlbMp8Qe5UchlzqRgiHa+f5gy1tc
kczYkza664d0Y05KNxojyBq0WyY6Xp1S4vf5s+E3Zr473E+shcNitOV+0W5jXhjbseGYWnmuq+i/
yarAtszFpSoHIod7Swre/4gZY27Qvow64GY0ttEC7s81JfwmTiYN4/mYayJeO7E3OMO+tS1+FPVU
tqyzYEBGsaNMjPcM4u5Iv3IewS/2CZzcLvWmZO+PFu/q+z1vWQutk3FHRHud91lxZdiXOIkLeKUn
uK2hlkwi7Ps+0/RXeoZAGWj1YNuHynvdvJgoINA4brZW2ENIlXxKVliysygCdRMDRTpc1hr+pQlm
sAF5S7sPply8aO6jAYhS/hmrgtl9xcNku31io6mrwJQ7Tb5zZKqw/a6BM6l+lrZAGNgwujqRWooP
V8hJYXdafZdAzfPNe31ePnnvH/0WEB62TzLMb9bigKzsDwnXJhSYIZ+Rc6zK2cDE9piXKmDz0paS
7or+On9JopN6HzRDcCfNZLmb/JY12zvic3GK6P5dDFaEUGVqX+TvdtpIt2YZbA/xCnvAGgVeYgkW
pyg66iw5oqiILnayTY8JZYTVerz/+uHI/AAm/oqWRxmDNDaFAserIO5eeWcW9f+z99N6ve4SWs5y
w7x7hfYFKCmZMhjpDbDPTYapjvwwSEzhzUkb+zTN8ejIMwEIyU2Ui8+jMcpZGQEpYwqynbc+POAb
cFAFL/drL6crENSY7zwjSXOo7g/soNVEgdvOaA1do35TZCGxi0QERy+GXiZtZOVHsj/K6vA5lF2h
ClyZE8UX+xNCyvomSFLocAoVmHucgNn9sEp95F1bW9p5I/jzo2FttcEVjn+aTAKN6gj9WnAxnmpl
OQ81Y7b4hHMPTJTiLvbQbr+Rjxzj/HG+cL86oapeKpeiTlbzyTqjb8FnlicP7wVMhpBA4+mYxTFJ
oIHppRaB2swifr+KIrXo64nT9JP6j/spqzLQsQBnFW4mCXxch0kVGqa/HmSjDFGKMW/ybEg25JfQ
9Q3/W8mZWJBu1yXywZz7TOOWP5gDgMLk75X57vo/VOOi0rHgXe6AB71/8J070X2fBeT8cJgkIfsH
XAb802O5GNaPaefgJpC8boCxNkZ+RxfEwov4u4Xi4fpWgJ4JrOpphbkBRB9P72p2YIgcRy11CTbd
z8hZmC97wJGkhnJ8AA+CEl6GIitgDIT6QN23Q4vO/UpkKfgMueAAn5G7rnK+dK6PxhYcdKdy6TM4
rVpXa1Yzpe1igBIh0G9/jmFU7Lhg4f+jI/rcxjg0+i04/MNOdzRufE5liQaP1qsH52xfrRHrLtyN
pvWYqxdha5iCBmCND8EF/Iu9xWD0eNKZ/A07et6TMx/3AixF0yrrAf8cbh8eiDT6Qqv0AFylZdtP
Vk5G38h3qRCpjBOQKGWeBI3h4QyEnnIoaxGz+wMy0A8daljsUCk/Qzy+LXMf8U2wYganPsbyFCyE
7QyS+PgkKu6HHV+ErzgQZi70w8Rz9nqVr7eaba3CjMfHN7EF2giK64SvGRMZcLo92yOzUPsHeaj7
NYkJUSMsVxxejTgWqoKr/Xr6bIDg/+3hJWTQ4XFzfLai4z4/58v/mWzoJFIU5CDrnxyANMnyaYSC
0QxtixFKJxuQA85lCDt+OcdpX91O4Luv26jsAI1q8ZJgl8UnUT3Dy3xbrLMV7upgW0UeDZUXLaGu
3TY+uKcfVKd6wEDCh1mWyEgy7XcrZb4ctQINAlgquEuntjAM7rMmQ+pgkCMjn+Fz1jtY8lEjJ5Pj
+6Tr4ibp70J1QAn0iKZtzWmWDtso9NjeIlfy+lKk4JFZCfHQWoD2UUDGPCfCOuHdKfIcRQq5s3pf
bBtKwVLGN6+hMO9xOeLl6fhBb2xrOQ1Epi9msIVYetiwoMw0Tf4AaFDL84LoAhnEyZ0ySR3PYwRP
B2HcWpUF6WRX6aiS61imMc6BCibAHZDEhT7o5qpn9Rdrk1JKd8A99w4OcKjJ0lZn0MRjGh3vPkO1
ho/+N2Dh02Y7Jqs0bh5jNmrRMzOS5yYguMBHj2CKxjp0wlw5VA74uWtI54DeNCqQzd810Mk3/iPS
zk1uyq53+5agRQIKAtHm0VCVc9dncqwhoKe4Qf4nPH+u8GP11C/7zZhJ8X2cML0DvQ6QhXIEsvOt
5XGg3scEC6I5VByVY9Cdv//WK/dxSTRyQHRoirHP9k+EzKrgNhzFYDE5Z3UtPCuzgpc6iwxChBnu
x/C53trvAE1fRUi2VyckMu6Y9acw7E9S5aGWR+VV/9Tx2Y3p6pi0PBjn0dPZpUhkPDMIT+WJbY1e
zFTbNyF+uerJj6pSnRlD/VeHqF4rXxlztjlGhWmTwj1h9G/Q0iy+5pYdjjPg0cGwp/Z7QBhu0UM9
7LffijQbI5PHvbSVyzc4079OejGw2z8iCe/Ia+0nfaAMGnbL7k7EcKw/QoAdDJ/yuZvFXzdMe6c+
5+Z1feTd4dO3ZARWjYcInZb5Nm2OIFV1VcY/jSjuGa9GxIemcAplVZEwcW2FmvdhH5295gBNxSRy
ohBpNOq2RRo7KopkOxLzk0jdBd2+0Xys3yNZ9aI2mJkiT8ooWeahElOegS1XAhaGPz1Z+ALKj6AR
Pyqa55swoCer/VKoSDQ1bv1racpz+rPzmrq8urg0vkOVWOeiVBlA0zPvY+cOQf7DhjzxS7FXwqFx
VAqRroQfDY23vtfPuk2UMZwg8rh18RUAS+nKQXrce9kQ8LlFiYNqH1NiEf6cPvIVx4lEcYGjLf9t
lilgMV+6/f/MS/e6Nftki31TOjDA+6RvZh9svxq7/MvCG0uvzHToWu+7S7rfbUnPUe1tEXL1vEiZ
l7UP8dnHEDlYrL9vgE5Bz6Pyv+Ll4kmYv3vG1+wrfsdjA3panlu25G4Nlwnpg2+C6vb0RHj8Ruly
XNwMepaKoPvYW6gWLwsnity/f8fApLqnNLRpQ1xcdTm4jPjjwqHne8RwvPMOb9dtHHj5GXqIZE/i
tI7bDubz+CsxjbqnRLOylfnq/lxgwYEG5HU+BC2vwSGMfVvegGqbjhvrp8FusKZuCNhVmCMKbtsh
eiRXEYQnlWTWbVECAdgPhEZ/GV8R3znVxAU7+5so7SZLm/KPmxVxfiIkn6KVZk2fm7Z37JTftX1P
+OJUyACX91DlZO5vgm/SFSd3MRZgpm5OPvHgo3lq5e0S4hAcvb5jPKuiK8FPkA3I2XzqiM18Dw+h
F5MGvlOoQBR/cSXu7EkUFCP6mRYFtFSqwPl7N6myQv5VPgcoF+xFV8ET6WVv2qC8PO/bg18TrKDf
K1GYhUxyN5jw6+YOhDtIrMS7zxNbQiP1+9Kr/MNXIBNuFuJRRp/yYprpMT6LJL4sGjzj125Pvb5Y
VfpUHEm+DVHG04F6u3/L4cBlwQccUxWUB6DFSiZGu8gcblSRogGHBticcwZ04SEN9NAi2gAXRC8v
marQv+RqKCiD39+UK39x2CwkVYX20vhnsMQjC9YkOEPDabulgGnDGPyTL8iGu8+j8vBTnGMps7/n
RuQFx6fs+DuY9nUEdPkF1utMyZWGaIrtBwwMkD1aTAYJEUdzickqAvvfXwn+SP1mVxOeUdGeogOw
LVDH7NH4oNdTz+mcQtPKVa0N9lL0kx+qQlJQM2hyajVWIp9bXbifsqLKvcayHc8LwzaDza+oa44E
WpNgyFPW4XTpayUw6EXyOM+nUdVEEvQnehgd0tOSG/RciaOQYzcDLDAQaKdVJU6iVwe8dye+OHB4
4aFqpGPbumP3ySdaUJShNNOBIVG8+erMsUSp8WJtfDNCUSnsiXCEbOFnsHOuVtDYUuzSd2AyEfYH
7rwzuuYFqFiT0U8km1Tc8HX9CSYEGf196Llr1do3El4pYKws94Z+zq7zNmopBiOHLOYCoD94ZH8l
GsTiiGY1mNcn4lSlUdEr/24T/kpufnEgocbmHtOCBnByQONSnA8FVRcuwmiTp2hfeCvTHTG7gAce
swyxMHmMuh2nYphaq3GlO3+O1qr51/4S8f1lPue/JjTa90fSS52oHtQbmePCRs+b6Zg2qTnHZY4p
354xQ+evJoSh6Y2LEHOxF4xrpMf1+GcVyOzgb1lc7wRKkyU+Ul1I0Jq3zS/0fDg/Q/vXuCyTDxKt
hKoO1oRKb4YeJuBZmvZ6GshVwSNbLFdRqhlx0JFjW754kAwV/J97u/pigu/e03ymapSZF6URvH8U
sPZ41AHfkSiiWaStZ+fVQMIYTzaNXtidSCugO6AskRubhgchnkpaR4O9FZeyu9NsmRR5w5lY5ryI
YLaqAFL4fdwWXdNXHcownUL4UeTSHvLpc9opjM79IGBXGNYCJFVM2ECL3CyUkPb5wyHCID42jSas
DkkgkEiLr/fTSCfOB7BFCthO/N86dPyF8VEL2us/S49+vEWRT0haAH2rZBIOItpGIqlw0tH7Ysu0
mVUmdYN7v6mvV+SeiKfswmhV+pHSRyxFSf6rcOHylgnxc8LZwq4a/E+lK3TtB1PAzwuX57H+aLxW
f+R8SDrzd/dOw9sDlzJSOTKUVDrAt5/FvNNVsUfOHWlvlvOJYH3wWsBU4Zhjpcf2qukomqhBsVb+
DbeS9cd/rj1quWjRXLX7RiB7XkoiqmYbMpnqBuZLzWvx+hBBnnKiEz5zbKD8eUZCDIbIbEa+b884
qUz/bFIfveVdR5F6eBDCInkrM+oojS+Xx38CbLQ720jWgIKdGiwsaxwhdOxg6k30GkO/hky8EcKh
dJ7hMZPlk7cshydpVbaK/NtxB5MMylz8GPAJlMAlf2wLiuYscxycAJk0Ibz4dsJekErbBiP2I9YA
nAHQe+uULYe3gi7MZen0/MHMH+ZxdUpyhEx7UNsT4yAE6/4ZDr7zVH8nMYO4KcJDM+Uakw9kmN0u
uZ3dkk/N7BaAUYCL24ar+apv3ovjDTw5e6mD24GQcqsta7TRUdPO6vz9PV6rcRMkkiTPw9Kefk/o
k6GXse8EHCywQvG++YpjqNBT7VIInagpwcsYmmxErompi/tlU7v8wFtgAsxN8jq63cUKoD3meGc0
ju1oyKdTg4mOLQHKvnngi82TdwaYDxVRLC5y1lY1BuPs86DP/r31XvnJt3jB6houVlM8UOOaaKib
qIU6tXO/f8cZe+Nk4Xa3Dl3YC1YDa56lA1X5ZiZ3fbiqe9dIOkzvNay4m4YZwva3stv+N5YbHjJK
0ySfgpxHBbXfZcq6zH5slTzpd+IvDW+EL/+joRSRFcS7zrwJNf18hnTFQbpRG4eqo0ysXJNz4KBR
aWwVa+lrQB8x28H5A9IsooX0LWJKCruXfGh315+T2Pks9hj3uDBO7BMvtWSccK+eySzH3f0fmUia
ef8U8zJAHS5vmhvCinV/8xjK2+uQLYRw0LnXUJCGu8sq0pkRAaWnI4FARnG9bCdXPXQ0nAXsy7zc
KdefeKmcGRDFDpFf4bnmIrW0zjIHUYy8T537RhTWqm0DeBKIsJN6llhNJZ9wsOzh0nnnZIn0Q3iG
PIthqFxy5Yfm1Ej6yipnHR2zMJDgFkudmqUvfEIzOc4iV0Q1P/V4tJC5EEgvh+wBbMgTOSPBKUXy
4c924ASa/rUgTxSi+HMdStSjCl5zHqQsWTMZ/qAQdodTILji2eFEUg2dlvFKYUqr1vLpFjcW9bdN
Z6w1DBowlRngRnjBuj2/uHzzuFsck4UKoD2w721ba79fhq9fAV4X7UaWne7vV4J++2LGJodKfwbK
/EJ1hJA53lt5yS3sHcBLeMqD5n5HnlQOpD5bWaLg8PPiDLCU7fQqouMVf1Jvm4x6LxASX3+Nij6l
Rf9nDzv0gE+4ySkEOC4btOOVfkE3nAAcR6rxlkPsxqjLcx3ahbJoBg6Qfh2RCQQ6PNAKpGHshMwK
MafVx68ru8qtHej41IPwl7jQf1X5N2wbg0XgJWGnCAyaDU5VmSJmSXmkeh0YJYYrj/JbVaTcuCDq
nQove/dLap1SF0q+X5JJDff79wPSYUft1P4yrkBjQcdfcnlXidDy/R0rwhH5fqlwbzPh0GlCj397
eyQbLv/8dBLiD0kPH1yJ5cuxn1EYAAq8oimXu7iU2SGGd7n00WYsJ7Pkc3l9hqxNmo9EO05froiW
7Pw6b4i88Nug7fbcKG1xzskdKfCf0yLIfupNSWr5B38cnrT9jK6zDIJepNd5qj+XWvWq7mX5U24/
V2AryfZdKYNHGWvSItBz4B2fQVVyvkwxkh5QW35OBdZ2kB82ReZMMV8f0NSjE17oR9EQ3a3kA6X7
wSqgzM34rLRTiP1dd5rGFzFQ6FQNEAkYvdr56oIknSVODvtTfodoesEbpB1KsaRj31XumiLIMIcP
waZkXbX0YobYAZo69YlQov2rEO/k1IGjHgX8fhCzRwaBntTmAwc3InDg6GX+I+daFviIpFT7wY6U
lRQb3YP0GuVufTbKHvlxf7YoyoZSGPPcZyCbN5lL/VTNnLdAvQDWV9BojI2VCtDrvtDKHEEHPjYG
Lt8pw34VU/+fjdLCCtPwaEXH/ELm+L7cbL1+gHjsG1k8Lz7jEcgJPlYkfIVDZSrSS23XZZ3KcAIo
ttQs0ElM4d389NkA89le5fKK1+J55JIx6pTG29i57pWt0mvdVgCfot11i/hozvJKwFGyWSedu+vG
2pL5YxqldrYgTCMV9/0e431IN7KZ4ERntcBiyCwDcCSx0jxU/XLSNFDHZPcV3bpEAMjDrUmNg25q
pPFvY2NW0AYKnyWV24FMNcAwGoU5OsC4JLkAml+pBn3OgiRVwQu6yNbGVaEqsel8vrqLSAr7fDiI
wBxJMxni3CK2q05USZ1/TEQaU9WQWpNfXoxvVcDMVHZvuLXX89oCZZHz1w4SEK6ICFMQYrzM1nsk
ZimXO7xsFIyxgsgXSt4sfbmQR4B0GsFGcL5Wf6aHp2ma+1LJ6zV4GN7VGkZZHr1CfvdnESxGSzpI
nxlm4G8NVGeOl9+kjhEjLotKwUa5PcYn8V34xuZpo9UGpPSQUYXT3Ux5ohzU0Z5Vq9GV2frMqrHV
UrTcdvKX2v8ozap3L11WZNPqCfg8H+ho9xlIp3t3HBEGC1K8mQEu5gwJcioeVow8RoYoIegmacMf
IxyvCrvX/BpsA6HIpyiOAP/AApwYortPpptx3rFbmyFYh6Ynd43Mfw+UwCPKdVEaM+YqVqsfQUbA
brjmtEhTD1VZxS4+pnPrPy9Hd+zKwMRn4lMhFr6N5X2kHYBa4CLszqWW3Zm2NWi8G9HWunLSDQHE
5SHNF5HCocjALK2LoXb5pA7BzuCK6tH/Aw+ik6Jt9VeQgmh3mTNtkLkBFpYmBw56KhjJNnrFSBRY
duACqOWBDkSGuTopGsJm3SaPdwf8/e+Qgq9nV7/fTrNczuKjYYc0bn9vzCwsXilZcwqv8OwPXzP9
NxgNk/qSdd44lBIqY6mG8BRnmhwmcZP/RC+2jOGMUDWSo5y+jNL2CRCMZNRLfHAfUoiQvnxzOpCQ
rOSknnrh8wHNXvJMWyFfP46E9pw3PAOBFuAhw7q+dzc8l3CB9QJRxk3DLqSJqQ6jr9INinI3rkV9
PekbiBqkFSZUv2JhvIRd/IloFd08KvB+xLgY9cIpAbueNaYTMIl8vSF7epTEySfAzC7yB1dC01QI
SRAhsb6MWx5Y1+SCsIkveCVzPlMU6KttUM0pJX7DTJ9wW2TmROvunALCqPuPOwlUx71h/xVFIUaG
2zsdDlk0k8ZDDcbqaX1xHP5WbdyXSX8DaWXrpDSAgbIkLHxM38oiJRgOUlrizIEr+lcOcaBQzf3y
7Tp/BRDKATDI+jFJLWqHfwKawoM8lDMssMERfZNO20vprSZpOuu6HCM7tCVX/wFV3ODUY3VtGsNW
pzbcUho7DhLi0pEqUsv7AF1da2MthaAPT/JcJn6Gi6WAYfRiIPc+Xx7dWk/gbV/qr3iTs+zgx0rd
hy3Grme2e3UBr97iQ6Fgoz7kKXVJxVQJ9DYN+iZPcOjzj/dvi3RjFqZrhtgImc1sL/WilwkU8Trv
7XU3nmOK9YhvjOAOxZTzVidvrkiL/JRdUradF9V4urL9tMa3vOGGEG7x6E9H8cCWLhMWLCpZFHME
n5Yskv6pPWorjnplVZ8y5v7jCu+eWcSAWOdPvj8Jb+ev+nwGewp5hB36zE1XH7Rmd35+MA24eqhl
eXGwc/eZEDAes3NTnWJtz9jPMth0H4bp1rWB+mHe8pYLT6BYwCwCPVOIM3FFe2SjogTcifMvmGlt
vkfjfSsoMdvxM2/Cxq6/a/dzEjSVcj4/4Mv4Vlg8lEQqLFS8hNoPr7GJg9jnUAaWfC5QYs2WW42u
CbsMQBhU/ATREWFaLuE5l8/L7XURIVyzLb4ThNRJ1TVpUpHEPNQsrLARaE7cNwt/7F+vkVXElLq+
WDCMclbH9R58GCMxYyxwg8r7WsKcQeBsY/hTrGwpEVnz6VMjB97DDWqX1cVdqc6TpXV6LNhdoK5G
+N2nWsfWN7XAHIOAEyajkjCL170KFIgBFlVTHt9qtzAGcv3pCeQleDy+N4W2i7Jo4l2PKR3Hew1j
5LFttSHh0hcs99Wc0LyiMvg0Ssu6FmPSUawN9GmMnY1dXr/BUnm4zrHh1jeRDDKwWxof47n0FSCl
45uMnJtZBFN2yXiY0jmfz6h9XAYsmMoc2szw9g4AfJTsu1iQCeMmlTrm41RRFSP+r+KvWRHcN4ir
MWyqB2oEcRRSUvtLkyrw/1GJim+m3veYj+eUSvQUmI8+G0wSjyQVpzG1bVWjSIyVdZER20kgO5yi
oqQIuBvUUqel544yBIkiCII4NDWtyndLTwhgCjObvLC75IpWEgYhEze2u6fxbo5EgYZa+W6E/Byb
OLcFhGNZrE40FmMJZz27yHPvNfPubrp527IVML1r4OK+jfTG39wCIuzDEcrHsWGzPQl+fQXGLw1p
WhWJivSHc3soufK92e5RUM4MKWK6FOrr6tRRr4Azxe3nmJQ0ojOc/D79z+ZXIb1Wc0uRdlIhwwIg
OsqXXBfFOBwHOUmeT8HocKy/osntdTobornHJVyc/WfXTsUAFtZeFjIwVExkOD4SsvxFqkpyflA0
2jkhA4ipvLzqNEEp+VKNdjRVXZzvqth5A2jIqcBZX1MP+FPxycFVQxpNfPu0penNMsyUYoqu/6mT
MRSqrmq7jO1vjjfJMlDUQCQuaekQxAXxgEndEodyBPovCG+ceYcz6b7p9nhhMYGTxb8PniuhYhfY
Hia9p/lUB7hFvyZsHXujOGat2x+QSlMCtCGhvsCJnMrJC4LFaJQxSGmMziAa5n56xsXPnjhZJlg6
N/ftq7+eWE5rOGuWAq13jGdei6iaMHrProvUDYM+P8vbz72kph8RC0sxY+FdgB4aW/EOPX12J0nJ
yI07+f+BSxRdIoCozvUFFabulrUk84jjQUmAnj7BnF9xZF7FOZNJrfrtRZ8m28h+/eUslxBmSQFI
IuoI6H81JlOdl3P5OckE0sj9f6bAtD6JD5FRXutICfY2Na4dG7Vd+obi0k7MlnsbrFppzJcqMSNp
j1n5FFpfYr2nbzESud6BwLKI6BGEx+vQUVDXwF2FPW7SJxYPcx5o5Htl3t9IbzR48lZ+Hfy49F5a
5dlzYI9RVCCAWYYr56hii/ETJQB9yo8+WSbresRRa8m6DzXtSCWXFt44t69otyzyMAINaikKY0rl
ZqkLPDhK78BRjOK/ocWGPYtwN+pX5lfrUNz5WzGIYMjq7eok8l4mEZTINRRO17TygWyuMqldH2Eb
qWnTt4wRJE/NK16IOfM44TmO9jnCrgDr+HZWB3jeR6MeMJnCrvdknU9f5qmhSGZfzlodpEJjNMIO
mIltQL8Zkn09es2Fzd0QS/Bgd0Os7zjiApP9XreBDdZsFK7iNKS0GTpZAOxwcQDJ2f1PY9HGg4RO
aUTIsf95heHcP72pSwrQAJRHDNTwmfm6geXVw/wXb/QDhJBzRDVoI4JvUpXx6Xo7GGIAQ7IvVLtQ
ahIPZmInJeZQAVKZ3rEczQbPg15/2h8QR7lFQig7R8HEm1TO4+lIURw53rBVEmZKezVRfkO+WYit
eKc5aOmQ4lD0aoMxRJHCBiimpR219fqWfIApfikDgVc3gSRWdoIdDVZzO/6d26ph1FcY5Qatjxbe
URMubmLQ3GAGsNYnD4lurjPPPCs8pSywBZKK2f+BkEC0qWPvvtDdLUc+vUP/QFxa+20anYKHJJZq
hiioOhSBbe0X+ebpAeYTgng3a+N9Lrl9Rqgm2rrDBZ+MeAh4i6s5A1x+AIB3xojRQVPPJMbykZpX
gBRV1BT+fwj2Xy0hrWlbrnpOZVXzcxaFIYQghObq1OFFMn0Zmfcj5Vz1t5+v+tMxFc9Mv592visG
0DuqJ65Zdy7mSIAnfbMT+DrKtz0mxt9zbY5jYU2Qaj8s/qkMX3VXA4GDk9OmIyF3lDrgxPPSk4og
sv3DVAurQsBL+8oI2h8NaPp+d1va8CE4vJ6zSQxOQ5r73HwL9MGyBpc7TYXFgeRvLJeoYq7N5cx1
PramiIcnu/q0zQ1h62rdcYqkChX37Hf+4Gg3ozcJTxWPOXREyVGyH+JpDwJWnoueqJ1wcgG7vOmP
i7Qcz9V44hZARN8FRhrp4NdYSRJU5vPQ7eoLxYxfuTsCzt+femdV6u4VPOAzwpixOov2JrVGFm7S
uSStqCzNa1eyfmU/84jGbDBLroTj3HApmBO4BD8DQzox1go9fCIRZojadcLtyu4LP2oXFlLe3YGk
3+PFN+ZVTJSz3AxbFo9I8sg2kgGobOtt9YFmxdudI2WwaD3YXzbCaRwv0JTsVhF2xOdGU4CGQMoq
MaJRwjxEselN0egpsrq3R5x9/q9Mh7WVnfHoPzuusk9ReL611183bD6W1wApEZ+GeQTqlMFN8SzB
hGj746iVfq/gPGmtazsOlBwgop5xwxTxeIeyF2UlDN2bc2ORLfHa2+7gAmWeNRYtW6Y2kqW533mT
DQapyIW8q5+X+tsOytiQwSZ2gROghSwMm9qejPh4OLhcM4d34mwtKnEJBSLNSqXEVTCdarj8k8+N
23vssID/L+Kv4fiI+Nwme3K0jomV9T0vUiznySxzF7+7dry9/s5N4jckUCu9L9PeROKCUpQ8mkKk
bR3MrAklCC8oAqsgG3fBNbbBywcCiUPjFYQOUpmgVoENgWsaAU90V1bkeni1XVnptylWg4NIp+eu
2jgHD3f3mw3c8b9XT+mdKeIHcXkd+gIAu4fLV2ZnJjDeSU0ImzUEKCGB5StjEtM/1RXN+IuCEQR5
DEK3hYPQLzJhuw6rmYAggZhdIxC7b5ZJkeB0WwGUfMrrIGM10U0wizbQ2FHse282k6z724YXAnoy
djgJTvR46TSSgM+6oG8Y5rfM5lOwBn7Bm/vTldtvzB4IyjNHVdTv0PZwpZYpT5RTTMJ/cgHvSbvP
vJOcEenCkkoIhf25Sj7ahooebgX6delILaVxt0DiHkLxvvfsVKBNHSl0twnbaRaPhXcpd0fQ0V1j
7ej1rXDjnaoDVQ+ZSQ3EYZY+CSg8fc7omRgRFCTPr0qA5mppHqwM1hZBEiOxO2WImy67D5lfM2GG
FjXmnZ6x+fo8TwBplACPykbnS8bK486aqvuQVbRaKRhPpOO0UyCHvTgZc4fILssb2ToZeXc/X01m
oXmlMUy9Z4NJ1dQe2KpkFzDpbHckJHz5ZtMFLCKrK0Fm5oDAxXbLyYooBKvkGEr7878G7I5YMTjp
ALTMNhrxV53MqKK/ZXbvLfONjrTqz53UkL8QVSRAKyMmPnxeE3JeulF+q8W75DFdtlQlkluZEMJn
YuGKCtbfshpY3s8sUANnhnAGd7xrEzb8n7m8jf5XiZzogXGAo8gJRreQ3ePhOI16Fea+VIRzUK7i
6sD2WpUeqUzG4kQi7ODkqmpe2tFcCNOu9fVLpleV+YSQ+EEdmDPbKnAX/sFh89MtfLs6mLVZEPXc
4vL3MSHUATYcwv8yakZ5FW+adCLu8GjmK2iHyBdfMkNhXFOKoORfZvQGdka3Ck48sLKV5aiIabDy
Xhg4ymgILPmkEalHKKNdOLXmZZAvoiLg29wzUh4IHRES3770CN4Rl63nBPhJ49hC3Hc3TiMS+2KD
M0Fr05vD8yKkwLjitAWbajLJSevHv/vlz/ccgI9Dd9a+HEOigP0ddbVEQfjxP2bQAqbSLKK06Ia+
M7viC1I7ceS3WTMi9Mlh0yFf0DiTdONhpn1xBaqzjBOGHCz3l3Tw/BqJ27j8qh0Ef/Evvr9cNlGZ
MGtXO2bA6fDjU4gz21E6dgn/LhfUWBGNVEAmKnpJ4fiVTHZ9IuPys2i7pj0r+SP5/Yny3W7prEeo
fm5nxBnSeZKvGkdZQ73yLzGLhxIieASvEH45NDBoQX2RbCbcK/hhEVU0Y3KFdWWZCF4Rngw3CVFC
OvdmfzZz1ErGlJulBjb1MfjtMP9uyJXgU6v2smzusuTg5H1wWQxFR0+6OiSrVnLQIMm7PYkaIw3K
UjftrtcBoJgibPOpDphnfai1O6fajnffwAUxEc02NNon6ctDRm1HnbPl8I9I9XkCwqq87Oprkale
fsB6BKxWyffSZPAaV/Tk3I9zcQjrajW0FqOBruDRg9EKEo8VdKcAoyx5AcBgpDieMxffye3FcBVm
OBj+dR+Q4WSHfLMHCNIdmVUtIkWCfajCyKIeUEygssulf+nJQw9UYAC8knn5NBOj+F24nW/hMyXa
PPT/1jiHVmMkimy+t9i/nXSO6xjbw7E1YuFxkePnEvhZ+MmtzwtczeJy5blVhBWr18QLNFyY1pE7
XGiJcsiJDpS4zbma+fK0WLG+WVAtW1T6E0CblsaWqqKGYv/6nn/cY0y7a+604MGFrQINJ3U69eIr
peCVwkVBcedTOe97QCrjmhUV5U4yMjj+ph6/oTTuoldHnOOHOKGnXqkG6/kCwwwzOAn+k5Cv1rWj
c6vP9HqSCSBHT71EcppRj40te+oh13CJRPTKH3rrcxUfzvmGgQcDSem61dFDK/axKo8Ou2eYJnok
boLT/OVQ+vFaP/4AvZarcTeg1UWL07p2ifCIvvK151QHNEOfZzNa4FVQLawnPhoBpj4zvAt3jnmQ
tLfMC++1YwJ7wckyV/J6QbZXkM8cc5iFCuJmkTNba/x6Yx0Jpgc/22j4+XrX/RSwifc5uo/z4C/s
mXCjGA9QCV9DdL/cT9aiyGi+GRNxmPsnUYJVK9l2CFQriY0U8wMKrsx/4gPFdBMyO4oZ0nZhSWed
3gvTOk6XE7K2gaHlQTHnji0Byvo3TNkIsGa8qEzdwUyXdBQI/rUUf7Nw8YbGGTM1AWEFgDsn89GA
CM9QHV3H0ohvHjXO+00LqlLMJjSKwBTiJk9Kmn+ACVv45czTI8WK/2aIWcJQDJ7B/7+bErO9/D68
xc2+/vkZEaZQpbA6SRIBI416DjUeSGq7vuxYTn64EX4y4s/iHUYeJLZqaeJLjqV+PkV+EbSM10VS
QwGb33KH+9DIZFzrKsPvKY4BxASFnR9G2RybnHMS+g8/FQEPxncKZYHZa0Pr/340W/N349Di4+u8
leSVsywLhq0gXF4Y10R1tJjjN6ycb+s75ywR7ShxctmEzs3K2d2pdV5lZujDEruj+3Ttvu/+xvnr
bt/YSl3dbryOBSxr+4ghfOytYtHGdGdprRE1FAN6EbaYu4Vp6yMFbM25OrC6EJbgZiELRvonioWS
23ZF522cwDneTE4TB0l0DZWK7Kih8U7Ne6Rx4iN+TTPgJVULrMRj2sev3X6LAFOTaE3Ipz3o2WC7
4gKX+WIRYzCJLot75l7lmNrFpOC5y4GMIVazVi5mj9+E7Wqf8eapPKTnXLzwyG0KTRPYQrDV+Z6r
3q9rpNescdTZEDzC2HFCLHCWeeMRWGHiyTA9QWr8kNJvI9f4EGe9UygZqXHpf/ulQS0bQ+YiDW4W
uSGATbze193ETDiqUIVctaw49lO+IpXWKNbPWxXYMqvHSy2KFGhvPzMQDK4p/5Q8Pm8omND2Ie1l
lM4sgcpf7D5MPm6iVakhV6dSGvw7dgbA8QkmlsIbeTaf/D6pr3xrLUBMK/LyVzMZVokuJHr3DXOh
ZguwRu0YFCC8L+Sweq66YeQIl5It1UkmSA5M1rWNdnuD2k4FLNLpyyjoOm2xYbsDE3747fU9Tjde
eZw/MJgKLJuIpq/bnoao8CN5myTjjLwlS6ZJAooR61+E1HUF2mzt5w3RH+ioLUZjzwpKM1vekzw7
Zpk/8DFhbWouOEi6Qio0VCjgqIAVcIQfnnycdoLqpXa/bXQ8jjhgwrTv6Lj7TWLd7te/xIVH1yCQ
q1IubZNw5/csNCFrLmavpCQ9ng/Bsb4iZsYUfE8WuJ69NmnyZJszrQPJfIWLVneR/pGl61UvVwai
oogrEce+70LvHxcoZRpMy5bZ/gqmqvRBpBHPv/Cks6OxAVmz6IH/YduKPQH0JUW+jeobiKkWF6lC
w2f3nFQceARKhQ+Rfs9Clm0yxBBsgSKbR2FlpeJpitSKVzvyEXT8VCBKuT5FfImT4hJoFgmLGToM
MOs//2y+JDy2NTUag4TiTYrQpRU7YIWHnO5T38Ao8mOZ0SZu0RT98vTFFQMmEVkEMU5VatrXAng/
TfiRBFVz/npFUO4+v0j9OfXJiFQbAWAjw1XuJvT6SFoX436R9+W2INn0057nGlsKQpM0UYwI5hNf
7tGn0mWptd9pNSbZNWqJvvwNJraOXGbxQfvpZuUWD2P1lPDsKZwJUngItizAC+FOQHSpePBtDBlk
jv8n1hEA8/VPnhMjn9lad48KWuJIXai1SyIKSAtQCwrY9kZu9cZUYe0SPew1p0b86W7xlUKA0JR+
Fs5GTuP25A1XhLLiivS0+mvpwV4RXiOT3YLt6tEf5uwEjOPfzPyj7vKpcv410urURiRW4+ew6vOV
nJnbQ5z40UEMQiu+HT7+1RMTPesI+xYeDMGum69k/LS0MfvgkuxdeY7Q3bjcx3ZwAsjDm7zxG3VQ
wE/1Ef4BsxDiSHsk0EbQXGrLye7sgkWGfyGsVzfQOV78Q8jshMuOloXVlpvDR6Vi0XaQHb/38FZs
bVmgtdYtRkYbo3lcEdMIjtJIrrFUtDkNzCjoGntWAVUW50QAFEUYbQ89HeWCjNcXRq8tzkaO8T2t
vbOR97aQ0Yn9Mop/fwJN8XYbINegyXkvGRfL+FuNldyuxJu29r01oqVeV/kZy1HhL+NTlDVrVFye
cA5eGoZGeomipES1o0Ph9fxnGJWMiPIFZIeEMDWfGFJ3U/HtVbvnaLmkbmmjaoLrj6TONsJoVf+F
ySqlcuvyRrcFW7VmDYtAmuGeAOhj15z3VV6AYw1+jzbr9Sfsff8Xno4agNwpIcVAekjc1sF92xdN
a0zRCrfof4qjq968Ir30wmv0F48xhkKSKSt6iQyB5l1JZAB8ZN1RQ21ejW8Sfe4mth+JhIhnotvv
igDby0ibwd68jJOFQU1n6zHZik3qxSTXmblj8okzYIMCLxktwkM1A3pAuFDGBFnQ02RKRop1EbH3
kl3jzv9CO8u6xVb0HSGqrAEW5yTxhpjkR8zsibGJbFUKwjmglYaDNbpy9qMWG3WZAt/GfHqcEIAH
pmvkfMHkQjcNWxnspSNILA8qC2xM/lrd8DXT+UFKlXQydiZP+qQ1da+mwFbWyx0IyqtTQC0jsqs6
mX4WjZw/RX4T9+LqxJbklNbrk8Z4eKlLs/DC3GMF0oDqWSLSGZKmfSHk9XZkLPy5YhhMhDxY2fTZ
+vIVh7/RRZWa/op3WRW8tuV75LeE7L0bERJV5+msyx/jUU6CCkHoEdkd7t5jb9tB9MLhlmavhJk9
uelQ9uSnbhLpCX2uIEc22Frc3n1XG6ji9HSPw1EJA/1BWOq/tDCSEyh6kNy9O+kpAlS/rzBZkxrQ
BGFoopp5SUC8xfzm/D2D5UTE6yY9VGfS3Z1TOVy2GEVZZkDtmnsGyusc04aS+dq39Droh2ub4MT3
N8znALlVWfTpx5jpGkwn+eoP4+JZ1UqrprjtXAHIlfNvFA8341QlKBiCinX/JXixJz+F20jpoOKp
kt11U4LbN+Vx7hWMbX55hyiQUI7AVTzgqxlV3eM1CHK5j4E4CcodYygxcJx7iZmuhGiFmCbENf9y
gA0dizN39djZzvTTU+yz1u37WV5WJe2FP2Ogzum+bXvbut8cPSYoHL2hKxU67YXjYre28vE7VXjA
SSDidBP5ILwMGVPonT4Wh5XT1PMiQtMB55JVdyojaBHcBcNDdG2/4QU3BKo0M3NlUVt5/hRN/nk+
io4yZrB5kttFBlzQhUdDMzpmrgVzNP1xPfurZngLBtU/GdXVWpIbdaWjkE7+zx/M4Dzywfx8mk4z
3ZeExciFGArAbbEbBqUHKnLs36sSdwAOLGePRbFrV9vMOexLzTWV/oS2H8Kf96NOC8CWCe49nQuE
XFLuGkFdTvA7usgXn4pBUadGLVeuQBfQHcBixZdWI5FDz5+LHlEJR6/u2+D3lZMZD2e8WzFRlPz2
Njy50OxvrPRqk2vkmXMWvPs1zbv8b6K/N57oupj3uEGxaXIWd1k33atPA71jkMvmWOe83Blot8Nj
3GDLsYsj3nikZnfAP9KIKeqUKycNEcvlIqCodJuTaaeYZikrPPpgPkZ2SBHMbC1CupqWvrZhYIzX
34y7xxBFK32yXfql5Tmmpe5NkM3ZiL/ZUGufmpt9WS5nHfeUxpKb36bE89/ZCazVwuWmyv47vGn9
kH+e2voU/vq+6zCfNrz+NIEjHvTJXD8gXYx/r2fzvOBsGvtG+YX98C5znhZvnGyhTRKXorLWX8AY
sxtpe4shJGLy+Q9aalFXXHMqo90UC4oreFdkUY60mYxg+OeyjGO/P/e1kO/wS8xjbqy1dHsXbSb/
kVM4kwpG/Vqseq4zXpM/jPyklPdFKCr3e3tA6xBoAiN4fhGjnVgDQFHPC4byYOC2msKQ8ZqeMC+0
NecJIzMDt1pDQngorWeW7RV3dyktPuyWz8Z7XMqX5sCgMJEh3sEClQGd6Sl1OMGu7/y19h6cwBUz
oBSf8Z/FndoRg7nWVOIC2N5RHtIYUkZBsS2X9swMRq29MpZn9AudRpHID2Y1rm8MyGx3gWBefijB
bXR0wIlT5kFtUVB/6Tqj4ImPW+XJ3f3Qu1W6MMfumP8J/yfF0PjXjk+gGCQ4SWviM+Hm8yXZ0gDn
YwO6BETCQg5d3XHB9RDi4ib7O/nKBKAt5haMlQxkoHlrYesbhPR2M7udDKtzB4Qk81lxpPxo/iMm
026XqfpbLvF80I7VZV76zw9c0DqBKWDUtpdm5y3kwboyXVFkzcHBxPKTNwuAauxrbF8gMyC12N81
0pG069S/yLQHSSwwtxTq4yOrSVZ//DK7hRCNkyYipRD1QHReQp8gE6uOxqbozTKcKce6YN9U6Ink
gbthu7w+jeGqX2WNmBOcNRbopsjExkficI/Xu4eeyzWTe9eEKE/Fx0JIwip4YKg5HIDOCLHMjyYM
PCTxfudVwrIRA3sPNXFQXfx8FjfIdCeAjSpmD8NNSqnF7JNxQvmBxrUIxA4kvIV9N84S3G4a1lsv
kuTYBLZgI0fuH61/TsJmYPzyVqIAf7g1E6slTO52vCInugFG/Cy3p8gaSlSP+FLe5XbjOlrvXTK/
Ag0qiopOA6/IKNwx1A8LxojTPkcFVCbTarmyaV7TyqMne9nY9Hkz4Vwb0Dv/o5Qz+yNjPbylIvA1
YIziIpvx9/mx+w0cCn/JtgXTO8uLlcgrNh5eodX459p+2bjAAmtFgGH93LYnNoh+dA4uuIamH7kf
1GqjTi4bIvrMWB2ClFCwDToSEyY520wZGqoY77FWnwvCzovNVRg9OybWJstXyoUmN17AKDz7YER8
l0faJyIFaXa/EhmVll6eCa6LNjPioDnBzD0qw8dl1Dy9WJrapxFYFvRkOmiJfZgncPluBr4aytsV
PVVBPkv+lhRLAV/hYITy5vJ4g1TlXUGOFIlPBi6YbqNvkbzZvTrMb5H5d1xO/Wqn9BtHMip9sCJX
oLvCV/Ml64fwnaLH6jXrtAFSfX6Mmw90zZPiaqyj/DQy9IEM5x6GTlkfHliDq5W5nIJqV3s/lVZy
Hw4mt2VhzZBX4M6TcDRRz4MCdn3q4LgwMlqL4o4U/UYOMrxTCDU+PSZ1BqJQc7NdTJeLo/b/GEpR
WYSNDlxedWqAj3z/8pBe8jUvmf5knB/Xi9XDEvsUcKiDVp5yEFYIhYLmOhG92ntn+fLH4+I3U07b
eqZ5IobSe2UNIpC7rFpwfvkN/CLUaf4AX3G/dUmQadPP5OSbjrQ/w2f0G80lb2Sq3L66ysxWuhA7
JqE/qzs990UMMDbkcadSnYCVF+bkWiWA/mbbdjspUlAhG/tZ1EkdH2zu/Nz4XBIlCT4FRb73ZDCn
8m4GNl/DisrcuVTGciikp4YSK+4vocV7qGCjjYbyCGBJZQ9R+CyUp6MPdAWOCsGNFADm36nF9T3v
YH330J2fLRx7XLkWuLO3+GW6XIUhRu7bAfNGoRNrj498z8yZNKPmTBA9Hc/VTG9KBL7GjIv73jXL
v/pK8On5hgzUrK6qFvaY0LU6Djws4VrkJXXo/eGTK3HA25iXa6BxMkqiP6mXlZmoTSp6tYvajRaW
xdIPR82AYz/Q7DWjFog5RX1U48xzlgczN80KDJZcF6FZ9NKxG0q+cM2zVpPLcfyutbF1qZYLvRrb
moc2hTv92GKOsCvGRldVuN8iazN1RjUv0MfW5NtMre88Iu/G6bCo7j/pbQuixHM79YRcrCFkRGwQ
H5QSec8FP7+lwoBCzEs+1k5JfANtbkJxK2wOm3xtYXQur9MUVhdnmc7X5hx3R3OLUygFuJ6Wosmo
cEq0il46UZSk2WQpLb3J7d6Z70+lGsSZbltBJ3GyduJPfuDilNn3iLdO4uEI7bowvvy37Hnv42a5
xSVB7+leusrgp8hR3zO23lJ5/FLWPuv2/Dg8LH5soqdR9GL9t508PoQ/M52mU/CcZAo+v3s8iAsf
6T67KUzQRAXwicLZcsh4Iw7avWcpE6wFZ4atjg+MhpORcqKx/2SnzyE/1Nfleg1R/eysz+QY4gTk
Yab5j8HTlhTWs8t3qRES3a/FJJE/Rgd7NkT4kwZ49+Mq3eikAFja1it8aBU1QYfB7wIHttQWnZcD
W6H1A5ec4pehbFnTheKKQ4MSVkO24SusaNNJW2EGzsrB/dXjlXDOUq1Pc8ZvRVw79A5VqMm6XDIZ
kA/XfUPwoWbnvu+j8xHesbTlydOUdGGy5oqLAuxtPCY1m7eeLFXh6McpGH+p9KM0dvxx/2Ue4d9h
Oo9wKCtcASiSG4794scmuh3dRkWvWISVgHCGlJqZFkva1VZiiD/Ba/NprFke0MCPYxrZ8lK42NWi
10XEBe4jeqeaF7GPvlpEYO+DQZMjeJj+PMd3Gp9DzcRJY9n9zJUoDgIGUTvx6QT1PQX7iA+E1dbC
0rAR1AP5WoVyFJGBHBy2jLuEiqXIg/HyTS3KvtMY55PtHtYRlSSI20phFd9EJI0gxyxkTk57Mbxc
46lLIF4cFVl5eJKlE65LUpFASTckJpp4nWJJvlROrZFk9/bVI3jcQjShZBakeMmUxsww877+Ljch
jE29fRqII0rddkPxDYLsCVEdxIHrOzxCCuC5TF0KkfZE4Zx5szVHf8jRIgYdiQki8kEf6E+2G99j
Gsy+Dv4gADsz2RqcA5BZlck+FHtdu6ma/uwkgGqr9b63RBJd/oWmnx/sK8P4mUMldE6LKTZWxZJu
poqWKgHdDS6pC7LrqhV8irOs2BZw6qiiX71d5cA3XaWWJOhfg0Szyk3cOZE7A6liU2hfqmgrCN7h
FFeZin5XObkPfYaoVwYBVyZQA/DN7EOk+7rjqQRJmjHeAis5lmCZPZUoa83sQ7tfezScihYR32ZY
9xZDKd0HwS49HQshiorRLWM8HF773sRXGoZGrjjWLROlwyJeoy7moEY/STOedoeEnmQXzd6qsI6m
dal3bMU9CVtyWNUwAz5AqSpM5/k6nyF8gGCDgoXxXo6ue2hfJ+6TMF+/5aEmIWq1v47LELR7VUHo
NKuwTh9WR6vKDHooksxG3uayrWtRZ4iGqmfHBiusjL9jJQ9LccZTbYMGW+v3FuBl9QyifwKqLCbN
w+rWQHGnDJIv7rsoqSgyeqXxZWnpc0nuAhlzvwD9yjAxcHQikD1JyMD+oMacHact/V7cPZxTa13y
vNzp16EEKf1/7jlsuV/bWyUpPgqOLcsGK6rgR8LCXm2D5zQanN7hD5YZdrlWW3ZETAVs0dQyYlCK
qIeSenDYaPux7b98Vkm5+NG5wNITBP/42BrodYINgzh1uGPRd9zA9hSht1z388XXmS0IxTKl+LZ5
oht9GA5yh+VgvI+Z9ClKAjIw550ycPIklC203QNylb9Y7xrgyJ93/pAD2ELMWIaXsKe6OGVGqFWw
1SA5PjVogyuCZ/UWsECPpKtaJXfmC7bMlCdVoWGfkgy9JRUs4EZobKmw9s2sUaXxWuVGF5SnfsUC
OIyUEJdtMyKKyK+obKuAMAEwIxGY/HwV5Xi7m0GbQhJZJJxvs2WXf9x9NtN/dpdvEgbDbY7mKCfS
W/EhnRmAmVrdAAKBtCi0wLlHEj1qeU/PCqQ7nVz1pc9uq+aFhd6pxlTP19u8eeJZbX1q9ugZ+/bX
aCJejgMNcdQY2rQcGr4U96YKN2z3CjdhmlHNKckI4h+rC/d5IxfwrMNuMKT9Yqj0y25Q1bneRAhT
ZahUnmCN6XKznDT8KdudZJnODAW73YFHla/cTlNeymanI9O4x/Yeo+6LYDY7PgTfz/mjrx/0gk+6
MFDpebUBl9CTvxDqjslWQzGk9rIIHvG0jjk9VQLSfOCmRwM0wuauNYlpZCJIjw62JMisWpjC6Q89
EHSZ1Gi5LUa4lU2zAlpZicXG8plC2iP6NB4cEfqjMj2VrafboYnOt5je1YZsjhe6o9f5j+mtzGSa
tzPpk2guyYWlYJBTE7h/IHbDynXWXpLekcxDhlTw+E9M/OQsy2+L6zgqFJEXiUaIE1l/poVCxzFM
y91c6DS4kwH7sgbOC/+AhzsF9STkupuq2qkTEvaGvH+bYSzNGVGc7rw6t46FgwsOuOYsTrc8oOKq
Tbr0E1ELzieLRZ3xDF6rK2y2YNeaIOsXys9dyYND/0ifIJFukYcb/rUoqy82X4m9IeE2IdZ64Nfh
pi2UhbLSejDnje+tZUzx/9mwU/Frk3J/hJ+G5GQ93Z6FDbga5NkUqrlQrSxv7BZVezklInTWzPWB
TJxSEhzbFT02okEvU3x0IStD+5pru0LWy48yysq/zIS1W2T7VFuNxaH5XxWG8yGUxrXzJHFxFV+s
mO7SbCuMC9Cw4cqeHNP7kOyknYVOV/zSjS5tWs8nBp32ptdVATMOoKgSBPimTqeEcP3SaY4euTbT
fDHp6OZQMH3H+0iVMni6q5EMH/yMVtur328xHMGEwGD8vSekSxKczhkfUkaonnaiUhiB7SeD3BLl
oLPbWuIfRBLjge2l8/xOQl2jEumCVlFPkwmVhW0FTr5P0VEbsjWbrg3DL/cRoViKLolW1ET2+nQ+
fqD/tUzDF9dCDCg2LyBNePQo6fHZKmFo4zx6fB/2LKy7RDwLj/IOrxicr36UC3lv1IcXjYKgDT3K
+h9qgZ/PpR7mdY1jvmkq7dWx07AIrR0LUF3ytRsgxRZC9iGTglezWeBM2FEPJrot7vd48vnwvuuj
FFRtb/tb/y9V0VmdZCgbklSNuh8FobgJHThipWPpw4FXdcrHNaDkFttlULZ2CVXI3D+6EfiMKfrP
JnPEWnktzNvdC0luZtiifcGx58harlzxvG9QNI2ScFV45Rfef/ojXSzKxJ7EylwzCYh1R9xZU3aJ
BKsJoWdeZx1QxI34Jtk6URvMGxD8YKzxjs9upolw3Dn0uUhpxfptbSwZtbBfpmHSClDyJyz5vzl4
w4La+FjfAd4L91eCCkNAoHVk84ogDx9rCL4xvVxDAP9APHXWZSJwk2yCJZGALVJ3eTi4JbR5aEjf
NWZVmjE9yzL7rVBTc/HY61t1rYTR2rez4T7RVog2ILKxpHzCa19lwDY9boKI5R7HpkVm0P2pzd8S
w2wbZ8im0QpbFe/lqrjvuhOqo8RzKq45uKB5Z6DI4ehnVFiLwAnQlU8aMGgyOJV2yErxswjmp38Y
3HV3J4qcHhJYv08T/0Npd47bjVlbagLwxdPMd3kAXp0saI5a1gbyDyJzP++ImKw4o4rVXk1Ml1ZR
HeKpfDG1Fo8Sklz1KhjbmPzmAZmWYirjQtYUV3jRmfuuaRPrAIi9joifP/quVtLfB7ZXxdF6B14h
RkS117rp9kBEdW7BF+cN+W0TL7kIkM+ApH1JeMQf6GtxFE/mvCzwBmfP9bSOXRph/DZijvRuPij1
H38NJAL9eef3L2XnUsBgGz+tVf7/K2rC4u4Wd/+b2j4wT1lIZcQxYlR2QYgquxQW/TbToLrKKWg6
F3cWistf3ZiCXiCrkYnIfYzLV2hkgOUA+46bhWWQoW1ElAxG2rSwYH0fVaoxLJ7WYu1v8hPgO2mo
NjlIdwVfhJutPwTjdNOe92vEhAJZ8qzHsdNPfCgm6hc2vAqbKiw3NQ+sGGn0pvw5UjYfpFNOv/VJ
y+pXuoG3LY4kV2X0Yq75WUR6yCtti7E0OIQ9PYGX0Ajwi9eQPITh4SjMvEQgtFkhntMsC4BMLsbQ
mxdqZm+xpBrkPo9wf4kpt0vSNY0rW70Y9+1ANG9XWACGMYt03NnL2YrIon5lQZc63L9M+Po7wX0R
KQoiIVEysqXG/xIpLRyqtKq1G82bZyy4EMOIhr514VemTy1gV/uhqoMv3KfZrjjbQcGtpIgh0LLo
otbv2xwapaz5DbhocHYYoZUwgUNYVujEPlf0MvLPNZbSrUci9czraguuXXyiYN6jMcAQXQ/0qdwH
Nh+l4/eP8gnKTt/aBUcId04prJy0h72b9jnxHJ+BT/zoFEYE1xW6Jkx5ItJ9UrOtGHBqsi88WTzv
FhXEInxYocFy6GQ+zBnNrYkh3RIvZTWCjUcYIir+7YiP847l3Dnz0ZtyIcGghQx8OEsbXNfj4Nwe
/B44RMLWtdWVWFmi9jcng/POQNpLsCcaDr47BsbDb1Qkb5fItwX4AB4t+5tmaVWWDp9Pkq9WkXdC
XXPbwapItCSzczjkLSgieAymM8DmWTjuVIIF0JqHdBUb2RnYj8qCTd0c8ne0l6jSS8uOFnqRfxtg
7H0JRFNeWF8COxRvIh40yuz1V2ITz57lbfC0ZeifnEbTMQHXqMiU07HQ+Uev6fG2sgEy8nVtsJzS
IrJsKQ5dFYPIeENIGdF5ymXhb/1p/i45Z7mxqDVgnOHm5VXo4HE2kixf0KDLw5NAP7a6r0CFUais
u/TSOqrbgAsNO5ddHp/PLVQBcjoZvnTBglJgLYHFpqAENS4pZ9R4kQGEX647zQIw3YCMEQHaQ1ND
rzBTKOJ5nDDUAgSv80IAnaKhQeog7Z7BCDvIypIzdFmMQsMUKLOqets5pjTsjz37VezsFpLl1NYq
M/Fl49MAwY7BqKyYdSHNio6F0QiHhGAz0JImj5JIPWqJ5ki85JDQ8gPTPZb7uWLbwpk8EodGsqrf
e6tYCG1aWp4ozBW8ypS5gFjIMkvq5W9uFmYDU6Zfr1Kxg+A4hIw4MVzmRR+bF9hXmWhAWulDpAk2
K6E+/GhdofQdY6OzKfBpSpLACMKe/Obw64bwCLBlsX7d88h7HDXCGml4NKz9IZob+2o5JIdahj8+
5dhnWNBvcdvjXFbbf80+epf7d66NJnEEtQBwJQ78Oveau8tjOerms5L7t8m3d3yf6X/oEYN5zeOy
aPoAHbeayRYtzunSEaGqhg1wlUZZjdtZvUjf1SCpqDAPudCLohE7x62t/aks+KR7rA3lgygZAM4E
/+j4ADf6HDb0nvKMMMBO/hwRRgdm929T+l1FWRl8ijuX6IVy25vrYhS9vGXSakFKtzvygBi20SZX
zAcw5FlH7FrLzx1OA17r64Opk0gGMVateqTomxhNR4HNoRtqsi4GcrnBl5ommVRFEky3S2qsSNyk
HI5ugxNRo/Yfc8ig4TgK/gmTRDjr5BEoEgDX0dn7QmA2XeJXDys9dOM6WuEymMXVpVA2YQ9YfsT3
r9Sglm5cr7ljhCYPknWt761cS0qd+zMm+UnoAwYNhqltgjGjeGfzmo9PgIK3Wx8XKn9v7ggtU8oP
PHvIRe2Dmo4NJXjD4jWrBNyZdGWSU2v95OI6roOMdogP0SvwifR6/keqjD79u185NvfXr4vIKlz9
Q+VFuxTB2moSpTwShW5+e5MwjUpXQ+ijsNNexHz3xipMhiM/81mFgnaBbKWBlRLgAvOzsWLAXHbw
LyS3NM87KF73xvExdlNz8yxAPEiVK0i/9846m3VPWgbvE9FMat3dK8yRXKGf7KxvRN1Sw8Lvd8uf
cBg8vutKzPy4UPQPxxP116wfDuoCOVDAXGLMlcYkGfSDGeEMu7sAB1M6PA3bhS7euUnQBrgJ7t5e
4DZ+ijpbeLddMW6wYNpBZB4B7qVzfsDp2ePb5oZ/GQeQIEhLGc3jOMVFq/wqhusWm7D59ks5OWd3
Weu3wRDYpH63XYfODFus6PNSeaf59ybgvamMP0pU3mfedvRo8cOhp9GTvFSosWouTG8qJysQzSGH
LGTQvLHLSxCwsw5WMrVjfw2PvEKxuM9OZXOwX9wFatILef2BwXM+MxrSlQQtVonxoF6JrGBpT++d
wA+DyluDuA0IR/JxuY3dxnqNcbxLdWyOenQJBxVG/PxZC97hixlV5z90ciWOFCLe8XtNwViJpRog
q/CSEKUkTdn7f5uRT4gp0EkSEYvDscXMZnTnRZ6qNHh6LZPHNKZx9KDqO49ao1dPErQ8AoljkxwE
bUgIDxvVwS9SOIiI0HpPR8OJ0zDmtxgSrujZo4+75BiIE+EwG5lEkiOBBx1G20HMBo4qcQmF2fRr
7d18LHmxkQxLyuG9WqroCw1hnmm0C9+EkI10yH+yiLxiIRqZ2pKUnCPGFpgmbGcTfVEwi42nX49Y
g3mGl/odjW/2XjOqoCzZn4/H5t7ZegMWOWinGsO07imdoXPoOMa53thWLTAusqAJAgR9K3ebh74g
Fyez+/VYqdHR0FiWY4PMfNg9IDNVDdbOJLOnboEW5aX8Eff/p2l7Nm76T3HKHVDhuqodgl0smSKC
mP6S138MMYe/OJttnYw2+kNaYp43de8hogijfZc0ITFH/ekxVNMEQr8hHtu7oyOuaT9Mq5Xz5CmR
ieRPkWPV0+6nUU4KCmD2EoSFTtT+ZhgJnHz2XqkxMKAvSwCuutW5YL79xYKT54ww8q9VVR60Xkop
aZAwVoVqhNczrQ8EPHZCR7yaHUV45l6SffI/c4dkrQwY9zE9fVSg8uU82IrkEmklGgbHkAyyV6A1
4TNZZ8+ulO/95XvipwodanCCjUzBgYrGmRfpgLkdnfJDIB33ax6Hkkt/+xrwSKPfvxGCDb9SPyt1
M/TozGSv3knHShf38X+Pb01dQc06tOy+crlydK5qL1pOrKpO1+XMExuRZdSsX9go5Q18YxJYBvOy
m1XqyG1/9qY8GQH/P6NjoWS+XLwtqIjn0buqloWsm672I3u82jt0RkV00RUbr0WNzSBdjBD7IwqK
uY+V4OWV8LV7L+R7+JIIrpFCOg9uE51U4RyrHZRFcO5EIassUg9acsV6CdEBr9mMJqzxqw32GwwD
5VHjuOpWX6TRcExaPMmkVsZ8vrK9R0j2IEZ0tYtv+xD4NZiacZrXXKpN/8yWM/Upv9CBcJGmoB8h
e1dtD2MZ+jmJ4NruCI0/7JasAm1KKBEJbgekAQIMDGFdqi6CP33+pgRgbsKv2APfFVPeeyYGI+JJ
G1yNY9eT/ijSosqAT4nXv1d/yFxJ+7IrLVIPr5StWdHqtbGNhfLswu33It60qApBnCwczGjsB1S5
UmyecxzFPV7wp/njNsPLhkeopkEbHlMBQlOUaNYs2+hpvp6bTVMqR7OSnN6bVvyJIdZYa7BsHtLO
31X8CqpdYYekX75GvVO+neEep9jtU4B3HJFXv4OE/GgsK3rZS4owyKTLmpbRw/RnkOSuVt/9LQoX
VqdU5yJKP7bPVJLrBFDA4IpKYx5p7+rjU1WQeLcWBps8a2hKNxhco9GDmgAvL4BtVT2AowNNYUDt
ZofXSoEBc2wnRZ0r843IAi/rUrb52dP7CKvM24ZKG0PEAr31Ol14iyYzjzktdg7ntH7mDpkiq9ZI
1CPkxvCASexP7Ur5FgDnmQvJ+i6G5F671D+ts1QPBfP3IePbsEXDoCXgv9CEYcgang0H4c+GUOYR
zb4AmASwDvOMqEGliwOfpplq5yFk/9Auia74xxV5IdF1pdjdgBi42x4iEY3K4rfxhPuBlu1CVnrw
CFqZUBh9x2Ukb6zE6liWdjpILeDrWJuJ3IqHjRXcZCsL2xOJ7EgOfpYVXvcSqIY9Hyq5iH1Fm7TQ
40LeVnnuQgs9dBHWAoTnqyShEicedv4LYAeJWSEkyk+ElqdBrQrTYvCp7+unjbys0U+uzJI3PtDO
7QmFQJR7scJa922wg4gMSEOkoR0r31vFdB8i/43D9WtSS8SfkMXLYdhu3ZvEDUYxjmQQfCNfKZlP
T+YjSYmcMsP/Pl/LRvZxYm+HeMS4n7fOvLTeFlPMgNWiZ7vqcR7W32A02IN7dL75d6fluItUnmO1
46wAN6kmj+TPdoJQ4Z+QbMCrOLiUlHmBqqpqrO8SCJH2pyZI3rs0ldAV0sbn3H/fiamvdS2M1Izx
9wcWEfJu2nLR+Se7kVAs2xOGkt/53P7TTsnjCQa90ZLkol5sBRN0mj3ijylUh9o6xLd0T6ZmodNM
h6+16YVq6amN0se++rycrqR5cb2gfZhGDJSVxyNHk2CzqEcJJxqKjFd1zi0JUl/vKgHKtcGoblxa
Uf/Dj8w5jmUNsgd6haWWJTuFpoQW5ulKEHwDryx01PCdKjz+wn67UdV3AYa8NGrokl4ZCapTSeT6
06nhhlYoFU4V6Zj8Ee3DVwmuzOtjSE+pXe0loaKFU/PtFq4ovmDjg53MygRSAkHeJz7RFl3gMpXi
c3qMMduuwJybBctS7hhtcAVQZPBIB6SxLjc0nChuXqMjkRhmyhD9xpdrlQ874rZqmnXWADIwd9FZ
ifd4OYa0Ed4P47Yx+QvgnQtJl50OqHmYQ+aLvc/UK5efbNSw8dAClkgLqv3IcuPuq6I867gDYAA5
nayZPtJFmvy0etmTI8LVztN4Luc6r0byEM7bTCVl7khld68JaRF75A7xD4Rr8TXROrqOrC0CrTBb
1yfZRqA/WrN7mRTjln0L3f1tEkACILWVmpDYobJEZQ91oNyAjfKz6b/4buGbFM7bQUFrbDjPTeWF
9Xc2iACAocwrzF8acQ95pxr3Eu52hs6vYVYl5H6USTskuCRs+rCu8heMoXEoLWoYeCA0iME6IXjh
HDjEE0o9HLlcX6NVJigqUHT5TskWiFcjQt0UypSuCHwy+mVJbIOegRp1HF0h/gmKXYtAq0B1Xrmr
s55ilv0JcR4EPqvuUSd+2KBla96QypfoLRJGaJuCZ0mS3RDxN4t7Ks/QsYnKr5bOQ7Ky6kRofJVx
/18szmgJZUz0lxG2BmzlnAJAVc94koVJs4youc5G7gXGUOMbA5pMJAJ9PLfdHX0QI0M4suaOw3jY
zRznD3wWLs2sByme/N/2yeAdHOUtRSUSztDPywV7Hn3mwZROp94yxhU5s4otinFj5vh5zM8aYLgp
YkEJLKGp0QGfTyI/TwlIH2DzQ0T9TqzBgc0anQaah+3gfvws9Lsd6dJpMA17e/4oaNf8LkhNWhmK
XpboF/mYNuEe2GufZPQ7QUkafhlM7TwnDBEkmugD41YqZiOZiAOo4RkTP4veo+zSY+Btw1GB/BZe
gn5HFDfvZU1bobnIp7GsGT49zMEMK4Way66xcuVuKNQGf6IeO0Dp7iDfGf2fGd3raBlEAu1Fir88
vZ+WWbM7w4/9mPhLDKfv9kbSlj0h34b0eQ9zftQocmvLw/pXYpM7p3SuAw8zg0tcvE2WdQZ7PfgX
XSpJhgWKXnQxV4iVs2hrq+MEti6MZ1qgBdcpSVIz0clYGumll5qTWim6go5GGynpqryxH7+kkx5X
A0i/C2vPhl2oRE6oXNQtB3jGwBg9BuHTKOKBsUaZYV3HUcqQDAFeO7+nE9KyTFZDMc1Eywf0xqeB
hD5PT3SBGNMW1MhoRyI5oqLM4TCPk7tL+hV7+Sm8RCgjcTRt4EkCFKEmVop2TU1S++xsVl2PHVsa
y/HswHxqIOZrz827egDPuch4MEMXExpyiN/xZVXJWhlsiW3hiQ2Y+j+jgh2X0gfC5rZt+PeoxjbP
L1atVd8vSNB0pdgOK5O+Z/PimfofL7w/hD8LYlbILe5qWDaO3zUxAWogj4qvJhGC1EwbBLhCuJhj
5eseIAxXn/SCHEqbSpxHLxaXrdjmjO0ad3rSL0lbOryD+bDvg9D+iONSjN84tAEMp4sgiq2XiYFL
aQU3wQbNx9rGAoJ63I4nM4u/GAfUQXFcCv8VAnA3nWKSy+2fgtoc8EuYyg3HONMievW0mSYAL1J9
AgwYA3/XS+IEQM625qyioSoHDMXyp5Krac1RSfpJhYNR0E7Lg9JVOrK/oWLmYjVsZi8mV2xweO9R
qJP38HPqChma/EafI459wdfW07J3NZj5G7va0uJR67vqZ3fqwHdcY07F0i4UC+iCkN0Cpb5aKMRr
nb8UZyBEBR5TLwTPlwol5jsyDox3pjEzoQRjO/Em9ANUkXUWVVDsg+kEnzPwCANGo03lmroOELx0
rsFwadfjiz0RjnUuJs71vaZWWo0C04MnmiN8oPaRu3g59d9uZSm1fy2npf2oahUJslvdEOOT/QOe
n+v2ShuUYz3SCOp9YENSamuuDmFCvgqiTlXl5Pnk0gVCl8ywHlyLV2WHTS1J81RRV1zrJvSVoqL/
1bfSsDWGyRyP4k/DG957FgkkmrDwPFEEJBzl5aQMS+efkHd+xntwxoPI4aY8dpVk81BpZL6/vT11
5l1J7h+q8trhDEkm8gHwQLlrEvYpLazEt5IXBTfMiAk7AjRlWwOIshPkGz511uqKfksa2A3JHwbt
FOBAML3FIVMEpL3BDbm3CnUU/yA65l12tg6jMkN3MOaCNK0+MXLEvOV4kXrUqQEDnTxxhIUkZN/D
5on3B5Ejkn9WajsIWisKrmB7n3QzMBD+M2diEvU/uuEhLT9Sc4oHA72popYKOEhXNXaql4nrcO+1
HzTV8XrvDrRdrLs+Qk6TufCy2MgIgcW2ZYWQGcUv2nVjHSQwj+W02fvIoNALJF9UcsbxHMZqCP/A
bD0OjIsypJFRfCGQar67mwWOWKLKmXA+Z8HmSRZdzGKz506I3uYOO7zR/woOCRc8mm1ZUkOOC36S
EOU0VXl55+XLdw5yj7RdYpXFwZbHUk+GhswBG6unBUTrLbWGC2NtXTUhVx6oJe9XDBtVqJxc+ZE+
5T9DDIDQD7ANk96JbPYBw5yP3eRwYON2MUrzSvTMlZtH9nt9nsQXHfmSGo/cu6HAHsYdGG24geRG
GvN2IYCPehecoN+da/q9IjqjKbaSvGvqwBunz/VlGvlQ2WZrEYHEkOvFwhwJbheHxZ1eUukGXWFJ
Ztcae8Mmmv/QGl0ZH6tS5EaoDZVkc+LcsVuPLO8nCegBb+l65mUD76wnrD2/mbb+VzfagBA4CjNl
viumsrKBI8oNy18mxvbeOJfxMZOUva2WOchzKPObcPkC+a08n00RJNXg9D796OYeBabAFaB2C3pF
LszlAo9J6Yk1sqITfZOIfUfD2rCFOkmwtwNgyVzkbwTvyG7KLzhF8djCv4STAvireFOAittt46bc
nfJQIwGFbOFutWAnU0jswe+7aMN4Hq6lmDHO1KRXNIGz6QafDdLJqeod1bHP+rVd6F7r7gfUItEL
5uTp0YZdN5VfCCS5BFoXrxhySqlsEO6kB3W+WfHr3Mp/2lD9ZXe85oc6E0ZoDolgow/AfK4wRraH
C/P6jRrBE1WnunHjmYdHeceI0JkGQncRnjEWUghHf7kgKGWnZYVeB07AQOGEhq/NW/eCxbiKjQDw
4a5VzRg991AMNccYn6gzMGg4FseAQXylSm4iTSWORQEr6SNtnrOv0t+S5DyXDTfV3dIY8Ve+eZCv
vWDCN1vHS1H/syMcShnNZTPd2IsLtv/Y/B2Ihgfe2JVGGnJYle5CUQamU/K3fHL0BxX1VQcTny9s
NKms7ijB1CUY1cztpRMGWimu/1mvkmXXN56agNBelnjubUFcga7ZUOawgROOuMBsrrs/bfL5Cfiv
M9TOSkmXYBJTTWe6a8hBbtphIgcXb7PhiqH+1wRuQXSoXfoV2924iUUNh/BIFcREeZkRSgKHXhC8
w5wbb+j7XvwzFV+twuUTYpCYuTtcKGQdKHxIj+KphlcpGiyw0yTX4E/qJQGhXCgP9mBy8ZFGUmFH
aBu24xjXT+wSVJyP7qClHNHuj6pClxYRV/Qswm2vqWYCQe311IOmW/rhHkxgZQXx7q+PajqAGywr
7s/Fo48Qv6S9zJIV9bBgBleSLb6s7mbiSidgHnR2vCHxRUgrWXpoiI8l1lSaJq2CFS9YdBGMFCLO
scJ6RfotPStwzBLtslXeJSDHWTAEV+OvUrK82ugMIcNE7pjBfNu5oFjfOX3RpJE3xXS/x/de9X1C
nOHuovFLVd/smyP/HuKiGBZ1q51n4Xc1rTREa5Am4H/7xBeVXnp0pJtt9Saevj4bSyloKBkZwgPb
dQ2YIIS+ZSmno593EDhzuvxKQHdxad8Dl+PTlSO8DnFmWHDtEnWkWfQiPOV9bIQXaaq7sPX9wHlc
T6utD7Y7U7hillJVyPbr9naXMsYpM8dNiSovjiHPM5BIwPUBpcJVdKfpFuoAlj+o9dWy9cvacOW0
7hDJkg/6/cW2C6KoTQXTomscuNMtyy3SVA/Vzf0QwcqJNFgpPSzJGcvquJ0CTro7m4x+sK09uZzS
2YnE11cYG8H1I4Gx/6M+dswEYEL/zl7rU362jjtptMz/sEKTmWdKyQ604tCSiN1OGELawH8CEcFp
VzzEgwuYWBt+f9MatPCDTVxRbww55904CoM7l4z4q9xM7oU3WYz6dvS+xd81W5J+xECmfISq00S9
x1SV8qcc8FfJJ3COZ12U3hWB+KIZ7KC1j2yPnT0xTqi/XHrvH36uDpdEsw1nBHBqKaLB6QkV8sYu
knuGtzPWFPr65jEiz5RVhspeJRhZV6YbV9upSXUGe+wnUKlXYRjSwEPWFb6xj+PZJav6nnIZtE4R
0bxQ6fxnoS6CfKkp6MN5dpU4n17BMaKa6LTE4jfGETY4DMxcwfsiip4zf6VEOVOIC1bbJ4I5SBMp
I53uNhuGqZDMw0UYCrDGXfleR/Fx7ku8DbyCPTXG0ou1UEdPD0Z8BdNkCF+FdO9FakUyBaLESd5K
+91qNBdp9pV8APmc2/GvwKRJpuRKIC1gFGrQon6ZEuw5vZ0WAwipOsm0jOZydXu2kbwv5RGg5LXb
4FVbRbMREFO5paAVQMejsU2NssNEg+DpPPHWeXq3xj9UXk4pOor/rKZUYOJZNZn5RQoVFF97Vp6p
kj7v//iOuLRy7/aRqxEwwMLklk/L4bENxVqebZOYIvuldTQLgpJ7WYpBqAKbBebm5zaj6BZyEk82
cSuM+4zFgSFRcwyYMPNOeC8NmpfImczuigGvq2KJz4190EGVeIdnTPvdKeVzxxkygHa165nGtCht
GChlk1hNk7WD85gqyShKgJU78PCqDPci9FFYKhAPexBCcwkMRIwHjX+31VZU20EptIEAQ5SYQM5q
VxLcSfdfjDdXEQZjXzFzmbxt/2m2IkCi7g/FnzcIio1390UKnF/zHH8g8O05OvQPQBOU5rysmgLf
DCDHA4SKNJiv7SHAT9l75XnqZO2vzPseCYXl3coywm+gFJrEIqQiIRsUA5C6MO4BfHqbvPYUCrju
3LQCgDfc/+JY7uvSyEFK9qiVnTv3Pid4d+ApsvzgDa1Pesul/Hrz637prk4HenMSzyiojPtStJ/s
u3R7viZdnHz06KxI3PQg5dYTBmUXu1NKh9ap2jlfWUA2AjFL8zASrfs6veaWCwm5mTB5ua9kh2Jr
jpj6GItUA6NqHZ74sk7k5IvCGYzYMoO5M9zJnWK9PeaXde5hNl2U+eHC5A23Dkyq/+rFECvlu8E4
GGsWoU39p0Q94YqgKX3VbrnsSrJH/HhQsnudLrloabm9b0+Bge9kRaue/1F3N7nyzZ9bMdh+C7jO
Lgou9h/4+mwD1vNMD2f8OPP4nG80d7ywPsCGw6Q95kkayUzMzedhhKJ0rBr4OUHiTNsEmpqcH+J3
tmmMpjcl6QQZk3Kgxq9LuMMacCr31a6QCO1x/N6QCBOV7ImbWmjGu65fJ8UA3P4w3A2u1b6jRsOv
2c2u3Yu+9sboYWa+t+hdvkUG+6+JlKgcsQAJvSTxhCx7pr6QILRGWDRmV5AucpE6pnyUgK7QQbLt
igUgvZeGXGckVTpbQgd3J1zCRaM5wEMd2Ol2MXYqRpamJR62ZYqFF0r/jnryMzdn9Ay6rVcNG3Ft
3UJ8OvtW/Vp1cfo6GaxU+fCw6SRqFzyBjy0Jc4u1bNmsGFsS7TZqtsJrxyz5fy3zZtejJHZd8tE5
epJ2wjfdSzIWF0bqkvIWRckalgRVDBaI67Pv/jMD5hiABMPL7TK/L5zMkjJETpPVtG8jaoMx6N6L
64f38JhHEUd6Kezo1fol4azYCAdCiAoJAqbAxJ63B7IPmKl7MioA2jkytLMBMDWGH9fJdwCg5mnh
YLiLHsv2b47gVIzlLqbF6cPKb1aayf1j81QKeXi3Yh14EOamwZLYRPKdg8kVoKaUB++tgQyn/fwu
Ji6dlU21wy40d9Go1X6+1688FlE2MMj2/KkkOwn3QzThxwO7pRNzFIPvSXR6ydGQll1vEcGCTRVG
MrrigLw5eKXbadHp/w37AHgpdkg4c3Tt6iI8t3ta2jOXVk1xe8RFsuDEb8PSlUEbH9d9di0bkOvD
Z2QYtc66SOPhPjiIw2EfqKC07yw2vqTrhsYRIIYT3ginsgFGthLP5cO1G6Kr61obVSxsyl5tzMEZ
Ni9LBrozZHFAVfN3NHoW0qChqSytxReHlXz3FY9AGLfUL3yE75RAVHfDVbzpMaVUVTpuFYR3Yv0C
DUh0TPlscBb5rLl5u/MyfZ/OVouQMxkirL+FFcWcVOMjsMkjp+i5pw4Ldtrq5dcDzsnUY/3yF/p+
DabWWvKopimm4LxtCXptWCiKBjRlepatndZ5EcnuRUtDRHsjp3ksccrVGT2ngfs/33YS6/fnFR6o
G02wLzZRtHJL2fEHEADhn4/Bo6zg4jmyC05eTGOezbRxngvV3Y7HAA5nKaXM1cRR7+faK0zSkB5/
IkAjJ+yMyZPFWfN03ao6tdgnjFGLzyxK18GVgGSM0/1mf9so99/fs5PrzykxLPIGYeQGA5dfpUUw
7wabdvzbVnTL31CrD41OP9ftjSxuoS9VJBUXbX18XU5nqEdh0tf20AJmF4Olfrp+FHId87Orj+WH
/0AUBTl5U1lWwhXVUHtfJsmmtWwV923S1FTeoAxValBX547y+dm6F9uh9oRBzhjBdNiL69NWHz/4
6rCukUj52iS1+T1DMIY4f+HIP9+PzeGkf4IE2Yxd5S3FELtHN/OZjy6bQpn6HQBFt747tB3Rav11
fFIYrYGIgSo5gFOlDkc5sGFiGrn2bLaGQOfzOdwUaBAiFFIsD9lpyBaUOxRBarA08JX7R04sReU2
jrkWNKNhuDh2sIE3ABegoyasUYa7AR+Q1C+pTp2vZabHh7xYyAT/PvfezcOVGweKtq1im3NEJOx7
Rftxpssee9KdtEOYhm+z7yb0adEVgIMWrUbfI45/eF1PvsdlFzY+B4d3K/DOl1pfqCVGzyQH0Npz
7QhQJ4xe+EduCWoqlkK9RoKwYcISc9CU5X/3d/KJnyhr4v6a8LFV36jUHGpGGYDRIfwQPhTAVTwL
02pBhiFMG6A3I0bR1vzlXpTWmeUwH+SmsJmiLEpY6XSaHhGx9IYyO1nMExTGF7n8EtT+MMnjHUFX
0udhdIG7CFMBuDieU45D0Aoo3QraYS+VlOMysdKU2cBGg29hcS9nKdFVOwKLZTZLOngHGz55NZwF
P5iJwLwydmdG5O/+cEQlqx8EFRak+oTeUUj9er5WBYlgiUEeILVw44mB7Q61RbT0V0AqXhLJvrAH
9T4atVbxwW4XNF46v96Li/lpoxyXCIp8yMxO+sU6ysspEoCsOZpN1qm48feXKUhLqjT1xDjz4J+m
im4GAk8KQ1yZy+0eIGidpKQC/uBlmPzzkmLdfaS6MLrqq4y7r3/WSAuUepJIni9tQQYN7oo9FJJs
ZH/15NEJJs65892luTtNFt/ezypTUoLZ+vncwQuDD+Gxk9GL1lm2SGsTuBs0NdDvIQ7p9W+ON/ug
p3KPfiU82l2DfDaw41ij5DWnyOJluINQhqxsrrDWrdU5JaX8CNHHd+zsNbUfC6LDrBKSsU/r6FCE
u0TrEgVWLVc0ozuhhI7NCH1cpT0ZfCBs4nLt3p1H2+v8Ghlr1/245RdNEK+aYrg4tlyLwWMyT/nc
swIcIWKuYUgs5O/fekbEN4D9b1v+YpyvwmWgQdWRjMPNY6OwwzifijTcRJxnflocrWZY3T//yhWt
/AULZc99kFZEKGmQV2MnAp6t+qmQ7P3w/wDRMft8G8s2UUgCYF3HfuY+nBaOXunc/4VJeVb5bCXv
zaqFpjW9kieLYEPdNmBW9OzpTOHUx82k56AS1OLsOglFJYBtt4D3gEs/b5nCtyJySX9kIWDpU583
dCjytnK7unsbVU2IWLeKGP4ltMrKOOTzjvp8rhLjzai4m34QR8amVo2P1Y5QFImM2MBk5qQ4v0FG
JGxAbcJcrkAo2QrclggLcRq3lkwLdSO6fLvkgksdT9vrBS4ln0FnYqYJLZl9kX07V9GecOZLUEKP
CGDA3LwI7+HHFxFpQOQ97EesznWhgQozBlFwPMQRbmYO867699UVwDLCSPiJjHNi8NgCwDmqL47X
goXYB+Iub1HsvPFwIOwuDMM1LkZBuaYt+tBiMltDdlgxAA1+rnWZRZUpjwwFjslmD62S2ch+Z1W4
pSMdkRbXqso7uagXWE6T6FgwrXcuUeTeouM+tRco/itj1UZht9Sjxlg6Rg+YsLKEU2CY8OnbhWMc
nzShQoPDGXTqiG585EEWYYXQ2ie1J6QWKA0IvHAz6zI64yWpjw9yjG1z0DLY0GhiYBL27OhuI6Bb
5DW8/uNO5P++TrodiV/w3Ud2fblbrNTlq6w2ksi62I7MW3ZeqpcD7r1feT5PJ6+TcTDqjCxmYxZ6
nwY049Bcrg1lm9vXQx0A1wwq7fl83VM9HewnDaugiQScnSCeKbb3p4VmoOXdcq99xenhOcZJztim
FtfaTobvu3kjWgGCEtaMne8efqJPnICGv4rZRGeSuWruGZgRUGeUDZyjCM9sPeCbYvtAB9pUICKJ
OmCeFt2Dx3lZnAO52tq+PjSlczbbSKMg1+4zORMG9AsCjR7rONFXnw8ebsAKbAoj+MQ5P+xHmoLL
zA8rYtumT59pGEowI10lZPTEpD/iLET7XmkpfwY8LJhGZzHANfAIj+ZRovv3Dk6TL75zZuT20ED4
afIfttTpgbJbouYd6X5XMmbBqezks2d1hto6lu6nbN02y8XHQcGtQ07k/TD/o/1eftv4Y2owXmyZ
hMOYOIFIaXkr8HtImCEjVm/0+1M3QMwueW1L6S1J++aUKfAbTC3+7RenHA34//AkfXWaTIppEgqP
+r9tLjVR4Nzc5QUA9Tl1hm4JBc6yZtDSaHdLzMzdW6KT5Tq58I4ds1oVKOuxfShQlJI3sz9G6mhZ
EhIivJGUtLZXYU5gvcfP0hsgLpyZl0U841R4TvEZ42BzYNDcs9g58gayK2+yyyTlIyKtDXech6VH
imEh+esPTKCM0BD+XPvUbugG/XFd7e7ox21/3fzXoaY0IjtwvQmH/FdDnL13GHKO3Iju7erv/iZX
GWS7zrXus8PQ2CsUyFxZeV0kLGohC4mvvw8Z3w+BIfsR3Qyj+IjyIu1t0id6FGqxFuukC6NlJT/N
ds2yeOslnx15qFiPFYt4SbJi7bHv231qD5aKEYucSVBxdwQoVECgKfRcW+d+W6yrXmVmb7E+zjoT
3G5ScIkzspWGMshnJVyGhjA2QhtzF/5DAiFYfz3BYof8ugLpz8LLU66uCsHP2HtLjcJ6Lefcd27Z
g+HvNz5gOgTIGO48A7zWOP9c46KEqBPFixmpw99a1fJ0/IJ9NyvGNyzwMjsB2cRz0BERo7cjZU7K
ryqG62H7KC7ud1N3BT6NBi/h+LM2gMineybOVYfsgok5DVRWzd819ike9kRpxD8osNB9b+sB1x2M
KZtsur9+fuQS2whXuVloSjsB2QokKkqzeSzntdMXFRdh/xUTqK+I0t/A/VK7xV6HkM92lN2IevGE
RJftkEDS4ixvtGZ8qM3VTycwRmuzmbzy+mE9WSiKL57aut/0plebJKip9fKvRMnNNEL+IwRTFy4h
S5jP6mgCprWkXQKhpgGjmbC6cAbwz5FZrFSwG4nas/ivlY+WItDXe9swBfnjeqQGY7PMAPmvsKOZ
8kCCHIZrJlMpctAHi4EFwvLxJEtDp1pLJyp1cj76sXcC00FAX/rH67zPNE5hfs5As8Y+6Xaz6Dek
o7pE3OuADgOtJs9Hrg+P3XYDoX8zWcqoOCDkXAIGT6DtsjpE5mnGl/MCfVb10aHj2eb/h5zv1SG8
+7EG61fM6LvenfdF5+GKyTI5JcVae5NtOgz8ljJo2B/K0I9y8wcdKsESzKiYD8eEgKCrVdEosEtW
VsIleitBkXTffWbPWeNZiXJMz6mIJL9EEjNQvMDlz6+DiF37Zwh8kOuzLdLFjgC9YNo9Xx6WZWba
CRWH5ky5aOLsvIs2kHgCj4X90IvzkRLw4bxIZpsloOlvAwd8z4kSaaflQe5RLbw6KQ4u0c+WNi04
CMEXacpPeoQOrZOT8aHvGQYmpGzgxjqrcett3quD1H0cK/GGfUr1V/yHORO65uESvlY8X+yyM5O1
fMHZtBqAmeSFLQcCqIy8/7rsyf+ikWMJhNJOp4SZX/2ucD4cYN2Mtygm3KRfV+WM7A7/5kdMUfL/
K2d/yd04qIprRjK8ChqUq6EcTT2hKIGP6/klPREjNos9FJijmg0cuFX0qhOqhP1o1aE/4EUvzDb2
099lD/eZqGhxSELzhPOzPxTS4Gx9zxtoMSXdqyT5+FNHZtAKTYAc4I/0jDwqKAdRGxEdQqlL0bg0
gBp51l8SrQEfmyDipEKdzRenDoOxR+r7O5XOsJDdJTRuH6o8REKTBBjBo1mn889zNqBxKgm4Zvrv
Ux0P9AZBPdaBN3K6CX19u4e4s38ejJy2+9S9Tk+AUYOp8IJxfF2R3N3RWVhLs/XgFUXUnpBRUjjR
XPMGTJIJtG6sYb7nX4mkM0CpU8wCURkyamK0Re6gUtvqBxqxwazBCqzgdRKjRI8oKRZqXsHTyPNv
129pbTxOq6Z52X7ttQeetfIBmTW5z/MEvdzd/ssLqJJfn4k6yxstlw26E2u0YBwpPSdK5SopCM5K
7TdwibI4UIWUzAHdEm6xr8MHt4hrVKrspcKw8nreQTzDz4Y8mSosNS8oDNMj/ofw64792e/Yv/mh
lpRECDo3jFFxCUxa1T1VF/eVbicvRH/uwkbMPerAUnd6d/C7DfA74NAvvJ0GUP9uCNcYw4QbgxOk
r+H59fFLizPfjtRCpNGTAt8nZU/EbQ//+PIvE9hKwXq3Rf4e3y73qM8/2+z9N5S97EZuyrSIu8Fo
sJzeN+cUNBUtYiyQbnPplPgHqvU535peQAMGrPBOe8wuiVnnO7aOgVb04dTom0VI7jzOwmJuB4/4
FENbo5N3m3ikjnnjv3jRRrbcOq0tcbLZbxOYEwgmZpZEE1mTNSvm2UgjX0CpYd9+JTOwIGdd12nL
lyezuMjF78u6fyFKXYPnPurHXztYMZS/RCvzpR6he9op7D18FpKVeLBYFMIeImqayrXnmYG7omB2
FL+EPsLzP1UWE6iPQuAGE69Q23+Zj2CnYaM3sSbk+Lvh1YO+V6rALk0XtG7PeEmKrDJ+oHgOEWX1
2fGVPoc36+vLI/j9o1mLSDfcDs7M3QegMTVBDl6zLbgD3Z7N5mlvE+XNTEjzDaervwzSyIZBHJgZ
RWQnbOipOe1R+pUWMbqqYtuhsUBo+oV0rR/DMA3Ulc/86EC+o9NzAVj3AhdhfNipQ2FZMmZUhMKN
PshO+D675kncDOWufzXrLWdChe2tu3dqnsWox84CgTeeyWgLeaVmZ1SzmBb6iKsJULv6KkEcuxcA
Ia0Qrm05qfVW26FG1bhEGuxtQaJ1Bc6wpH9o18IPZTg6ZcDphW6hCPFQG8ZZyC7IJkvJbpjZDJAc
qITUJxG0F+uziDb3sjbjZk+9m+89URDMoaE3mKYNYC/3mi88dKA2mu4fLg57N+OO95WlzPxV9HTg
Dj5YrKFW85NWUgf1jSG44BQgROXrw+Zmr2qhrDRVvn58JT+xR1t/emajoajwa7E4RXbiY+wIZKmx
D0D0mIy+7jkiP7FgfrrSfh5SYuJ2gd/pOyEAJ00HF1s7kWLltDlDas0ZAtagiJN3PYy5uc9J7JOX
el9rzXH4g19FHCI2Sf9xdugWZifgSamzrUQWye6bEmLqlUVxeLZjhPNEd0qqAwl1NQBtZRbRmRH0
V2JTCZbo+f1JxV4aKHZMO+KBrBN3lXGgtR3iZHMwo1bqZntIPk6PDceP4BfYUPcvYYNKzwH25RaU
BXccyjUiC0Om7oLnbj3Shg7MkealnMMMVngIm9De3le6kxNXk3ZS6n0fexHPUuyeqXo1BkFK87Yv
/wKqlW87jJ2dVA1FJIJTQC7Cuxb4EPcQ16Ix8lwrZkRWC+z7UkdlKivLzmufOmDPrekkH6TaYAIo
1+Ksx6BoPo1JIazZHPU2n6ORobeYfKTO0SI1P2djgl6fhhmyE+Bv5PNWmN9bQfF1e/mkGO1/oGR8
+Za2muZ405thd9l+isd+3YLi9nBCkwp+NSVXgwb66w6fgjFNKUByAhgmgbtH4huE/n3sVA1nZCcl
jlxPgpaWAex3jg9MtX/bpAA80Dr6xoG5BcFzne6qKN/JOhO8xHFKvAzzD3vJJeJjvj+NfFw5PpsE
ct3Y4G1ricxFyGdRSO/djnvHz9tlKkaRRI4V2bnwdmdSNhYhFKV3jQ8zCmVAZKkfkIdrcjlg80XX
kFXpUPOOCw8Czm9LTz3l2wpEBaN1eiTD3vCZgjX6OFAI/5nNIAJ0orse1cc9rJ55mWS+UoRWL+cd
pUEWV39DhAEH2eKYRHm8nkZDSKFyKeUbKJK2LYG0+C8m9795j8D5CsqVQFJAgPSaMs7Dym14kO0p
SC6e3G4U4ZPdy3TR2pl8Wfy+VpX8gI3dhjRZP9uKrcaeKnCX1Tyq9SrynY1XsIfp5DWmOK2TJh4d
8plBMsgI9tGqpBC8eK6R0W6C+FjRC8nU9JyO1GYLNL+R0vLZztDvESg2CL3Zp9CLzWR+cL0tWKre
CqAQ/G36j/ApRloC3ZAJ1IrrVGTXeywFzjaGI7b7ks+CgbY0aF/zz/6pI7tGhqB6wvZQOVwE0Dd2
kJyt672kkZNHvh51dpZvJ7nU3eQj0FedKEwnCunQstybQI13knHDJ1GJ4y3Hv+40w4IWjjh89suc
PHCVBWYmcBtK51ycZFP8/29b4VMn1HqAnFFrQKdj/fRr2H2Aj73w29n7lDuTQnzysoWTHAKqVtWo
irNhj15z5CB+DOW4VT/JysZkcOQjFWh7EwcEcgkrkSg3SxdJSEG+w/e9pGEfS2qFRcg11w2955Zu
MdSh+Uj3D2EO/BnFNkhMWsM9xZav0GqAeZchHLO3LicRVI+kiI9ni+cl939Ht0Y5XYquoTYk3njb
CWeOIm8luQqbbF9o4ARXoqREDKUEjPq6QcmX0/kaZF+HBCYobwqzHlEh1waoBEaGZdTBadybudIy
b3TsnAvkTX0DNWqrNBuxij+ETnQ69edzapOdJHXMGSxxMueJc0vGEX7QURm1JSuK6LRKofX96UEY
aZEyc6mE3Gx2qjDznaGEpBy6fFyuYjSzxDmZ1Sanp3TfyjjOqn7cnOVLWZzMIxc7k4y+ooQCX/VN
nyX03OzReVBfLphejumXzdi8SkhM0coqA20e6Hgp5R0yGWjzwdzCTq34nObQynF+NyxLHTxIgLle
JgjJch2MLAC5ch2oNvDhEPAxkAMowonarTopi6G32c3Qe0yVLTPOxbqU0Bu3GgLk0hEdsuu8dcfR
tJ/Xg7h/+t1tHdMnoSKQdFtcKpn3x7URcM1dD4PLcWmZs2wCVYvU/uuFjnqCAsiVRjNpExW9roTu
JmU3OU0HqbkdWDzxsZPpF63qo1Zp8UznvUYooDBfjTAqzwokWp8kVjfGDucjfSkD8zzAtObCkIIf
QiyjHEkUFnfVRZcrmeK1pEUuHAdpH0365mCmYCwlKDYcQfRfIiyWD3x+Pm7wGPWOIXQrVKt4LLlO
rD9gXDDEJw91Uid0Qt5FQL2gJZYNGhRVpssCdcn3sWD9KQkqh1YmoLy86UbPdF9YRO53nOzhgQ1y
TuRi67uswP8gCHXIYwpz3zrbNhoMEGG3k3x7nyOpy+/CS6F0VDdNNNhWWTIpUpmVydf9BzkIx3La
NSR5oZZhmpAllWXEOmVaEQuDw6/5Wx7cbTEGciFlNT393+wXvS+AKQSEzYxjkdNR57PrAhvqWsID
lOd4G7d+699sqKiz0Kig0z8hhGC+AnczvKR0Fwg9V5AindTKRUUSfv2Yiw6Mv8hLdjbhYuIzU4l3
BlsY8QZFs9RQ57EGfvJqtygBYkbS1GNXGp8d+MOmxm/HCl3QLDe0pHrU3E+kz/MrXqQUGDeWZwqx
IKWr2IW28MMZX2YOs8fs3x3vtBOHL79u4IscxB6VOe/smhHUBZhK8qQAJT8NeSWHQHsvWxkCAky/
Qq/4XcWtN9EsrWBtG605uh43R+IjWPEEwvKuV4qK1XuLrQPD9gcY/nXeL3qR/eH7Z+g9abH/Ey2+
i11f88farJu3N/YjCIDfk2fgkujWv8awK9vYsNMfg+VUhZTLn+IgOa0wrqtX5+U8NNqWuVZVGt4s
FjCxQ6AT2W+xh/83f1LY/CQiElD2q79GKQcKO7kXCmrl2OhuQN9M/VglI+tJMs6goRxNYqxyvIQn
xlMe26aASVP7FyDnrZiJbdf9bYHgWS+NKzT9Ea6Q2KXZSEztdecXZpY+MRX6FDsNNfKBtMWDplni
/RDVA9+UcLiw+kDfQCHZNpYowVBV2aK6g1z+MWO3ogIx0x8Zf5T1+NZjWEqgpFy6MVfD6DsDwz4t
nyQdOZqwgdbQrMad6Pv88Fc0UyINC5YfvM1eI9ujRTAJoTS58v9yOvIfK6w1U+LcYbzivtgMzF6W
heiUBryLrp8iw7glXCbsMqe/eXceDJDPQUa1xA40GkHZS/Z7F1w715E7WuQMPS/0HREPfTvUHEik
htvMiz7r72xQBXxbzJwd+cWDLntSJspA3Eb1w3DjKBI6sSVomKpRruQO0jML7h6BU2OzsY9zAFaq
AS/yZfWQIEdFgXcHG8ehSy1Yb6wyZR/kcFz7YtnHxXQWLZDNlgcM3XWsYoIPPAqpclzl21YhUyWp
dG4H0JL1WDny3oemSAHM3dRZTZscIed8f0KiN4O5Bd6mKpytoc2AXtO/55j4v+zuCRakkvQQEcNs
cdY6PN7qjgbqiGznDlCqqEaaGLaAMMzXjvxJiu8LibMuyJKgzt9xGWltaUK2SK0s+aJeE22sdiHR
GmeZi3+gMzxk+I0S7K4nw8ckMkjmxfmsVO6Y4hGD3BB+u+UZCYdqyict7/qV3d06mT3Zffpe1OeW
Olny1nTRdOmTdTY8KAUK4oXfsZXHE6fNgdIN3gtCcnMB3lVZ14j54zG/fGncqsqDA97Ljkw0GZ0/
S3T5ajuh0cOiYBInWu1LtcGs9zeTne/RifQ7CDEjXmfExJKvk+hzmBYRI4m+F3NLuWtREiEBUELQ
mxyvzKPqqzhRuluPSf9BZZrY08k68eYGmqFHmpj6D+Mn3Jg2sxIlmJdE6/RWBGjueaS+Vy6wk3NP
90TH/GPmtTr1vQyIRgf8Ehw0oEPpYTedh4m2vmceOr4Sip2bRAaXRc849UjjUxh3iJSCwmH+OvbJ
QTpBJJ7nlmNZvDHQ+2zhT3zuD3XHL/5cAGDagsAd7ScQTG+STUJKcRNJCYFEGAvXL67TWkCCzwXv
sbdRaJOggte3YhEBXGzthPp3M1EUT1YEAvJYpbrQRdqnKUYlTcOtiULXenvBRogvxS19TMEo686S
p5wqrlffGBjAV28jISoJJPElN9QR1y/B59/5blPWBQz685n9sVjraNVBy7If5NLIYwmWnL1ywGVw
K3Vd5QcAROILyfpVFWvmqci/p0Lt2aYSAzZUlw60SQI2/WmHbOJ/NA4AbuBQ9hmXGXZzZFHyWUvT
GF8Ucz5ngrMTZh3oT3nxBnR2uAJ70XotKA0RMwZHegFiXJC/n9zbHZibM8Xr3GuPJzSGbNvx2Gqw
xtxBZStjFeNP/+CchI03fjywEOU06lTVUSurvR2LEFtoFHgd21JG6qtqFFvEcZiTJaxRMgNzrQQn
2MJ4TevlpdWirQZh0JiMwS8dZLjoi/KGfLaNkdzXofESm5rx0WqtwSmWUsfJ6ch++8BBNLLcfMdf
M2qdvqmBs6+05KMcRoMMqWs431UoA3I19pp4PnIbqzoTbi6HfIeBVxMb6qfrmRILt0MOx049T5kB
EXyYWiJLcFNI506cKq7lVmcjcZ+BcqyGsVZ8HNE3QALXBrEZw5VMqKw5D2jDsSBH2Z77P5TvUHaz
YZwn8hIZjl2TrNLDp9jHGfmEE9gGAe7ZJ1WFU2Gd/5LGPszPnmY1czF9LKuD2+vViVurDAGa/ayl
qDllE9ISrzPV9PnRus98CME+SxCshrQVwvpSnVFu3PHEAX8hVbzuYwdU5xBJyLW/nEhBDmQfMkds
J7u1H6SaqMdRw195y+Uh2AFAlmv8U90NT4aJ86RPx0FeuNfccEjetVmbLYoFKQBnUACSEVmY62Rj
u78Z5XEvuUsMI2vxPaFxufTZDyzJXCEV0nUqX3xlagiy1K+oesH1j33vray4ebie0KQuxqQOCFi2
vUqc9btZFidpyJ/Akv6nCwhe6tW/7aA07YNmKtZYK4tQxC5UCbpvGEXyYKeripPX4fTzriOcyJkP
AD0NvOnT+4A394NgCzsqSx95UsrCbK86b1UKTx4ifzgKIOvzjc3msmMOQCeqgy+BKFjf3ww1Kp+B
16CF/XKdi9Bc9FLARmLe9nPJTOrxvCuc3YuwMnzFUCAs9FflV51Jp+d8PXYtcnBlAMLBw1aUd3Rd
PSBYbFDt5CqCx0Rfwe0tTiVUGBSPAR6GXyUtvn/ejQgup2/5PTL4QyMWx3cvFARHN3cbW+c46KeF
HsiNTWmxIWqa/L6Cyq2grPB2J+QjBRk/gGDghDJEo78GXZdrUkUvdzc7hdcoSrrocmZyBdmhWjQV
3gVdbFK88Z4aC1Qx3LUKOzMhFYGjtCRI4YOemmK4pHBPmRPpnGwiT4+zs2BovhM3DUS968OsRsH9
C8Uaz10kiMLiS4Lt30MGp2fFfmgeW2nqS6JrLq+OY2zcjVxM25cJoriSXe4gwiK1HAMNZQtGVwk9
zA7aQ7Lwq5ml+7Rx5d3EccH3EfG5JDJUjALYgXb3BLiWBzMZq2rlZyA9Be+SbD0UZjjlKBqMewp8
CAJF/8ux+O8XZSdL4C2T9/sHM6U2djaEC6BK5ArgIJPM6phgeRLy/TfSf5UqzQkWE4CBwA+euQWG
oR8xm02p6uRnzD+9Rgh7/ko6ARetms9wY2YNWFsejvB1L1RUD2pVOSaKaHFracWV87qpyfnjLqNX
aw/wT7iB32SNUHuOfO364nVSt01Yo1+HTgFr9mHm/HZyrbiwA/I6MtBQTn5z8IhRxAdjHptwb155
6G1ce0aN+Kxryh33VmYNWsyaDPz4vOChFaFVpeFtZdemutR7AWWW05Sh+1BVFpg5wn9HIyDSw7bG
dzC4G05xc83ufXUMN1tTa+IAKgfJQ9MGCXfUCyvRQCCLZZdNPZaV2erLG/6yuNmAn7qie0HRTafj
UtG1Zigflc7NP+edxhWSOzqboSAvFJO1gF4yh00Gvok65+lN6O8b79ZKnv1Wg3pehu32mmTCuj0+
h9rz7W644ZTd/sdzDr9bllAt+NMo7QKA8bDKyTHtX60bHyyUcAxvqa+cHydl18USg89n2dvXipqu
darPk3p6iTO5RJZNR+JoOs5lsWiGYD+ssRAF5zILAYtGQuxFoG5T0fQJFguNSGoxr/qDwlxd8ohL
Vdi8DPpk/JEC4lmqLeaqDQtjMBNprS+w4U48n0EmX6k/nipD2mJlER3SwjWUADXVmG0EB2ja78II
9oPQqtg+mvyXQ2bovsBOFwvUJQUTO8ejh5dk7MnECe8uMWYyTk/i91ES2HEbtDvuWwR6j4VRS2bA
mASMsQdLrPBjKA+/oHU+uFL7zwN6225U0WLXxWgA8AIFNHEFqx0dJKNKe4zcdaGuBADh5saMKIg6
KA+QYuyLUD1mbQ0Wn6iD6Df2WO11xgGbXqeEAycbHOkkPsIQHJeUyKtyMytVyq5H3qWHiYzCXJ2/
i4GBCQA9T32TvSzuNwyLD0LEJ2UnBFg7yRxAKOQFJ1dJSyrQijr6FkqobYKvubOR+z+RQGxQI9zk
MlZzx3WH1Tr3YiQ5AZ0ITRi2HcN8sysPuh7NL0UoCs9hGUKd9N1cMuiyUPq26pcFHnWuX2Wz/BIa
A4qZAQydfIugZ8s3K0AtUckdLnJmQbQV+blGWYaj/9DAXo6PvimHIsmDzKzmCf6n0Aws9N8uegEF
BNRmBXUSKaGcWrM0XBK9RJLUmoLi8wiw62J7ZGkpdgc1GL3AoC5SW0FDKh24jSjjn1o0I+2n/uhl
q5//g4n2Z9htwJoH3fr+SK7vsr0xKWpfBeo414hQejpg0vmGu4VZWEbBynVrsFZaVEfUPoQXHksH
SBjqJ0cDS7RJy3fZwcMpGq6QmYTz19tdb3KvNIoP4jUNE94sDAEdwgjPEJAAnRclO2DvTy4nd8g+
yl9F02hN/okC0e0Lxc6ozy+KsVI6UU9ipmZzaVIyd5dlPjKV1pjq6y596/PAZtKl4yR/J+LarqmR
EUajb7MoMo50BbiOFDyvJmGNtZngjKDgM1PsYtJqy+1sCE16BOY+gBOyH46wtF9H5eYVAkc1QU0V
KJeSyzarSBg6eYAgmWZua5aZk/5BFnW4/q67WUi27tkMiq/vGEMwVkiCkojW5Ba1b7ASqHdE5yyw
ri0QWt9nxl/DufiSn3PLZlFiWhiboiyzE0mLFZYc5EIKOv1hdkByGvBvz42z6Vx/hT5KGbh23E/D
NPHY8WWLJ0zwfYmWphEQucjZpqIiLa45MzorcgYEkkcCYRQCUHPerf+UwffBx63bIDlESLNB3oXw
fpDTkDJ60Hq2FcqnFPpMuh9LQygd62Hb1PDri0tyzLYh1n/gYeFHLc5EJ+kUXawx6KPfDBx3HgpA
522eDLjohR5qcwRVbHLz/cWC+6V8H+ZK48VkKdLhQuA/h2xVBk5oswHSRWygHEqOKjWYssGMSMDp
mNhBjjLUUPXwEeqQn0bQgqnFxMBbksSJKTiMSEi7JELlDbcrw2KSsoIC63cX2GNxmNuV/buOzxVk
CKYsjxe34ZorCjwSM266wGwN+M9zVvid32/ALO/+3NTaJ8sz0YFf0WQwugGbseRo2FDJezGJFwMt
XsDjt2auJG1RNgUX4P+epwNqAhZ2ZlyJtMSwzcJvyscuY0vp2VARCo8Fa+q2QcEaAy9Wt+BjrEse
9f3oDWTCMXlm0e5ABmsPadf+dPllitTbI7KkgIAyqHGZDfjp5EVoI0lBN2UPILfBZM/svvL+mdoI
hia007KKr+7mLI5rpas35CcSFuCHVGHA+446wJ8wRIkuksYqPusBJDT6Ws8h1XdBC5ry6V9Ypvyh
vhNwlxV+KeYdECbX7/KJK5fHmnkaSkyvxicpS4d5ftEBs+QqH/bCEeLCFXAJrEWH74NY+EoSV/DO
WxOk8j07HJ/twzNBLT/3qfLTCDROgMJd0oULo8v0jSuLzjzXKjyYh2MbY1kL30OEFG9OSDUJ7pfx
kdcjwVF9hqu2bqRNlmLftjTnFiWNQlsTl9eCVFQYOK59sxIIKDwDEJPlCyD5Gt01KAzHhh0pYP5M
GUmZv8uKHkgI7ttr7BgIxjlaCL/eUQaZU2U9RP/QbE+W7/Slg/l6I10oX3EuLE+N++qQofkZ2uC7
jb/qVNQYqnPZdCIf96h3qt6FRyrEORvSgH+ht5N/6zkFQS9lXdcLCMTvtPsTJ070ZvzB9yVySA7H
ECuIbVRTtjXfOk0yfn4IL4hgLOkj+phYMWGqEFVqFfc+94xrS845BWOlM16Uymn8JOMw9iyvFqh3
0fWIzYjENrcY7unFN4WWNBzoMfVXrc/ZFgIbWZRXq61ZKDnUeaQ/G6Arv5gaKwGTx2yLdw8KixU0
XMSQTXtfJW6JCjtpbZrQA1WzMCzfVYWmC1d7h9StrWotTbRiWBgGkOOo5gYt5Q/yBSfUje4o4npW
NClKPrP9GRQ805++ezfV5Gfp3q6bfBO02E20zjuAEwjZMuZBE0/t/XgGR/nvmFHZkoD6tbgSZsEw
iGNyHgaWfrwMdlcKTGZmLPlyHYNFI7pnL0+b8E7/xLhOMN9j3OUQL7VVK7oTkqxxPJrhIgtW/D60
FXX0cYY046Bhe/ajoLRcY+8tzG7d2M5+9bJNUQlE/16Q2PAnV6HkBhFskTCIQDRASfoD5XPzNksY
WjOP9rc8XOgAR3YoMXZn8LLtfrSetZuovsYcfEA5igZD/nhV8PUVH4JCndvpXnnxWJ3xNme0LSOc
p/kJf5AQvztGYcQNq7OYSdXhQHy7MfAMcXNI26uo8EYwyXZANnPhc5QjE8zfT5d3oR2OEdSPqHjA
Pj2I69zDrwd0qTrnMsEAPexLpDPbGcm6GXlJKztltuD/nPnPZ+wMiAXnordQnxKZcsOF96VCf3M0
aBnOtNxDDw6RYgcP8arltJNc8hnzX/1OEY4mSTvWpOnTtnEM83+IVP+AQsSyIPA3Q4YDKl9SdIeW
78LgsJahJpMACFNrRKJOCZyOcezONmesv8s852HnBOT3FmPI1XvJOvgerKbLMzccs1sikyk+3Yde
oqEzfRoN0E3Y1DKN+y1tP5JKuwTOTWYUShppMxKNVoBgvM+Oow+9YXPWYdk4ZeWzJsq+GQ+AsZXR
hL8oBncnTJDTsOOydKgyH3MMbaPcycl7TZU0RpFWJac57ZH9GQOBENv0gMNVKry0hJquWXIWaSLA
ZPPkUuxfskvJmRqWj7GBqXnuKpkWiM98o48BqD4oj/3QIyPy1MxOVAUL7sW4S+5M5OeaTvlxcBTR
A54hFLXXvVczCLEc4DIXZ2uh8p0Wr2xZRXT5msnP27G1z8uYyLAcDkgtbHElTsx/Le0cyikuelzY
2wtGUi+NvXY3zzCWgP3AZagWkYuclOxtR0VFepAdaGkxkyz5lzqYQCdzave0vTeZhmLSBtMcRPjO
7TZSILl/RqMDtkq5McM2yJ4KiFV38At8s6RcQS++k/ubnbLapO0MP6hX+vYmfz3e9lqfOtKncZEZ
90v5JlgGx6jAcau1xy3TwLc4hhZaeiVkm/iXPNzM0G99r4pvL3rThfhPQJw2LJM518cZGE4htRPp
ySCO6ZlbuA7B9r1tBB1rIsMINSGWpSnYuAWc9XsmAFuUTRomX22mqruRrU9WksWnHU4O6i+kMWfc
/pKC5f8TMDMVgBNsEUpeyvH8H8WFC5tlOKJAWUV6pOI7OD6kK990bqkb8k5ixP1zex3vHx62BVyM
4a3QEf09l9lytvVKEijzeGyp6lXy+hPTxHjbxMWB3ej2PJM3nYvYvKYUnFYzikP67739AX6zr12I
QS9zvta7362SSDikjZYf8ThZssj2GxRDSMBgAAFlg8lIc8Wj/w6ZzBOk91vub+jp2DxxLSvhDJf9
cwul2GbjGBK7sH3DN2S6YC195sLzCoA4CAPmWZEBf4uKufFNEJXCCKFejS05zH4oGUI6btdQ1Bny
AyhSgWYA6onHdicGsKA9HjT9C+gdTZ+A4FjpukQl6Bt1nzcwjnukumeFThCpULgQroETUCdIMMzj
/wl5o9hp7gJP+Hw+PbHnVfBgmKtpWdPq5Uv/crUez5EKr0ykco4KDUKPW1tfm7MrJEalAEMLpYNn
FxmmiXHNLiommYhFsqAFYLyT6QElCpic9j42j0JKVrCCqLwpahkxy69iExzGilJphIYppMjKOO10
B7ThapczbrdWDEpV9vfXDiWLuXq7aOaYj8dzWXpDlv0aVJpwWxjK2tgvPP7QKv6EeRDCSW5cByPS
EWM5XooJf8DIDP5zFmP5CbIid00iJ2NdQkUfI3Y0m+RVjmMECur1G8DKQvpU/seZexUYiv3WaYNY
k+dzKohmsG5PJU0xsGI2/1sKi8ND7wbr1keU7SS6V9NkftXQ+IuwikhI3GF/oQINF03BcoUh150A
BSox6TYUwULKxvV5Ulmz1U7XXuBUn1jySJ6kstVaE8fpTLXPUC5CHbRqWFLmgqahBhiZt07TD/9k
KqCeSr5ip5mW1rBA0/ufraRLYFF7SudRxGwTU8h+tJQAQJOjN/kbZPb4OvHMTEqtaRJ5btrW2xAI
ckJR/FvOq6BVbNkIm0LLXIFh6QYAQ6YnM67CX178fbl+8nW1WCp0LWSkWf5ag7+c173CccI3RaEA
hAPqegtZUO4g+Yx6ER/YxNOpVX4oFWykbSLYB4EbeGbfECgzarYCbkEKGXUp9WEEmmTVdiKwt5X1
WOeoAclFV4ZJcTKC3FupdemO+PP20wOsC1WrsjH6rDQ60/S+iBVe3SZIYt9HRSPsVHpb2G1i7n3q
0Y87mlgW8o3C0GYwMc02e0r140fn/GXx8LWkapI1RqjH0RtCANAx4Dpa0h+j7kbZgdqvcu//L1rd
zB/MU4yMWwhLS/9zqcvR0j+11uZR0HprgbvCAaDo8KAydpXY0TMKspoLBczkWXYV6a6MvFLd6KEa
rdq5gXyff20rAKI800fbH/aVAgyTX6WAKSHkMCnzzpl7yZ8UMuPqnnMNeuk3/XpHCcv6po6f5yO4
+srlCGUahZOpw/mIPUk074TJcfCgatpeM86Eyypx//na+YaBZllz4ieL4TKSX8gEOjjqY8r0tRty
JIEwUSU5ZMvN71iUPnOxN+1xe8pCVKEFSDCEk9a+WFIxIG9847us5aQyYZ//Gi59uP32jd2QZDtz
E94xIyLly+YwyesIApu48Je891wWc7dJuDpqMxQt9x0cHGEh+kw0L2RBHCbnxPvdfKR3dXhNpXDZ
adAuVI3VTgyhZZJqyTD7cUZw/H8wX3hkDwF2hXcfHSBuie8PVQuAMl/YzSIj63aKc45FrQWQ/WbT
fsxLwj/V4OrltLjx1ib8t/FWy65yRsBANU0uPGsVVXT5FSoAJe8TXi/dy9QWm4JEipDDtDAnwKzr
5lKVz0JmGEIUx36HbV9LGluOx2gslOzLn/s8fnhmlud3DgRas/jpOGvMADeN/EryhYt9QMej5Wsl
pSxZtxQnFMnyi7gaPPGOjPIkjdpDR6DIW/fXprIhe8S2lm7XG45cI0cTVRhLBzoGA0YHyWkJ0SG7
EuNsryasdGUbk177KYBblr/qHjY7zESuNOFg9e0vbRGUZrND6oYqNUjogquo61UuYrnXq0TSzN3Z
71PkopOZc1zqp2wZAfEFJ9ZxIeIjsVTCMIbs2iUKO+fAOELKbc7js3QVwFcyqBPNqPMva6tjlJKK
QMUK2SZzCFFBvC3qoHyslWV5ZsxSqFHjL/5OJFGQuUJsdUAG0g+DHKOPywZN4mb9lISoaI87U1PS
EI5/WcxY8OlVnCTetO4zI7yBEIN2802ojzkHBxNiB+D64fM8LY6Wy8h6FTHs25oij6C1HwG//sh2
35zRnROv6E1xVV14+MJn8EvguUzXWAQDY5tf8VhNC03UZJk4DwwpVNM98V46eryI1mtEpISFmFXC
fIetmowZiHOKJtMTAPRMXmjCXq8JiXtXyREmnJYD0q0va0l4tiXAwZ/05JaJ5jywtwmQaX2cMrlC
+xFw56GgzAyT9eNEdX6hOkem1Znt5ZEEiyYkURfkl2VUyIqnPnYQxNzOf2e9wrqhPfaMXTV0d4Yu
OxkvKNPPamM8Y5g1QNt7MHHbNR3nQQXawW5oRA6/rgRqL1St40wJj0SWNFBvcXcXaB/BE0XCWMIL
LBOnwXQ9kHRPFhHJyn6OdfGA1lgBqubevkFhEKx0P8+mt6EdQoFQMDUBgNtvmQvVDfMzCB1GBlrX
lfCKNCiaTFpYm8tnML8/GF8VFV0sjk5v5bJ1HSbDX7qD8bHjXFTBIdPJmjZnz8tVtqkpWeKV5idN
Z+fct0zGY3J4cAjy7HEXpb+Kf6LY2d4PESGQE6LVxB1uqlr8HvrrlPPs/AqWy5+2y1h7/KtitcrN
MuPEOL6vYrC9mZqzJmw91fDaei8Cm3pZLSEnApv8Wz4MZUk/MrsTkbGp1RrvVl66JaWfmXgsarpt
VzMCsPmRRjtKX/d+sKei8k2PxNYqfQCoWrKA3D4W19My8nd5DJLKyOQmQl8MLpGiWGRLzjhzfQ9H
9yQQu5KqXX8f5kL27/Ywl3kPzIssTjuNyiQs1HafeBwPo9mcqYfqBnlVLzj3FJBUP2GXgKkG7qeR
LQao7MomaTnDqOXMW3zOJ/+06tOuJnSfIHNTERqj8NkEhiMovQhNkgATbwZK16R0kehkAcOJGC6s
1ic0yHOrOkgjJMz3IvuLswYYn/YEBRsg+M718p2wKkF2OhwrKutF3Gkimur+GE/GzePRBX99FUiT
m+rSrsNnnNkF2mCUywyjwww0ToOZn6+DweeGSps2sU3GH5HM1ZvJ1Ipy+oVL/+m3yOdPNbfTOhif
eafqCyd81gb+G+rsQzQIEeZBEZdRVQte7aBRBS2m6aRZk2vtJLEXi7+aYhRBw1HDu3iWg9VI549U
LHwuvyZJOCw+OOGKMBdgNr6h8FZpbNKLtuowEO/jDWvyLE/kQz39mQXnKo10W84kTGCK8NC6DQoe
n0tNmE1IxUF2JRdlcbgTSLvFW0N2cVQAGjQADFR0cg3KHg0Yy5HB1ARCxc0gJwZWVLfSs1hZjT3z
pEgiZxezQI9N71GrfaY10U7L4/rRnF2I9mIgkG3KAjUECS47IsPrG8+qlCeJopNOAPANPOISu8EO
Po4DJILmTm3vrWY5Ebndo84FHzWdfZ86CEP+sEkmnfdpcVpp0IXzKQQzapSOYmlLxF9bVvMUfMrL
ZNRArWdHE9tBNMp4GF4N47hlfm4i+4pF3lSEMNIdO8LH6H74Jv7x/8ytHObd8Iyq/qRdsofPwAPF
7YVZ0Q5vgPlbBUlTGPX3LNL/Bnc6Jb7mNoO1AGofSS+jWMK286Vmb1FEI76BCxebzbGjTDv4/6Gp
xzdpp+XnZqjNIt9cNjiVpx188XXGeapUf5ANjzjYn3b0W0zJ5dl1pYAWuOYVhuq6+B7cocH+j+YW
tDkPNzhSbzzSsKjuuA+l4u4wSIG+SvAM5aJ5kn6s34166AZ394Vp+HwGYyTFWSL9hJaGdji/7u0/
y67vHYU5EeHY758fv+9deffRV3TSOO5/RkknP2ExOr7drZSvMP3zqP4X5iVCIdp/AMEngN+PKTB7
LVVbxuYChE0KpuOYqvVCVeEQAEYlXL3+jOn5RYEtURGKqyl8E+KZN3U+gQBCqmqDe6CgYVWsWVmL
YLFJTgRVVo1i+drNh6s1f7nXSb+nG2eOe3720WLEVtMf6mA3bnVkhflQ8K3myIlYpUkCyskD2H7E
3hNqZke8zfr9ux73CGcBpw5kI7PQNgYZCVXUwNkh4KBrwkHbk1kNULe2jo0NWHyJyfgDU4w6GdT6
mbPxx0dlzqB6LEU0YF9lQuea2PkPJvksJ1LZKUbzCvoMETOCadnHt0VYUB1UaRni/6MDcwQiCjRr
FBJcTtZgL5WFt8yysPCyKbA/egy+HLDNkJolF8/jBRDAXTSgrMuDddJzRaeWlzpBWO+YvhYr86kh
CzBTEBbYc4irTGNmLf8SyBEc/6jhUs/pRlOIGtAntC/HNlGANPisOWoQzvKaospQIx8W/lCAddDT
IND8+Ggg/Iq1arZN53+HqwsqCYPvTM7A9v//aC2eTbapzrSPRiTM4dfWIU4TQ3WijfKt/Jas5XVh
ivaUYCJFSPqGoojzZnUTQXk4oGQS4HmXD2/+hG5eKJv+Qv8u5NcI0YkbXObqflAJDwbjpLIed1OR
yxBbBex5MyO4NQd782bNAC2Msmao2nWCpjopfRx0qGAl/3yrauhy65Wf54FmO4EEJwX3J0mGkxKN
AlN57VsujjFNuxhn+TRvdgutOQn2+pSZVki/sklwTCazUhFjxKbB/mpWDcyvLFtu8HD2DRnUaWRZ
E9YDmCZZsToBYmI94+EsnYMsH51RvnmzYUB92uejmz6kAJderojTpompn8U8o2Sq+LLyNg8MrVQQ
g3BZqmwjO5HTsbd/YS4m0dUKYsa+h8lLyu90puujDbXrIY21pa+8+85vrLGf3oZciJO0RAydkZcX
dkZVRnc6dKJafAVWACUEWNb1h8R3QtcyTDDWZ1LhV4O4Jkr2kQqFldJ79I3f5whc+U+wMQbyS9n3
bPEIIoU+FY1YyhU9VVkPj9pHoaxP+36IxlHlAbSn8WQHHJAe9fq8SoSeBWsynzyD6HQvtGD1I2a+
iNFahpaJTiS/zh8sYbF6hDk9m4wqR6VtRhG0jmkcVcx1YYaRvY9Z4an+gyyGjgGDAaMsesAqDN50
tLziDRMJkHUXIqI0z6jEOi29NfIx6eu+St+FPNAt2HTuGHeppcKDhOxNN2cuUiiBaq7jfgj55vkJ
B8hmgdeAIiwhDbCv3BXMk+9JuB8cu8qaxhfq7JK8UXoh0TNugPh9WjkjTLGEqWzjwfhBnXSaMDOF
okwFKnVQ+7eUohZVBLaP0Ww2GdlgW2afQz+2ybVMtc2Dlc0AbDtod0kWSFK5HNUURJFr62M9jQCv
Nkng0zxh9UYrOlVyFcK5c4O49DxZgbRoh7mVWhYfOarRtRcueMjHe997lvNh2ucLPVOayUv4XPjb
9HuWRgj8FjVexpAePofTg+oUC9BnHGBEdO1iNDXMojvSGVo4QNP8rdvTIl8M/AMGhNH7nDUbo0qK
T13u+3Tv8S/0hWgaAzzufY5KR6lAzPPARk7iXGf0tg0kvNX8j0F9JxBfzkhhYR0mE4FYKwFdAyjl
EMDYosqy4Lty++UIKk7fjLc2fT3t615qJuRMQFF7M+sFEPhVulWkRfOssImSKpEBeHUSZcYU7Tda
T/lWAM2UyWaRl3dctGTRiudztSbTjYH5Za6C128Uko2pDRAOP5fWYgNSh7jZvSaUF6PqgAPQ2cQg
PWf+2bIoX1jn6O7ms1QDfLqLoye/jYZUt+51ZclJDrAx1+mv7UxqKdPcd9c7uzenykJZLThO6T0K
OeWYqOaOl6zUj/fdLbPjvcYn+EfI+7KGh6pjw8eOcVn3d5zJd50E0xS4I+GHwDmsbrSJO9sYlXvw
1ts2szTOnMgybDQDMLwURUr1PVB73SY0JI4BOuZYHbwAl11GW8OGNULb5utWRlp7Z3jVn97hupBr
jONCdYueNd5M3CYrWY924U0R8Fr4IK5QMvdOWbRdoKOyLB57Lt0QTe7XeEQvL+6xD/Xn+dTOKzAD
Bh2CYx8yMeN4XUwGrG6QzFcwR5NVs56LKXI1TxTL1ud58FqHJNoTFlwRSiENvc/uha+37M61VawN
cs8wskjC3DJPm59T1MO+yhqEyQShg1U5aloXvzhJZJoIc8hN6qQdv2wbCLgYmpQ/R2LqfmgGnpf4
RaFJMu5eAN9iItUzWU+seY+3TpWScLNbqfZVRPP+1Qxlu76nYuMxJHpMH5Rij1OgP6wtfrCbmJhl
Gz3trWTcKSy9FUf9FcWK7zcXrvEjeg70PxmRSnnstxz6uRDZL90/S9tzh2b+ALq/UvhNcJxFqopr
crgd2lUBoveYZOhN14j3DRWpO9+pPpAEnZqhemzspbCwUcj/w9XGV/U3oSn1dBuSBAK6EN69oM1m
nHz8sUxzcOzTzlYZO1TwoYiHj9ZFVLdJabGQpWSI9zm53vk19bXxhLQb2VquAGoDOFLmGFtLwICF
VqLrpThhhQZxokDxFmU4JhaXIWmDudY85LalWMMN0f83x+yGKk3hQBk2sqEhNyxJ8gIFL62xQd5U
6FucBIEQ11JdorI1i2y0g/aG8apYEZBy/DGE7q1cECL1ljDnpAcb66AdUaEhkGwJq8V9RLSaRq4F
i/p3Wj9T9nzFDQSndMPxOkLP43g6SuWvpMfoy85nj3f0muujWElneojgr8NKChFYq+/epsqGW1un
OnKsOtC4va047XOuntY4b1RJiostT9tDfvuy/Qm/H55LcWj/ZKJnIYBxY19d2OeqPbf9GKO0wz44
XE5Ocx/f+d+lLCEmFyv0u4ski5LPZdKAXb7jR36vjro7P++S7FKD261vMIRwJ8Wiv8UBG5MZ4emk
wVPOAXHhfCCilXnujCKfqC8JaeUwN+3tCvThpRAmaQ0LNYJqUiwRDOo/cNQEiBoMEiqu7nusPhLq
2gjmPGxD8JtaVjcUNTvwYfugAvb0XGGouwRabWcsI8V+S11BLH06fkoHIciwwo4m3wOTJ5b2FodW
mvrBSpRsiYioJsd4s53CGQK1Z+nyPk2w4bO2aSicxD0WW5O9oOGtmNYXIbmqk740TkDZ3+7lyElM
VYNsrSDw+5U7rDrGlDNQNr2b5cIirMMq7MCaCiuWKgFeE/u+mnoiS1DF3KJOLOQEg40hNnTAJ941
8oLkNqD6GtL4/r1IlkSvpLLukRVLLrnMhFLavg+BK42fhYpr4jwX5qvRTrQKm76MEKEA5LnlIzfK
izm4+Iz5AEbFbmH14silOXM+V7Ro2Sg+a8aHTCrWza1rNVKe/5OG0Ld2PxOZyoVBqBk87lQbJix0
IHM5cpZ6QKpCqhbA12SpaRoiS3K9+sKn58KV0+oGDyA/xnC42Tb1XIJTzcgaDZFGhTo5i1uK+oL+
vSDjdmVFJso9qaz2jkoKPpXnwlmLiPEX+RxBcm4J7SgaWBP9l0/nF41T6iX5GtmCT+nYVawlwhPY
ikY+HfukgRCk8Iwhm3LgO5KPbHg44wBMLaIiHT825cC2V7kbWqkZo7a4kIeXGaSQb6pJplbJOm6I
Conf5yCgosKZzDA0omjNfTj1OriHDR/l2R9PkIjXqbdG3M7wgKSpm3t60HZlEO+OigrII7FW4wNU
prJRkGNr4CuMm5ohZBza0cXTHq8kkrTsGgW7SqdV4dmxrUzC6aMqYiunQJhRaIYnhK+hB18CYHkI
YDxrECarsMo/f9HbFoYaZ6ZurGnUdBrZk3jjx57MR9nJlIp7OQZeZWSvHtwQxIk+fb3ZaW+Ya4b/
fYCBDwisdvUnEvMy/qA55tU20oRcx7d3S2R2u2tIAH6bXUAw2ECM8fe9gwtpMwkRPGMBrgqfkS7Y
+r+ngm9IpNpw2vWmsugaypbDWjr90/hjOJNwOdaZqM2t9gmkhGKB/B/x4dfUiN/EqFPgHwRCxVIu
4U/9QEbrkepLM1/AMgZrCcw5PuplWq+E8DGyc7nIXSDmp9y0xYMy/bCiARMgP8VUl9CeML4/toMH
XTVD08E3SkpzNb6ctVV5vZoyS0Gh2R+87zGj7FvOJow2OiMD0gKt7tv8Jy6Sbb/E7Osl37teg9Mj
2GoTd3MXu/Yz2YOEoQFqt8COuQiJlwjxr/GMZK42Lg2s1KlsrAj21w/P2PgZLSy3SlQ2v9cby7XK
uHsI0KwNX2V3MLdK3AYRe40JNvyT8mUpC7XtyZA+giH8ujGDObPZRBObrCyoimka9Scy8xXERL7L
ShGUbX2LomS836HKBLrAuFDhnA2WKuRHTV/dzWu0AVPCoE89wQzlgpt2iUyS1zztwOJoDdty1WBq
Wo7ygjJD4Cp2yAteWcTS3McgYPuhToWpxQOxIPR+3aSWtEeSUc10uG2gAPdWRM+eAHVtdA4wNO7H
dt2JuomVQTtRMmJOg7HkVQWJfLZBT4n5Udw+4UvDqJZfvuybxSOJXRTQh2THmCc5ji0PA8pDAgyD
beQ05b3oUurhWm3e5Crqt7RM0rPZyHiYv49v8TH1Uerk5I2UY7qnbUTSrJtuKeTZahEHIPRYbXSS
ZmTwcp3W2upSAihNtDKRRweZavtL3sDOGgoifdvHacLhy/1klhHWw4UFAtgcYHUoxyyGJVjMfP5H
JZXrELGgmm7jIpgezXRLJvhwZqvFA+KT4tg9n2G4nHpCfaBoVTRw6gF3frSV7J+k5xuUSmLX5mfB
59uGQJFWKyAG7PJ6U4gm+4sYFyuBhvKlVjxlyyyBuUvKNO+vRPCqZ5Nt2kosMM8eSUKOXl6rE+tH
cPXvLdmgnvbf6nhsAnF6ERswx2ddRsdpHsu9mYVuu1URXKY33Hzk94lz4SZCBFwwpwMnRAFOgyH+
0z4mBFA3IJ/5/NgkIsDdRKoSFIyhgQy3aeKby9MwnoeEYbZPLYHQ10pSLM0yUHHDT0OkIWGjCKlM
riEl6sqMPSlwycl8/dKw0cCfwkKRDQ18y7wkRLVZKrzE4Kl/xEZrWz4RITf9D3DQGXOthX2aJ68E
70Ji4KzmhPHJrvPOJH9mduTcICC8AJAHXqCHYb1sSuSjnqqY8QraJqhd3JsKjYXoFI7JSzmnEiQq
auXMzN6NWcWdkx6QEYL1WUnl1QfKbmPWGPBMADFZ4Z21omGJDVrESKMeu7N12C8LKti1BxkrjxEn
JoBTv1KO7GwjsPbUyOjnk4kWUQDHo4sduwwLZD8S6B26Czb47ks6LMCZcKd1UcVfHtC3Uyyt0UFn
wp6Z2eu2p2y9njKS5ufaBoTP2i91BfKZmDelnxeeEklGOT7KIcmVhQOW6zogid5YTm+DEuLLW/uF
6fA9K6Muzj4S3Qr4nFk1ejGBhQxgjO1sjLtOwll2Ft0uygvNM5YISrLDq3MpHmIfL29tV3ASTE6n
hXH0kgL4xhOX7P7cXbPiXflhfS/W1cVSyOMkHCCf4OyhXf9AsoDaXuxJTQqOFN8t7SNx8foD0pdb
dmAdOJ7mrDtKkO8S6s9x1U35rsys1KwWrepGnP3N7br4TJptpAUXpZPeAoPOCqjvztnIXANWl+dL
n3ua5LPZV1MHxRpDU6fIhtZYy2nnu0GouL6iyERtwYJPZDvFmnjdNyvlAmADjFpn2ql4lU+H8WDg
mFi0FrnNml9Km+05GuAn9DxuOVtUwnDftOQnOday9RJZeTlViznG0AEXkmdPYuAn8aN62Q477yW4
7luR9qPR38WF3Zf6zs0t1px4IvZX9GRGrXKcPjHUzXNPSKeWyfFA3Fxe5o2RjbzSAcLBgvuh54od
vd6wca/5B3xaXxLPSFQ1e3UkdAZN3JEvt8DD3bPVLQVswFBTC5+t/N3nuiBH84KVfl8Z2prsSstR
lfV/GyllcpwujJatdeIFz+NbOWEi8pmh0NAH7K6pFg6aRztlGHwqkStgWG3L6xHYAjovGM8JDubq
X3RUZCWS8C0qQMSlcbau4kGmBAfuVG1ioM0z/bNoStPAUcr2Ezj8i6jhGw8wvCXB8beXLt5w3vH0
PqBuqydo3okVXSu/jM2WkUc+XI9ohpMGD9dcyjpeBr61JS9geyXEPWOafecsiMMhl3r52mPj1n/m
0jPM8iehgZotV0SS7xRFRa3jgJo5nlnR6T2uQejJd9kwqrK9JubfoTzw+XoWQz2lxVSy1WOQWYfG
cK+TzOCGUEDo8y/Rtr5dGAzDoCCVjXxQKzSjN3IcZV9hCIe5p372TmbDJSnnUQyEwxdBLi0RCZFh
udV1D9eqH4pEDJdGIUhmSIaWt1nk4ftr/7h17as5pNl3orIkd/T4aC8/Cz3TvbfAMvx76waKLuHv
DX1tapr4bA4SGautMbQLeJjGp15xA7siFo0NNvszAaLtXCAh2WLDo374U886OwRBTT5uFkgnF2d2
ge+3A85mR8Xq0/m/fwYT40l6ZwQLPW9JSQUB1M+oE1f1KmerXqRBmbsexWynhtICSJdZFoHhOQnV
+Nt/OcOG3dbPHIsJIGTykMRSpe61l8VNvkwgdtUnSJvfctOHAVsKxh3EFmuUn6CxrQXPKfcGHLIf
03Lm1w0YQK1yY9IuMayLUjb97fd41fYgf3Hy1XvkwX7t45ZtSPNZdsf8GKL/8xsjd1Zb5mseFVqC
BUr0VeCE/JWx5HGmef4AnizFik8F+wsUum6MG3vjCBz5SlMGFHtA6sNdXWpBdXXcChdkUr3U55VJ
fHLD8TK4oPiwLA6s1mUckNt16QdNFXyKbxs3/FUEg/K8a/nSw0RS3Ov432dievlJV3Z56LdSdIDx
msiIE0xIRVJKJSB+aKQQH4Xmy59w0trCZJ1Xe7M+36FzP1F/yW+NrGcn1gCspsjMJTMziJ5a37Az
kTVv3oobwtHCkTvaorYEN6CvFnYvahrsF3Dbel+xtHCBxPugDqJlKLgN7akMLcXWA9bJ2mltcWoQ
VI64iUSCkOW5/OmKbc+z5Bxz0MhQpqfi03KCVvJqGSGvmVwOx9oNV2tvO98sNcS6Z66na42pI8a1
whaSAZyuTA+6FhBhws4ci3zJ4Zccuq0XreVXa81w1Mv9HNi1phTOtGg8J39RyHd249nKAtPPNUon
BOmKxdVs/OxeGWKjQvJc2cxvNbUOu/6Drma5iI3yMsHt2DAtMFGlGVU6GjAoCBS97Rp77AUXR/MB
cLLzepG+vY47JTM1Iv50rGWNURZ3+e4dFqNaAe7y3URa/NtcJoxJYqDemJPVmsfzdbOJpQ7X2ik8
2ipPhvH8pOjiufzCBBdbTXVoPZ7cgfTFgi7l8ud6rUT7MqUoGvqgLUbNxDxx8NRSyGQoyGcvsQUj
GtLGAQSu1UY3TY9i/VEf5xJUXrGe0SaxROnOWq5MpcKl6ciCzOd7AGb1OBtoW/hLtonAHVUIk1um
E8NAC5B1Tq2tlzlVmYV1ErYFVr8Qeb39TWETw3msMlnZnCEJBaQZaade/+dRTyXqIHxcBGK8UFpH
LBj4AF1qTFgREq4ew3O5urQsPosQCQexa8xM22qaxG/tZY+rFbkPpQ+WOmH9ZBBllFMWLEggTZz2
sPUwc5Ut/mNFbiQSkGqYBx50Vcam21Pnt+3X7j+21Vs6sXfwcYpLqsePmOe4o0Jhlqq2K3kBLhcL
g84iW2tjSkcj3YMLvjCmlVo0/S7iGnLBUtCbPIOiCdTWnKh4XQEHZGlofoLgIZDzLCwM/lP1fzWW
YNRbv5+8q0DR8g5RwjdBzaTlDt6gW3iVN3VrG4GdkcuN97f483uvr6+P3Cjbi3w6CU60ZfpE2qd9
8XBAKhMDOyfV1/KXTKHCWeGwQl/PJiDXq9DLftExIUv1N9DW7xzXAzYg8e6SzHQCffa2jdtk3EzY
xyEwwJ0njt5MDAinpxtDQoHe/ioc+IUjwlH9eL63Wx1+JskQPNp0WOWlaVMngB9cJ5v/7Nc7jQNr
dDUklPk8qtF4HFOHJx38OuornDPLizZuAi201lBRODrQP6WWcYz7cXtuJI6mKepb3qPJ3t4vHqRq
DMYpF8mNP84rbC90F+AUrgzhZhcVxGEmiONMHwkEW7COf3y1s7yyqdu5CJcJ47dTAYJf73qmacfT
mbM99BQewJLewGKDuznl23lRRrUoaNHHhkes9ZF6R6T9XWn1VRk/aR+rAjFGdBKhpcxnrYL9NNgW
w68MSy6Z/PHUAd68JXE2T07Syaxm3Lr9X+jCrrHwVwYDFffg2BmmFl/rsse6vqWc0xJqxIkZrScn
ts7Q0TM5ccCS6Hf+QAkAJJxKO1Yb+98/37dMFqD9azMJoxgzeUQrAYN7rDWr0gipkNSuGp2/LMzW
YaQBK6uH10ue4k+tQS2QVKGVCQYui0+N5Ot0uSg0iMoBvgk+J0CbOKHktEXm9H177MTZeJnnzILz
Pp5iDPVtBBoC/aqdzI2vEogrfahvfi38fb3yOP8Ycc9fpi4vfe4b15Mu0aVTI43VXkYWRQhHKM31
v9pmlC85h+k5n5qeFsRaL7goEsAg/rDjI5feUj62Z5aWIu6uHslO+u0tePtEkwiuW10xGJBHy14w
4RvAxR0mfCusCwXipm5viiRUN2GH4YeO9srXORvD3OpskXOAOQHLxTEfFVXIeIXFACsE5eCi3b9G
D8ZBBj1ccFnlMoDCieQnpehDJoWgUO7AvcecqoZBYL7dSJS+uPZvSp69aAR+52lLBKKiHEwhjX41
uYi7GhZq8G6uPVPo+VtBjxGw/JV2kfwgfvuV+3O8A90T6ebADZiclStE2LEfEZIBBVmLLjePp067
UzEARPW0KljDhLLyH1wqAcVoSMPo2/yTfVILml4AzBonor54BEacTLyGjX0UKbYmr0/fTeBNUQ5y
DzV3oNygcK/Q1SK/ncb04IS5AQ5qfqWHChpgAuesnPaknKB2eKGtJh8KITV6Zy1vjHCgw4CmOnBb
A1vl9E2q+5ZnGUYaEPflp1W9NNLuVdGXQZXYSWVjbrEYJHCfLmhj9gQ7rn1MymrPoXreJ2nlTAe2
1KHDPNP0OqJpNZ3rTtST1clInwjFg2ERAoGZ85OZoMtRwqatMUbM4z2xSYsrwQGZK5t1wPMmtPvG
szVYh3pzIouD0nPhMyVMQ86kGm9FsQBk5dyFL9jJKyu17dRyI7iomllEeJ+111pS7sXOeAKoyBTr
+MIqh3QTa+xIRjv/BDY5OFnoMB6OIPWzqhAXur6ieUBTs9GwhaQeV6xFOJhwpyx+UYZ0E3s97PfO
tuuDn78u4QQc33u//FdrZwswjtk92ceYF8R03DTf7soICGksZaI95ghRdVznVhU3MT//bE6U+3hd
EfDWypf/BB1FtYTLJBMy+E992VDU47ftsNTuqFN70QV4awIs/ykMTrnLHqePSGqZYoLYJ+s2dqto
R0KfwFLJaSxPde4eHYA3WaHGap7FFHAU+3k/qyOQ6aI35MmVJuTNYh7/QVyizizKnP6vPhDWnhMm
N7xCGDJSXJgH1Vwt+RQBVcZb63GIrF/uhwPba39BXhODdpNchS0yQ0f4l9ShNl44mWtxAadYR2sO
PytyiUJWXIOlMWLLy51nip1HsqniQkEzD0QZkmmERX8uD/bm0t0ttWCWJGfnQL22G3y8VfV25MUK
M81kmvbynMSnduJ93Jgus2iASlzKX3VfMa9iQs3xcIn2PYDW50EjHntyhBTn9xW27hry55ffGBxD
ZglW1BP3aAUNGi6oqrbNgF4Pj2L/N/KoePWdhICwaaW5ZhwG03B52roemOiZlXnQOhu+fCsf1b7E
XOc2aZhwxMTeJ9z6zRFOYxcsoR7ostX2LKaZ5X5ijk1O+PCnFceczhtIbBnSxybHAbivUUDNElrw
8uxf8VE5hG7/teiclPQORxN1EqISw6L/C/c6Lmvz5nctQOKlMDMUBHEyl8RxKEryaPiyoCMR9t0d
XrndZBj2cc4PwuJzlCCl6kMtYQC+k7OFdA6wSYAVNk7dvzTZ++AuQ2MepAnWBOGfYDtreBDkLbPk
3Ay41V+exO7ZJMruwRy7BCOGvL/if8U2pHKt/mbkpVhzQJ/Q0BwkaGYZzFzZuILM2CTWBhnyU2UO
sdbfF2dfJz666VKNW4Pw3zNRssXcy65HaVCcxjCEZT5GxsPz+7I1s/dSi2rUbMdU8zFq/27Mdh0j
PzPoDQXM/V74QXYdyVk7zww2AF7TSv0j8DjEcCd8NWTB8CJZu9DNtqW7HPY8i0MgTp4aKzxvOCzb
Q+Jgsbxgl29IjJL430ajKIDtDyU47+u7FPMDFxZqGzzh29u6GtMDgt7uOzheZuFPT+nhJ514RnmJ
R9YGanfynVgXbI5kwohVr3ODwBLr9ki431nBfPSc48DvKdwxORTpswzjRBDJ46iTXSG4I/6U6slA
yXKOZRN6YenBjIhV7sv+64B4MwSFoDJFz1797tb5UqRHGJ1o91IlHcVRrnyTCtTJHXSxONgsFtEQ
/YANB3j4OM1Eq2IK9rETxbfl2kIP9cl1ZhSj5W2IA+Dd8OZYrbNFeA4jck5aOKWoM3Y25ZNO3gOO
iXkMi2IjnQIwZJkns2sqxD9y+kYeahwUrGi5v0yr6TClYwyageadThu9ZhqXZQlQj9XTAdvUm6Qi
AzvvN12DNk2plK+37dioJFsO+f7avWxIWiHk0KoOu7QSXSn0aGd9Sp/YNqSPy6Grf/9WMx9naMdY
5XdmWli5P6h0qmPiTsLRSmPsG6cZyyQ5vTb2HHCiu1hgKSQXDnlSrWDxW0XIsa1iL55Armfirykg
DbmvQTz+6poB+2GU1j7gaN/dCj5eOV2CxLmuPK2rcv0qqi81wZi0xUF2g61osX2u/Avg5Cf/hutX
ayp0afKN8SAgLJreGksVX6EGg9b25P+zKEE/xWph4zo8RrBzhoqDIjKPjlyDiHddci5TzUFsYyYg
DsahAAAn75VjfiEbd5ttQ8xjt6rkMCzqxs3LO5C+OoMmpmRP6ud62/1sK57J+B26IDvK+fxSmquU
0QAowyyUOpcQ1+gpWJOVEaSOULidSQcZ67YAQVCIrCEekoGZ5C4KXBLEF5dYafj6kfwRlhcsGFcj
XGvNqSC7hz+/wlK63+WrNxXOE9kuUOJi6u8FKcS9hkxXX6Eu8KdCaljzTHUsYWwGR59yoxN4xLEA
Kh+MQm4IveA9Xg+vmaE+AOdUcKG2Ap8VB5CJ6lVFbS1dbvi5sUnME6XiH3tjQGVwXP+VXn2gPHSH
fytxjtT132K2JHLOwVQfLzY9HMX+YJc33nUjVrGhIlLFWue9R/exfMt7nm4ljc20IKDFm6epc8i/
WcXDwjE7DHAqnJ5BJXSPFpx3a7OLGJgl2pAfFL+v6Lk9htw0D9S0XT5PPL+Z1sP5XoQWf+81IFlR
nVUavXPeMvTzoouQev0w9zttrOBnWkqJKqTSp8ERy0djZbBcDneXc7wbGggP9ulM2qMdPmJNs2kr
nr1Druz2YrOIrbcZCwgsviKNNy/qu7KJpa5pW0U/qCml2ENwdrnHWVVXtaaPF0f0YytAdeb28cv1
PbMJvJA0VmxmUDsIjkyZhrytTXEIBTyczES2f+PqNv9aKtN/Rn5z2CAolXQYE/ZhIqq0xcsfBmZx
CdZ0ReuedxLj7p5/2QHODgG/GY64ClwuxQOQZ6RyObZIXjUBrl+4RuhxN7m+FIGwg3rRPdshxEF4
oL/mYCMlgz6Qw6NjK+0RCPm5a8wKbE/jke4ZnVxF+Y5k+6wZDnGA78qSU34VNwYiRjYfcxh7u6dq
OBte5Ic1U2M7XJlsM4uU0at4d3FONSHgtVZCt4+LLztOZgYYvqir99dceMCEYSzMV9dAElCzM5ON
mHQTsu+VNCdCfwC5ZLmxWCzQsPoRZBRWCZbbK3P/5U2/FjjRVnCS9Nkk8X6/PIpK+nwzNjrKW0wk
je1+CWto7BiYBEZAon1q6MUr4SQHI7JzdBgIdNo8twOK55dvJj7GI0mbKJpLLMdBMROyJCoymBGP
PiEb3loZYePtXCIl4XfLPlXfLApwFf22aFvY7NlLD1capKrep0kBnDkZQWC7uVaku4zBXmtDOjNq
viGyiT7WaCEk07cNaYUAyNTNJM38+r1YifFKlMuWBTRRiO/5cepDZbFwjzLjFCiJgWoB7nwLTVas
z+M1zjw7FMboviwluzpJ7+kPNZ0OJgY8MDobJR/XSlTT0ngua/nZAFspwCfyNTuaEAFXF69Ry8aM
/DB6vb/MHc/A3nvxnuqROiT1XrY6/GAnBd26iJ758DaRqgZ6a3KgTFWWIjU/xE+q7MunulvqWJzW
yDkufV4w68WNuDP6TS9UUBgYr2dht0qqO4l69ZUF6Ww21jj7LXNiMgDg7XN2VPHyQ0nYiPqN3Et7
x9rgvjo3+CM4vkm6e1ipGiY5kEYhsthUAxLi+9kC219f6FEJAPzt04U1cXlUxgvND1ODIzH+CAFr
87RnXaz+BESxIb8HhpErxIcRRTmyEWm7zsztnOVz8ZpRKxe6ZY+B/IW4rk4Mejy/ghkNZORQNSVo
2TsKe1N3Y7qhnQzhnhkiWhyIDVTwC1JhhKeX89wuDvyKXecCHoiiByr38K40k1EpQNm5n1BOIx+C
fgKVSkKWs6wU7M7NAZXyUo2yRBCH1muCapfRbX6SQsvuG6mHzXKh5smf2BQVsd29hpAZRANiW6Ge
NqB3sfFFJI4Br1ccl+lmZle9OHj5CMU7P967AePXsuSKrWx7iHW4PD9Y71eX0A3/Yg0aWsoFiMO6
cT0i4ggR69X3V6NJ4R6ap9H9DQgdcBUjDd4axC+9n7Vjpc4IvrFegUUViRngOoKjQOgqAey2pKqq
aMD/5hncPzBPjykux98cClTsBsM+GGVWIN+sw5YMTPSplwe6oJQLY/0b7Bd8l9kITJssZmArZUvF
YoO8yDADTPwptn7Pwpk2Qugew0N6V5DLUgOROo2+hxAGV6rF/YuYpev7aCoxT3bmxW5eSw9jOuq/
hRv19bZBtigZyyCC72mNLeqF02yWq5gOcdPbs2SqOJ1vwRq9zXcRZM+vS3mqTODZNBCqi6iZM1h3
0qhBfAl3dCWB3Noozc18RdovULWywnH4BsnRqRQ9CktSfxnsFdYXUnD/vngFprH7RJJW+weXJ9/e
ladPBpZIeONwf6ITCBUu9Rxyb4gDPlPxJsNGvPs+RNBqzVlCmJXEipGo9rteO7yAXY7+HmKbXB4S
Qqelb77D61xZ3nm4LIau40u+hZT8t3KbQxNKwqwjAAo/EirsyCvzXY1SSKLBs9wlROJU3AjR3Gp4
1IGllnQj+E1fqgLsEPJYppbudCQVCbx5PQEHc3/btYj8j5/dmp2KxJH8DeXMfm1yMw3w04WoejXf
0e5D2IFltfusEynmJuZa1/0AVKDPBAtQsCQv0Ml9kE+IKjZkLjyN43mxmzYIcl3Drl+uJp3drWfw
rtC3/jwe7m32+NHtUVnSSYjEtOtvlPHMCRiNALcpe0NEd93R3LInqxcDxPPlu6YGlUwyjuO5YaYn
B1HQdKbXxa+nGNjDzxaafUhhdzjhrI+B7Im7F7MlU+zWbQJnZu1htz4IpH+1yO7cA/T0ICCOB/MU
99B/6LgfVvQJ4eegrmjR35PseyBOhppkkLiEQ8Rsd1MM/PkHgro1RHbRZTBYgOMfLHld2qznhlxw
6bc9BA0OSLt/Yd8Gfn/WH/pXdcN5IsLqmSMVFquYtJs/qcdQVR7nTO2H8XDd6UAkErg8WT9YRqL9
g7uSsrkP+IAo59GgepW6xoMv0N9d5J2wcrQweQ+pQLRyDnmqkzFr9iU9ugZ32yOkmS6Q2IeGG4JY
vqQP7bFyLMUCKM7wWJMRyDmIedFfPguhuVHCCWYUEXaBBuoMjUJudnHP9Jrq+WSUcQBzE7y/9C7g
klXCiskTBWFWuanwodjnUmxJMEpfkuBhazdjkdv6o/z+B0Eygrvi/Z4/JSoHBWQGqKidhLHEBtWe
0k95jS6Pwj7weNpMnEkHi9WoX22Noqnrv93Z/s3QMa9nYJNQsZN7JPtuW0g7+PjN0Qlt7jvX0ohz
Vb9M7r1gkDYUq/gUJSX5UgRojlJ1X6tCAUV8rOaCKMTbtxyEwjL2VL8rdlbWk2pvpmwgHsX41QGU
S8JtcQDb9I+dfKFiMwvmsGl3PXDQ17hs1n0GCAHAua4M+oVvP1GMsVViB2OLiyL8ADO9bdEEkMIl
+fGJFkkhhS50PdsYTHL1ytiaTk8TrIG0rfFfinDvi5JlBpfJCaiYVmY9d5QpJhWs+1LaB/5iJUl+
+uEZ7MYDi/M9Z3QipYKlxNBNEN5zX1YlRrOtYvGL+dr195DN52h6tuaGwdqjGJXPvy6Uj3Rz7hX4
H3b42/sf/mIyOR8f+uQXg/OkkDlFfU1SnpahCIGJx2nb6A9tqYhIbPV5DTqosGfowm6DdLHnFTKz
5a/yq1vX97g0MT/IlHCAtweoXGvz70Mk3RY2LYMUB4Q+1FkJ1ul2iz20aMsWkwNEgH5CBQZZb13j
7R5vaibXLulc0y5Nd7fj+a5yFHwvVqgT4nCD4Eh9GK1TKayhuu0eagRM2My/QI7iOI1Oc+KnmbLQ
Oq+6eOXVEnq8nHyRdv0PovLV/TRxCnHAU+CKjzYPBkT3hGWOldZ1s37eDqMlAl04rPAhPL2wHkNL
vkC06Zv+jFhMuhXxEPX9c1rBf9ThcFqq7YpULJL2WZjm8fKJ+Q71QCCpg4Wv+en/pj2Azqc38Dk6
SJfQwg3JzFUuSXtO3KCpfBuJW/piTCpNV+XXjZjrAtOm8g0fSrnRo1QqGa0U/k8KpxzpUF1G3Bp1
BmAOW47ytjJ6R3Du9zhMUqlXqLvLNmIQ0lbvynyLagg/ik+ckDw6/2nNWRsFvnBNfd4vzVLLj810
Mt8JnzkluesASNa7IRZQneNnBoDBmgvbwB3zkqH1zn4Ta24u+HFsa9C9PCMEAkfceWXyKp9Xuvr+
ksoJMYoc07URUBQlOeNMLR2cjBOotba6DhHtwwG6IhU/VJJuSTSOr37hoSmo9Ud473vcdBtoIUC0
Fv6SKR10phmTucx2nRJyR5AdLXes7z943XR7+QEXiomyU2/J2Na6RNjR77t3YyGAC0L68BRZR+oQ
EvWu9uoxH9J+cY+/ifnQkqxB9rRRRV+5xVeSg6YrCVjQgjOOzIs5h8WMptuqolYPC/NtGbHcqlFa
dEvfkfepih3L2negZmAgCWGLXxqCcdlohfNGjGHApHJW1pTsxRXGa6UOzQYQfbWFf5Hfyw2kBYYO
QeREDnCeIgpEs3ylv74HRakfHDfWFcpUOk9P6alRnfMmKvAAHujk0oJU9EmgsF7FD7acgxpnPB3p
QCWIgomoB3YoABcFUfS/tGoqVo69ehA7w7/xtTjRheSLb/bo3/9k0YmF0kECbFmFpYQodf9sylHE
kU5MNcrINCaohoWSdIISj7CCNqpxsKVUBRLAKLw9dHizr/w1cbhwKhvjEfnVpZ8WzpjUv7Wu2Vnz
ztOuBH1yTMgAJgQXRd4Xc4/zXTaS6h/pdjRdgS8qZ3NOZ+H2hmv5dyzglD0mWoCdqNYQMj8qPcZz
qIWDn+6Aaq52Fz/I/uLs54rAuGreHkgfOLPbvGPfIHkiOPWylyxpQeRY46k7ioBKz+nifs3mdHkA
w0mn4P9GgVwKbr1tfZ9dcZH2hGefS/WRsRFRUhfJLBye94AhhemJkBLxjDQjFa+wCafasmN1S252
mOSH/P3sj37UiSXbLeZ4q+ZK8GxEEjSzM70sEOtfT1uNJvR+Jo/1nR4/h/qjAj1G6ZC0sF4azIpV
dz3/9c3TJJ9D7VZStuIk3EAsjxxSIn9WxWvNn5hmTc/nEf3PCFoJuzVBIdc7Y+ZHt2XbHpI87gjZ
PpTe+bJ+z4WoIfed0r+PhhGIZh+ypavKlGaT9EOodzZfx82VYDP23bEJSm0P7TdDoAFRtQb9ZCw7
VpxHXoGkQIaCyhdkS1RzGWLWE8N3yKxPqsXYxrTX37MX8KyT/FKVHAxDzoTvg6LC1RgoSzUKuuvt
n/iKwvMmxKgqFztIQ+mJYxvLEHhp4Uy10DeAaG3rxdLeSmMlOeRFOMIosN1ss8IzCeWaBsOFlzsa
4h0Z+SKU1kCabJjdhVHSUvsHBz1/dCuNpAZyxMsB3QLAh5F0O9Gzcjnunh5FFCry2p4relTTUOaA
hJ2JaTYIaRG6kGPAoGzg7RFIuZkpqbu09TVgQZztGWIFhvEOgmruYjlaAqXaPx9kxaZfTo5BclyP
s4h/aLysq7xTrYQnoOcm73nnjCWiMvzgxTPMKKxOOBfQq7lJgGSrolouqWTIkCed50wG2TKnnUc/
MKyHxiAmR219XScL9bZypL9xRWWVHbZA1St+a294HZZDYXIQ0phphc3OWQOm3cRqlxuO6Q6J0cKA
aKO2Xsr1U0uhNcleHIuOqCMevLXnTHfrKQaQigHb8o9negK54K2UfxvIOMewCF53CPyuLbL+Juis
QbhWqFHqSsnCclNse9HK9aYa0AL6gZjDsrOZ91PUj5mxFG9McQbpuZSdzpKD+HDFhW+LuffD/IPI
5N1dMamBUDdGIlu6BKpcSfo2DZbp8EunnwF19ir/0F1gJJfsLEROCOUr9pPV6mihuIwOwaWCHFG9
yp4ar5p2/R57Ra7e2MAPVtPAK7+C6LHh3+c2b4PrqudgHaBt95qiegPU47vj8Ir+f1bPIXkAkM1j
tlbWGFskvEn9N4m04XaT2bUgwzuRo7eyzpj5V6AzVvq4Xaoz9QP3XvCInY7Jj7JJxRTwFJMx8HEI
dd+EwBofmpDk57BqvLKqxSzS9UVOu6FvElSO+OP2YjXbUfMwAClUImJnoWgATkjBmCEj9uYkEeZ5
g89RD6Wqk7uSb36cZ8iTre/OdLE4el6Q/rY7uS2tWuyRYmE2usQysBctlYdWaXcZIEQoa8Hbzxwr
23jZ7AkoOm+HOoYn//Gy1B+MtgudDf/ZX1PrmXIOXncWt538Jl4OYt7sz+Mm/Ud6dxA6AF5bVLxN
xNr6ZwpJDxRwvSdBYs7yDzLzEmPXwgvEHGcWj/yamd8UGyb3eOexxOsO1PPsYCPykTKI9/LKdc0o
KvLZlxoGMTBlIktcrfgWoyDXSTjYvEVRhDO+/PqwoeRwi6JNZ4++/iqHCLdF/GVH58ddPBJN8Qyb
nx8NceUpYqAAN8xY3qZvKuK/dUAOCwMA51/WgUeEOgOQfG5pTzK66JAeB+kUtiOmpcBnS+ww5/E6
ba47UygLz55XB/xZKV7CGB/q+F1rbC7/z2xU0vtt0BMmH9wsQL7sOqC8SFY3fTTMZbbVnJx3mva3
/oTa6bUx7dOnaMBWAgz2F6X367aVn6jzMBkRqyTUpdKwFCEau3NO1xaZ8lgNDohSV7mrOcS7MbpD
m6qkNFEO8/E66MOXbwxYgDC9+veui5TDTvJEMOcBeGRBiHUW9gTFbrPKLdN41aZGFIS+qNbXr0uV
gpFnFofND3k/CW8HDNDkbIZSgWlU/lDliUr+G8RwIzWUSyc8Ay0xVpGI0Odfa2/q5gJTetuW9ULK
/+3pfakCBv431ninmYwFsL+lWZL4HWYNgHwUXqGm90+lMmwKKH+voz1Zf37TrU6W/ayvNFjSvJls
MpvTZyXhdnCV+oaqR0ATI5L8AbFgbYl99nhntwm0uRxQwQuUiv36D6Ue7yU6bnZLMYkuUwUkUFv2
Fea/E/n+ypTkIpmZ/i+9lyjS2bGiS0oZEbdE7RF2IJ91gHVZQne7WMlclLoeYQ3CMUazakCe5Au6
OX1sDYRHHaMho0M6ys0GvDY+m5b73/Aw7aNI/YAdSmy0R1yuCo7CyDkAi4u7S5yOXUjJjuLByODl
8JezIVyZITDj3G5/50xeFwAG7BK4NQZ/M535SqmOvtit1mf1IB3gYG4mOJ9XMDzExj26wl+tVoZp
EiNeXXEgFQA2yjkaNzj0tioRhJb6KppE2dY5jkGhTyLQBSQfXaEfEps72V3pfGvw613idDvaXpCf
11yAMAMGOo+5Bw/YONo9eVtL4xWW2x+v1IuizH8NXbdsf6E5YBOSg5Xv8w8Vq6qCIP5beSnfIiFb
jjHeahi23O2/s1WFbszf2rKZjtPto2VDVXANqX54FbqgOTnDf0eFv0exhlHTkAgn3GT98Lmi9afq
4HrORTeIw0ClQW14u52+F9+EBg3wiIItinrg05JQ9Q2yovfZFtGhnhVj3+dUTnYqUk6uqIY8EfsW
E+AOHN+hEEBVD9smnpY6YC12D0RUK0RuS2JPklSeL1yFgbrPJZguM0XyuK8W31rxIE/jugvrq6Nd
jFzpf+58XEQ0t6dClDR3INewG2JDUUIVC2ddS5R9tWyloIRVrpBPqqqWxkMBlNkdMA7CuXOvJAbE
hAoZKmjCHZjKYhkZG9xy0dYB7wftbluRuhDBoklhhF/bfkHUjpH7G5oybIuURrfBANc0AFwIqwyA
yB8LLMwKGcY3UEUSN8RmjtfKbga6O2lOwq8DECtdYDjPX6RYabz1fD2FwOFwoIpmZJwHqlMBTG/v
aTRmYrTbIJVPKzQWGTkZQFD9D1xtTH0EMMWhYZXdp+Yjn6CRVmVkG2VysD69lBlkA4x48+HpPy69
l83FXvinsPESQsD8de8lWKlAZv6e/n7ayNaV+AtNNCUB9jl30aZCMKAWlbfG7frxjyHFX8UWC0/A
pmHRzwS2z8jOMDYC6HcH3b8sFCxX85AMsGucef1eGjnyUpR9Fjn1aw83Gs6SJLJkJi0dtWFOP7Dp
qU5GSA89wpk/klHDN/dIlnEMvhezcaXJWwlVoHhGa/F+JFPMzVeu0/tRuf1KXxE8LCEw0DlZ4okk
E008vdamn7wVJ3ty33DNCKB4gddFObAY3qVpH3e8sm+huAe6TpvOOePUH7Vxonx4At9TO7mpmQlF
VpkzuwvoMJa+pFJiSyElTgv//7YZzBSmBcTxvdSTVeGWs9lJvxp6D8hrDgsocSlyabKLVshppaIg
c5EFkz11tFGXBeVOyMPAgXqZytwMVrhnS3z5ohKlE8+vVpCBfwzWfCMgwPsDctyli4h9IO73BNZN
8d+UG+xuOxQbCmc4C+tW05xNXz4E4sFuucleX/AU43BySHWej4LDXJpAr+DxMlfO1h924aE9AO0V
4oq2L43jiUFsLBLKR0nWpktwS4suUo2c4AnNHd/g5WPmQgSjd1aQoCvHMCsySuCFyPLb5a9KdMdc
Y1r3v8QNluTjgwkZ33zcWs051/AXL+jzkKSNxmxY2FsZbWqiEbnSHAy6fj2vZHaqQz8hne6/E7Ab
H0+oFsh0As+Roq5cmEXO9IPh16T1voOZmRJmgwksB4pZXSZGbU8d4cQb2iurMEjWwt0UJT4ceAD/
7sdOib4ArZsPMHlwUFNzKdPym7bHFUF6pt34ekgqmBl3oj+Ju+ulsiDjDluheL195w92oa2VN0Qn
3ClfFWZ8Rk0WfTZzGLKDk2Wd/nzq1S3tRsEjwY040n25FjA7ZUGeEmr3makFwvxephriRMlVnmYJ
VMhllDN/lS9OPgCGywKXJOfUBY9BRrcP5qnzCDwArNtJaFGedn2aX5LeE3yoCATCsRksiW8+xLoI
XpELmnVHMULe+EsfmKLfV1AgX4i9gEwmNwi3v0+gayxkHt1XH7Zqt79xUwotrpO0J1xtPBiob68L
iKuLJn86yAd6hq656lS9bgqWHDMkyfek42uTs4/yuAapLrnYHV5AHUKtEjQnW7IHbHpbELPrwDC/
oAHr/nqTnZKSeX1bJg2Zm4u/OiLnxbzj7qCkVxBJbEuKTESCWVuxve3Wg41NPQ7zFvH0IpqpATwf
90NWCy47Cm2yYli8cRg+A5Ib3nnyYaysG59CN2nnZQcl6sQsjiEP+jAspZVjzN5HhGT7Ews7zUDD
jBqxOE2s5pze+7R+Do0AQU1m6IiEOwm3XRUZN9j2j9y1J5AFANLHclM/2aJg+HECqXXJb2u45skT
O4P7eMqx1CRRqPJtvIQQNScdtL8K4MoKHCoaIU0DdMmkArshp8I6lOcfFSxlYSbmubdVuj2V93Jb
6JagoEN0VkxnB9NpGtpiUSoS6E3kz2R3NvrON4FPvg2cyrY04KRR6nGxWtukES7/lsDvN4O40f25
XIz+fDiORaiScI1WaPElBkYp9x4LWCXFQP+RrYmS9+AR9eiVsx31XLo2VLHuK9EAn4ycz9kfTFAs
vvNjYIKhR43zGeqomJ2lwFvDIpQ2CM7V//tbxES7/nMujq53+UzjKLqiBjFuBen5M2CdSiRx3f2S
18Lw2p8Xe1URTXV9hKY3bZpbQiE+wdiCexfNLfLflOWsesrpfZ26XM9Q1eJN9lq+QD7Wk736I2C4
VZrnfT0itEwo2O0rFmynHB6ey0lxaY16c48/bYkS2HZ7O3iqi6Jxaxu9ygJ7sXXhOs758K9hmBux
IJsz0BwHCOBd+hoajcVC0M4WkVqrchmH4rd1od7ZRP4njRAOVS/aFu2B7N25FvB4JnEXjtbYXLK2
Io+xiPjg5vzMqAclmKUdFIJxbZ1TYePjPvM9JZqEWSHxkPvnNhFSOaIBSgGdLJXDnETWlXSGOD26
l5ZhGKCvJKh6IN4VCrQRJdgTHtdB4WeVsE4WDgBYNP7FwNQcziAnyagLTOYLi/vJacVnDRh6W7gW
3DRIFhATeGn0gf7TDcCNdVLuWTXqEi4a14gX5inTXeURXFMTXun8bW6J918wQRLC6QsiCXhQEd/z
OdJUw24fYdS4X0VyZz3a0OxhMoPjKO3zUv06Vmb03+/IR4WrarfMwvtFpUBnKEhhDaKx91ZFnDaq
l1UiE+55CS1Z4DtiuylEq2sLug2kJYx1TfXkOhYD39z5djfhhw9VAEtN7MYg6NPvP1mocEq6r1ZB
1iyWpuDenuQRj69/EIFOjpsMVkkQupq2q3KyMk+KjOf+shYlAtnY9MBQBhgR53ktEieCFVBQBJ6R
MFDamOUYvcIE5v27vaiNpNTKcghuvGWVr3x2Zc/fDZ9Mn4Knc2Q7I8aFKUm2wTGhYPMoXsvEOu9q
DYrZVdBAvdwj5a0/ZLHme5KDEb7Tj8T5zM7TUxhrXVvhXWCBbLiTybEIz3sSESFizcjd6gvVfWJl
n0wWDG42xuqWQccVFzRPeejeHe6fGicmrig19dxzc1f0vEfE0+Ful7e8yghTvbZZbbpWrRMuajF6
+cttAuN7+RKdRyAAYMqFphdJC44ii3Kz8Sr0StVHhdM/ftJcwMWroR15ogrYPtGUOMB6awAlT9fc
8kr1EqSiM6h31k3/heyDgaJgVH1Jz8/tFmycXoHwKH2jyfXdmdG4ZzciQ9N6ZlgRdhDymgrSzyVg
9iNDJEAdCbBlnLmSJo28+8skFUtNlzUzusxVwZiLJlYe5eIwyeXEElSgATc/Axu+vrjifGVKAHZb
ipub+10N/OftT6wsAAxg42B9tgY/vfjz+op6nMriflkSfyXJ9L3IIZECpDD2dMt6zwDB4K7QSZKV
xCsOJZdtwcOXbqiD/iGUldW91T/pB+l8XxiQzyHTBtGXcLX6hifeCRqwuN5W5sifOpqMJrRI2Aod
N3JFKh7/OenMRQydPtFbm/OH2nyrPS3qP6AiMG90wg0wlgjYsvSZo5Qjq/A2UMQQyfWctqV120hS
ezJ8ZvomEDsXCPgG8ewglUgJN0iSNQrlQOTAqbfN4pOEgGQZmRVZ5i46iqDLlPig7o+NXXKzAW1A
qhkVoozGt8/36/bG7XTtVbTMwZglkjhcHSUSDTKoaPYDIx6lYKYX6pR2wqbR1We/WM1Ebh43VlAz
BuuoksJ8YaIB2wCf5an8bjJLXNEDW+kIptxHUINGOCV3P/gR0c9xT9Xv96gAfmX3RTVT17EWVwEw
Ypd1EWPEHf+ijXK3R4Qvist+Z+odLqQaZtsfVK9bcUsYnoOYmqgVIlQSJ0Bm03RIDtpqvNdhABFd
6JRnGxUJKZx63nr7jFL0DGo1HRDTYw4OoI/NUF3aV10oYMrEoT9mdrHMJp6ivmyhQTpOPLEs/Iai
i38Krs+21FlKsEngdKIPp8o8GO1rOpqojdf0Hv/+ckzt2zHqMnd4EQ+EQuxMPVcTv8GI0vwXqqD6
38wXFUK35oAeIrtJJiFw6t89RF/r89mBfdXZPeOG8C2muPgBlx/ZC1t/8mGzuF0MLGKT642JbKAM
azaoiO5xYNCCwy0WsyWUb3MCwEF7LAZH7rIo8VjUsTmDjfmAvjHGgLVef4aJLt3RHJwpfb1D5qU6
QN6k7USnismjDJsm14qXsYOZ0JPRRSOzDMy86jSKw63fqrywnSLFaKl+8W9pKFg79uNrpyyYr/QV
b3O9mE8K/WHPjUwf/hCGSnhWZems02MZkd1bqGsmU1NhWWC1xRVWha6eRASf2rqhLs3Lm5tvXKi+
5vyQkH1bxQfJvwab+LosNAynXajqWZehINAFfI/ZdziX+QCZgWMV/8fozmxhS4Y/x2iuMMaKtOum
kEDDmd8cL7ONqBsQJB6nQn7lfJUfD2c/VbflzkhuwTCwUu/8F37Q9ak0umI8VhAz8jmhYBtUHFJ3
EHjDmGxWhYWq0mbkRP2ppg1iQ6+vK1mWvAEjxe+sOtnVjX/Gn0GFe+cCBiQ7k2TnLgnXG6BAWKeL
tfNb8qdrzkBO0EJFfOiYnQq+B3k+ohcLONlurt06CDm5dHjDG6oliG1Y1y0IkeUgdKsIDC+Cczc7
KKbDfP6ktvTyto/Xo+VZT4rkMBcTezfvegTmyxShE5trdSiEbYLvf8zaCEPaF/U46RUbhkUr+4zR
+FNoUjrAmi5LwCMSxSoO6UON48pGyFpAuK1oQT5CmyiI3vAI0gATXGaFPa0k7BStQC15j7jlFQsE
X/Qg2R8In/MK6PUeKvr3ujXfgKpTn7yKHK0iR4mNOXvTpTUSdiY4HlQ5Ibnv1jKvypN/HatgOIuD
0VxvoucLVgWSdtnR9kyIGzCGrYMRdDTx5oxuBkBO5o6Z5hDd+lqw8xD/fTMV33kO+gkKwe7K51XP
hj98baRgjwyMkUBgSGnysljezdDIQqbz53Y5w41nPeWSYm9Xt4YHzZ0J766QbAci90xV+pFyn6s2
iMGAyRmSTsVq6AwRv2XjFnY5ylkuLHZ69DbJOpVQupQ90GA5eDKy/kDrsBfAuBAoASTdLRicpHsQ
okhneciBOS4ZnCDZ9HPnSPeywpuV5/0FIyMraUHxH7wcWE7BJlF5rvLvqNzyB6Pb+LJbmQkk4mbD
XZQlwT/juLwTeRga5GIdy+7qvCbRnOAqQRjEySMCdnJITg/W5Ep/G49/XwbCfNUAvccpiss5Ncid
byXHNppiGuh2IGuJGDdzjQMJh/p7XljU8rMCyFOW0bJhE4txTR7d4ky0YK8HW4SDAO2WBDUUTgIb
L6/zA0nIQIneooaPR+zGA/WD6O00gp/hKknDbJfLR+39soHiAn39gL4AXdDjIj/qPqpoSmUOkxJo
Rzw74vpDyDkEiR3SR9hSYGkA3goiyDyHBkeh0lWDM78kYt3UVwW3WLGh+CfLC46HDQ6NNfkHQKJ3
cO1L6P+4miZrCu4lkeTPrsXaujAHtXEqBvkz5s6vnQRiiIVseGa+2c4F6AVoTuGOEUVsqCFlpHSk
Ac455OlKE8pGVxZEUX8Fw83ELOKbmAafsMpp3w47oEenpn2dvo42q48Q65rvgvtRRvDEveVopw8i
Gm3pT4pYH1yaFSzwoj1cgTEzG9rJRckgBy8Huv6JCzjqBq2sALRxo+SnBGs/RWfM58GdS02jTGA0
rPKESTKtNq1GQWfGJs6/iLVzXjOHqs0uOYuS5DJkVnR75q9XwiqFBnVY58z6gpLK2FxSbFSaGzj1
WpiBEXQix1KaF9NQ844YzLjLX6bT9wF4diZaPEtn3MCYZxVX08xN0/BzaXGjfS9cDZMzCgTAIIry
oW+TnL2visCYtbNHc/Q3X+t1DB0XVHer4b7CTzSo3bJLeLTw0jGhBo6w85H90ZStkgP9ZbAmLLY+
ctq8dopwA+OI5/0w7+FOBMzCYq+KHxkY46Dc3w1s9C59V8pECjER+Do5cEqlMcyiLTytDyBmRVtZ
qYyvIAZiDB8vLKRpRAId61cC00vMFU6Y2y0v4fEcw7RWUA+f34qvwvzIjz2JBVlAhnK/Loj1MltM
u/RRknZ1rYxl4Ug8U4gb/Mtf940RYuC1MLw/s/OGYKjDoKpxpW5/qzxeQa20S63j3LYRb3Tr+0Zm
0ixZKo78/sJlzlVFHHSUEdleiSF4Lm2EiWPn+sGoleJShFTcbTP+s2LcbHkrLunaUiBqNPSbcu3o
N7/ScmASsyoHXxrOEm80MM0kyOopA8I7WvCD7JkZ+gXKmh+dmbwuv4GcuXRn2428R9cOpxlkbwqd
I3SuLImhebYIRwwzmvf4xwgk5hOImLnlnn/X4QIyDaosyDwlTGf2Dvkn5nV/adJITeSulZHAKtVJ
JLTKmCerK3hIjgNRFC+OYsYGKdtDfOGrYmTTMtZGYoDXtwcRDKBffIT7/EOrkOsvytPFOktZRHSG
wcuzUkSXyYBmANy15mj9c0VijTIGzKD/DbfROKEQhMX/9M6bhqO/jS5gOq9CHGYBf0r9Oia6zCaO
fisNF4Ye4IZA3BsdhS84/MihvE1Wsy4FddWVjDPDmcld78F0jdet2s4WO9azIl+9EUKynGwgi18Z
nq+iyAN+nz0pqQEsbsp54EgU7oht2BHD6yrWj5Zz2bGdE3EgE7/euqvGWaDhHpccxJpFP9pdxEOi
5s9nGvnHo6CREf9Q4MBON/LnPSIZy4TBr5140AWXyml6Q1KHRzPRioy83F42qVOjES+ynS/3GaT1
Fz/dCLX2MkYTduXgEOt2YtwZN6rCevXjBn2zh17xgoXS7GQ4J5D0SD9cJW350brDg15qdBYaWsP6
biirVzl15X0sdPV2BwqBnFKCktdPzfkhQ0Tk+HFEFDVSex+zevkmCCNOc2g7qFRAywqkUFhK7Ws/
FMSSyeZ0QFi9rj0v/vyROSCIG/REz4k/Jh/gOLeXw3Ws94vg84FLkPMTfKiucKBYnr9I2114b6/M
chmnWX8UWTnhkAvvGaAHxc4LmYy7xlQNcXmmzkHvbQb5RpTz9sgims8z9Y6XSou4+xEbMMYn1+Yb
gDtjXc+mdOE1QAdPbmPylgvdXrxhm0OEJCrnyP7VIffVY6tzBj/vJv1qph51SIodtuYs2kH6arF3
/Hn75oCjHIvX4vwEREquo/StkOMkCDdnXePMCQdU93eCobbjnGNovCLQ15AY36dmLOppBy/bbmxC
O9iYyQeEN3VCjcPGgGuydurtmZN82N54o4veDe9YmepWJKYjJPPpLfueKZEuyUdOV4BID5gt8/mi
z5sv6UNk05sw2s52Snt4GrbOknzns67VSANTYGD+Yxu0alABwDQ7P6VPh8QbwH12SP1sD8sQknh3
9w/2UBxYPvdiK+xaENHV9ymam5AiYeEkhSUVxVDsJ+VRQ4jGrDBzQE9MG4wcWLITHaDqrAVzi1fe
2JpWZSY2Clhjd50GGvvX0req10Sgfr3sZL4LwCH11hw6hN7Ulsq+SZhR0tUVHXbljHfAg/2yxnlu
X9GtlBmJcCtlzx/83oe0DTITpo+oDtDgtVKfTx+p0z9Fbv23agCZ6rFY+HlaKC5PpFDFw8WZNATW
95zXTkhK29aHej9Jojme2FlXYgqOGeO79ABGQDvmS1bgy79CHl20sCkcjM2jN5spm0OVoDbUwaY9
dqdd6QW8iO8v1L5RpGeuXX74kgdSpecpZvlz+51RaW67EzsE6khYBeNcMExkzfu6zGdxX4iQydpJ
zit2VGyMkOT5U9/P9vfIwKfd3hOUlPdcNa1a09z3btO16Nd4eXnGTVnnQsw1MdlWMhbVkLr+yFI2
XfNQIsEOOqEC4LO09UQrtEvaPqYSBEAYP/GZUOMg2yFqe6gjFetosIrGb9p/WjQgnbdKCUMMnOVj
gM3qscrxoBk/rBAXGmWRnROZHrduZPh4UMMES1uzWu2HGVqBUFWC6iwoT7KMvjeYitAjci4g2j7h
TlivC2f58OPLY175GeFu6Poq2Y8E9qn93sgjx157AlNyVc8Rz9+6WS5adwj0QleXxrLRT10JMdfr
49YL+hP4JDn73WWYv6q7TN2RYLEDrZ3pBB5eE6TiYmebDC0p/cSSQg2iu1ZOuIx56E7P1ruvKQJ+
0gXgUIhmB8FP+xhm86RWJDx8zdXDD8I8mmxV6ZcYfZXBFAhBGZNbBqsure+mZjgFu4KJp0lHchP3
vC2ha/XW2Zm+DV9+HXDvCvrTI1/gIJ+iBVXPlroEfO8F8LmMJ6OjnEph/ZkQfdrrP1KKmnaLL3wc
1B9BDN+9Sou54e15urJdzQAzmYeyBuU+1hVuONV4Alb02ZOjyeThhjnQpVpvfJ5M9Gfg0hrhhRCw
+h7rbu9SX5eRwTOJMLWOueePCaCZ3zRyB5fHNYbCrPDDJ+ejlKqAPzs2BsCq7NQ2GJB0sovGX/2K
MkbEJEiTwtwKRs3Ka7hV2apBdtexkNGXyxdRrV/5FUlaAOKN4nyeJEv58GhYCh3QlUWtrlYntr0j
FIe7KK13zLnCPinQcStgctq1z93rNSzzJghVe1Ek5ttFcJ4+3/FnDrdpf84A3KKURVV02ePpqHvO
45h2AbFziGNAlJegmFCm45C6vhtYV8nnaeAN2zavkWfv5y+bKFnsinuDKdbSrhqRfIGkn0vYuEnb
6w610UVcro1PyRvznD/ti3VbZzZi5WOT61IfQescB//99D3yE+q6aWCC+VM/Bh+vfbAiFqgfpzmF
pny+iPPN1LFKnLZygKajuvPp9gwwR/+uDYBw1wHh/RqbTTj/m+nPzSeBgwtgf8z8aV2nwrJi8xqO
kM6URwIKLFy1ZD/dr80QZU+z7rxgVfvbeb/hZ1OLP0byL4BQM+TovWZnq8EOgmNjbHfsZ6DjzC5H
E9iu9I0WTZQkKhD7aRMbu7TNeEgPfqNZtb/Yfx5Xkf03VYXhpm55EmloF8WgBkaEyTAJTkizwUY8
LXRjzRGQXsvjK7O/vrdfGRSLLtLALXD4TXhXrXBIUqPzACc3GiOwP2B8G1m7FJ7bkV2/MEVpWapR
Pu9n6zTeBwyNPqIeaMv9Mvkx1hsFXas80ooxaggtIck7bBf66dXdLDIdJ+WQsIi61DmXhTQBeE17
y1sl/RRmsTxnsMIcp+varNaeegOORLgwLOg+l4/IyswxnKXJAbp1GuPlIES/KZgt3ho1R4mrzrnh
eKZwo2mgWOK3XI+IdfxpB+udT0KWhaODbLWE8ouIRsWJekFz7UAl5J6fYqWB5lV5cD46jilZ3TdR
S6caThJQSbi4ZvhL5B6ICjZ/3zfOQ63piCu4yzH8+FJ0DlSgxfcq9+is+XI5Utqs/uTgPkcOW1FN
9iKbVLkNiFtlPCll6e2QmFzYIWY8qA+fMvqS/COwNKgut0/BHFDK/v6zV7ng28B+GS/AvhA4/CXs
SiNLAZeRzgULgOL2UJdvMG3BbJr9ejBsNOnCy1e0IXpXCVGOdFNO0bZJFF5g4uhNG5cP3jOXc8wL
noR3MVd2n+pQgKPRg0v7HJgeEwqXyWd/YEFjGidod0XBgo5B9voBV2kwpMk0h8vW73jOVhH+p9qq
igeJPZLV9SiDIzBY+vFX9nnFnw3iYY3LvJUe1jdxsRBfvcZCZowmIU0arI3IQnIUvOdT/nlCdYSF
OwMVuFV+rC8SekBb710I0RDOE0HuTkl44SGls56su0zGEptTGjFnsbXZWF/rVBpkH+MvSUGVfoHc
fImOhuHM/t9WUubjviizGEfWVZDX5/Yp2eYjQBdKEr2qjALXayEFDf/+29T/rLkgZMsq+61DUXcV
GVI7WfsEM10B9YU92yomuTaVwk1Y5lU9ip/pcsmF9qIQAZUvfie2EI46CWwX9MRj7bNx/cQb2eki
9iHJDzMGZ/90pNYggGxtbxe48xu9S8m4+IBNWjxd5RBOGyK6YMNp4bozfzTogEXNjlvVjjjkNBcQ
nwl6Euq9F3mZvM/7BYFyNo6c6dVBVSLmMKKIvHw6baFWda+v8hB0hEsgFu8Jy3uw/CwHDQ3dGMaL
zLBmaXeKMF/H/MHK0GKOlFHRmLNxT8S3oWOXW5ZHiLEttabL0QegL2h3VPgqEkUHRdM8hISc2SrU
TS9b144xatPLE/vwyc7HbSoVLhXGotuEaQaj4wuKbENBddnYP2bLmWZlx6hqqJz9UtUll3YYWH94
S0B+QLBeD7e1QSo4/wp3M/0s4Zdan62giN9Yw4sOV0Bt54se243wlGpU4FmRYlZYPdiIsXv6QO6/
X5dO918bsg3WOQQQfxoS7Vw1tOKTBV6axm0wQH7nvikNE4EuoaNSUp6I792asbpTu9O19qVvyNVP
xB4OR9PULUQtWNBAsw25SsaglJzgZqshmhuhcr6Uarc92kzdqPbg1SoltP8+ypx77hchYgDQpfuC
i7nEl3+6WbSbkL05Ax/ocr+yx7qJ/06GYdcrTbVk1vB6Pr0BrxAzdNi33/ZA4AXAX0oaNt0l/WNL
MJxZs0XT5qfok4seT1x7xHt/WAc9EfspiKZ6EJ74C+lTGtK8O/zFysyB/6gwYo74u79Gs8X9iydp
fCOZ4jcM1EwexrdFjvqZo58oceHujsxfkQ5Und00s8c44JQo62na1S1cmCOwb8CPZIT5QCved8NJ
628vC9iboP+/sCa2oiEBa+Su7mhGdp20ZOKisyqPKUFv48R+SP3B1O+nkN/PuWmeov+BKJH68M/v
pKhA+6DkARDfugV/rIQXjCiwW3CDFNeBwq9+jcqYo2Y0JXxfrtAcht7dPk7DR6w9hE8t3/xlGnPK
Da4zR46eigAWbQ7lSPMgv/RechVedcTxt/HLDFxihlUd/9gdxPjjqjD60bt7wuPHw2cSNaJJlY0j
HQGHOek/1ddw4kaOtSHtXpeEftbNg3joDJL6vU7JYD+Spq8hKI/cEKWc2ApIGfCCCB0DxtXjE2IS
Tj6cObpSwf2be0A4ElSHP3qiEIVzCm2lxv8nNdOiN8PFBeW7/VoLIIuR9C0VUyRRaEFpGgJE/hC0
scCx8qogymKGXavVPTpLGTCOcOJrj5/dMXCGO4k9XSBIOF3URSMa9sq2c06gDsaCeSCTbcXy5krs
4gZpuDRBfcwKE9Stbs3z6yXi9/yU/oOC07qnce6ZEG1ubJBsB69nfeomIWsLtvl9x5A9mtLlmQGc
0LSnzpXOZKIGOsaebx+gHgssyimyeFv08NGLl0FlmoJgHSd/Y64clcSG63bDYUoJFQ5DJc86lSjQ
RsMdUA9Rn8EGRnBBMNV1BKae12zSx8YRRPUGFxw1CVPKzK3sC5aXdwAMoC/XqNn0spORD+z8aBI1
8n4rqKcxaaDwA/aPAENGNGcwRP3vDYiyP64uX2UwZaHj0WKC2pUZlvC4H1gM0bldzJCB0GEvR8R7
wDvpitM6Z7cufNs+RgfrUD3NoLgKQ93bQBvlKl4iS8hd0uM8U3rU1zdGq6b+StQAAl/1JWiL55uU
bn2vlmfVuFbItQrqEY1pQvGXJYONcsyBtFEXuNZydXsIuXzOxbRW3H27bHCbUlzTRPeDkyrJ4baH
UWs/I9SJmn4hdfJ3Y0UfqbOoAxoTPqHX7KIx9ME0yNWqctj5cldUbQyohuwMEWkjKuppR13RnKMr
Kz7vVezidJjRjplmsRerhWCQ1MueM5Q1ZxBsiUXVvtgxo7ICBQBVjdLt8fA6JIzcS2GPywvVe5ir
U6hrtSR/R4fGOpuIv9gM1SqGpffri6DiBTHPChWlvP4j979vsU4dwAzpVStMLG2nsC5TSJwKYwlN
cMSbO+3/XwzIVPVPFvZ0UR04vsc7M0eHveWD+PyUefiau154IwuGDjbqc25rNsu+vKlB6w/bIGxx
5ySePMgUoh27/ZniJ2vPsuVB/fapDrK/caYSMt+O9qZDJz30b82/D7jeruDFxjEKxpC2lAY5/nFK
vXKnkDSGL7d/33ZNS6Gxh166AOieljFAf1CnPkcW7XmzBYYVyRnrFPCkz9sFdFMB1+cYTRILNsJ+
m/I10f8ltO4GXRkdVvWTuBIo4PoAAgk7fJT579N7McUqiNSng7Di/Ujhhx1Krx+uUtzLRnTBn6Gp
G1jeW0VtiQmc1bNfgjx0ywXyiJMwJDNBLaaCDV4j9v9HjmgJACdzI/bGgc1iGfaUPQxcjvgrKCIy
6N7F7Q3whi57FKfOHwaG3SdrISanfVzUYNcanWE1zTansvJlRAXrfeZuiKGMi6dEKMB7ITrYjDFt
DQ5+wj7XQP/7hiFDez2HYhIV/WqLXa+yudts9h68DAYsmSVS8iOxVazI61Q0S+Ih0W+1YPesXRkl
KPl2hvYb5NBIu06xxqWU6TFmtHWtr3+Am+h0PqPZylNNU4z5NqYomVxFX9NdaQw8j2hZksQmGoGp
YfHLtBy7kmJx+sc5Tf14ulXz8Y544PUoXlsye6q0vX+k5lVCppJsjPsVFDxdgozP48UUCsPiuVco
RyG1e1PRq/gA2cVidVcWvnPkXxevydxYva9aDWgoZgOhoi8GXUsYv2lSKJJpaXWKK6y5rR1TGMv+
71PeLMrjhB1DRDnfH82pG+Es24qymRZ81pAGp8N/K4fVfpnSiBcMxPpqxfP1Kqb7Bj3FIVtxfcqC
2h1DIIuH6+khEjIICu8oZAJbEZYL6MYCJihZZnuVGAr1kWKQGALWRpPFrwf0BKIq2lnPvdvEGHji
J35RRXB8TZjds63+XLwQrd45OL5pfYlgmJKQtZK8qhRqjVZ+d/8iDFVnSFXgJdL9iIZ561s3MZj5
DxE9OD4GFztCF03/bUX9xPC8CbAA69GozeW6HKX47/TpVQeFR+Wv2aDmBq9CQRfyN67NWGijxvRc
P6Ud740vJZXOYbYu/mo83YRMS8GtKCiTdyM6EIeVPHzhkGYZ5SGabuYxWigMGOZjV2dh7+H4/dyE
VB6vbEOSVyRDvhYDc/Wpl01TnmrduPhwOZ8NJZZJi+wNs3L8bfxCjSJknDgLkocOsUaDFd7XzkHo
cnpdb9k1vCsIgjr3U4e+1Fg+99chscS6QLV41l/Oy2LyEF+Yz/PP86DnyP8kEiNWqO7FFMMG+mip
8Ailpne0COa7rb6JY61nA+emUGUwaQfuzOjDcQZsHj1D/DRilrDA3gnfwwYfsjPYlRJdwq8xWZrK
17z4CDkRIg1JQEIko5ymUkzrshwqGWvOeyJ7f8OqkVopZkfLauVXv8Z0QyRNST+OTH5LKh3/zzUt
Z5XawRJsvpF4xHN3FZJmgMtzPEtQ69uB1QP2eGGoxHHiQpjHL68IcAuVFN0M6LuUIKZ3HmwpPJJE
KEKNwjXrBcH+8jonuSzBCrvvM2IoTSE9Vxypil8o4nsxhxGHRpIszvs4eq6h9uJB0/X8GNyorcqk
6PmaDb6dM8vc4yD2tkPpVftaOGudGp2USEKeYPSqyrPIEkPL0wrKy1wKIgFVE+As7TS/L/wsukJh
QLepq7IL9l0/ppUw+vCrwlrYzIrS8QLixi0MQdhVEu5Dma6waWJP4mf4OjMfJma4kgmegu6coTgO
fBt4uubHmnBmceEjEAHPGjejYhacnrnSTutbzvXq7R/ZXXMKOybWVrVY3ZNgIOtkT9pU1SNE1hbP
DPA//p1ejHbjFujqywxH0ym5ucx5qoVCO2HSGNKHERAaLjijpaapO+HvPkW24mcDsLwOkOi5heDS
98dvF84oJD+x5aTYvgIvBDNqJjKL1B+CueQUSP/pwe1qaBg4nZEeE3RUQoS6NDTV0JC0tCed7ti7
o9Nan0VdDCfuHf7KbTKsXlBqPiHQ71iHNNjXFatGN5ZCeKehZT4dajj50AmnZLSVENutCzG2V5qa
4b0dB1skI20lsl9NNUIvS3IfPakVB+TCcJVEYKdUDhGXGOC9yd+WrWJeBGjBYpy3fMlNqbrR2QF4
Q/sFzux10hvLJ9o2Jv3s3/WO4ioeLf9nJEzbUPMYL6Ap5dkzXbQEzuzzvHZ5graK9mLijDq7Et/9
dJ915wmvleYO7Zw9Txe/2CeC5fkXdEXk89DzynxtVUA0/ok3qXBUJse9Zlkw7nKcJM27ZCzx34/3
EO4Pi3aG5i5oM0xk1jKhe35kE8ZrIpMgDLzMvn9kglkzD7zInuo6PCm1k5zHqK8wfm8rdTl06kPw
z/Ch79RrtniYp6SbtVq24qQwN0qVBFutYkTmkUv3Mcn/KPmDkBGGpzenyfXFOs2DpV/sWau/EoDG
PC92tIXZX9wcqLdD4Sjkh4jvLi2G5DCvA2cUdstxAjduMhi9wkUXNCSYyWdJDkOyme4MqOww8hEL
/H20sYiLr8BQ/pKTX2XBMXpUT8qO5jQyDmLYK7aqruzjKZUPSwq4neWsBTAfmtPkXuYukRkCTrHQ
GmqlrXWb2MItDGSaL9ip1Q+dGIB7gm+FodbbNIJGCpJQ3cWGevpLvTlfQSCrQg3L6JlAV/lKib3K
cRom1SvmQh4EV1+S7OHFfit6IwrSyny1LoCS/jcP2ND6a2KEfzimyb/3o7Z5mqOfE2RwLm699BcP
2YITQTakidNH0isCY1svxuC4TbK3uvbpWPxILRnkxHnoU1sB8ah7UveQ9GTNm6XA4MiGaNw28IG9
uWAGOjvBdwLXeT8KJ2AVD1FbFXvh7rrJBG/AP+0++qsur3GCtWGToGEzpOXUQ3e+P3ATjLi+r5+x
MbQTT541zJseAfzkylqxfaBPXla+Usavrt0JDmRvkx/0R0rINAST3nfrA8MDJR4wQStalc7PJt+L
MwOwmEmh8esHlNLneE5Kk+sQT1yWwlv1mpuD5VmJSnorLZEtOlXOiRSPXrJYhY5m3La4mKdLX9TD
Oc37ZJo6104YpEbulOV9ss2/Nyx825bRjcM0U6Eb43FwASmCfpPyhyfKz3bn7CgeQdlvosAiBSYh
UY8beS9BEJ9+CdVTq7l5lQfMEKdxU2hqq94r092deBECosZ9Sz8NuC6jjqAbsmNOf5yDgUm2ysc0
CpIt3WQJO6aaSEbO5I6Qp4bIBxOmaIwzayRPycLyuF3PhvKmFc8oqwkXypJrwAUc3snwwu8D3qks
LOyOL+yi++viocVIetQ7e1T3jMzHc4asnrtFKQh3fAHozh+iFaPAd8t+Vw+NuE3z0IhG01uGnsXB
66LAtZlLtd2kEP4Nh7264atw9BlrTmACJ7cD7q04x/kIvHBwkb8NUTCTtdLWw4my8kpLbsGLHVlr
tEIJOJQJnqkDJJx1n6dtL49xBhTwUkOqmpQXxi4rpwToDqgAGWTOZ+i4fpEiN0xiyNwSvB0tCeFu
m6qMMLNg6I3KtFGxss4TDPIH6xr5thgllDRJ8SClEvvgQ1gChEBBPv6feXHM/986m84J/FLRJ5uo
+pVAi8NpC47Yu5OYTezM1zDoM6cXGwUQn6pEwzG9YOaYezbWiHKOmeBOWAsQ7EReuAJo2oHT7erN
hYYVfMUltN+fq3zGkKS7Rqk1j3KD9ZSBn9XuaQWJQmnVLVateDhYfbEoNnSyG15tuW5YGqn8MFHx
TTOn9PwZ1M6/K8uOV/KIdArqtKbBNNYaXdUEGG0kV/0y376enuEtE+hYsj35mT9uAPIbnL5DwTbK
ydV3KxPfB2CGye7IVRbahpsBxU4nhfzwkW/BuzW8EJwmNONofb0LsGQTv0levwaAU5KISFhVG1bf
QeUrDjYbzm7qBqvMI87tOU0xR3YE5Nbe/wDzivXhmi3wcafx+G+Rfyy6lWKridp9UYzswUdpoY/y
Ij7scO8sCsne+AXOe+erMfjsFLbePACbwLIZtjMSJW9ipBrGWTXC1YNFUiRZRNIh67iD5FDDh5BD
gm/wy2Xg4M20qQ3ijgJfaSBshFBT5gOpiQL2m2B0j8pW8jpsMk4cXQFmg7V0+XxQnmt0QqyT8bPf
d0hak/dFYQhQSdwhdyrr6PiRRkQUqhyxfcElU+Ix3/Kvqq7weqdMrhF6ymDSYaGhoQgW5Nrw0Kl+
/KOEt8MLb90kbJc+nkUkPHslv047046Ex4oHQlw6fvYdQ6OWovW6mfxCMqLtj427GJoBYz7cscZB
P2+CFyzrdihqMCuL2zvhreI3+kz5OKHZTGsLj0DPTvPDK28676AEoAWN1dKpfTcs4OlxP6WxmGdR
ECptdSFCDB+ycgl2dVVO9a04arSBZUqfWIAptm66C5rOr98dhlQAWFy4GrmCsQDxYP6IBCNdBLMj
qQk2UW4kNTVlj+rTVnLIqP2CSeGTHSaHHPbsAi04gfU7ZmJa8woj8tUwAr5hzVzclHCWfMoiTsR5
btRzlxdK5wQaoeKnszfp279AWrJUZLTMsY9A8P1b+8BpDhM5AhWnvG8hSC9yJgvJ3rhsEwwys0gu
TPzz5ikQT3clvLzvrBZXb2+sTCF2Kd8NqFgZCe4GAOKP37HAVc404I0PtCt4EUW1lXjfRp6T/8Iy
wVnPYcKfZdMq6CjmKmu1L3DxCtiwHxO2oZopK2eH3EB2VKDlom95wR7QSk4RumNiIExq++P9SlNk
Z6xRc8W0YnyAQEn/yC7evSys3USZQ2L0O2e1DCf5fTJnslyED3CK+653tqD19iMIhy4WeL0vmAud
tiYFjFlEdQf1Y0gHG6ICw7v/chkbKr+IZlxQMVl4BIKwfmZq+JihgM5kY1XzvE/SxkB0fXK8i196
E9RaS6jQwD7Dh3vatY45HFkqR1qlt680nXKmBTqtBwgK7EEKh+xSjjhfaLhv5KMhF1gXncyNamKv
GtVea8vdCe42RMe4yH9vm0NTRKfVRK1+FZTb5mh4a7YitFElhPm4sJnrLOxygrDSNVZ45ft9ClvA
Vmzt6T9Bj7L8LDtYAWqT56nxD8QhyDw9pMv+nabDjO+qQuLDx1ivSIy8uQVb1HO2GGZif+mIJa2H
QjpGIrqV7U90zPBX5C+urmClUGNArVCAmjR3SKFLuYfSEFxUxyBiDfZ+SRARRJC9e3xGAysWyN4T
N6KPbRSx/hy8l3KT7CxZIJgvTcvn0BmYRM6Jhlqjkls1lC4MAvz9ll7BQWEyDYF/JjfsvPptehD8
AFw14CYUaBS11AfPDa03PVIwvS9K4+u4a1XriGp5ZNVD3sxqMbRs3GZSKy9G5DUerAb5iayt+nOX
r8NlPq9BOoMtpZVJRIZA5VTo0611vibWwK3+lHqMDYRVmVLF/NP5Cee2QXoXdjDTSadF5DG7qHVS
RY+7RIl1zMT3qp5CzrF5JvUTBM3yVT8RbH3nbubV5Ngu/Q5ukqNBJnP3mUT18nmCpWO3hnw8KL75
t+VRW2FbAYGbiwhBIY/cjfBCl3Wp/pxy0de78dPXHhr3audTGNWFtoQgWZTpRgS7mZiZsLCfl0ph
cjnueCkogRdFdEcDeYsN2xdUSlvrC22ojBZ6CLXNAfr8riG/i4cRXVV+vLLgFxwUY2ogeerWlE7S
Wj0jY42057JzIeDf0WFZCfSW/31XT9WB5gWSkgx+Io1C/lt5NsD9kSuTCuKg7ZpzKI1DwnaUIsKF
BeictFqqc1rRAwfjmMiMpvvrXgqkOdGMzeoANk5jLWD2J27zskMJWnl9YbPDN3MEQ0N/JE/RlOoc
J+5b+rbY6HyB14WFmisGXNvwTZx8hHf/gk/gg+BQ2P2EhzQ718qwRZ2ktv44ZA7HnoKFCdtOKDgH
2TbCx4Buz4oeGcgC0u7eCFEnGX10ObTa7oX5XW3Is2Up6WDf43g3zzoRmjQ7WpvrbO1EA+UtKWn/
QgcEGRuKeA20KERvTdpAtH6rWD7UyfRHk/CBDy6jDJHOmtnlrV3lnj8VUtNmxpivUGhPvpRhJgOI
Vm6XpgKdG1AuDwVkmnvSFv4LM8sV2GduSijodlAwjl/zrbBBn7BjJTbIoWb2sk3zyRTkx/F7nYWA
MceMyiFfpl140drutPaPbsZmWXJ40+bO4M43Cl3l7U+9YUfno6CAetySBqH/CVMADOcmpM/ZJPaw
gMjVAf5I3ZwcLUw5ioLDPinXZ20lq9jG3ZOTCpdauFTwQ/AYXiE3W062mUzCkKpOlY03zmQHw3/L
5TRvZ5Jr94JNqMrTAZlf8ADu6Auue8LBCD/PH5RhtSVha2JV8pvJBG92ENgomcier01YUpOAj93m
uU8WuxEQ7kwBoi3y258MKVjXX3ZLdZsP4nx0qjmsICLZEOfnCKYXFaGJDBc8CqCqtRPz7YyYZSxs
mpMpxYs7orpeViexjanPP2eClOdTQRWU6qyhpPRVMF1UfIU2FDbIULsDoR4PdV045iu2m9BilqNd
9N09lmbCy9KH/iBDyRz35D5u9/nsdDvwFTIubBKCjxXwifUbcK+MTKq+4z+MhWBr1w+Fxvptc2LO
p01DxGGkomwVW4sfVyIfVeQu8O2Tsi1pTPMfSOD+4IAVcauE1FGV1DtV6/i6M6luodnZUCAI/aAZ
87GS1p9RZtXKnd4liMcEAHvxqjqo0B6VMqS8WdGAW+vjg5Xx/CAnNsJniciXzEPS4vl+Y+RYeueq
oVBVs7gyFIWjz98/wUGJ5f+Ojb6UlH1s2lZl8DhwDa+1Vpim2SBRx4MsHLIaFWpvWVL2XHCDQOHJ
34U06edYZ6PEPR1Tm8pKlRzl7zTToburP+6tc/8xX51O/ku+MWR+mPxqnzbHU+pdqRJV9WPtnFo9
0QatYYlysxZoPHGV06PXtLRmd4QaauIUHYtDKnNDzYDgupGnWbzSJbmcZDRPcQHgIK273PlOjThP
aKjv5Kx2CLWKHa63sg9Z0ametTX6IlCH4EKItI8w+Y0CR2Qw7ypZXgE0fxlT3tcEoBVmPODiAoBe
noCwPxjiEp9Fp6iwcGYpyQKTDinb8lF0G/hMegtYe47e5CjLmLqMtjxeBZ5DwMmCwP2kG30ZBeEN
OtRvFSrvlf1wI5156AWunxw3JE0QNwkeSwgxYKozsUi9YtX3FoxJAjRNzBYUOpGxRjfgaX/jKgvq
VSyAzbtT7ESlSBolb2OVQiLODND1bTciN62lsu1AB0QdhBqMNVMmBzDdipJOXriSzzqAPM03etKb
pzfhhm5nsiRr5Lii9Rq+/Z0kVQJAaHi243vGNgTMRQ3RnDU3+paYhUyYDXGhJewQ3QmEtK6h6uk9
fLirVitmwJ0+C/sWbsht0NSWtih/SKzu5dEnfmpziLR6kkYH/bjwyNSprblmiJVB4SJB98vUnLFz
itamfoCKWmBpTHuemfKuYRVe5FwXa0MHo1L9DvLjAbBgdnBkdRAvM5dM6R/wWruKuz4FfhcWFjbK
OS0sscK1JT5qozRKCg5/F97K6PSZuW8IhoJgTTDpN7bQIwhGToAgmZxLBHZycY/MaHq+Dd2iycTF
JQee342l8qqc3dWdekW7qWIvWgEApBTCe51ODYOZ+XYEPCGrOoQ18k+Sdzx6RPn+ee3WFDphp6fK
glWLsXPntlaOoZPL5EnsDpuz6mZekyorPON4Fj7LNGZWNjqPaxHX7pD/cwnI6txk4Za4D5ekaDw3
n9IfANj0jASENWTyidO8PDWMelVUURGgs1T7t6FzGlgNVPuhDM6ZggUyTkkBgvrr6P5NfKcAfp4z
wgkEHVkGCynk0vtu+jO9RNYWvV4mbeAGrTXGf3FhYpc4bfXhp7EbRg5DOUXYX3mZUou+g+0UxMOb
3hoEkoYw3oQdJhAyceyY5sAqx+g08kt3t7YMU1Mvto4hohDDmPxYtzsumuv30zmSqOZHG+4NRZWJ
15HVhUHjrDUlTuorqv5JN1IMx5QNQFwxjDV7jv8AXM51+F1zRboLSAEH+kuG7j9NfIyHqiKTwvAU
VEzO2oDFgjcwm/u9SFFPJhmS+ng+9w4AHeLYNpT4rdeynt8/yfxTXhP19cCLp2McTovXzr/Fn12E
l+Ymkgu7THmSsqmiJpzeUsny9lYJq1hU9O6WlJFyCMw2UWYiSfawXcDNX8agmGxHA0dfsuiGDvYf
O9DS5qo1vg8ut1ZgIOZ+A8R6Ec0Fz9X97t0dX3xfWXzHdP30sED6YhZPiKFiCQUjiPCeXYX7zUXS
Ic70F8V0Nb5ZFml/sG2kIsvWsGQ2nRM7C1QoqXZddjwUkmsNPIpbcNZo8gqjpLCDKFCVRJRHItk/
ubL7ES8s87k0yJRaswozkwi5A6pv9BVrIRrAf/8vKu461zYBdw3wguY7kRLbJ8zNzFaTdkBWj8pe
nhgR9+EqLa0RdRdi950kiwLH5mb56oe5fwPmUxP74BU1/Fbx0sOlnHnAn3SW00C/M+AyO5kJWpJU
EkKNSFWG6UlJEJlX29Spt15iAEaDl0v0jMP4prWj9odRLE+XGf1FIKMMC5G0WXThcA3BSY7Xw5Tu
6eczqFCM3JdregqdlxRzqJi57HDDJdIFM4SazWnU5wPU5pfGCFhRkhJP+fmkWomVfPYO6vl5+s0s
bT6zcvIDyPBE02mH9HkRrUOO/SQSTRzqNkyv4tSFJYuAxKM249nHAVWMQ+ObbuhiBIpDVb0NPMbj
ss9QYtZuRIq+qFtj8tG1DRx55FVf8Mo2P0jaiCRgudYfuv9/sQt+e032Knqb6Huc2YyjSo61UWTY
RUwBqorQKco5Kol3wFfQupIsSLS+AiWAUAYymNKavadGA6TsHeoHFoXBnd1hhef4SOzwdH2Waw13
RD5KnFRSKOR7RLyaILsjpELWUByqzXN+mfrfJKBObUgZlCniTlwNFB+3pMa01C+HCwwX+BwBs3Ad
Gkm9bvsZxiWPVlEYUulFMkAu+aXLJbt4gc+TCalay3vfog8RjbVGwZJrK5UeYB2qm7+RPxYAs1ux
AFOI8ySrRQlJOI1M/8RF6XKpkgWQhqEKmGXsW2JG06rOKS1bfnWuF9KYvT7EiXcmNdr2rRw2UesV
5vGUbM2w9lOA1nkREVECfMtq/DzxaXPeuyIqY/ktqaf6JUVVBGKqNy8p0zoNQPx8xRj2hzUb9ffN
tYp2mUzyCnSOZor54EtxrXFweAD/tglj4jPcXGw8EmQ09x/pdyxUEgt4IdtdFRAMLr8lsQy/yQsa
hCPyD/1l9JLrwjqsfj0KnF/5Dnd4LedN/ngol6NkcqddxXumydP17mqaPCQFfbqV4vVhYbSdVtAy
UHmRAf3GUJFlOezzRP54k7dQJjZnulfb4agwC1GNYrpJnSpi9KhboREtdEK4NgNfyl7fM25eZ3HY
+hNp/F1wTap+XoxXgllD9t5aD/Dwc74gOPEqcEOGDGkulSRuSKqaIIYU4atoYzPJKSu3FFrgMl0t
xuIJNh4PHqQ/PoJiJJRXm0Jj+sErIHswV1g28Pt9MntTn1PFkheR/gKd4ig18bFe4iNgLWDfESLL
s7nJK0+AEAeP6+Le14vsaTqsI9QJpmvEzPVUD9J+cNdPcJWLNLz1dQvY/YTYJjwiaxHUZvXz7VD6
itnZBgwBg6J1E1i8aEtV0LEOZKjmIawxf6jvvniiIuYNAlXtOKG2ypaYjvQuLUFtwFoBKQ/GMqyJ
tIHQQhufI1pQlyTLkLw7hoBUu2lEGALP2RHYWlarNAodbtEd/QYFenDAZmj4H25x4ynqNOURzN+M
CXzUf9SszRTcHwuKAsfZ8t4lpBKCf16QVTinWUrFiyA8TffY5rfaIfXXMg/sOUkU0no5qX4y7tyW
slT1ge93gs7SlZCWLPO5T4W2ODlR+57BdBcVra0jxo5DY+OF1aP98UCa2p6/P11VNUBwbm6Qb+o0
jzpJVJg/BJeP+vgnL9oR14DlxmmGq6GShECmPlLgVBTR8SqL59RUo8C+kVmf+7+y9cAaEFl/gyQR
M5RF0cOgsf/rDCqyfq7AVZ1PSuB3JeXNgsd7HqKE4HdSKTEiE7fnviIXBiaPgsFdPvPfbxd+tAgG
ZfYiqi2QXuFOe+wW86L6XpaJbFD8WrxJOIX7tAo6dmKRJZogx9PBLt7B/66XAnRoggYo7wviwkJJ
phse3KX6zy5yGsyf5dKhFs05LtK5NZhmiHzEaL9TeACAbS4IY+Qaeae9tLQB47ddreV4OSR/qSTW
/NTIsyswJDsAGJ3aD/I7UzFjoDmySfaqFyaCDG3Dya3lP+7B0uJftpBOiq/Ql+CnixdSbEboCZhp
qzimsmzZQxneusT/RgxxOD2iIStn9NKxDvO5Z/K/jNbKwbUR9ePFW3Y7yuy7imCbQF4OE7hT0SZx
VxLKzP/wv/4ZRx/V26+06RKQkBWUMFixJx0xhIRC9Pj6HPQUD77dgnr3mvfYSxZL/jwCiJoe22Ja
IiV58hmmOohhoOAVK4zzx6PWyklqZq9VHXAG+JyCOouyoJM9PNmCkEG3BsuqkehAHLAJx1+sR6ky
XzFUFGqcTAXuWaRyZopAb5SXSB3zWhtvs0ZGzn95h3wWC8GdvBD8gMKk9MvO2hJDMXNMO0EITsX8
7C2fFZEKBQvSrXLrgJYH6Q165ydQ1zvaDKBA3/9EYoZK7UeVPETdW95EQXHlqRL1kqb1yD3uYMUo
azIkfbIV1MMDhbGaREHmT98vg9N2nm+bFH8uPIXO/nigeoXf6/NZ1TFkkVtrkxFzlpsA+EadxF4G
3DESG2sHN9i1qpZvuxBC2joDb8a2fPjQ2RwsqQfiNHn20UqR63L5SKT98IMZnfvcTds4zAtrlJep
Ns21w4iEF7iLflaXRHlT60Z1/TtH6bSydUDNhftsAvbFAmDdsUL0YcTH9TJyrV+88PFLhf37RczX
UMD6U9DkMH8o+rQvhoa3tkbZDpXuEg6NUDDBTKOicsEmkoCDjNgfVehGy+tMtGIv6SxLYXfrTNIx
UTyCkx5+RbuCF14tLHiuXM4nSdEANEBDY6E10KIFP8xbFN1bDHBhqg6LFCLXFh8WOE9JlqWpZOYi
/sXsPhydKl95Pm6XbbFDppabQMUzwChDo5gfv+yBrcmr5Rrf/DinwdyExPwNs9Gjj94Mq8+PGVkY
wcH4ajnr+ghgO9SkdfS0eA2EZrN600QXdD3k3gRMv82P9hZCSPBjcwluc29WinaRpMM7bfy/ATlT
QVQ4n6XOhRxM246zsrTqoQje8E6Zq/tQ9yCNUlmvrOb4OhAO0DYblYV+jgekfcHlEE1MsWTTR/mj
yxQT5LKrwsNPme8C9gdq2d4fg3V2uhB5GMTo7E4cRPIoAfB84cvnzhmqXBB/5YIXDe9FcJlPvrbM
bJ8/3D7bWLkSLplAM426JcLZLrPOItXbVCZ/+ioawd9cepOjY+dg8rtW1PuRSFJzh5ProfLT2Vsu
bm+6VMtGQVcxUS2tWNM0aPEn3L/H0OfC/rtqLEUQjxm7eb9vIh5XwqGNagAVmheQmcl5EBpu5FkB
aX08A3bcRppQnxq2HdwvMEwpWh3mD2Kf4ytzYy1LJpM5e+vQjYt474FuyI0jm4pxjAzPZkvWOQle
uujivIgUmVnD2947vQFtIm7oMDv9oU1d0dM2w6ndArbdDPBtF2Y0gX7aKAKwaRJrfXKsxlSweAZu
F/eTtvwhnamcnPi1FbyhhyeS+K3T+68cfbJCi35XEfUaZfkqijQ621rTOST70Ii9rtRv44gO62AL
2NQa0IquQ4fFPk25w9f2uNHc6dD6YSbwzcH6dd8K9tQWX4khuXVu+eoWc2mHjJibB5pfAr6wRYDA
H4eNHH9A3jTERyObFd2PDv/ILuAL3/9WIZKovN/69JSG6Td5vTFV5ojrSUuN3FiHPyr47l/bn8/N
qlBTdzH3dF6ZOLZ71T7htG1ZfwsRUUX6mwwea/jEjF3TyZqxw5IF3Ur+FizDz1tnbJPtUBw1NXGg
VV7I7TGhiCLxP681lgqKKz8OUO5z2zNli2xURvQA+sJKthKRCORxNG59iJJ2kEA//kdxLIbGCuSQ
9+n1CZEU3Nr1egUjHdX/yQALNYOf+h5AtHHVfr2iyT052ciYTDGda2h6Ni/DHLZTW9hCnW8aubiS
zc0rsbc1uCNsot7+Ygq4NcTTcmgLuch7dI5vTi7URbJOGt22tDM4ByU25/pvB6v3+/6A2W54dFfg
a7Q05rp6oVUkRneax4cZSivCqFOTPZoM8urhT67XOM9cFLP/Yb5TMKWHfpSL4WNck6rVUFFFYF82
AxFOH90wO+DM0X+5CMGSrDt2MugjcZ5Net+4EYbAuPjfJszfyP7uamrGL5whHpffK17lTDC5Bt0N
5OPUZLl7Bsnd19vZRI9Mr2geC0CdM3FwPyrDatnD9OiamhIKIMzlsMoo5PV0UCQVdebKvnhwt1Yb
lI9w7xGYi38AmwphhCaaLghgkPge9tVhzcJUXvyGbP1cGd/xukjkBVFgazkw6O4mRneNMPHN/S1o
+ynf5ARm+/279lHsT06pfHjQmrIrRtLuehH7U7PZMqOu9hZlvBKDzvxTd5QGW9kDLwpcs2At7/0x
QZ74kpDDnXzDXbs/BEXt0olF93f1ptRg9xNyAYyEDYtb4IjTMXaoaaHSoGOwbA/ld0Zm48hISXiw
UEI9ai7NR26AbFpZfaB5omOkohOFHAr51tNARc7CrqukqyzUKb/+1bjfVBXWIEIKuU97js5dHkFW
lxCqYaJ99gj09PyLeIMLaRAkvsGGBmnJE7E//wfztE742RKAaaPrFuecl2fo74IsWHQPu5MvGT3w
RzHWKgbkvtQIrgebCoFhGtpbYOXlDw618C2o6Uw1LIa0jo7yTD9+PMzdiEzjI1b/yl6RqYaY/ttd
NouI2rFz/QQOX7CVG2hYZYMVRPaLOzsqQId1eg8jWpK8q9aYUQ95BkjYr4VnTEvE50uFTqNiOZa6
2Akl6B4xdxIsodiR6RgUFytYHP2tSIGNy4aqtaKLMpIRyVlVUTNLQXTKZNTqhferG3/fODKAep2o
aCmOyDhdxLzbBgOnONQVJlKVAnizsR/HAlYgzOo/i7u/F6LtJpPdBqdZ8YLm+5NahsLFYVO59wjK
C8vo2/hv3V5B3SBvHnWMeNbToc4Actxhsd/6vAGHx7lgdp00DCtQ/nEtLCqery+lDPySxDHq7XnC
6bpmyt0/8jVwmGju/d6Sl/pXsivVNxOTyXPem5nQsN2LjkcqUpRxL9Rgv1Dft05CGuij5fZW7h8r
K3hRHya3mf5NiAo+sNqvRTwF94fG7pQyKHQv9PyLNc995NrRib12BIgWRaytzswKduQF/xeEb72U
Wmc7jYpUmr6uVo8uBkyb3bcgCj+wg3yPxJ3Xhfdadc2XdNVKIDO48J/WCPN7lUXHLN+bgrOlu1bz
h8ZJb8weFhpkOCPT4Oc5PR88jeJ1N7J3eGUiX+BEGzOryykRr/U0HyGagDgxEyFBMMJA2UztE9Jv
gp7lmX1Tt28a5+wvd+NrBB67kJivxRf/mWFJAKhluYfjV5ZWoP1/A/qzShcrKEyb4xqn1Y+2z6/j
5i9AZ30cow9XPGhltkyI0c9XKMRwEWMG5ND9v93m71jtm8KlWnS/4AG5t59Be5q7B6TiPA+y6oZs
bjvuOwAWCGfWuQlwr7/MFGHdgWjwIbObdAIdqQx7QGEPqU/6hkT8WqTM0GrK3laUSPDcZRrNgV/2
RXDFKUOzRp3/BUh7juc6ubzYU8CZnexYdfWhnRbEl+qS9amt0nqgQGd0xFnGxw1hM5gsSdI3C2wB
qDvDqzVb2OYnafvwUZXWZsRcAIDDayByThrmkfp35Vto285hTPk+mTiuxLQtwKlC/Rst1xxLOkIH
jHDNMVoJtRW8H3mmT1acL1vvTQTs1d6/cCIL6xTyjZEtogEImeKgI6GzJg7OhKgNU2RJubxIjGds
YRj3yB8PmN8UgE1pim3jrOus7TNGMs/0sI0ygpESHtK/A55V+7a1AuiKF/mc/PUoKIWEvR8UsIXm
Hrbsg01AtksyrbZFCWPzNSWt/FkvJgRRFaNZLQNwqw/7l9YEyEbCVs8KbvjfWbPz2PrBWYUuMeeJ
Zg3SKKWi+BOE83lpoE/zSTqwpVucVV4PWgLQSThKCOp+ih+1E97b4ASmKNB15CCc3zfp4ICsJqqq
h/W+BT38blVJ1/X+pnrFP4oJeOCaufAZ/WPlfA94Z4MSZSTrLK4M9FyLMbaAY0gAOCpoXIqwV++I
1xnFAEK8SqnaV6oOuEkyPAFxMRZeAN4E6/kCM+U/aGcKemsmYu7sTs3gIiND8Xfcg7HH0Bfba5M3
QYo+1zXz+v6X/SP24ts8nOI/tyycNKYA4mBCb1MlUVrrUzLalX+K9kMPsOh8tYl0dMmgwGZxYFtH
VC0wEgpw7S1kujvW5Dieo/56DDu5L9ugJGrGrnV/AWVmfJePf8NOFv1zPClMTCJdizw/FCsjjK6A
EBaJESs7HzgK1PHCg7c/oE+CtiHwQyDQUmTmWyzDehFgstOINDHb0LwAvidLczmyKt5dh3nFoiVN
XZg3yJj1XTjpinXmEFV6AJvb/25zpaGZpqbo+u2JBczTI4tA4WDiLFJHZRYe905SnW7S2CAlneCH
HmQmSeKX3ZMvoD7ti3oQ2G8PIvwCkM8WzuLyU4yWIRL8Z04ot8GZo17CGzsYUsaGUTw+TwHkW2ag
s7F5HenxsWyioI9XfreuO0gGux9rwPpRwA5Fbx2F9u1q09I2xCq0B7L4HxzFyd1bVi3y5lDtiCh6
uW+QQu8DjnXiFQs1BiGzS9TLx1iIuyhb94cR/MYoOh+6FQjw7DjUIAuYzHxiXDZQYvK2I63vmGHf
YszBlloOzLyOQwc0wFmeDJbyom5KG38C85UiCptv8gPHRm/hLDsZIsoXxPOAGx3v0Ji2MaZzJ1HI
jVKolHLmqTOJhE7b495wGvcOIGdzFC7/kaFrCYNIdEHFOP04B8IbRxLdJ0F4oWzmB+Q0ah0GUD6c
JeHtAwUR/fOW1YPRlHqJKSqw14jZaMyIDookjA5MKeDsz8c34e9EoyYoPkD9eD+yBIoCELnr3zkX
hWAppBZnNsAU3C79hzmt6FfFn5PIqmQ43GyaM4+ZVLZEsaGjzDk0m0eXmZFjoVsuzjZ0eYU0xbcZ
ZjrjkGmRwyzO6e7mN5F0lRnkcrkn0N5O+AZqG+evlqT8E4DEiD/le5FGqz/IfDQEzW5tDq8goxqB
Mcl47HSoHi26Vp0SQlSAxfuM+HlF6/r1rzIZPzhqDb36apDyWdmLKpjrnTZRhSWdJogMiSMvZP2x
gOVjg1khOdgXrqgKmJHGdx9uFtEsLayTGNQg/C9Oaaff9ZyczA1VRGUM65txRiZ7D8OYLg7mHrpa
tZKJFIl9lI1lnd1yw5w8ro6mSSpzAcO7SzMHCOQZ2xDpVJe0quxUWNBcjY5BGDOnHaJZMicRbhWw
GA2kQ9z7X3v0xqPMVMzF6vavXwwLV+Tl0LBemS/nswZGW0RgqNTo5lsIVRYopr0wdDge/J9h7QVH
WwH7Np1a/l2QGQrOiddASlJvVZvVyaGNUdrjKTFrd+eJUQ2eb/QWQ/+BCDCBH/9baWBtobFygK1U
6YPMYchudzekOcwpi7mfcUqkK0r219Cx343jSgM2zbUAVLOI5JDQ0HVZI2Z/Qhu0qEn+RHuutadk
ciLclwxPRf+bd1smi3PMuSB2TT6jPavQnQ+UxVAsXOx53HJ2mD5K+O62zxanFkbrC+7T3hX/h+cw
lb/Od27q9qlaZ0CjK/eCo2hZFqiu/RPAcj8J89Xp2/Z1c6C3m3l2bQB2G4qqcWNNv783rjj2MDMj
YrX9rxMgjzk9TgDfneL49tiyHAG1OjFm2WdeXU05EH0tXcLZ1DwD3GP6KvEL46+Uj0t91ice0AwZ
oeIk+RmLh34w7SksDy9f9xODEsCOkVMsvye1AyxNfZbQqMWUAj5Ov8b+yIMM9brMraZ324Kv9FQy
1FJzvD2/aujASGvgDksZz4eNM16BxcYWJhUWwGRTtMHvZztEJXqMgdrkmDcmSRXLU739/x8XiFYy
HyxTjaIpDETV7Vc1Lt3f6HqrAG1F9I1CLRm7f4zLbhTyYF/xuLNJx95ebpQi2HkdqjFvdCI3Wof4
zPklGja7kQGKhgGsxO8vmIlQammy3MRklZjGrIFSKFPbGV++gceDIjaeSX1x33w9NBwGPHuDipui
Ac+7usvunygjMRU6zmiTeaiXoXwfoI0ScPFYrjPtUMvfUFPyAK7+Xm1T1KwIYVKh5ZHMe9V80WaY
SATt0eCng6FZ2YltyaZ2pfEHQoYlicordXXvwPso+6iLTZT/b34i9Ff7DFK7mt3cE+hOA/j1Nu7d
b6R8SJ8O3OdMVxtcZzNrGfdcYbicOvH7fOumfDINpc3bpva+AGJIv0kNkCuJswctxPf5hJ3OK+PP
tl61Glvz9hzmCtMmkngZxqLBe7Hay1WVqu0xpH2EhC3hrbCEd7F3zBx6lMtb7yStmDExDQTZC7kF
0I7J3v8qLAZ85gWyEzQ9TVbLYWHzbTYHvGIHEk5rhVbNDkbEJzGXt2UhwRUWh8xhyfHI7zXj/CMF
zDvT79+XxBRvFtHibv+zkd1TLODNTI97GnpMFusnpWET4JsFX7ZooD/QMG59SDrs6pwC2nA+234/
BjDc8xoi/bdoXl3HRvn2pKwasFPc2F20vJbe6IiwjX6ADxPyBja5sM2WuWiOUqVtgzBZBeYjlYcv
Fe9dP6Q8lXmghUzzYBPHo8h01WiYgwUJ1ZKbw0OBn926UYOI/P9R/T0rDkM5+06Iz8quQj36ZxAS
zfwtAYAJvXfZUAyYYNwpxCAf+9LlAdcSyH/u38Xu1mXqEzMUldwI5JaOH5DVL4XMFBJHfmya7aUA
55wpieMohUFXJeMKPqQCzKHt38IyQnOZA24Jo439woKXIZqmCQX9abOF0yhgsphZ2nDXMk5vqz2Q
GajpL/HN7rFWztqXMWV0dgJLvfnHZt+yQMp1fEKlD3YnYtQWVk/gfqCCFZ3ZXk7W/7yiltz59hQe
M0o1XgFLuvt22zKXP3xHnZdKqVO8G2hNdreqxV9WhBwp5Frk6/+bbJo2p45MkRmCpN98eEjJ8GbL
n+oDGxx1LEzkzRQhQvviqPVyb25L2XdPSNnHjl/zEa+oK+3JEBTc6JK3aD2pXDS63vTzDCOiv5Cs
dc+muenADQtAaXsKQYH2Llsod5ef97DmotmanuYsJmGXGx5BjwEtVbnDE5WP3mx4/ayizwS52jbj
RN069OzZ4V5dMKmhMEKNjXHxFArj8Rh6I5T87rKJ4uoI5iV4taAiR2qeHucUzHbj3LamtSg7UpU0
BdwITw/08qcvZZJqzJch6kspOD8FqkM/7l+IYPspnOkUht0QS/yopATNtYGZzXAnQuxUt+X25LW3
C3/mq9zXe+HT5jKT4zcqgNbTxIKourHJr2ydA1e7opHzFQ07d/0+h5J02wCg7FB91KukrWNNIwyW
9IV1hJo5hc1UJzwofnY/VkVA4jytpnlVGnnQ+Av28NUjdDQcsPZhsryaZpVeQ03NnaED0kSFRQob
0rb9uj/QWCYtv13UQRTFr0yXCLIzUUzVtoZj8P0XeKPxc4Ew4dJ3s1Z3TAVMU9+Xc5H9IFgewsC1
ODPujS0kJ62w1n25UEQ3gvE1mBkZ+W+ZLEeN8AVw08oSEwreajfV5oRmEjUuyjQU7CFwhd+8le5e
9//DctowmkC82bhzQagh4sal5OxZS5gzgT8sqipiP5wskbrYecblzkBuzWqobzIyVTIUtcGPv0Vn
sfGr5qu5yC1xgZUaTbJb5uUGwFez6q3xj4lP8lMOgk8yPtFv0BJUQ2J0C0v5n/DHK/Idku8A80ld
ERRZdu/hQag+Ds6E9dAFAOGytFyGNYxzfJmKOervLJGntp1g01FXkBSvfd+n9tOwEM8h76hXG937
WpyJMA3iR407M2ZFLwrqTHS/WauNCG7LMKu7H1Z+Qn8hYAn8a6PJDLfFMwC1Mv2SqykyxbRqeeuQ
u3MVYLYkvaIUCd85J/VvIS+I27gzxAPURuqiWdzfzEMxaHpBWfACL0UtRV8d8HJojtlOpYWjIsV6
utLz5tSvYrgA5yy9psu6EFnoSdDYXfYER5PegGGuJAaN15LjeS4vKrzOmY1xKya14a74lmhfaLHa
HzZlyxrBoOA0SJm+v6yi185voK/e7SRl4yPqBAeb3ede5m4Ev95zk/LTOiTlrk0FPpGeJ9DNLAAp
AJlAWHb56jstSni6KmhYPIEuZ2uetAfQW/IPCKWTlpvJpq2cPsps8KXwiSCrv64LiDeZ/7n8uHn5
vmj29kpcfg7P/8RhH6msgx2DSgtCkObq+6X5afcPLuONdKnptfl844to9F95ikvuOgvnKHkBMY5t
RK81Hj5IfCh7+5e3m6ttVlTVoYT+oQLgnzC2BxdDlhBmJIjtSPsjCWYwEZLQZELOofSZ/BWRbMoP
g0KTKqP6UqcMtIbs5GHLw7jili6oxC6QbfGf4exRhfXkj3jwomy7wrMoxMzMVStpc1RcQNfFRqeA
WsVYTVXyCUJRsS5FcKr7OTkRTBbz+SyBGrkwvi+iTGUvR3Rn7nI+azu/KVZ1flSXD8oxAsPraIKm
vvxx0ANYsU0yfJLOn0hEMire0Qoc+UpEN+Cynx8nARr99fW7MHtNEXqOEk4zrW1O0xZWkD4q/KvK
/Cj6eMqO574+QGlwL9+3aomDBJE0a2Dhl/yagMUlHrXNC89QRsmYqg9MmcZm+lPCFsc+VMVb7yzP
/Fcwk0jmC9aggLFxPmyBFSabWN2v2EYHQL6tCXkF6aXxgc80VRdEZkEe9RzapDl4jqaHvWOtwdfR
c3/VWKVAnropDAftAvVB7+NlSl3c6rNr3WQFdeI0Ir86kzbI/HrWbDZZr1FUuyOyfe3KuJ57g4T0
7PRlmX6VdCaQReqZ23oHAB6VlhlUPUVRJIs50q1qXuvX1NRH4T9OS1ULpFIhgWW0ooBDx7rzThvM
PZ6+1YNkQqJUoLZEOP5/JKohUrGy7khLG4jK+IYoFtaT0VC/OCsivlWHJsQzm4Fh8a0g4IvLeE6/
DKv5TYVvn0xNKBudK7PQrn19KPgcHvGBs8gw+OGf9NNl8Gkja5Pfe12e8ffn5jiQxLb7xYgCw7q5
RDxcpE500/rBZQ5a8ohYI19llrT/ad+PfOPqpr8oYK+P0DIvKH98XNAAeyUWF/hRdhUHSKRdHK/F
PB3/QW6LT7pUgdIepvOIb5Addj3F9QpUigbX2FeNvQfFh3k953uScdHV8QeTxPDQPpzrVtFZqdSd
wRueU8BA/AdTPsxXuV6h4PIO9Znen9bnQhJn1WLacASmURO6AtCMIJ8knOEyN1y0Y/s8gh7AAa4L
o45z8ho4/vEFVZ+eOg5oZ6im/6GurZ91HSJvB3+0e7zNN+0dGgeEt+mrAu1mI5orsEcibKgnHCxu
mOHM6da7mcSDu2vPta24RuXDP84g/cD46rjHAIPT/7KTPdGLl6tMJliNb8peekWgwxQ/IuAuP8BR
eWDxGdg1JLQoNFEgjkuthONn9F1zUeqmxeknFYamwvz8xKQ/4/M67SoYTpHQ7uGvTRIEuiP+fNBT
PXfee7+8JZKI6FqSIwvxKAI5ivJ+iAPMXz5L2BT+MwoBm/Zjw3ZomwDr9tyXLi5RSo6r4XHnH17T
H/P5HQ5ooMXo/iUBq+/+69ROzQXnZQDYZbc8H5opR2jykiZHhzqawhU8I9SJGfMO9PTKG5ttqnNy
ugWV5GdqMsiqPJ3kpdR732SkAj6Li0neVNp5JVNparMvLXoVb8VsEXsM344ytXvP5Hcy880UbaRz
D89FtuSqvefYdUFb4JIMNtfhL6PUKoPLxwjwe6G2Wuz51nQil/DMja6CNxllKX/ttW9pwkRbt+nU
vD5GCNYNGZA6qe3U403B7Cx9H7i7qaQZZ8zbCBhlXShCdXrn0Hh2HhAhPqEry2b696+aufwcmrOp
IW+nQlKRcTv6HjfAEAVGufsfcYJ8pRA2hq6pHkEIOBi2L+IazQFBSDzvPjb4dwHGamOB75V9FWfN
oemVu3dMOcoApZA7FZ7cZJcfPoErQZFkX+rQs4ZK62HHDZMFvn2Jmaxh1Uza381H7cSe2TZABl07
cU/M44SDu6VLn+ZMbUcBqWR24x/LETF1eppCsjXSL6PiqrKBhpDQVPW0dmO3Ro82Bg5RbjX2exfD
gDBnCI++zXOB3s1zD4S0uPYQef8YPOVkVTYyBgBL0EYtgv3iHRPhUeG9hB0kMc87+Aj8KY1zDQnx
OSeynn8z8SxvbG20d7oH87bI7LgnWLAIl/Ic56BS9/zDdm1MEg8YLAVIFGCLgGrSeP7ZClZeXxSG
Td4wJniQtJ3si/Fe5w1J+DL24djtZ/nD2dt9mq/P+QRtYglT0wgZWG0AHFSrEDd3Y1quXxSw5e3G
eTPjeRli7vkMVQF12Vu/a5FrM/8vyFzfrAjWr43uk57uX/WV2qhC478b/j+JqIs8b8s3aD/CNeQq
jun+iIiGJnKpAX6d0STHMjAwu202gfCW/iRMqucvR2osRRtkBdRJNREGaoQLty9MnAME5lD1TX3G
3GDlvmNfAV+aTxZGmqXh2vjt+2iU+6oi3pJ6AXFuMu5FEsu4UQQB1sTkfYcfiDYKhEYAcoIfySC2
WPJ82KG3gXuJ2kwRkkOJkYdY4B8yS5pgwJZzVgBv7cCLMfb0CJPmmBU67ls1dSw111g+UOs94jhd
yr7kXe4bfurxiPmTtm4ToH1olgKGOmVspYy/H6lcK6dCWrXvMiPKjJFZH18iAzF0ATVJFkniFq/G
hrgsTSYjiGcj1dplVMESOC7FQK46T+DTqSqEqHFiD1zwG2PqnTi3+VE8nwiY8GUltpdKooZL6x/d
RwRMotWx12olZMFq1W6s+oymDBJBW/FLMJy4ty4iTEGMq6X4r3r1BRJO0iM2qVzyD0MlDmJEMlrb
aHNZ183T0JkHJXZXEyHz+Ao8wvR+WLCmLEft+fa+tnZME8yLE8Bg1KANI62+h59TjS3y0nK2y00C
LDUID4T/svXpOOCbP+5DtA/NYRfDutmuQI1T6UQgNwlpjUvk1/RTdlZlVO+iyEX9mnteb5HuXtHk
uVaaQJzr9kD9lg+6Wsr05m9UX4sRFQgmBbYASPdczgszSyM+UxJVqpop8bgFS0e/+yEjQhtimHXl
S9Y4ploHIhJSS5wGIOZrYsSUj7aydkLZjOR/1dIn4veupO6JLfNIxuQ9Zk6bRu73m6At2SK/s6Ha
cnIb8P4s/nyU+Zx2D88tnTfJ8i7JUCzv6aufD/nQ/W2pomCsqOJbj/Ze6EL0ouE6p2yiEYxsuNWV
R0YNDa9lmWN1NeJanJv9+YT8B2dDfdcHVlDySva/kfigkzg+Flr1lMMaXJo+VHE9qzBRhZcWVBZo
O+ss9cnPZEygOFz/RgZqioid2cLX2qxghDr1frgd+S+TiX5pPPFmFoSQH0YsJ9iHfdw+QNyhWZMb
srJHTIoAEAZ1EIP+Fga2vTJ4WNZgKLDMXCfqMvjdBj6CA0wzrJ8WJxxjye5bUiA4UnJCqpX540oU
zBAiSW90EN89D7BJWd3sD4QZp9Lb0qLXdPfJ3Ndw2BCT5OjGRls422X9oNDQHUOsxwsXkNgY6JrY
yJFry7V770CWYH5vW1+LtsBi92JoZ87ZomH+x/QY1mqaYYBs5U8v16eHYzwK1ZmQFzGAOBaAaYc0
4rWmszXQF3jsgaPJ/+Qurp6M/suosCU/ccQfZgmhM3eFd54vAPYnw2J8+GqVr7vJaC5cFrGugIC/
iTv9Y1bDX9Heo7Q3uzVb10g/086UAh0aYBtdRYnkuQ20cASIIs+ExtDgVUZIIeclLm6Gpr62ec0H
K4UOPt8qA4H3TLKj8K2Jw7AdqVv+JxLrXkMfMO0CIXfzG+/kWfM+CJDEXIJX2vIbzBGR03+ZwQ7l
PE+asAm14n/BZUl/JArVeE63Ie9Gj+PKg0ZTy4rmilelwp+fF8pDggWxtYZnm+0vjaRSqp87Ug5m
cl/oTnOSZ4B+0e6P7pUjXmwSB46/cy6/2uWvNBmsLbiczFYUSvgxYeORQcHP4BPVC2tqMxY5REZj
pydn07REl9dRWqqZR2bjAdOXLSzi0VAdKrkE7luuC3HDw8TnQG5Qg41D4EbWX8z9TMrXFygvC+RY
8GIZISw5Z94kem+sda8z5LI/fYoJLGowKFObl6sQhyW2PMazX+EPLNPb4DnMjyaBwEPoR3rQ4wcv
mwy2KvtySRJlHLkFnIjXnOBkmizUFFkVM1DNhCZhno/hLUkuNkAi6cS7xmO1c/e351oUQShmWNpy
t1hi1UBf5gbWp0pKA5KBoNDxjPQ5a7s6ylSuEVNYcCzQZvqinwEIX+YkCvaPklWZP4SyUCRKSXo6
K4V2dJvvci+Zcv/PvFtpjCS71OEpA8kS0hr7rkJfUr3G8UFiGn3PW//yTiZLEeklaWcWEl8RTWnD
WVH8lRYLxTrLDShLmyVjqfCl3FmwSjykASuGfF8EGpjWdRwG+MS0tjljFwMfHht5KPXb+Xsom4vo
0K2CjWn7ph0meRz2VVzyaNauzmnAHXTf7cL9y0EWkuU9xOectYKXQQi29MaJYmKQ6aG7404IV2pz
YPbzXjSFfrwOWIKGONkRvlzmuOXRCVx4pR+c0VhBxDYl3fmTcNCvLy8dauJsbsHTTXOFA+UwEk6u
pjbqmfuSs99ue2lkrju18hbBNpPA/OK9ZqiyyHhERBjaiTEz6DiMH4SkeWg6DQRMGIYWOjeXVttI
kwmiIFFkzlRZvRI1diJKLUmWtx3aU+UyZMKqMBHXyl/aTnQQjuHji4/IHEB8nGQ1LpzLDdx31jn0
WRbngrEt19tDeiI+5PTwSc6iRfGPjT5WX4k559heRagoyrtZKHiSA8sMOlOckdknDMro6b9nLzYJ
Ecqt4yTZ/6LfP/QUDBykznmOzIkYhXMC1sYeZJoqom9fQUw/vzU3oYkSayIdby2TaQlGyD7hdpEN
hBOdDUBdoBtqPKU10xWuSrZJOnETMZDSWmuiNXMEpa3TV7AiMuqC4CmfWEGqPk471II2hndSjYZO
MMh4nPnuyOa/z25w1ztS34Q1Dah5qncepDO2qsfPEkANlY04y0PfGdPPn3j77RfWKepQuRgckG4I
KRVtdCLwQPVWVRX5wXagoXP8bYHsQM6HB0N+omPHQLYqYWfdW4/WANCmEx54L8FmIoRGqKj1lqkC
New4oXGJk1nnSjskmiOXUvO+doHWwESAevQlOQ6De3HAFrNp+1uNm9DH5Ptm7jGOjENVkB8COBh3
/SqMJDm9og49PkZZE5FhQoZMSN+LaKfQ7wsLYgq0HS5cbxhkKHjO+C5hHAJCHEPEBJpxyb1Q/kMC
zrJEtpSi3MG3eDNJ3LTDg0NreNdfcKKNm7FiTBDYpI+1iYRZLgr7QZRXo6ckTv9XkXgv+hSe672d
o5yr5YPc7VUtArU18pB6ss2mOxf8jmWDAhEOukdvwDprXwRdSDhkwmoJ35Cz110GgrSYzvQGdd6U
QoSYy2dyeNtFhxwuK2vPlV1tPbRGRjd3Yu2BVHX2jS5KhEqyIZPHJQY0RYTiX9Z2PzNRtK6Q1yVk
/1fOy1Vnp8OLwOdrDNmrdl95zaGxvxnRaCZZNtKObH8oRkrihFCQYSR/hrJylyIhqk0LH+0bSlZW
l93qEeAsm8MSxwq+Vs7negGe6O9GRRsfGQl/AyiWMLb385K46V9OT3eeDQpw9nRlKTBtY8AedLbC
DDmNI/7+blwbqyyYN3DM6lq0GEOxIzqwNJHjypGsuWuqizDwQ666YIrc+wVNk18EXhTK4QpX2/XE
DTZhIuTR8l4kOozO3ElYN0hi4IbgQPeO4uEIqlNirzJyJ7zK00KV6miJ1MlR3hyl6P71koL4yL/G
JZzoR/ZFQsx7MPN2RfcCPOBPsqubwa59F1N7qbqmp95QHZ/OoK5Z+POCUcWPxWg84vHu6GDfSfXk
l8aASTEVrSwAZo2szPpISYGh68+IolM8YQxNBM9xjCBdLx2s2kFf7s4ScQmKDPPcJOJipxD+RtQk
O8cKoD0hMJEXvs4zFogaqGxbtRMUEPMiAa1tKoui0WT6R5Bm0HN3uFWilGG2JXhVbzz0hYuZQbTM
La7S2rimyqD9CBj0zb3/UGioCuWe4Rz9thmT3L/3e/DWSW4fB40ioz3iovhZSBG/kmMPhlziUkLi
cqLGzudy5EuM95YsnhIWA8JihCjlzhSa192yVdMRvWJSp+dAc7+o75QjTwZqXdzUKUXEj0860iun
mqkWVJQADlLeC8rXIP1AAqBeLHNjJAeM7LgqJesU5AUQkcwpzTdTBe7PRXiHWenqKnwR+0h0G2QX
nkMVGXtp1ADZAX8/1SAKils13UfJhxppYNJSpKKFtxiStYluBL8A0S1uBJO7k8AINfR0VwIdMByE
klCnaT7OhfxIRrN/zKNhEIZ9wyVySpLcWe5pcm1AmD4RdJSuQ8tZ+oehpw+6mQAqFuyax+5wNyW+
CEDoG58QB0vfI2P2TpZKoLG46PW7BSEA1VaD9a9VTY8P+VKjSBd8k8g968Nezjic3AqtGKGINWuz
5LP+kWxk8E3F4gWNPv65fWkbf/N53vrAeXFyxjFlstZRMvDi6PeBR39gpy1nqcP2UXM5Mt7op8SG
QC605K3bvUj7p4MrOnMoVdylnvOzZC2CwO5jewXauVraPPtWrI/j899rPltsX3+f+WKbxmTqBeAZ
JAoCNqusgKPCsTGilmfJc4x6WZPOzf13o7uMX7ZtEkfCAUXxHfGn5MAFeXvAZQJ1dARq6DU8YCwt
a3KilxA8DBI7cmf69A9yI5AyYKFx6fb9d8URdOB8973aiCcbR5FCwuD6AcLnRSLU8AcEjfz1/cDP
bzxFpZs4oHHu1VpTSsn6vq6bVFSr5j4zqXL5DZUEuzQBa+dd7vvxmcAAAXvW3OcfJ/RD7kXFFrtf
pP44kgdD8JzE1TVuYntLkDx5U3L53iqEOCbqxm+ctPVqqXjCjmgyGAnxTkgp/hD2AsoP/TbzhIQv
gs3Ob/t9qLkzcK+3Fg/lHCsZn6bRUZskwlzmnMKEW/zJn/Z8RN+Ro+Rki6eLDyzzzp4Is1Y6wM5q
qQb6wUARTB9fHF+1irIv5GAZdk6laapY3QYrwA3P/2z5qsXgxq8r0J63MdY/cYnO/55ouJWnLZtO
RSQusG8p7qds++pd+HejZtJZyC7EaxzFi+KHOm/Rt/p7Hs1g80B5yeNGzLY05syPsNGpkkEbFQz9
pAD2cCsMAwDsMg61EI9g648hozh/hE9U74orHxdiWQH+seFxl56tDI+zrG9lufF1Rtc8RNYiKVd5
MIbv/3UU+oO/ZcUAXTMjJC6JLSPkZW1QN8UNhpcuvPBJHUgcAc7bdydShMuSa3y59LcDbK9fG0Cy
HwpzKgWEbEgrlofycQRLYyH+xOuoPD/NKvJTKo81JdPbaQUqod5HnnO2ZVstMqEycD+pEpWnm/TA
S1l4l1y+N+o4gHtNygwgIxNNBaTLkloFA9c1Cvs3dEpaX+3+6R9VNUwB+RRhyEFOu5qIMkDywfma
DsEAixMmWdpzk55OTosqwOmwuQZyL//SsIvaucIo6kuuumJn1m3Zoi9eXtauxTwdhg7rLBspKRwK
t774OCEJKdoXRxcMWQiL4WhDYoPNrr8p2rdq9D7gEjgJlDunE2XkBLvfB59urLboQ32eLXdAy6SY
+IZ0fbRKdvn4CAkHqwmC9syRYNzwVh/K0xd7at9Q0SSDHzfayt4Gd6VhQTzDhrFkKFJQirr4chit
15kUFKQTFD8wfXMRPkF0FgXLboNxJe/K0BpekXEDElQ5MRqeQ3FbuXX92dKZPpmG34berw0olkho
AUmbNb1FfjkSyTYAKgzgaCoqo5axzpYnl+lPP5KMRayF9ouEX4qHvGWsW3K3horDowgda8pizk6f
QtdD9MprirpsgNHnHqIUNwHusiAmo7cIn9glJB550i8g018JK92NdrRQXY0aaLLX7r9QkOr0CtuI
GfzOtJ4ZtAfMGb7E4qeP/Qp7BTImUOIe/2BY1OeLnMkbmUdinR6PYU1f+qagJ0IUP+1wL23Wg9h9
RPaj7fKiBK3T0Sg6xsnyuX7KGWeDRlsouGmpN8r0IVFxpCcNx1e/egByTEY3SwULkO2Z2+W2TKVP
6JhV/qkDPTBzBlLObH+PD1bt/P0POtHBYLD57f37CFV8hLkAa2hpc4VvVdNkku5QuwLF2aK/K2bo
1ov47W9mdqphIZkIhZ554rV9gLxCLy9HE0ew4R0x7VC+3FJngHYKIsETfRBuYYK6CPUqMOCHx2oc
hd0MnQNELPMsryJ/oFE7+91ixZ89z5BQalXdVRn0wKfMNzx17J5FQFNlpJqoTBT+LFwUhgydhMA/
Hd+RSt/leq5bjkFZ/wMVN70S5dTgf1GMixgbpk6ZJ2FxAVf1E4ihpVrN6yEPZWkefjsYzdB9Rm25
CXmUA8ueLHEdOX1VPWHIGpg77hFPYRNGTV93JvxpZB7I/RAlfWP83E0q7qy/+Kb3ou5WUOc9vxwK
CCGwKuN4Su60wO55VvW0h2pn7iCoGgqWi+qYaqK/ilDNViEBBKOqDxYZf9aixbhArBBG0d0GQrcm
MmYM9Jdj2GeqTiNxx/l14v5lW6mwiaLeqTbsXe8/DTWMGcAV1cE4kac3YV5evW2+kwATxJvqGaM9
eCfg4iFHye6rtwW61WTQ/zeV3PxdqcrVzfjdRpAB23kHI5pR1x8ByY2+pZY7wRQ3S9vcG1ixAurM
JsRDVsFoe+BKQ4vsPOEeOpA04gBu5bqAZaqKElrNwE/BsMlTO3zVIO2U9likgwCC1bnCKSfcfVbn
v0zZe/mOuwy0FHc9OHazdQCZoUGV1X++JSLKViCn/ENkQ8mu0nQvJAMVIjrr8ukcTFIk0qynW56k
/jsywrA6uEKgsQ2R09kra9mtVw7Pqd7u3tK69iTnI168Ts3hTSBMGM/6o2RPTMEL/UJr8JiJgEli
+LPUM/xaCjlURpa5tsAXtoCnoCW39kAx015U+Jl7c7mnjgxS/Z6SzF7m1TQo+rqscvQBLv97UHn+
uHnUIHIxVcBttAK7G0XrpAP7EKMjnWlrZJjcainkw1+qBsuRe00hnp0vGxmsrsaArhTLw6b/ZZWL
YqJySI72TxitWPlfvGSMjnHBPM7bO+e/jm5tcumf92Qf7JzA7G26iON3N3HUz9bye/LJAVWZB7IS
bYn7hCafo3vednFQ+dUOOHKS4lDuF1uVQeL5WVvkc1bqGnulKNJENdw12rkJ7gAgS95vtA52NAH3
kngK5ToQ4YCTzi7TlvGF/vxgKe0amchLC/nAtQffyVJQ1QQYD9cB3sOmT14Tivqz+urppcY3b9ZS
QZI82nnmF81oUBHGumiz+JGISPt651806DSYSPv1v+wBottL11JUve1YmaEMbEAhUuQ8cMkIWcHO
5tWG3nLNujNztsM20zCDrx1xmDHjMGRsYtCRD3mT3yjh56gcVqXPv3+BIrWr+qzFaWMFN1hYrLZa
1om7CIZBAIO3IbrjXrON4FZwSRDrYoyjvsOyESk0Iegn4YzeEIiyUH+E5A6aBZYNVC3ZIwmOZxnk
/J9obzmcXnDoWekmmu9cxcpIy6qocZhSEP0EZhGsi+HQUp/p8FsQrilqLPEsKsUqXE/G8GaM4Kqs
LFkcoeb0886hnPmiJZkgw1FbzDl3/xgdoqG6guyArLrGxi0iOw1TM1Zrj4k0ek0nyetsscRK6Scd
j2titH3zbVx7aZOGYNhA1FXliHWX0owrCl1u+uo51CO9uWoJ1O4mqfYAnUzo+44d+3Irs3OTIT/9
BZ6KnF/uTPhlhYCk4KZOCu0iz5th5efVPYKzQx0aWt+usrI0K5NwE+3LBP3bbbrWb1w0/EMZyd6b
0amHBQCVr2fd1fsBfzg9qr54kKd6mitMQrpW8HEi7PTe7+j6g8zUm8f3cihcnR91wEFxh6TgWxnL
tYIu7tofxAZzJVCvbCYPzNnvMgIbTSchKgb7TJc0UWtdXRiT402U/oV5Q+S/XZUuW+IfqWhOLafY
nzxDkfWXYyuPMtnG7uJ1iqpspj/6rRgdDke+DFbgTfvocxBsPYLbO3ouylx2daJykMLlO1NT1Qpr
ih2BZJvtQ8hCm4LW/jngaXU8Odut55jXUfpNe8a/XxJc4nphi6BCxrA64yfPMBvlG4KmSHDukLnO
tnA1ghkkl1icY8olNtrjPS/Br3P3pBAwtFLYf3/b/70iDbO4rFKGXIqHk7rjWK/yp1fLY7t74qcl
he3v+jqIUmuDIs1kcrUbaP+W8igpwZWiGu9xDIRLriWGbyBRkbdn7tQBLsMr1RBwifxQsJ4ted1S
EFWZXjTZoGgf7L3FvX5iv0KeDE2np8UFAXGw4stYfo494NmfuyndMZjdWIqCvD+xsKE1OEdNHQAe
62w9mvZxLcZbcyUqlCvT4SrvcuJrOh4IPZ3py/K4Al2nTAm+343WqSnxbTi6zxHZIrRGrmfl2qbb
ZiOZ78XtYK7glpfODr4GVpy8cAa6/Ho9hstYJ0SNTo/x8/hFNEhCsMCC+i9Xdh77kCOWe3qdW7TX
1mdtBdhjOnbZDInwgVbB/msJWdtdRve1I/jodSYktDacbSZi1L9c1lpvWlDWS30iAjeYe7i3Acbg
Svmz3Uwm9uBhjRFmd1w8R20VRT6t2ZkIQMUP7daPyxxGldt/6y1ZPZDKAELxDS6skrF8HVig6cXD
Bx4B01TS7ugupIVUX2SstJbWbD08r9QwbtShIV5n8ia2D0Erdn4cLgVskSpMONzaRIR2/NJ1PDIS
wMTNw4pq4bdgdA1ApjgzfFPOgo5Qnc4kafpHh+lg4DG5rj3FEDInqFPTnESJedN96des9Bc2YZfZ
1DwFcQOITvi8/qdT99lkt/3LlkZG+LNIemqefZr48SRnBxFviY8MtgEHL20biOykBFmBP+7IFmdm
F4D+lXlpgyKAxoG/d4UcL7HIyj6AAFhxwJe4TrFJ3ELLka35+ijv5Sj7p4YP6GCNRUI6qQq4gXZR
9UiEJ+eSpbJVfMtRcuTB/PXDdRiF3rpvJM2WDlloQC+b09J0/VzLxLs2+Se1bBD4gYWas5EmdqRX
zGm5EchCdDftulPaHd9on3ViwmKo6vN2fnRKkZTnFQsaET2aNlGN5kURGNejNUrW9/euV5hgGvLu
xkZrCdxRXnNcWVn3qo7dTmQtb+nHl5/dRs2VlV6Vo8JMWPJ9ZZlN8pyIW4WdYDFVwxUiZtHXCIJ7
9qfxXb6f7q5yTLuEFL75wJkI/2i2Qg6f8wZx2rbcOksd2Wab7nq86nhlUQDTBya5qx10N3MCa//Q
1g0x5R3+nmLaNZiXLvCKOZFpty3C1qwXvjv5AZoR3vqd+0aMXsa5cUoyHpgPbhoV6vMs3t99gluh
gvUJSvCjGIvC0SYuwIWlnuN1223Pn166Fl8kU+55zCe/LwWZACpaK1bE3HZM9jjQvkwJ+KFgwfgh
JbHfTI1e1agu738uqWJDOdZK91xReHadn9I+jGDiG0hsvcZOBIhXiwJBXAECMtWdW2rGhkBLJHwP
rE8Ihs6asSF4heuQbUFUCSDg7Xq49uSU7z5/rSgHRnsQ1V7XdfsnvEhHrdvE2ZoeIHI8jSJufCCg
uNU1UZYk4nj1N347MDw/jU9XNFATRpkDCKYtBRqeWoCBOcYAkQA8s30j4Ec22tD2b/LJU2K4iZQo
+jaNpXuiXs3D9ZRMOUcgtdHKdbJWHVdOvot375V70fZ5t/c4ESmjPE8EkhssgEeXyvB1E61EyWp3
qv1iS3eXiGdehAHeLgArE0M0WKnH48kVyZsVdMG/hoAbkq1oAJWiW5djCZgPW8kRy9QHj9/7JS9C
gPm+zeHa1lKVO+Q+l710eHARHhr+6to6DjmL/WtdnyTOqhUtsvItEOCY0IvWwpEsy0EPxuerhyo+
1lUoAaudmiwQxfnBPHSyusLEALkRPAkUXTR2gyIqP8NjgV5HvE65xquh55lundAMLg042riDE6iz
I0H148BzYF8w2US3EPd31R69zsGi1xDxRtUkrWH90xcYakKe4cgj2NRhyubSKq5i4YxD0zm3k07P
o/Tnd4ok9VypmeU1JUMgARSfYAWl7EqALRlinQOhDjzq8Fk2aL8z4BMhKHLCtVMZEQ/0cjqo9Xzu
ta1uNdI05h6OBEjzsyxE+oJclWUKS8fUJET6+Uhakp//Q9DpNV6nyxI/T5dTE4OTnxtjaYIfh5mk
+d/ToRUzKxetzh25tt3z26z38rCWbov94QGqpUjsDSBarO0EogvqmrQJwXA2udjusiRWd96vSei/
X9W25g5X3CowShUsBl9ZkYcwggDIUCfrOqAq2B+G3yhTACwtTUQTmisFSiJz+T16fZPD9xze7G8i
aFLn4LMtu2yJC90ZxVakBGdAQ5cZdS0wd4+VT1rdmfgnipOzS0uBnry6zK5p/Q49gE0gjKrO4haA
JJCAG5r18IclIc8JfG1l1FyayxxP7kkKd9lcsUklUSBr/dlbNs9isDdPqy0vpydItzl24j5nAW/x
KRcZr9mASLn7fdPFLaokCWvYv3gR6Cwvn007Bw5WMhNjiz22sgdvQeqPVoAlWY5EbtzULML2pUXK
C/cVQXupM694dfctHpI2jIFdpgPTV7qVyXC0EcLrpHdRdy1EU3y5rHa4sDPs3JcIaiY4k+Vhk2yN
og6gLLOq7pd8jCqXwVJyfIvzzv7aMRS76tri+fgFxP9SI3Oq0IAs0Y3XanvofavV516u2K/1o3hl
NgUlvio8OesVsrC76P5D2bFTkR40gR4iw4QOXRLNeHq9iiwEq+Tdd1+y0PcryfYUzed4QyHA1idA
j3KzYQaZdJTlvml0kWOnHOEVt9DnwEwU3A9AoNWx+bhF1gfQx4dIjP/NaFIh/BsEq0aWEFJVkdtW
JJ75AF/9x6veQFS9I4jmThM1VX4i1uMibGTGTsUdhmHK53OzgrSzqwO+nXn4m5TFeu5vEBqvpaMD
cBG9QXL/fMX3iJy0l9FM5kVKheB5bn8ZcZYVDNbV9vnc41coD3tIiPkiRlu4cXwhYEkF14y8sygF
a5pBZUTOhcYsP562gHacmSjBeXVp1YEY0Bg9c/5jEdsslHB2dmoR6SULrw72XMJSkm/0Jl7KNlOW
V5BpiSLguVD3RtxwWpVu0SRlfj5yeTwUg7E4bLYq19iFAY7/JoCrjZ90GViZg+G+8KVrucHGGj9P
0xnHwrYthJ41vkUTapm2kfY+Vvr3mD4dUDe7iwNs6Nz2e92sHQoTEbvJ6LJ87r9zk2QJ7FeoIa3m
S/KFPycMySEObubaAXxXgLeBp8pwF2CQsUA2riluvKWMKQbdiaoO8U08Qk3q+2+e9N2n/8dr2s89
c8szZVk6dnGrnZPayL51yI7+75DxgV8tcc0NRIECntvQp+DAL2x+O9ChHRR9ZhpD8x9n/GjDIXZ8
ycFEPYsSe4h8EeBYL0Wvzxalu7PoOtjxvqxtGr1ITgTxXWww/2yqFUH+1gbV33/vMVym9lKBnEKz
p6DDB+9a11zx5eYWXoTHjjd2+hZt9gCk2Ba3vQiNPSsBOs0q/QEc7Vm8DDw4ZuEnEriCe8q88FCt
PNtmwB7tzjHeXsymkP8vWisC6j7Ho+JYFkSszGeiSKCdsxBrKTPeQVZ6cGP40GAP/fY3yPAM+d2F
TWRU8j+RXrEWwaKWMYTBK1Ox9kPTfY6yYgA5unLn0czQxH7J30ahHO/KSoIRBU/kF/PQ+Fa2t2pe
oTc2MYp3q+sMnllLwTvUEQue4m4N029eM7Zb5Dlqbdrau2rE9VipKbMuXbNKn/VRB+Hs7OiuzCPA
DTm8LREl+ppMcCgBfqngEEKNAMrckXpV30QN3tWVwmgT65pWGd87dCHEbo4ANY1PWxoF1cWnApG5
2i9N5jrwPiERjdVrnEy8P9Mg9p7a0/z27YhEBRjPpmze8rfU4M6s3edA6sTKh4QJN4v3mod6xU4j
x9BRLe6dCTiZMZ9Xm94yWL4/6JzYycLVxjGp4FXgK3d5IR6FJPC0WSP31fizclEu11hcYrD6LYP7
/Vmqzb6KfnqxDKbcyMpAOrIC9ffRUnZX76jmiDcJsc1yCLdxw7On+RgMwG4++bJNl9m4X9+dolF3
tgK7wUZ5zSGlwvF6sSodv3Fnib70Gg87wduhZRSdh5E51PQ34IYCQ2svE3J2OnMrU/f4JZqOVhfs
4p/xuwK8avd/GbkoSMBKCkatG/y26IZ80bAP/BZTc5Xgmf4yz4GemHVgj1z7oyg13I1C2/RNfdP9
zT9RaZHYDavIocLvIh5aS3bOTVXGYYZ+7OGV/rxXM1x0IBsm+s5TjssBxgfCc4woGGAxYhaHZUjW
kO49YxsPJdkm4d0SjvrdxMVUhL+d7330+tOmcUi7Jv44Pkrs/Mcjk9Hv5QaynndDwD2+Eweo/+ld
2Rxo1ve+MwFBj8tkkMR2KIiYAxXDwLjPH6o0KE7e9CDaYX3ER8q3Ixq0A23j2B3iB6xlZHMgzfSl
ANS7pgMwdk3E2IwGZoyyJcZI2Q2ukPzkIgLom7Udm1E1Mz8q3AtAMiD4J+KHim0Lq1Bynn2JoX4B
8MseZLGfIb6hoDGtBnBzLXazxrbdIXi2DFgvZmaZcw+pmoo2fmHFeY6QiX9clVCMJZgTr7/zui/R
lZGIEOqeWa5HoS5P4kjn0Rp19d5hXo3qFJ+vzwPyH1O/abxBRInJvDQn+d+2ohxqvcqlpTURgFCY
gOGKgxSxWG9UduaYQSl//X1je0hRlzaOfMsiCOLpKBz5zCh8nbxyjFw9P6ns1CbL8fqBJ1FekUC3
QfHg7zRC9t5fn4e9xb4qyXHX7a1uFq/sUSamEY4MPfkv43rL2nvhVLXvV9YA5bCNjpLnvzPq94ML
tdZUl/oAoBW+1jEY3cHwCHFofNYJPs8IOziZzFILYIy+GbZdO7Gy5qg0ENQvKNLm5HuBkoL+CNU+
stCisLaGkE7XSBwKIN8+uxIAr/Tx+gAvlm6OKn3C+6ZXCh1OIQCQyw7SzjyK9LOMQfBN22F6ulT7
n5tWvr0AbxIJGLoBvxszBJa+QjiyWDycydkUNYVmG32voF2im5eW1MviMmJCnnRiLsAnyCjYAYlZ
xuCl6aeocxR5pq6kGJHGSQnMp6rfulSjE0hE9fNMM0Vsjp6jFLD8n6uYFP4XPKUwhaRjgce6Pu9T
Dx9EWxAyGwna7vnfV6v+yPzHikqDeQg9YZyGM0XTFg5PsbFuaWzmJWrH91gqFeFqd2f86eig89Dt
NKWGxMJwS7u4pr6maNas9rxQ0SqD9zffh5TDX9G0zl3pVIY7g9MSVm25iDKkIkBNDK2qGG9ARZJJ
TP7Z2Mpza4zg3q7m7AxgihcPKubOvcJ+EDxmp4vTcHCowJGgN9Za9kAaY+e3kNEJkuQZ9Sb+zGjW
O/LCj8kKEtyoCaIg0eFbu/85UNcttQUWf4RXegDcO9aBG3RApQFuYB9hWoBcLEgnKqGA/mRV+czb
GOCXZKv5jeSYDa+D5Fl4rDOoj9WEyiwo3G94kz0uvIfUSO21Ul3jB0zJ99XsREOgM08LE8BYCidJ
9Xh9cSyG//zoGzQ+Xci4kcJn80MmJajDS+UDjG0BKPBAyONTeG700olFcWsM2qJC/oODscwJAyDR
lcdtYRY7MEhafb1zyEwTqtB381z4s09Q6dZP4sKZpRe7XpUIcK3ZEv4JWiyqbBAqfbZyUYuQZuZN
p88qiA56z73hXF80R1/RM4ha0JZFa+CL/m0QdKNWJ2WW0RnYZyQ1IAACzwZbWk+PwXqnbFYwdJHh
CF+nCM9hbmPsLQ9CarkZJ1HchQU60LOu7TBV+CmQnleto/heoBDWhnFOBg1rwwaw97cF4y+2JqUo
t2I8XxkaK7IETU8OAZ2didr6g0gc0Bt1dNoy86B8ycsURVukPW/6nTS3xaRvodMXVjorSicpqhMH
phzIttLYtlbknGiiWdUYMOY2XaDt5ApyI7joKCW+s63gVObSzUr5kQ/Gx5JgBrPr34nkMbxulvcz
Evkiq7pYqEsPzMZKjvUCzum/WWyMZtAPgqL85NRz2P37PuAmaqtXLpfY6WPb1aTRl7dBwAYXiUBj
WajtuQjZaIwNLZZokudM4Juga8I0RpJ8FyS6ESbQLUJ0iSYYpmqoMN5rXwFt9imk/R6zDzcDl1x4
R68F3AQcRiYvPBjsvfYl8IaK3/9kequqpA+fb0h4T6jSvAcnps7r/BZTaRk1+mBMShJOmsPXmDpC
yVWQLUwdqOC0NVJ6QX7+QqpMBjb43F2DIXyQGhEy8i+dluQYNr1bKnDx01985NA4fL0n4yrwK+Ij
L3QO7CujDpRyC2XQXkLasSU/ZavL1H/HvaXU0tjT9XKSokeGTGqW4OHeHPHMVmE7fG9fPgK99YFU
TQcVZrTR7JEHX71/QQPLBG48UC5oLEPbY8c+PBq2isR10K/AWQLlIz+SmcI9o4oLGZNgtOiNK/u9
dkvsPh1tZpnvwlW/D/KtGUXCdhslPW8O2058BeNJ5nHpL0ll32ewGDqN13Uf+lmdSJ3Fl88qGceu
lRuHcPr0/6OGHteKQyHGRyao3xTPosBCNjPBddkKZ8y7/R97+l5tNdpHP7uNVIcENibwkWpFcevW
96wKW3wifiualf4Mvx2M+ge2yG+S1hnIz6b7zglCzI5/2t7Ia1OArQGN4M1n/Com7Mw72zLAqhnM
ZI9LKR1RU0mGFKNm0MuLxhHtmdbK/ljFDs/GKK+hIgOig0jqlICmR70OCBbNBcX/Mfmr2PwITbzt
IZnmDeNxTuCDmGXaVbO0qY4G/syHCnpIZuS9kfRcwOCYqV/SeMVYBOPE57KpUTqQPsAH2VtNnmec
A2UdASEZec3qQDhr3eB+3aRRuLZ53lfivpDio+MTLDf1NL9B2icApI2oeSW5RHJxfGMvw8mDwmKZ
QVozScJb60ai5L33GArc4HKLVCAQ/GmuK4cSB67fk4NwOpQa4wStslWdmLJIOtmrOtKnWAtcqBOk
n5aaeXnmbFzxQ8F3mcGDPdehE6SZVwwX1ztJFGKdrUGpYHw1y/ffcflYaIKjHUxl2xqrJVZ37ZnA
0D5OJG6lhin9yUWqQs+/bCfzYQ8AnKu5sD6zTMcEMSj2/fDyjlTqo35isbtiC8VhCju+Jo4/qpGS
1WH3e2oBbh2Wzg5blwo6OgW6PwICp7VJouVTvomO6mJK0v6WnXMlyl06wlFhTRK0HyudijW6O0nc
tL+wuX7emMulQvY8tXBbuS+GX83tqahd55ClDo4rFqmGhg/vmlohPS06EyqchW9ZV/Bgts1EWImS
A6UMaCZSTLRwwpQIqU/8h+5Mb0NmMzsMj8Y3OLKDf0zUdClc4nxn3pkeP7AhBYY45HBTr/yzp2M8
XIVCeF/tRN88ujusJFqQY7J/ioY134mrlMXSPinQCxFwIeWDZvJtqvrKU37XyUccvR9HfuyMrGrq
Bvdrun5QhPJh26nVjjGC8D2GTbsde31Qq7ywOlzuIvMoQDggSX20GgIsc7N3sARcNv09Ob1XHLYU
oxzOS7Bt8yYYo/nIr58q3ZNZGzES7CH7TQ0tazfDdM9O+klXcPRx/2O14T0hS6c7GjzWkiG5qbtA
oJgtz4emSBQgqcJvQc2lrb4Hie+pl0pKGf+tQHf2WKb5LBt1Pfwuw0Bl+K3DwZveFtTVlW64sMoW
8q6kVINOqmEkBQ8ac7QKToJpI+dSXiCrj9CtstCAftE9GZZtYYLXz/uPAZQ9KWI91lCXcV1hIR8O
JZwXQTS4/zHAE709/+B9TTfWdzFXhs7yU8qOeSFSLcn90vuOhrQv+XkMeOHueoaVgd60uCWlkkct
R2YFcL8dJOi/VmK5TxZzDvm6Pjo8URUJD87ZhRzIjvTctVxjqBaDKV8M18eTMaSxGy7ULTLAZdwz
kuHWpYN1Ce3G0sARm9xxuSeRMiUJH/8Rnvx6gFWIQ7CUrmpm3JpOchaa8nvvkC8OE31Sh3QPPHIn
yO6sHum7LRptZeZWdcSVyU+zzdOFn+4eO7mHfuZEhCsuIauvqoqFnqG2SLb+t3sKgzueECjpyiRh
9tCJcomCIuHsTp4w9Pzb2Vf1wOZX3cUP7br0xeKxSmW5dIDTS8a+f43r5K/zyJqcFR42aUc8lvGZ
Of1YfpXIyXuGw3uON/lktdy8kPzWsAToD8d9NSedAtk2Sfx9sjch3OjmwvGYG7jj0gBig7FXSgMU
ABKfWJNvr8y7FPV+JBJat1UA7AIjmNAeylL6F/d0mlLMSc1A4weyIZEWq0kaozdjJApstd5BmVDT
myz3xB6gFVQm4vU9U9EGeJN/hln/J2aHXC9f/PduNvZccmsmXJQU5oukNWsMP2AfS/Z5h+YMPBhS
KhXbwwGvvh33Wd6PoAJhaF8XlIXFIXVpnNl+dvKq8a0ahUQJWfptwzgBhnpIyjxNTlJz94Qr1u6M
SaWHTvS42YTlgqgfWreINu/5ObEznLeG8K1vOhcq63SoW6mBIq1Nf6gNiOzFjEGy/QpdiEtnDylB
VkuxlW/3BvKe1HoxlHW5f8Rg2eJ7p61n9uaU0VL7Ajw96kNSSVOZBacw9grXdRlnvZg4k1ubMVqD
frf01Il6UmTpWdC/ndR8xXsjqKpDhOGB4UbpwMLdoK1IWKW4jPfD6/rvnV/S7TmtB++2Y9gcsXnp
zswmnpb7e0eOxdXILQ+yiOl9jFj9Mt72wmlGoWm/n6HQbhMi0uUw84cCEDXKD9VZvQ4PNl+2xiUR
R8vyWfhQ7Nudt2i45vaNnKZg1AJGvCe2KEJVP0z5P5lB+9AnucCEZ0VEITcWybzqHZ09zkjTNge1
EHcpCIJ6bKIb5dYjQyV9RTib7GIVrEgmWPKlblXaUsh3dvgtYBloBw1FchqhwwCm9AAqlQq9H3H2
KsRC/7ep9bwofE7A77/XCA085dWdiNGAwXmL2XaBxK2P70VVQgjv8U032nKVNeP/SMUFn/yMMOpB
CmXInvgu1BsDkCNcbHI85CykWnPC02dW8dSNbGZmZwNEd0y1f0iuCBthxcY+TkRKhleOxmnMOBDY
kK3YUQzjGQe0Ij4v/yK7a68agWC5Khi2pxERdFz6TCYb/BIzuJD3oOYyt2h0x8zSyMGclBTr9IB/
cH/I6n3E7kCumUAIiJ/zdOiaE3BPHdL+7G8egUuzSRHQY/bPL63J2OZu9nLvIVKvU7q2AXMXVXOH
qbvYvzrwyqgsYI2y/Qyp6VjCBhFnJ9DdnMckUrKOQHs2Hgh9IYkLbt+SuwzGdVuEVZHmFNHjh0Ef
QPsujlU9C9/H5nxIw5HUqh9QQQ4jyKcwHMi/uBWc1m0p9GNhYeom1Jevq7iwFossNpZmz0gwC9/n
4s9giqHerxAheOGKVnZqTrY0UuBtUWQp3tzO7RLwn4DaX28AtBCyHj39hAigWUYNbI7oYDw6aqfi
6JzX8A9XcvxmyqmxDQ2A+ukrjhnM78pWIjMneUQ60fhjVnMAFfRi/yfQoNChY5+Qgd15rMSS4Lll
zv3+pW/8evdvBcgTjy/kIJHSYUA6TI6BjESbysHKbEj3oLoRPQxn3MYgM8GlSbFm8G3If4p2BR2G
aVmhOxvRJea8pjV1F/iIweMGXVsOlsye+a2mdkOwe3IQScSooLzBQKL6alRuwciP6EV7gPhMX88S
GQHPmSANtKVJgyGGki90p/8oCfJ+moGPwDbGDkBZu9HXw6SBXYTmARToqOs0sn48JNeVm4kVQqEg
8znIi6vKvoTHbDT1C+DcWP1X5zprGOJrugROUfo2pcD2/OBRuLFWhS/H2FWTFFwOfxDf32kn3R+g
QJapq8hBNrL0WUaSedkpuIrjG6yOEJKILwFFtIgPOXG+8bL0HaNqArEOXcPcCbR/tG3qxULls1lN
+Zo/D7CJQDT3zVgWD0Q6DSsUp0bJkTc/OnEXr42Jx/AIxiRb9GLCD2BF6rKHSfY+AjqGnAJstL3n
/MZIemGnxLyqHxHoku7IEd9L+CTQXfNe/aLiU+pumSzzogjSD/71PzgpOzPZksKj/BhJZJggTiGC
nE/Ew2D4Mn5AUF2cQm0FjLgK8Ujx/Wa0oiIw0sp+y5Hm3kNL1e9MBqwZ6lxgwCczzrYy1ab96CSS
BsowDWUmKFp5nYI6W0dXaD6IgTRKrNwKmmYWkxvkBqAIfB1zcJAaE0F2AhgHJffgpUM6nii38sJI
Vkicxsoz6ybokzueIKWjHivDhszt8eL2xF1MdAysMiwck9u69Bs6/IONgPK++i+4JCiRWbWSthDW
MG869M3XIaQlKKg8ExRaXBNWBbBxn89bbszAVeGhpX5IpOXXCQ4qcS3jisX4UT0LIKeRUmRGGlRC
FTwGcIgSkdLfet4BO4hMMx/9d6eM0RNiSmEqe269KlVgm1/mRkX7daTSC8+paYMUUX+lQNwYjMqc
eWr0uSateM+R9OfOdddGNAjyiH7b5SzFE7hbByOGiiZBzECnv76PsTt71Pox0uBdfeVs0QI634Tb
bzaiLp+1VCLJokmxO2TVoaNJdkEdQaCDKYxenwHiKlD51doFvDUMQkDZWIULGYdBr9jbgw1mjZIz
v0t+8oJkF8gtXYPZDpdpJB13Vw0201iAoWHEEsGzC5EJJmer/i2zQeIg4IUoobv82S84URgicwBI
mi3H7JG0wKJq/pPXZBKRdvUpt41WHVVnclkEDIwuM0Rr4/o+OSsOmIiZ1eHrxS2l+0geIHmuyphS
PjE/4IYTdb6Ks/np7j5ZrHgAPqAPehsVcoYjSVYoA8cDJ9fCNd69ixzVDpiO7yvigIkv/4MLxQ+w
aKv/NgPmlggNdjM7Cbg/+6mdEicYh7YZ9T1RiNaveQ4YyMsneVhx9BaskQpeg+jN8Y43Fs7aTuCb
i0jKfUy1qBf+A4nKcrUOvRoZhlFhD2Ivy/wNARFrYQyclY8DgGvZlPsGq5/tsSoS25KcCRcDvkn8
3LmFnLdSdnNKSzAeM/+tAiETNFA1YPPyU516AVzeeDy3vKZxRUhH2jHhCX8vIaevUX1m8il0Lrwj
GTTg5dgZvlFzT1KNdHK9p4bXWgTaK8SwTytw5wAnLWY1ubRNJnKDGqM8hOW7OdPDbNRQkntjjm61
rsK5v1ZzggGPcapL2D2afRzptAsKa9PN1WRkkcRqVgW/8+rPvYdrTnwpepueW5cCbPc22vDoQTTc
uhVhYflydXPpyCUhnwsCgrOzriJsev2FUzuNwjeIS06nVk9M+K9HzG7rdGb66D76IJYkgJkPyNk1
SlD2KLsNpUUsIz/180ZTM8QR8fpTb3opuXWAnkv8DVdf5TQ4LphL81I+ezgEabsmP6jrjBG3v+hA
Lh25y8YwSo6K+uepynR/0rShaP8kzUEq0J2zUlBnxwP3klO/SwoxT4HjQZN3X0CMjVgoKIgahSqn
8DwF8Butl0e88aAvpdwDPz1spOQDvHMrlExfUSOyUYEevHUJOmRYCtp+KzzVnzl93xFGUed5nEZX
s7PDLeGXhwP9Ti69seaPDL4/AgMJT0V1txu1nBuV3N+6rvOZjPTULrpolaDXb0llTEuYbH4Sd2g8
cfrTth2SoH04Evs1Tfb/+nAwgROd204egk01XhirElYSqFmSFq6FYmYXKqGEyU4v4LHSb47TAeuu
aAAxoSgSoDgp7uv9tKtBCdyNaWITAviJ3J2s1KAXDlwUUCSdNo7fCef2wSS0Nxl8KBz4poMnNWQa
kTKfU/YRvFefGG2LifjZXGHvO8Gw+AhV6dbWW3pSSkAPLbnyf4noe5RgFCI01t+rQPm/CYd4TEEZ
4sM64Offlkk0gnnq5fkXpTjKc+yz0E2yo/fTIJ9K6xTl70wZCzqvHzC5IRPP4WxmzcYswSKmx55Y
k2AEZRciv768eKSMVnasBnYc6OpLb1T2eVhf2Ni/L66nS758/JlOyYX+Eal9JrwW/4qNU4iMG/nU
VK+derTlj5MJZm2c/nNb8qOm+MQuxVXryF+ARk70az5VoZcUJyALjQRwSXyHDKiV+Wgr+TnqelTt
7Msyl4+d+TlPWcZGX13CbqS6lM3t6dbH1aLjZm9/IplgwNs/r94xwJxSHPOmayAb39OzRcUCW/eo
77qkxN3TMRTqXRYqurPRcK8HPECjaUhED6XdJqdUuFPK6YiQ/c9D2x6Bnpz5afxCN9s9PpJ+6LDS
nZ200YR+ls7NnM5M9ZX0jp3to8vWg9kKPOKxvrzVE3EE5lrNydEzFreG8eBX+XZZaWyjHTLod//Z
wJ8CfqXpK5vOVeAKQe8RQnFKe9ZnyZgtDHUENiD7DJU0s14bolfMtY2RccIse96VZAr5bclbj8d0
Q+s9HX68FfL5rpaM80NEXoVw+BsYANdZnTu0snmCZ/WS3+iuVhfbBeEWHVZlNeuiScoUqaxa5RLA
K7W8BSQ1+44TRp7xFdQ1wYeQ8oGG1I+uhYBZpJa/xaxLDzeTCK/Gn6SHEXr3hPTG/yeJ4kSF09IB
QF6CqPU8KW1QL1GmItA4oCvlD+bsl8kslMc1er+cGs9v3Upek7mc7B2b09DFSdquzZcaEL8bvLGa
7svrZFcfWJ2Tmv6yQSpEBMe4h0eYY79EEw0Xn6STIeT4cD/Q/LxTpGoMRVKh1c+hYxVJAJP8fQZj
00ADMM/AddX8jFX1fkBrIL+Wvif58tLZkzHI3UDbO79T7IyjQYcJoSzN2N0UR0PH9SbQAOKiWwAx
w7Y5pq+NmZZplyyEa1GjJ9zdn3B+GWzSy/8UMakSf05k28QBiR71E3WLPJ1yREqYPxA5j89igouj
c1p9/Pej1VQj6i/Jt3Ip68AN7g2wxb2MouPjMOgT84Kpq2agiTjLWTLgPkS4/TPb+fGzO6Y9qgyP
bCSVC37s86aWJjA+rtGpxYXxBo3GzVlCrsjNqD/XDNljIhBqGa9rZ42CYsoKBA1l1XqlbXBvLYmv
tH/7pbvwP6qw8VqFVbmR1De+J7vK11DytCKF4daGFhr3MLs+elok3+u1JLGVr1NLMLFCKsWxsXTc
oFFO+/YdsbEfTb7E+9V5XDfSd3SI8fd2ys4QSZq4wu5Jhy31f8u1Q12N49ENfyx7mxajDnmSpd2g
shDYLfOI6vD5Z5AZucW88TmJYl39mB+Nri3f5dp8jyIa4B7tnc/XroMdieI+z8wrXjmxlW+OH4fw
OBtMGTl42B+PlxD1B6ykCvBLfMIPaGWEuC3J3PI9DlKJIz6n6AynWYVCqK9tuqejyzrxbZwKmNqn
QQ4w/RJEtRyWzSFolFBTHDMLi8ERyd8Tce/t8aCZdUOeLSXzX7vdjnzTyjNP5FL8/xJP1+uAAvnH
fp+skGSKD5DaDhdzo/HW2grMPg3sS1+dKTIwunqYj/wQW8G9IIJKcp/xjno7hDMq1JrBrPWBDZsN
TjCE36MGBdrPnOVIPKtQXhZiAVCAfPj5qNMVTTPfSLc9XBhNLjAJ1jVysULb4SrLVDnoXj5Z17Il
45deK5yXRrgt1HAyW8+wKeQ5Jd6jhU2GFWJEa3iwciN3dDOdBMxT9WeaYitQNN84bg7rKVFj7nJR
2PtQiEgPdKZdBzB4nYJ2118ZgokNMXqT1ZblRtKSlQhVfOwEw/LKPyr61oHL2n15zDqn17K4Esdk
SoNROD9IytI3mJPR8oXgg8k77IetvcAlWhM3GXTVXDaRVhNKtH/WUOf4oDdwlLfYCKKBbmglBNTr
H+RZGZ9LbmSqgFfkQR2DakpXR84tvXsZGXqgF9CamwtWfKjNATbZI8W8AdVz7QQVpWGaLjr2be4R
bW9X/TOhP5ByhwpZoV3lpDDEfND9SDrq3I3JLFL3voOI80KIZ+47FdXYJNtxcyYVJvvp6Fn9cj1E
T0xWObCsyNhZhVpEdpN97WPAWitCcNLip5QrlbkSxeshjuo3/Oc2juPAX1ixBjv7vkE9m4mlQ2LW
ThfVerZtgAqRwFk1BLSI1XlkYL0+dxHvMOdMk0PG33Kgcf6QmgjULi1Fi0oWM1t89NvNpH4h6COe
6uGzl9KA44rLWzfUG8m6xrkTKmxtl5zCMqlqoFLUcXBrorlm1fUs2cgXuN7/2mqP3piNsxwXGY97
D/fYZXgTXt9Vyg/F+QU4ZvWZZJXhAs+odZ5pbHVicUdLODPoLQ6QPTQnCcjpfQ8WqpcXrzMh55dS
M9AK0JM/zH0ARuRqTVd8+V1Nph4w8SPtI3gOig0p73XbHN0/wWVcugJrNaTfUF0Fy/5WFxTEHmPD
XeJX9lnHqhqw3pYdg9w8ReOht7fTdFBhm1/ZuBMZCJr8+9y4QzhX+XRoa2rM/hzOPc92P9Jp5Lg7
R5us2TcN+LABwXUk5Frx2rQnXhIKoEthqaSVzHnYnSGYM3lUs1nmYOhTIco8ayHXPNzKnuoh0eoA
TXIXXtJe9cF/ZO1LIwnXHRkCaaqssADybgTP+zW/9o45M9cPKZq20RmL76ZjLlQ7FajTTfKvUbSe
Qu/5ArrMOZKfqsfSsBVkhMGHjYYT/EkWeDvf8pTeqClEuvc1TNKlksFrkOcvVGqiUKUVoqGrvosC
URNb6Jzcu0mUpWwCFGv6SPSz50ONYt7qCtnVLk+eWJF6FhLp6D51wIwMoXXu4nmz+hNoF5P/xUZW
5uylXzaE/qubtFsoB4ILxuNHvrhiSSegDjjLTPJ4KnajGlPPJCMxlhWbYic3msiPe9H6y5Ila3Xw
twLxcjX+1QrVSfGT3MOR9ih3Gus3FV7XKvz7nz1hMrSCAt7lR26zK5T5iCm556oAPGp7y7gRp6J/
0Mrk+L8/gjKkEz9iDW+7DguZgozEtBizATOsooqqo+B1vMKxQu/7AenA7NX17TkHSdZ6yF2UFXG0
rdZW1PSoQP5S5kMcEu1NlWLm9WbkdRFF92uDFVNgigHJ7EX0EpJOEOGakG+Br/SshklfzVQSBlbP
TT9S0VRbbb4sMOI9oG4avLH8C/5yZLDqia3SX7tsRZcazasE5/Py+7YCCH0sqFbjfbEweJrrP5fR
05DNrZf1U8Z55bdROBiQvgaS+Wzjcy9ikj2vZbzj/2/cy0dSzij5Kkdi62a0Z988KPoDdCEVAlBg
IP0E0ItvnZjlpvVPIZAAYpanB/6wIXTqkINEY6PFpuLBzHzA25ACcp7JyywNLhQNkgpz5UWyC+8O
x0Hu3PXfFTswGRZrYJEGbqBYEk8TuGZippgZWU2goegHAJYmanu8aXiDDg5F19F579wCKK2FpL8B
xvQB4jKQPo8fAJNCVNJndjchEg41mD1Z3fqehGX9bkt1+pdkycdS7yi6BgaoPg9h95lfd8Swbzi4
pmbnwvv2EUB/mtJ09ELTIMw8kyj/2QMvcqSDeCDDtf1gEXPKoXyNcfa1gJZ0NtDzVqniJnVkbZmb
LlJs7gl2X1JHvfbPLZRh5aqNXObhVz1vErmZ/bhVhsenRGM1zhwnqiMsPa1XhNrRP1jva7APZLEX
dqVITXhd7c4EZ69jGEJmMT8hdh/hxVvAQAy57qem4AVerYUKV+1unoZd+TYhW2LpO5m++CyHXO/5
WNTrLWuwKKy0uArViVMFQjiFrozZA2Td9HjQb5w18VUYbaatOSz5ejMlDbdp9DbkWc5hsKpb3F0g
UpcMJ0dBDwBPp1xTqEoagPtW0pPAK6clWNivzDloZu5LcUrzber2ElKrEMfIcJ/MWUIB4FwaRdBD
iteglu8en24POnBc0hySNh9p4vbOgxe4zcZik5QzRTL9IZKSgCEITgId6D39qZMfjolnTSCSd1BU
wExwDSm7/vv/xpZfUtWSiN9M4ZPfVpb2QvEYjpH19hPM5M963mrZDOW3/i3jdstlX8DrOpAugo21
dYWTHksXoTNpplbZt/Xp5Q32at0W39zvjAdPubQgm6yNtD33GqLrW8UhyHfVHReKKoTkm/IkqXiW
eKchLl1xRzpcQDQrotD2lbjbdfVxpWeoJboa+wVTB6YMiMRf02XPWSVXGCl0kbvJJD90dIPH5M9Q
rDmw8KdJH+BRkFxD7N9uLB4Boi96zaWJRebK/CqhNu3z+fIR+MPuMKg2dusNECCYyh2miYAAti76
CQyXZjDOEexnqVEGrc2M++L1VAF6v5I4HzR2/HF3FllLlePTQCJml5Aj0QJ+nBLbYrEKtoL1rF0h
Qt0tyDfp/GH6jJqv4fFvrS95JWSyJv/1g4rCyHT0H59GVEENlLti37HW/vXQd+kFAgCTTEsyXk7I
oxHxhwh+VPATrQHEdR4/tB3Ql43jFWBVEjFFf0qMZzjIDeUxlKkIDk8hjCQQp5HHI8PEoRNj16tQ
aecAvR1nb8aj0pCd5lk88x6AqmI7kQDeVSpFWzNXx4ktXcQX857ILUTI/GIEcDWyZXJva9sF3xPT
S91zzdJpYGU9Qs8tcjJ84s+vZes6l5DyEIEYhBM0kIsdxxn6wrQ9oZrxlc7jWJC1UrtzJDWElzFL
umEG/y58SL2vz2dwuSdKw/8VvGUnln6Imhyw+Wttg413TOy0uiJJD3ipW/tAl4bA8o58W9+Leb1z
ffzej0dfs6CCOJKKSGgYefrQ6+9x4IbHMzw48join5YIhcVsKT1AD3ajLiORfTfzqrTu+11xoEmE
lHcibNGzbfzRNC9dBE1IK2RvUYyAFP6hSFFaMHfTGxlkRT3IeP1lQOzt7Msd1hx89i6mT6bAuucv
FfzyTJOma2Ik0mH2KpF9LhrdObI2XGCUtl5D4L/wdbRAgKWLa+t4gGO+KJFTX8LNvSObEX2693jW
REHpv91cA5wNvAZ2oY9N845+PV87KJ6bXbX1r7M+gEhg7hNdYjOWzyUTOlbhHfSPTfMXDXNzTjQ2
D+/3YgbB9DM3KhZzfot1C/YZZpcJjPgUpVzUCI8bmPmN/4EZ2peWPRBL8uaa9zkzz+Mt6M0u8esx
RNqEfPa2zSEUQP4YM4XvDnGgurvbJsYizLWmHWuRxVe8yBp7U0qggPNSEyHGzkuvmEOeoMUUX7LB
mPRIxWwSFfvnzmzGQnVT3KBvkCtRTfWkP069MlZoVCwf6U/EleHOHcz5PHCYQW4AY1aQ/Usvk0Ru
8g3s1EZiSM9dSRymk/raVTn400dgivzIZdalyHBSoBgrGrQWIDzb3lDAZeFYtjfruRGa4z4VnMHE
Gl3DYWFiwz4pQ/O6sSYh5lDeS4puIVcSxIpamFRN/46NZqycYpQD0DwmVGcJ4UpGnj9A+mfwL0gU
SF5KoBmxVSA+Yiif8R1btb3baBx+C5QtXG0CpRrUQgp7soDa9ZXaqZwaXGqhMnay4iV/fjMnwoCe
xQAobYEKrZ8NGjPaOI1vEt1zNOfEun6WU37O/deM1Xg3CZPAB1E/UhSC/erlUbICkIcd0g6mHVjG
ZQqQ7zd438byH/ec4Nhl4uq4m3KkSfoYDoQMOz41T1LfCnb/1+4HZe/RqEVD9zMg6drVNL/qz6Hd
daqxrm+pumcc0zYWei1/yKCn5BfYgUgdTDXmrz5+we67u2QCsA9ucUHzN162ZfJhLpZGWW5ro5EA
i+5Yhva/991eH7BJOCIMFmbJUlFrxlqSoYqFQoFxC+7LaHTgV13tSAqDNEDgVAVKnChcJzXuIdYe
i/t9nSnu0pzCcylK+N8bLkpm4aDtCuKOtcU2Mkqj00yDagqj6GVAb0uE8CVkd4SFllQR6zqRM69L
WJvCVLGomsDjyO4MPRbpaOcrfYEo0BvFYwFOXZfXPShdQwXDSb/BhFQfyneQBKOJ0ey+IUd2q77n
8+5KijIJWAXrhANcYIk5lax6nPjdVqt5dygSTs1/PdPuECyopyBs009yUuu4YZgUH7TzBXI+6Me2
TBKGTHtTU6E5wioT1DYf9ouNpH65i5e9eFI2wWBG2xKuXfxhdf+B69YqUjd6q6JKx2OqWUaJqUXY
tIiOa6lMYp62v4T1eQBhW/ThEpp31ypQNdbPs5g3C9/LZNgmnr5/U44aWJF44DK0WK5v7tKACywo
KfOExbK7zdAhpHe9T5e1f1ec0n25pUMSjgkfRxGvXy8jGTXCw4R4WEqNu7EA2lYiAKLPEVnKsEKr
dMXT7+TetsXbwXvuSkLg8HiLLEIRK4+YgEW35LSTu+HLybvvVGBcZyjUwbAIfBLu5DMB3U4Vlc+e
fvGRTXW62ZImpKxpvGonLpYFWnrCFSDk1IsA1UpLDjKJcJ6UP1il0+pv/nBnJ6pVPcMao2vP7iE7
UMlqMDppmgKe7iuKYV937PZxEmEyDISmlVG4z+x556jtOjVNs2njq854gXtMD6ROKB0SX8Quz1VX
V3WaOTRJptfSy3KnpB4JQ4LmyWbVaTtnRXSvdKYdNuuortmhOtjsRYnn1gNU5q+/SqhFwLlwJp0z
8qdM/SPtfoUkSlanExfsNuXZNllFnt5nJ9p+oayYGAJmX/AaMpa16xl6+VKE+s2Ym4zWscF0IeTd
D9YZXqF/EGV9SkevspWlFXTD+kk01+Q9Lfxr1yGiW32nCU1nkKUUBSkB0ToIX3EVV0ce7ESlorwW
L+oF8TrZQnGz9gdNJVcZbe6Hsv77sJ+u7qPjwfgF4psderKUa4LaHIDk32vvttDMQHIuh1HSHbDp
YiVOE1wnKZEnMJaORAj2dGBuV+ijd2C+n1sUxjQizOYl++hGpF8YSS3gMf0i5LwVTWh4pCCN97N3
mHvM/BYLUCt8nelrHifqXwzhE5llwRNnGhVSLYYb/cKef1SOUBJdITiGsupXqtRm5sbXViCDXqbo
Nfx4LDBPDdiks71HazlcQFq/Rx1NPqJdbGq0u3RIgzJoFCq0Z1P8x7jnmrVJMchI3Iu8KGvsUWkN
A08wotihrF8prEnKybJ4xgnkzU1QNd4Q4Yr3Iidc4uIoKJtDvll4WsrIFcgt4V2zwYAWIpdPNwBK
E//ELND0vTs/ZSfGA3zVQERZm7WOKzJcRuBpNrTiuN+jHTRLfpvM9d7AZNw8otmCSaxXZ75NgBUn
tKO1I3dYruGc5UO8/KkAk38xKZWDOsuPzdYXCb01PLXrtaOtJiwMMxhdBK6/DZ+4eWJJ0KvBAjvc
WKo3sPkzD69xxVskmE007zsRvkTVDXP7gYUjOo81S+7mA4lGY67sh+Nm7Sa2Sy8vgmr7NCZDSY6S
WBO/ap1soH3sgppgKqrA5zrZblpO4TAkGPA59NbxQ7sl0OLV/PU2vfoAa03e93RaDMMeptjctArt
W8WJLhQ263yzeWzrh5lpJax8zlgP/x/HOGAd4mA95dza2+swz81j+7aJaFhmUZrGV8Gc8X5NvGX4
t1C24d16lErBVQmFVmB/DffRDdk5bTmk2sinEkHph8D91coFTtssQ/WdyqGxgviBG7cZK1bueSU8
8OG9cEIbWFdlrhv75CyhC1xEXuHflI1jlT94h+uJvB67eFcV1OmZWHQ4/wVUuLyVHMqUF7EmTQE9
gT2SMBWWNIfz6Z9qSmUNHXtEvYw8FDe7bzY349KQizIhMrKQi3MhPyVazfHji+ADMVtK/cjznJRg
4Uj6lINgqCifI9ZeXef9EHU8zn3dedMpxY1ZuuLPra2fk6vOnyyRWXythOU2ed283OZgtUC5AFSd
M74z18euc0wTsoVT0Xn5HDZPhMCvc06fuI2NXIa2Wo7kydBGbP9gXmbWerT0qzkFIvvxCStb5FvR
tx/Qiez/2LxsXI5CsO8aaFfXuBlVqOenFwj89Q1F85Nsc80UjdsId4BK0S2YJIfNQ+RnaNuTiUMY
s688WFP1AG9lM25+P4Dj7EKQE7euav7+nTuSm1zc+t0FH5uC2O56K9z91t84ahmZ3n5WasM86umN
GVyK3Q4OYfecIYUZg3G7aBhx4QHUd7JYsejPXRN2FuYppNKutVU1F0TwLDfw41urJqfOqK2sonYN
WruaHGEUQZwtknuRs+sW7OxOSZJwYcLouCzAtZOk2yMWNB7aK7aqqdlqM54jlH1/VblvetzZUNLH
zDvaoONksYgE4+RuRKnmltzcQR9vn6WKUlW0PFAxvZ8dnFoG0h03Q43PdIFemgWaPHP+AVPJ2tsk
z3XkMlgU2lCSC0MeOHMAkow90vGXfCqNHdjvSLkBV1n0OKnMIa57NguCrsvAbB4DdbTvF7/tbA2p
7KSxeAijeDTElvqPLYEeIE7saUu14BXpPN/OFTi2eErWU4s6SyDVq/GiTW9qGWCFmvbu+JgkFU8/
D84pV+gV/pF3GN0DF/ctDXFcHXkWutmtpsz/Q1qcQj+s8Ecsma7KE86rCEoT6dsUDG8gdB6o9LFU
KMp49ER9S1ijurCV9MnM8z7kUtELZnFr7/1WUlp8GntnWq0QD1mJPLvMHbeTD1vXlV7FVFKA91Cf
j5Q+8dAdZB4tSqgi+4tlhmyFToZwsqr2GU3Db5Jl+Qzq2gLIbPbL0oOrPl3ZNHeqVE8RvIWJ6uUS
kr/Hylqd8xvwGOCo8nin4LgWRX0YNkc15VPD8jeXIpwqmqDe3qLKsw5WMy2fXcjiqtoWaMnYSovY
zMTO/O2wtODKY8PQQod7/6fcHGQvTqk1O6oz6KXCSkOXZ9vrjuN6Ez5Xnm0qGQBKHC979VJ6DQ7j
MnBHPZNtzBXV45pxJUR4ZO7oa/XOHDRB4IWfrH7sElufv7zD7MR9fXocUpv2O1sqOmr3iU8r1qRn
aKlmnVxEy0EO/vmFRuokgrsH1M8acvsyw1AUMGrNs4w4d9Lraff8YHgFE8PB7JeQwCedXl2anEeO
AjfLKNIdbdo94oyou/FKNOHdaNLtlVXXy2+OILuIs2EEYGt0OfzQQJCCYHF9sIiBGwL7DQLvnPoW
GxiPOqLR9AtM3wOC/8aCluhtI6HvLVpX/b8kyR6P8aaEKs9LsJAo01xwXx23N4HzF5in7zD4Pvex
QUv41r6QxTLKKotz9I62GDem+voBtU9qt2Slh8/XSN8GMRU/CwC4u+0Cpks3eWoZWFCMs/qCa80I
S5/aIdQBJJoLY96TFlbLK5gAQwEfDyDTC3yH2tmdbVNwyKrNMziYOmTig8wxG9z9MysY3Fz8Yqu1
ENKJdHMkxSUn23nlKelgr94q71Eaz2CKN+Q/wFmexJOrCvcolvziympCQw9/xzbqCrAbyPnyQEp9
Te2+8HcjjDbJ2IejNYgylD00kGIX17Uiw2m1HOJhHd/FYOl/gblTEeKYYqIJp85ovDziEES6rbSm
7FHjp7DcXFAgs3fAqGpWf7/ioD0rVPpTSH1vFO8ZTINQwIvip6ln4vWjXgEpILmoy/RBDEG0i6jq
xQHpigafoeQVfvKgb8/U5792Yb9YefNar3Ikh+zP0MDjXFCZokyz3jo7Hgc0ednjnZixQaI7vKRd
U6FFDqVUUPN/4e58u9YcYenrD2kguP3McKgsZyqfD/h3/jrjSloHYQNkHccg6K8ijAjImyVDjT5M
c5vztqXsFw2L+rdnal0B0LT0Wi4v0QwHp8Oe8X6nUDUNxg/OTfj46hSVA5AV1/nJQCL3+CZI9OjR
9j7LWPDVurFiR95zqH3FsfRuF3d81tYKev5elfSIvxHoQ/j4wGVOeRbvwnw7wz0hhy7h+hk0/3Lg
i5BlDaXmoMN5F9/RETEMDpEMTVlzrTyiaBrkaeHF9KvCCLpT7z/iCiiYw6kS5MXWuIX9W6mE8G5K
z6eS4gE1LVd5KP9eXJu6xcr4laRvUpe8TXxsyROmJ6NnxHOCgZGzTwXeOJmT5IOdDUP2WYMykqSR
LSoLy+qMP4x9PDpvx+eAiVpGahMegeD8EK5JOHiwlmQq5ZqeKobxwQm4jb2QzgIsbIlA7r8NhwZM
PDJmEf9ZxUo4bPA0R8hmWb1gFv7qOXpreShSXLym27GjiKQASC2YOTl0pB8RoLLeKxqVq+UFpooU
/HzfL8ZZbYLxaAxsAV5/CjaY6zyBd18oq4BpWG8MgXgwg4CNFXeq5N0BHWzjqvNR18xDiovgfOrN
qv5N/zNLPkU6Ctgd3kO2IJ9zEc6WV8vy+ZqE2rN3jJcet/yfLKyI5+h+wUHaOXHiy5K9xjKk4b65
7tnZwQzMUuQizB9Ps0AU7Kf+J3dj+lLup5f0wZgacdVatVi782NNWEBqnGdlB1G3TBORgJG1G312
Y0v1Vp0VSSjZ/z+vPtZVx3t86gqDeEOxojx+4R5Ml0NfX8F/rzNRqyy0o6SVaWflZ49b0zDocPsF
gprrQnWjsrD0LoeXd7gBrPZHFs5+PDW5r5SKxbVvfrUG7dqEyxs49mxXYb4qG8f1yffeyc47zPCc
Ewy4bXsbIRyXBagiOtvfElP8mE16Fq7B7JcFN/mfmn6qA9A7e0JGF57OPnx+nIuRqOi3dIremt0F
dEIJ7Kt1PPP0ba1ijp5cJSGyv3MeC+I7uQ5gzRS+qR2CRwNRYbMod7nuKcz28ARanYqzYt/HZai6
bVNoyqNwgoOLVgnjeMXzVjO/muc358+Hn3V6t19m+dTzA6xkzrXrIALcJH2gig9KigTQO1Zxny1s
Tet2/Av2TFmUTdlguJkHQsTmpI2JxL/DSrDeJrauTgU6fgUUXv3P0QVpP8yxIkb0T5WkCo6wtMK1
cFMOwwXOMDuviZSvGB1K5DFXJhvgGD4LhofrjOPXaCHy+7rELKCvoO6QIs/VEueOxKWqjXBnPrn9
JgtbuuXsffMJFwpaKBoc7JxmoxsUPqwIn4iSpLLPG9YxtrKtHVmcw/kqSH5lw/dxHVql4ibSSu6T
ZsoIK6lzzI89ORp3GQncCZ5FHOlQBnokUw0Je6BLVgPOP4KDP6HkJJI59BQ5W1hBXKUVlmljIevp
AZTdlHgW2D3rR76yWfdCFl6RYiU9pwNjkzeeQYxviCp1BRtHg2e32CFXMcuH9SmM3bk/XRHkNG/l
VcFdbBPcFy1aZQEaxNwr2l4FD/fcnFG7G6bcyVpdd/7cuJPO0yNFl2kjZoDTkZaELjbTtOGdrxmi
IejrsJWFmQUmeuRW7r7/fuL6UAZ6iroHVvk4LwSREsQAZvh8LS6gI+Ba9j7JN5OazZBKTTKhhK/e
WKl9AhpnBpSgz83x0LqnwAIfhcefVBJpOn2XpfCUQgErmOPm10w+ZMViJT1U6urahh7GuHO6MJQW
StSUfRq6edvO6+7fBGRkN7QIUGWCPDkqmAEvcuQGww6lLjwDL8yywqKXl5kXhXp8W3YWL7pIgTLj
U/JW2qixIQ7vcW7DEU42++DQM9ML8PEq1UZDyA8+ognwraeErk4NutLN+8xE1G18DUV81JMwJ0D5
TjPX1xt8ViD6gPb9uZt5ckcE76dhXs1yi8wjHV5Vg1lsiefBQhJ4yo2293uvpKn36p7Iqjddj894
x2LetuAsh7SMjzpOLPydnAcbGmi45p4lorYrPyT4kyY26vuIzH0Kwlnx/ULQb3YLaavrKPYqsTnF
neI4N7sBPTBvBawC5NH5wfotFKVpyy0iE24HU5MHqSh3EnUptNWQowT8rAMZE9P6AQQltZw5iLHs
N8jTp8yBlAwHDRM9UjjXKi5OPxgiy7NYVYWftaEXiZLJjT5PaZIvl/Adx0kLShMmRc8bFHO16jul
T8SSggTat2CGFIxievWlGJ/TqAU6V9HmGHdgylKRlsAudkT6qTnP+klIvdT0ydsNx+Hjkoy4dsae
IdGcqCcrWtOzpaSRRVpJxWrTWQCOdRdxIfI1/q8D9naeAGCz+5eHMJWTO//L6/WSGomaILBL81Z1
aYGcfvuC0oeJsJS8/zudLS06hVAw1q+kXxSyArriQgniVEkMdJjIepNI+NONkj8j/j3Ot3FfktJH
zV2rQcpsC51fY3WuWrMWg9WR7t4mArhFABfOan1mXBR9pRUqyltpt+p+AyFDL60D3GhOZmJEHtXm
PbT17h/Hxy8gfqjzW/4xgOcxeHXoXej2yjEwnxJj2vFdCquus8T+PPn55LehrwPKdFopP3sMDK6y
8E40Jkjru30YUIY0jrv3fXy+KPjpf5HyxdKis7eXKpRzfr11DEJUzD937MyMGotQkkS8M8hTkFrw
gZSza3wPkPdzsuXVQg8zRBu6yRcRrB8cuMW0OYZ/hPg4GUFpUYLI3NOyVEYFL1fsnSa5Pbn0VbD9
BhxYIwlFKRgpW6B8KfNCt+KNjpsr1x/kkKQuIHcYBp+ZYIWekqVPus7oJWPKeaDm/lPoJMckR/tb
uSd9bFwYsf6UJmwiQ/gDUe9t5Ey97K8S/RCX1QEnglSfQAtOT0n1+oVTFeBi7R4z6KUjNKpea/m1
C6eZ+SwNgmeMnC5HiAslpt/ovlQZdeiwBKAJkoFCSQFJBXH0tFYImgpDLltPYWlEnRDkLxZJjmw4
kpfNTrdqF+oNkHAnEZTY5kDh64qQJi95GyNikONv3KDsQlxxIg7cnm0Ftlh0pT+lFM2nLvdqGjmu
7TkSB5xthpULfDYHcG2l4NC6ECb+OEkLATgWPjYbypyuce9bnyROfDwLm18uaMdUZAp+RHthW9sm
wh5R/4uEaBCI6JrtuLvC3EY7ENiTaVzjNEFpkF8yC++7IZzHXCRkSVGrWjmu73ox7fRNjX310d+u
KxjLMG4gqLrUV25jy8p5eJaPt6MklRIQ1JSrCMUPKYQ+2R1fuJwRWyIUMMhGDDeaA4Ud98jvqKr0
KDjEOhgEbfqGDQMTF0cpPJZBybqbnwc1ygGxzoWnj6QFnt/ljUGCUKm/14YH/1vYwR0mvZyiMGsL
mkykHbYurcjmohehbGoau2aetUZfVHTKa3vo162TP2mPN0BoABY4oaft8aiAirGXIDzeCS9eCmUI
K4JE2D36/30SJ5+X9NlMbmO6jx6SmcRyH63cjslWFup632BwBGzx4Cg7WC7u8INPSOfqDLKH0XXS
fqb8Exza7Wp7PomsbcSWjHUBymQjYO7KuJ8VTeTeOyzuyHEFXA0aqQMxKxrEUhPpnjymE47UAbU0
mZQj4TigJY/VCjA9AM6JACIwnbNd2Gl/Jel1Qhu6oHlgYk4yoHAR/enkdBI0/NrJBEoLOt8qN3Si
NwmPJRHXH0Jd0DLsakVF4FHEWzIUhHJdBOLSuLhQD9qmRtzX6O43w46s2q4y8LJ7YWGizt8SUz+v
LDL0qbQ2GsYWJsuf/loZuCCMNhY9hF9qnOGrhpNrMSfT/YJdvoY8YNCw+TdUr2qCNGkzWmS3GxvF
cgothxX4nKMXIUsltd8awnwkhr2ENMjboUoP7Q2UKGj3B8uIGO96mhbWP9CrReWg0O49YTGTnyAp
7sb6idnQbyXt010+Omq/N/SPtLhK4TnzB5KwGGpzjujJfzOHShNL1LuekkiansJW3WzdYVWMgXmY
rRGyn6wXsHmI2sdkNs+CWrv4xXsPyT+y4JHnuzlzHq77LJNq/K2eNXb8cishqQf03/fKWnBOGKjg
DiI+9yqOnkAqvI1+5lVyU2pqJJiLX3+FbBqTRpzZqk8OmW8cM1RXtTrvrw64THk+ozeaHuhHtLGW
2bhXMK2LZOMoQAxKm7FfCJVZWdRPvUPqtm6xtBd+S/+zEB/gL00+ZMZBTNeSAXA0AnQVTpfc+mkD
IxygPtl6cobN4BmPOBt/QZj2IwHkfm0s4EexaLz1dfVmCYc0zN58sN5h/Kaft94gz7Kac5F2ejbT
YarlDy0E95BzEnjBxuQUoB2O/Fi59TFdbHgo5N1lze9z4WjXv7fIgEypryJfd6N9ie1HijHHyAkx
S+f5qrlGrociITRxfPCZ0mTv4U2AHJrAphqqxbbTH9OLT/gBq4SzOGpvz/ouWJrsR6fph6gbNP79
0PRogh/1JAspGMYq1pg7wKFQKdTrBVUitBCkoWhpRpDk4LtP5yejZ9F7Xwpg5awO+67lkZO7DTTt
QKKqp68P+lzDBjdPadMEiM/gHP3wmVPpOe4EcqCIFjgrRrecoxbNUiGv6OO5R+yxU0CabojtBo5C
fmEMT4GsyMAMhmesgHcnUZPYSxgFojC5rBXb5lBO2XJDtUOF9KfpNvOYq65Exap0L0rKjnO2H/Bd
82TKbLHgdSy1ebhr11cEu2oAOYnSi3nDsxA0DMlyipjqob2K6HQ4CSKw6GMeKod7mPMeSJ0MqBgh
MT56xwhvBmW9IKHb9GHtffUYwrnG6CtJlW31ywl/QnSOVf7IfuRFhyZu218Futwx6Q4PmEY2zw1G
m6Wk9EAsAWx/YsnxKDzZKo1iFKDkYRgXptChL9ctZV+aOQFjwRBxTll50mVNf3pW93NZzYNI+2MS
dlhkQGDCdb80pcf1Xpc0tGDX1PmClWc6blZfLzFCUYquAdhu0J/MrMKFunRh0OPiAyWcZAESymr4
fjUvbW/HejjBzEfWNGn/dJPAzIRRkUSIXZL/CynPPb2xarFOJWL4qDguaw1jOhQ0+Vetg+jqo7Jz
q8sJRR3K4WxsRqB5g3nPB37kflVGdtk4LpnZBKolBxWXxYln2t42Vc4rC9FExKcpY7v2cN5Yp5sR
Q3hclb5X227sPDRz6t8BBVt5OhkrJ9hWfAH/nES7Es6uPs21NRw40KmD9TSAqdQFe0bC37spyh1j
trGOjihA+muX4djXb9KxFv2gDgNj/ubkxM78EEnsXFBFgoBCMscwwn4Rv4VFwiBLZbfpCXhXsvVk
P+ZASaupEexITemeV35DqMR7ZbIGnmqfnejCSbnXV1BRqwrUEnWxQKld3wP2WytqiZlhlkKmNnkM
oHOW2JG0fkFVrtUkrVopuhEiBtQpGg4zQ69HXrOlxf9VU4X/ZVEjz9Rg/rIppN8zHhPKeO5kt+5S
LXacsE7N3mZTLMcx1XUeH6VyWYhTgcDDY7s1LKpKx3EgkThsQyqeBmoamt5tBg8Dkwu3EmNvaXNZ
251zGDi3Evri/LuJOPvAT4LOawYF90Rdl1c9fITdJiufB4fnySsvBBXmq/Nm25NBUxCwheGkvdzj
VtyZ5KAa7QAkvYI0mJx2I+vhwCzlVNXHZ7afXoSrOqw8Bn69taky25QdKN3yMaX92ivC/eq2dkJe
x0dVUUbf9rlCDgut7gUDOfKCxnweVM6Q81hvmOFg43g4hyHxKkDCL73w9dqIl1CgEO1UN1kFvEuw
lSb/1AAiPjg5E/aLH5kAhbc+9RvqAntcDbdyh+oweDXVD+9ty2wba5E/XyQBEs9P9M0e3jUbHheW
ojm6IlYgyVayFC0T/NaMPXLVitPJQrfC3P9P+ofLMmbbgwWjrVFCLoy7F30zV3/tgavCibGNcAF0
vYoYvLi4E9ZweUwjzaoxgV6+TlMRgxUb4DNe3lR0hQnnrpIagAcGD3+zCb811SkwoK6UXj5cqGg9
8g/mM9x6V6k0vkwO5w/ynd/+FO9S1BP28ueTvadh8ZOR1Rz5ijNioX78CPVGLvyN7oAR/2cjxgsd
qK9OQeASKDfqZJBMsdDi1KVO/UERpm8FgZ1Dc8Um5vxMCOUF4h56N4B7/HT1BjekNkwbxvPuuv7E
YgdyX1cHGRV7/9SY2cz9IXIC7UmvF5JieR5Tay0RaJ8SIFvEatrdfPRgeTFOTkY94DCFaQT7nB1h
EJo0rfcXU6QdCmZks9qZv+yiO0bRFu2AupqqfnCcnaT4cAmiNvFraVnbuuZVzRFapaFv3cnXC0Mg
gRFZnO5bfSZadS+CgyNYiMrT8xk6gxvDPHGAp53QCc79QJm84Ek3iN3t/eyyPFyn4bwXiYQN7sYS
cirm4PtiGLXxuBwUQHuvRzWdbY57hjPSiDNOpW/YAZmcUrM8vPqhyY/JgTj3mZAhPwM2QIjJjSw0
UFCfB7yLdJ4v45kdalEmYu3zM7vDgwJeAvKlfHrG12uOi5s1njwhPbln8cB2QjACtx4PTJEgLkVI
DIaxT87fwdwBz/mdSG4YtcBqukz2oq1xsQpxTUkc6tJSIH5QXVh2Wl/HLBBDUk8Tu9QXPEst0V8m
Vw/uPV2HVBWHZDsRZUyneFrVW8b7Pz63gGq+NvzXKq5DRa80L9T0/5wDfuC1ioBB+DGGP3alVHsY
sNhkDztREh9Jt7pkv7WaQYodhTbBvmAP6aN6sb90BaTbotC0zCwKWu5wAfVAQPZhAaQkk3/lpJzM
TKQuPu9rb7SLMzH8/TmDKN0BD8jGp1PLOuL1Y/VwinrdYk8k3uH5FhbseBOZj9YimnRNNoCCcQns
UVduCvoCw93zWkwuofN2sa0fmrUYxTtOa25zjWT1W3uux4CA5k/AGqizmDq19H97+/mWYSCDYvks
LvzCxf4ikWf+45Yc3Vo2KTxXgnNekIKByAb04xNJgPwJ9u5qCEKHxxBHb9u3ijKYvvULXjZPkYPw
cVAn3dWa/z7pUeTEm6mlvv+BA1BS+pNMpeiPLoZxEZ29U535ep8vBcjziUQDb25Km4lANPvitw9l
QTS+lSotOArrn4T3otBH+Q0CqM5/6U6JclTKh1iAmQ8uYKC6RaVfPR+raeC8YB5iXWJkwj2ZXPBH
F8O5BjXxsRXfPv4VvLNshb5FdQBu1whBW9zyH/H8Q0fFxwNppWxnFze/aGmS3u+sBkR5w2oV3kQq
XWkGlWfbuDD/YFDATM/hvXPtS5zPr9YAqJZr8XTfuPpKwn9GQYB9/Wt7hdtJ2RWL+/qD7BVDR0Iv
de79mtLdm0mYt3nCSwlmMGOcCCVMrFK7CHfHrW/gPUpd65HzX4gN9qHzkzW2bCZblHZMEFqM9qsB
ndvi4VCmfdAfy8ea6lXB4Pj6f1uvY6e6S/KmqXYiXZAYSHximMuseVEf9HcKqMlYSOwRRpxXUxgX
d/R/1XkUKlP9nWKzgHIjss/E0gB+bzYGx3vUjDIhfnMJsWnTk797SaIrtAWa60S5WunJLGJpEG0I
VbQ9i5zsjARbyprnYeNFT8+p23iCsnRAzAsADE4ZpHELFS6g1R7Mgt4jhUvXHpQfIWvKxZWfkuW+
qrA2BBQBX9mW7zcR6VSQFddQzft24cKSyaz63/YazAad3UgVnG0JnYMrkjV0fqgXQ8dpqNRPNxZr
o6QQX1VQrLYtre2KXkhvdstGsvj+qQ79WD/CTNkq2v3H8vrKnAeSWPgeK/qrSvczu4fQXW1PCV5E
MKkK91p5zqxbrwoGna9z7WJh5kHOwfkcgd7FbiVYlYCXDJEsIUGSvUsvZHhs2HjDKSpccN8AizRE
bukxk63unn9ZYb7hjUtDGAh8/zzrBK5ngTHiW8thZGFAIB/h+oyxdfnfFZc8V+2myB9Z8BV+FNsZ
Fnwu00KKAZ+QrZAOUSMZfPZ+n5XCMUn+Eq4E19e10ZKsHiXKaPVPvay2rExmga9eVsofyiMlxwlV
zGwOzvDL09ji6QZmdQdyGpBo4zrrxHjd2A0dB4WcXGfiHyo0VmUpd9jiISlQZUzuMljnytP9vKpS
yXtkb9KyBBaX4wth1dtpuiLu04DWmWG4lkp7j3kir7PYNu1nAIoDEKnc2WYYiThQ4HtnoLnEH6eW
PdaVs+pEv7uxV+V0qRR8zmoVS1l3xH+IJd3NWvrx/uveSHaCEJ2FDQw5h/R6svwKeb45m7Ma7u6s
cxKvfQFTcDvz4qHvf1BUVJgOFv7OEBZ+rYAQmzQ/7agah7b23kR9RzQvpxsg+u2ZbxsoP42qjn2t
H4QdzJDXUcpOxW7m1+J6FlVOw5yjuFJeF63fomtNhbkFT6a6Yf4FpD5fxczXJT4NsNxqzUHWgL5z
VYTmFvLaMozWVFtHofEa3ACRQ4i1TKYpvshYFPlWRTAeQuv5TvWhgnpPfxV0y29O1iUO2eOkzVqR
qgYlzM5uRNhLiKNVmL1bpniYwAcVg6egFphma7ufgamyNT8VLd2cU/5tDtVJ4zuMWfl5OCQ9hYUb
6I19iZtgdKEEWwmGRYseY4bnrVtEL5QhLqh3ggkyMlOw+LyEziKxSTzUDE6n+U5ekhtcVvfOmUp6
BZhVYeusA/6CsBHazcFqk7kUXKW9AZuOtibYhOGeMPNpCw9Sl3lsksD+/fhEtq8mIvF499cBqje/
ZTozmtQ9X7u7kxYwLmK1SEPxbb1vSRUkPaqY7ZRfUc42lWgHNFTsfHxPXTaoNORl9BD5y8xZdW1z
MGdj10K8NSCeC8OKhqEQkZdCB9xGLOLDWsu48jMK5B0dwlqgr5bp7SKwueSvyku/mXtnzkQi7beu
KNVMEafhhIXjgll0/h55Vttz4J6juQtnmaUGRqEqM5cZvRUxaLEKrXbmQ+1pZVXLpgcZoZrJmlzu
nsPFqOu6T7FthLJDpgeNZ1gp6qO9AUKoZZg9dpjmDuBG4njkdf4gZpVNCbAcFzLejATnMGJtRORk
UX8P6ntmYk0GzQDwGIwt6aC+p/Ur7f4atN16zusNXkwTO1N4Itv4cL0TV0GLqQmJ9tW9qRK/1mRY
8hSvD7VfheTh9ADLr14XbfxmgK3XyUFr/mqaxmVPxdN1ArR3Wkvv6v917a4GexT3wsEPMJWivzpL
1WR0GC05QVus3UfQ/FSMX9MFtjFGwfTAvU5kdMEP8pqyemJioNmEJ4RmutD5V6daN8pQxvP7iZXG
ZexOFxHyTGwC7rRuzb4mwMqKlFRwY4GeW7KtwcfL80LM/nruJ+gvtKNOXWLXRyHvJe0n+JbAbPRb
sykNcr/o57f+QR11QlDXtsmUX1QaLxelBIpVlM9tiQ0O23LVvx8QjlgWYE2u1LP33Yv7u7Wk3Xm/
EbGgkIW/PagmIGEx24Wp8s1jyNujtFD8w3d8tJuPkKGPYCqvZpKdifyeB9pLuNS8lZBTMA3Rh75X
crnyeGgLyzaip1gdGiuU1pGPbZnNRHywXV3FphxRPLN7PMjXO9XW0X9ewWCAxC2C1yIlTXH/GDPV
gAp/oL5PaBVwdb0ikvAB61W7lD3wCu0ixkjobzocLcqmm++RLqLyatev1T/GCM/SSCSiTnhQQ2MZ
hN8T+aGi2W/63pP1Eq5sv2+2P1EBvbs/wR43syzKDqSgh4vwzKml5uyOWzB2weMtWJni1KL/WW88
3t0uxd84IaXbe2zNof9MVjsAlPk8Qn7vJt+yFGl2ZLoGBXxFNeKhz75LZwhpaYq4KtwHPGXQR0uE
r9Jpygh0mTrkYqMcMCKbhYrwKbbEgPdhMtgHe+yzGQHAoUzOb3wxJiO3RT63x5E6qGNb6TtRIaXd
O/pBD1WXHSuNxBd9AcUGJYf9JiRJFFMuK1aF1dGvb1GP1Yq1KaRztZhIgJEFQWy2ZfNQw7j+ebFK
wR/+rupUb8z6S7HYZk3pXJMuveApI0qess4ul/88pOqXnQH5vPBw5sgNJ0eTGFDO+41QnfN5OC/k
MUel/p83SF7BZVktuztsMx9eUIv7U3rPgbc0HOw44xds5SjrcH1x0xFEoTD7PK723w/yXJxj2TEc
oRm6eAdo+Chle127nONBq1ULORt24q7VjF187V4m4dxfY643Whu/sF3bKDjKhJhuQMqMa2BuFkci
PE7auH4VcImwXkwD03dwTZa7gVTxvDTiEMOUFByYAsrtzHmtJWKpAZQMo0caXZ72OdJwzNtmHkqH
ncTdZFlbGLBktmDie6V4ktaBzAPUb/u8C1aomd1WtwULkb/+tIBpXbEFbtjN55fpdAeh/rJpdWf9
G9/c4lzq2M7t43Z9Z88G8rUD5i+vM7heeoKXOtnLIGdbszxarrqp0I3wbkliEZqemwv9d8AdBrAs
Z7qHRWrnXf3WTXGI4S9v7G/ANSMZ/HLjZ9QQervCeqm0KA4UzkE7v/F+KwrdG2Ueyxtdlz1d3hnr
wWBX3EXOzNHQVWjsJy8BNm9wMTQK7JsCms6BIrNEIN75Ti0WCl7ziqoxi7Ax5LfGSgeXuh8u5dch
dxH+okTbbEFJVfGUzTuZIKWIWAM8lBOSfGZZVym+k9PGoA+TYrHfsZNJ4Fx2P3wbkTxW79Vjw4j0
Su9Yx4/HuEiztZq8zEijilkzx3lXYtzoPJSCSYutWb0TCINlFBEkxrnWSmf9ZCGeutmVHjucpLwe
pU6dZvMPI2lMFKveCjeiUPFy8UKw/W1inrZBLFKlNsVtBsf8GqYoEGP34ltgjFVQrIJM0OiT5Clv
FhbiKTJWm+yvZb0JTZiTLde45sUKIzcjwcp63WF7hWS95YQZOYQzP7sP2uMv1pAzse5Gj8suJm91
q0cLA5AwjExiJcGkQa08E0taSH+X+XKvejtBT95mGHdYsD9/ePYV8IKD5HZsbvIgX4ZI7Ks7bFeU
i/32NRE+6a8SqKlKzCdCDLbMBBAJO9Nnv+zTtY3WqCf2Wf7YSEwcROfHfKmSMpFQHU3EqPL3/kDX
dP5eWazYyeY1t3mpYQgzCUq1V64YdtnIU0fv9G0n6hn3kpZg1b8vwwmplI9zjJFRqQLoR40JwRFh
1YjvG7lKZDV7jUT8iFQNnxJxYralYHgbLAZ8YJSVm/JV6MjFO/xB4eYAeRKnZ+lDNOBxka+ToP9d
JFnTNx35Oj7iCPs46cDzduBnNCVRuc/Xxk6LOh/0qN6nSRoEEgJWB31bGroFWgARas/PahG8hRN6
uMRzGqjL4NmLHWhujYZlvl5DoT9YG3du/ukFhMavMld+7hgUzRiZWZV9N9y9aovtIHvxh1SkmmU/
nVdZQ38vTlH8YSeXJ/kYd8W9cFGiO6vhuTfFPAtkM8qZb9OO7hZ80w6bbWxNhEQANOjOZ4IlCr26
cyzyQ3IJrDfHx+vDW3e+SeguUJc+sr51/YINpWaT/1S2cmu8nMbL3OlxWBSlv7SHJeZgBKC5hfyC
jFLED5f4lFjzihS6zp816EfviO4dhL05ctPEGZtJOjeJYx34+cbXaLxiHjbeDj7+U5Mm4Mn05tL/
6X7n3FP6IJMW9DMI33eLvVpMgw+Zr00u4EA74ttMOToXmzrTrGLsMpbz4pBWF6l742Q269zMC+K6
YDoAZ78yOwtfoVhtNGtQ/L1azYdW8q2MfrHH9F3tczZDxuKNiH35jblS3r3jF4E0LrjDKeB2zAIP
IlYRwpYcD38ux33J4eMbJksEKx5F2VY66rgbbP4qe48J2N5MAMKGQzDTWUqwIzmujB69VvWCqWSQ
RU11OFB9SI6wfwEip/XVCQXzLMABJA8m11RUOiDmt+7mHvP9M8Z3SOKssmEhXlCXRT4pINq3TA4o
n2i2lifI963tfMwlUsXYM/PP3qc9tbe2tHfCbU5cybtA9tWJDkODlvWKyM0CSPjr2w/4kU7vI3tQ
cHszCOVsVSArKkNSX8WOkVOItT3WI4eH/NgVQDDeGZ5Fkp84yGDLvT10o+Z50So2ycTV0Er2zi4l
w/QzkK2ZGMxh2fskcoTVdIgrHM7EBFI6IqvGFFuJijfAJpeQgAXXlqMjDOwK3doLS60KAkD5qoHc
jwBUxo+zHw38qzG8NXp1u0G4skPBX29JFsJoL7l5QLaIfKQMc6fACDOipmoZCj3Nh9T00xQAiDCo
U4HmetAytVNqYnwiL+Xxo2DHjNlR0YznKwG8c/Pncev1xAtqDJ7OYT4bZ6NTuOPiuRo4JuLBe5SZ
tpyvqlXaSJ40lOW65VkhV1nj0kycOd7SweayQGsKsIRWtLRw9jvLsnU7CQyrOge/EpgbSPTOpuk2
FAuMzHT2tcwTkPnp6625M76pmotcaxBAVOeLxPSbte/jVRge0KcslxpAKnM5OreALlkF2+OQcnDg
fPLUrrBAJpLWMjN07+ZNQ+UbP4MWtIrl5F6XYXZTnDTY2WuqniXRWJOTZH1zgL/Qstue1DC0F82B
bsG/+zuOg1bFfaW7WF4mkyeS1xzCIazIexqHLPX8jT0ansd/hPukhHfkgElRAOyf6C7FsbEnUXmJ
w4eFiJXsfQEl6kNlM20SJVYtS70m5j/ZqnYb0vixjrBYwIFr09wrJqV2cYq/7TcG/oGH48eor2Ug
0Z+TP3DKzyZCIYcrO4RXc6RHRrikgVBVZtkmp/RTkSipzlbJR3OnIILv8mdEGyUhQMlxymcaQyjZ
FVJuNLghiTSY9yx5tPoPzOK/7fwvGxqCBw5whPnTn8OyfoRAcEX7f4nXSrUKdPJz3lcoXeIt8+x1
JLgozGa8SoJQA4Qbc2YGO9Rp2l+mMTqJ30WNzZ4zjCp4RHF546gyfo72IazU0AKlvgqfyechosGG
0sOzi5wb2q+Tywd4CNZ1BX7TQDASIqSRCY3fIB/OnqWNmbguW/5D62+z98R04aDiRzaVfmMjf9ou
CgtPYpUlCg2INv9XnICWoWKGBor9tLsVWv/i8pfsMuSjLwK9vMJEXPG3R4YDE0xlPEGCgIlCHmQj
JNppSfvpisnheAT6bCmKvEQUAInI9ZNDjyq74z0yx+hYTdPkIiwHBWcpSWtTwjRxDlW6VA8DMsMe
+vVDaCem8uaz5RvKSu9FOpKfV5xYzGpRgFSZXk9qT+j0CAGrruiZZtA75hxiL2YO+4QrDD1OQIfE
WH5Q50tirGAk9oHAJ8XbGC4htzfsIOVO58bY6FdJQfqZ+YbS+MLp/l6YfmtNiKv+Dphda4cz2n/S
lG72acIVNomutsxHj/kubj7IqR5jRob/iH9tjWPZgJSA9gTvi8v4TawJtENq8Itd4qhS5MvxlHyo
Gm/fiShbm91/yCY2LEXWT7OQl0G+XA603yRS9BI19iNEdJvkQqXEZpdYAYToIMbyZFmrwu9axkvs
DXG4XiX5g+RE6YsVB/6ipZsnDQ9eHeqS8Gvz08IxxnKDaRxfTsfyTV0+EFvXbg/KUr7ZReJUFSXg
ddLF0qAy535O9OtFvMgah42UuDfoZd7IHYd4vi2Q9ZQAy97MYs9xnFONm3bh7vO8LySsfS8T+G8p
HfcZZjDO7x7+gnI9D5JhIeKW85tw//ARnNzTkiYul4zVTLF/iMJ85Jk9CQhPEOYCTzq+liB8A+x6
bc2DZmitp92nJAKmO6XIpHLn7+t+09Yt/H5cJjpu5kGm4+v023tvD8koR00ts+sIPW7GM8FxzjkH
b30EXBSCSAtIjJEr77e08tax6tZpU+DwkDQ8JwnY7eLG/1Uuu+TCWL1LlYcwPyR3GSMgXEq7sCcY
3fpyrwMLWiwuiTi/ENxwDwwd9bw/o6VDrbU3sfxKi9HK+BDDAPVb7+KnPOMCfKgVgLa+RfBYysvP
rTBROs7KVWvhwY140c15qkKgwG1NtVKN8ykIQDK+2Xr4MsSzfA2EqFJ3nlOjDtyvJP0UfbeRHOX7
XZc8aYMKg7y1vwRVSI+WangtNMRGgNh1R1wg6QM3QS4uIcpepruE6upzbHqYxXnOBbkvnxgzcZrv
9tXlnNqz1NLcHGQhaELTSY/deGs0jjx6+fNFYJ1gLYptAdpXgp0hq5YxRGVxMZ4Ph4RTi+0dkNd8
q+kR2bqJj5zjeUg6jxDg+HoKoY2mo5F6STrF1pIyuVxmCtCYdu+5Q5GHucn11WgAr01G/srQkkFr
aAgSCCYfqGC18KcYwTUxCzUQVTHE4qnCfu1+VKY92MutmVFXnerBXc3rAKXzzop1a0QMaVdlEn7p
Kea08DyibE87+p3EKNsstMTOeId3usWP03TIIGb0+Bb6HwdrnbpfFlCa3TAhhy0o+laywhVH5+fi
P5GS5WY+gp3hYUtmvAXCu30HCOt01HL6rho7gi2gnBS1tsPqmUjGXBq5vIEpUDZcUiEagqZH5dIW
l2zSghmfVSGes+XwTCY+78clmuHLCvW3aFrRfpQP1RQys51RMI8fIlAMemUs1V3h7n80hbDqnQxX
CWvD9Oq8V8FhT3xxysmUeeZDryNwsJTXv2jgbVk+Pu7/LluurRYRTAwJUVKtHpAgPD1/CaDzOODt
cGiyL3Zs2gQ2NlWbkv6RO4U8nlf/fsS00BZmOLiDMtqgUHDpSRpfEInW8KeF3/u86LdHulzObVOp
boO47GFUzYwe+qiswBhA7jgIL8oiUsNZSNoHt3536lvJR+xnZv6BSxMawQn6zT+miIa4OX+uc8Ur
Rg68EIgwjWmFBk93Bjne6tArIK+CTAAeqs5YMEikPQ+PqovbNExcBK/0tqTj0O1N2qZqB3be1sdt
4+9VNuWEdDg2UrsHmxfMYHkKqxkaNIVsH8Br2e9yznQ5d+8jdpKX10yXuiXqA0HXzao3NoRyztqD
JFPr4E5BpuZl28oZgaXquthevfC4Cne1gBmNXTFpOxmeH0NtGyXlwTWZjc7p9ZlNxBGNV3zBG0sn
bivnhOXL50zLQeq8XM1/9FnRdi2iGOkT6HY/OhX+D1nGYnsMN9qG+Km+J8Y7bFQZRZ3le9gqZzkq
2jOHVfO3pi50BKuVkqi1t0ZjBO0aShdbEv2LRQqJMbWR3mAlb5PEOxNMklACO1p3XobYZLAFC2RJ
PNfQWeHfJ4LR6gJJIpCMpBp6If0eRpM/ZWvZMJMyThBLe2rAsWBzYlxJvlMdrV39sBRcBBJX+0T1
rz7PKJaGlXQUkx3u7ClyGAH+rH0bDINrQB3no3B5VjRKeEwVXKkdEDODSynIcA0eh/g3T1Jl9mHZ
9GjAunJCDzZavU31pgW2iUAYXxd9qvTZHWRWTAHfcgBFzwBjxjvaAnCOOR1NqGROQQTYshsxp9Ei
D0XxnfrUUHWCkGwdkAzYk0XaML1cWihM25NEnlmBduwASVHxuKLwS9YdM2TRsQmgWMCCWnBsz6EA
kNWZ1CXHJIApT4tCqmgiXdKkw4v+80lChyasJY1PImVAYldZGoALBhQ4iFBJbmsvzoP5QZzApNt7
utHJxNCTswt9mfwdqO5ycL2wS2T1JZ6wIszlyCTXUBoowY1s/iEgKoOvqxapnsbbee95W4gLWrjq
J/YaevDT4AXuRVFqGiBlFKyRHR6/kTHazeIUgryXw1aaDWwbRhz5hVKbjH0PXU6EJhA7W08c9RDY
esFh2TgiiKTs3yc2tL6xfcpn1+9sKxGMOWTuM3Fh0T0ibNFi8vsSuXS/n8zKsZ4++YQNcj0+BoYu
zXXNDSoUN18n4D1X4ItZGTsC41qIss4PHXFb5Zjmg0WU7+9umkwopFaxzaQ4irqayijbn2NR8m1c
hHLmSTS4BS3BurhxSCQJ1H7yHr1iv/jmzZ/Tr0qC574ZZzhTgTVJHUSEn+wg5lcoGi0/i0lriYEv
MpDsaGaIy9bTZiF6j/YZSbJQrcxcMU1FmgeZ6KzbtrlQbW26VbpY/erJtOXO2XAu3cIXvz7rb/Il
7e9SSY17/HoQgr1KTcvy0Pb17traJGDEv2pENUftYevDXFHk6pqlm2P7ZSb2KrUbNFt7F4Wb9NvV
h5Z1xlHKidYMoIYe9/zAqOu20CsBpkEl1OWh3ASxpT2XnnoHU4CFAHAqrCWgsiOZOJT6SIq0cMWC
52dfTahFgIbLD09HDXQplXWfgZH2FRMoXExUDFw3F08N95tX5cb8XfOPu+bzrbeCXNztDuuNBg6z
N1GC0N6U4KjfLMKJ8/09htw7bFGTKbJ5T/DGpMqy3F9pYD2llBjGeClt9sa3URv48iSyY6/xb/9i
FrZM/WNxKG093asDW4WsxoWC+l6htNK8sBrNoWorBkW9ktrzO9RWOAoBGjFEA5lKUpM3EilILyz4
1XhFsU5NpZRJlyXP4SxQwC02m2BkyBkPI4JI+hzNcEnPUW7i5nTTDs8DHRiKfLhhl9oFK/KaBTfy
ILmZhMOXOibGE52Mb0u6gNa/2N1h9j6wUlqN0FUJ6ZchBx0oJuPTrCZ+ZBRtVaMdvk+Dglp4HWui
WeM4Ar3f7YwIuso3eePv+tJJvauNfikwuVb9V69Rug0D3Z6N1khyDZhuNa4KQnv8X1DTFtdIU+m5
YpjJa75tIjuMN3Xzi892hrvM/BwIs8TzLiyDz6m7uiaCF9N9VIzORUxMGUokLzNu22dCCRIeO/B7
DYmCVAahhCxFsVLrXfEfQHoVzxwohvJnjag/8aHHAVpy2uj8Z38lVw9hEXRR8gSEoQf8m68Nuv0j
zstTAM72kLRjHvHbA8sJaJwWwpbBkzz/hxGTdZSArZolE6oGXCU6K6rlcxMUWUIDELyjPdOOwYZV
nBsB8AJqAFWJeRdELtW1tPVv/5nyT3FZsz83wrpRlb+anQibUQvXM/SsC32Lm/vKpdI+JQw2SiCc
utl/XsYaN1FHoGHVWV6pq1/jl3Mcc03m/uIGRyoC/iG1kixEOMTY2aZS3RNddsX8NhF2HY4EbQ0H
3Ym7lsZBwownO1gxYFpSVXkoPmPu5mjYmX//BdboRvLyh2n+Pqk0bg5+fmCm/wxgksTfM7mbMxJw
nENEWqeDTxPgLLXRxRs7VoNJdzfY3tXMD1tWuuTbfEPM1asCwPsgjBYOHsai+j5QeL+iJVk4Scy9
w03vWyt14Ny5WYAmXrt+GWccGI/UYttgbg2s55iXi35g9kShPoJyWNb0awGOrrH2KvLXUzQ6iJO5
3ECH5TpVTKxEQLozKQww3unYbDlx/CDxUTP0B1y4LP+Z1Nt/Z67NBcUBOvU5u41DcwB//h3M/xQR
ebIEuoLoYEtwOrGyhwsZVM4OKH6QYp8JqqdqADPYj67r69O7Dk3GMqrceqV+iU3a+ZOqcQJzbzhf
1874MM/Yxop9+ed5aw/eipIiW2q+6nos1R7vUdXN/zAhEBcNBin/q90srLgpo8Tq2tOLsxl/1K+6
/bKlEwERAN1mTC4LzUh41GNMfuDl8MJr7L5buYI+MpAyoJLoekbe/6CTPPST2j5rqo3FPgsdfqk5
vKJbMZaaMSxW55KkqwXP8f4xZOuBH7RpDSN5FOtvSm2PBjq+qKthzFRxwHFwRv7hIRDQ9h2/vG0r
T9REQWb49F9Q3rXO/hd0W1RtLX+1eDWtopJ6Xix1nTccoY4m1qwKxSnsnMlkYg2APQIvw54SUfTn
UNzZJw+DCrEsThjkC6qlVt5qSmHJ93YgMEj1uHvBn7Ao6Yrgp7+aNqtNm9poeN8/vdmeKe5/Q8S8
xQryPRWIAbieMLeCX/LLWEV0SN5FbEBAIZ+c+00iDtD0CR7yEKNdQ3XBJ7R72sFGN+YPI90ZZn/x
MI8EVouaI3t0Gon2LwA7uLrHbOTeW1/4ZPU/nelF7TvXPWRyjcSLT9C8yWlEkMv3utLTDT01K1BD
Rq0/7HHcmGN6CJKbGBg/AGRsmMstyatEotVYX15DbRvhkAyEDsSME0c0+fm+uibo1ASMdg7y7pq+
GHcQExwHd1cURuyRaUZ6saRK3CTJmttRDyeuplS3KUMRJOcWqnsTBr6Z8pIKZ+GxLqTm47mNkbik
IMA3RdSBF2LcxfcdVpDg0++piWs5nPB/xrQyjMgUP/6oIQ4PmfD7FAY80TedVV+Zod4zgYCyWucO
BTlDHTSQPduy1QLpjfn4G8O68uQ9RgLySCtbXf9g0v38q+qpmJoLkfwaDkXeUqb//pTUyM4i4kSE
DDAh42bElvjmtrICbPxSgbpP+m3383v28S2PKTSERTdz5UH2iSJGJePDBIE1o8/kBzDWgD4B7b8m
LYV0R/JYDZq+NZtLrOuNdorrTclJWzSp9s8e30rS0oFy39+YlU7DBaPOInppgV13rsAUbPQNPd0j
zgaM3G02Ccel7AeQ0HNopp/4oz4mEFOr064OgaHpvuY7Bw956eUbAKO6AbBwjvwSlJhJiJwNIV8B
dD7otC4WYKLN5YFFZT7zakz7LaGH6ncLjjg7y2xFMJCLQJTdCLnBRK3gWuBosDAFXTgNXg3JQc1r
Ha853Etb+3nQjrvRtu9WYnriluo7VQhIcZS91+7zu2Bqg2lekrnX6vUmyHpda3nYS9YfUKxwHB02
sg0XwuuX2ClqF6qNdS7uYCdcCAnwmKDHO5wIpiM1UaY6t9yrF/ZdpnDyPeT9dl/ErDHhRfKQW+V7
74xx5P3A5blF16CWT9xqyoOsTs8acTrxxXt+MFG66Q1oen/gWs91FNfNJDLM8u/puvAakaQc6Aja
0cGuKcdsi+QQ51WQAmkSRok8/YMHujLbbDS6eNrjZu9wYBZunOx71cGU0Vyp0r3rofzlTXqADoOc
EWG79Eyx+B65PpxYvgKrWSeyv30LhhcKl3KDLptZdE6cvKsLIPANH6TWK5SNHpVVEfAru3VZAaYw
SnNmgzgYa0bqCL70i04SVCI8UQJ3veq2FNI0d1p/zJkKY6rVbkv6Q+Msva5BPweWauvMatEkkFhj
7ORCw9G2KuLd8v3JnLEmiNcMrVkALT5hr9AiLmUBsMw95Rzq1dXdZEqyl6ItmcoxvtvzFh+Fd2VV
LNx9srVMv77fKzA7tcS6I5B02plgWLBl8t0BsiyeG6MGtQ9Jo4VDHs2rX9/tLFUNunme8F6XID1c
x2EiCiextQa88GUuSk40yOtThveglhsGootRwKcm3jUTZhb1BYGw5itXo+Y3UBMHNLpzA7+Oqw5j
P3wpcrAXZEv/Mf4VXmiv6b46jMmJOYlshXQECM0Xq5GBRmVgRwYS3Z+Z7cJCGGDNzmFnLtqqyDUV
80S3j4bfLQPeXDSQx5bQmkuTA5VwfN+zNs9KKuCLLRS/3KpJ+GOcU7uRIqGnz0sid/R3UMbtWp+j
4T0ENwI9S0v2And5ToKDP0K5uH9UOgxEJpNxeSjtZ6+n6kCKGndP3PhxnUOfCk0HVIi3knX3aFQ+
CVxkL/d0E62JeooQs0xAkK8vWA9li2AruPhfdw1TPWMTU5fOXbeITJzJOoj5a2RAO0f6W9TqwE0h
dsolWwLvp+iwKWnjAScsIewAnVK8GE5q5SKVDIBJPbphDbvak39YFWAjUm9jtEoZaS6P4ihhieC4
fjSO6Wd1cCgfzf0nvD3mLg2i8ll6e8QgEJeJDh2vskafq+XbswYWcCThgatXF7tT1UfS7UpBoSc+
kvFAP6D7eaqTPDaMGmy+ugpsETWGlDRffupQivlcffq/RG2nVZ3Hl8kYrf76MWJcSTeQXyN2jlfJ
SyaDOPAaQ+nhyp5DQy8kTEVIFyudLkyFGvUFamwiwkvbB99kfM5w46il8bwUH0mVNt1rFPweJwa0
Ooq0tcvn+psvBEa7BrRPivMAnIFA7vwV8uTENi8N27iBhVp0lK+10vxLU+X5Tx5GrBfsD1AYWHbo
smJsCxbRauImnQ5w5VqlMaXBeCZ6yx0Qv1ZEsHjRcOpoHoleO4e+RUkGyePi/ZQea6wIAPoRu45p
HLqdnuHJMI/+saRWIFuFuFv0kD2AdOpv2ZDjkYqOxexr6LU1muTmZxYvl0wVzEWzFnmaX+YCGurj
2YiLCVbhmTtclkWSEIr/tJ27Pj1FwpwJW+j50FGRhhyPEo3Y1z9zkBC+lJLCYd6QkH2EQid+Hsat
7FXFel/d7xB9wIbQ4Gbg6N8TrZsSvZRQagCHah+eAR9W/Fqc6gaGnUPiS0hoV3M74LiBIGcsOlhq
XRVBQ4IiXn9hGReV+Lo7GB+lNWo6evrNt4HwFDk/YoatYxbtMtFqhNuYJduWPOQ7lybIxHOr8e2x
L+gyPq2PFMlBKJHymTjg6zRg932qhl8P4TTWfL/CuDCTxbPTxVZcD7/9fVpe9EtQ/Yih3SBwBSGP
FbgoUTAmyRK3WNYk28p2MeCD0BMruLB75ooL5wV06mKb3p3h2SMfE8MGqrHl1vNZW+4hPPaRrXV8
tuZlkJ1ePpXsIGdxYf65+NdaCROZ+Z+Z5Rxx0eCo2YXRPApGy0P10c/TRZb8QGGHDbt+o/N7w9hg
mXKLv3FSj82Hy8OL6gVrvsVIWCrQ1DkXCQ83/YS7DHTIQ34S7kp/r6XBnTxZv4M4CY1AL7WLsPZu
k837SRfzT0J0sroKAm4TFShOIeb/WfTszIQEimevuWuMFzvWXkFz6ToY8nDd6+2FXAMi8bJI/06c
xHCmJA2s9Gde5sTWSzjKu3BEzmRih8GxklBBUtmwF2MET5CI2pSEqxzWM/U69ixQLWR7VH4hpXNo
IlcLvkZ/tLIiR7m4eJn+GRlzF9PDhVqNpF+O5avF62ZzsdFIDUW20aAORyjLA4TVp4e3eOK3bSPT
1uvo+wv+AR+Pz4abh9unkzWs52pAFaohrG7BrutlAijI1OLTQCODZMCFhoYUIcd/nvL9RyGaP2KB
eL7FC/HKdwFmPId3aoQUbjlfgPaINjnEJksF0Cgd1uu3ep7sS9ERA48zVbFLz+yJmvRb7KUmmajT
LhXVrd6PRbwS5my3ipOEVf1EHRt+LKsB8Wr9M4xu8dx6JpGjZVN64m2ddMQPP8TTxrpm1cAQWOy/
CAYb+NkwqFz5U4SyoLAhNTFRaRNOlxXQXFe1tw6fCXS7e6sAOGrfBFlD6g7PFLBJ3UlKNbBpxOul
lnRgwFUiQj7laK3/tbZ3XCKCSoyp4BWmH018E+Wf/WZUe15jklRCwVYiG2oAw8R4KD+d95yi3EVF
dgjU7gH40iJOgQoyprGA1G2vPle27RRmHAjtMfRr/gDIqi0qRXkD5w8V3WqcRD49rkIaHEbRuAjj
8qvYcl1/5gY015wBlILGYiDKFPgXu2Hreb8E0yi8Kixlukr7MUD6gRsux1fVpdODPkLi3UPrLWmB
MT/ZvV54a2FVes7N+SswkG4B0n1T6BB4bURdDIiQdyPD3dX03UNcDLmjiVKA0LDiMA10rgFyvJsm
7gXls7l+uPHpZYFPUT4BicpfpYYyWIpPANQ2Vq46e1pJpUwRGt4ezmUCQdQ4geH54JTrZghBXetO
ftNQkjxSgtPvjUtoBBR3uHpC+VcX2tX9mSnwuXGR+hS9Zcb48JuRgopQ91yeaA/E+dMk6xsMu9Qw
cjwgmiXNxhkBE6L3bEpuI0DhIDiBPdbk7DuqLa2SMA1MmpfDr/5NdH7vDdIpEESwLv95ZwuD229P
vSrbyF080JZrbZLKmsNjjqbV0s2VsWDGFcgOWZMzUtTyf8gAd8vcU+Wgo1/A8qavoUUHK2W65mVs
e3PyoOlUPAAxFpdIfFGP/q4g1GzhxNM+bDggTPOtL8ssnd6xaTKMIMAbcDJ1IWW2z+x6JXGgYgI9
1LNV7WyGrEbweQXJVnmOe9n2AWdcHg5mIr2dZNYMSQPftXU/hihBACV57XhlNAGYkzoYa9ie2zBb
njH5olFBa3c1wfyK1D0VtqGwi9sLgjYMTKyW2fTLlTgl2DUjZHnITjis4kx0xFjYG5xOR0EQyldI
gqhy+q5CWJtiTjl1/c4Qf98oV0fMw/0vUrAcSGt5PtfvT/3C+ZGUry2/p4yEvKPBD5iV1O959e0g
dmOQYEfPtinz/lCVsree+tCDHMKb2OqMHP44STJQXfOF/FkNOvnkeHzeXmb+TSzi7Cx8/Qd9Xmpk
eR1IaVb3xr4E0zcwpv6kgB50jLGWPrJX8rqiTYhkcDMTjv2mqoULYtZdtkw6hrPP3kbNWZobBVSq
wBludginAlsGzybcyUKr1+GsBBsvLjlrf8vtFEZxMp4zv0cVPCms/vZ8oyYY4FZQsdoIILcraVGl
uogdr/o9iQ+YS1dJ7siS4+260VN5z6Rq4MAYxVzpU1l49JlcxgCurhmMnSS+gz5q/1mJr3x4kSWo
0gLf7/CqpdOJd9B22z7uP1XIlWm8MWR6SAoWbse9MYLQG5IxeJy99eSXj/vIjaCArNayXy5xAfyx
yH7V7Tur8AZcJ2OLN7XpzEJbbY6dnk06n678WwBFQEyiskEEamvHFgd1XqsN3YjWB+eVYz0FH/2q
F3WFqXvDqH1u4e4tnVO+qMna8vRYSO3y+nRRWaErI9lAymZCPWewldZQ2bl7T6AIr3iT/YbcKdT3
l2ktvurLsrxbt8fPCwSoTP6V+pJmLSrC3U+miv0DV16wj9AArsC/iUP14YOsWfGnJWGTJ5zevb8q
ECFTvxotJGuYAPnmrOzr8X0jm4mE9hZBUhpeZ5o57WwpG7ql3LkvcQoGthDse7xPbO3XxcOXitcz
ZPTWVTnEpDLj0PKfSELlcLETbWr6GTjTvhZAZ4ew1AB+KCD4/4cYXQqZO9Ob84PfAr4utD+4JvHi
RgYUESv8yGt6vebifBSx19p1WwZPPG1/l4cBUehK+4UoPlYRKppNOrBY3OrODKJvgDku7Zx8hENM
ZToonF2Dh8tsn2QujEqgcZucnM7bjrz5A4i7Je34SUCX7y2LYGWWhxnUC2GpRv+ncQMrBaBIfxOa
IJZOkkmA0kEHgtfUgTQJmaX4aq/FpUxbBE6Bf/qoo7K/c5zkD1IIqR0yvrX/6JeZUnOufcOsJT9D
EPdDWrNOG5vUicbxVQQUsd1SpmUkHQWCmc2A+KGXUgStL3GkiSJC9uChZS2Dr1uYktnZpf3yS8W0
1CON7MUxWrmO86JXPuFYFx8ay4nkMKIdazWNV0E98Eb6tChJt9KZF9oN7S73Eba1TuGHzoqxUj/G
mzPjcZYPFHsgNsm1tRWgqbd5uupuEQJkNjBitwrf+1fFO30dd0O3SWcgbfD4W4mc6wR/GOECb6ne
V2A/Np+UPuBiPC6WNuGRR6YqovzQxYxp2gqTql9Rn0tqIJRh2fFwOj23b8lwRYLu9dgVb+fbJu1n
/5TKI6p9Ur2V2mC47kwAK85auX82M+/liJYBek5umzpeYH3o4O3DDkYomnq3T6ar4BnF8Iy4TWYL
jxBcgcySOxbSFaQQA8GQW42l8kEVQDCHaPoze5AUVzWDIleZvCMLaizqC7+7cntARCaDIJLGbGWj
J/A097ygjpCHUkL2N81C96PDM6eS/uxGpQFkbIjH9qVaNrvslXlV9yj5/PTs7hP1WMDFGjWpGidb
/dtzXnJElXNQaDibO26K+QsEwHg0fhOjvFhckUbmHjG+RYyeoBCINOB97PRR0bdjMuhwq1KdO71U
L4Mf4F5W8deGF+XoHmpHc0G0+Zo06uJ9qRoaC5zSlowHKug4VJxOzTQvdgEkCUQiwB7uMLMZqy/X
KL1xFy2lf6JNZgrAugamDJqMGdA7Xv5alr4RE7b/DXHQo2ARa7hHN8CKXiomHsSCvrO06GXvaHoX
QJh+okXZQCKpaTw6jQAZllfznZcH/ymCiVYnu2nmeUA9XrifwBlA3+egrGaDLXtHixnkp3hIu4cP
xsheHKzt6TW14Pr8bchh6DciVQrMbPwwv+CW+0tm2qLx1EcicwuaKfmXhInjeQEg8JHOc5EPxJIb
ShJhNSuHk8a7GzoX/dd+l1RK957OPVj2z8ArDKKTFQi/gmLi2YxvtCMi0kFxvJbQQX3ohYk2u0Kw
HAh8zmzhyxZz1EA5sm32l7NV3g6DfHwMjvk39nYEnOfz1hWUZqBIaeJClkYuReXEszi7fChsVXjx
Afk+Z7REcM+kI5EMXvzUJ+FhEMZ4wRgrcDB/jkbWYK7cEzee1dongcI9B17yDvQ4UqSpA2AJp6hn
pS20zKRlKBcvPD0DODOtNlN8XlbYZxroOkAP1Ur02uHVdBs7YrOUzcT4gRgHHVQGzuL6nDqtKO0w
SAL5uYnPqp+dLEIJmdrx1u6PpxaQQl0WA3QwFlHu+axoc8EdQ8t2op1qJMPKH30NCA6MdocI0+wk
E2nbVKyJYTRm7zXxWiotC673eRe3dTINPmFVB7LYwaNVKN7OS+NqxOzHNkgrZ/M4047BLUKgP+N6
BMAAFYo4OF2IyC0itCezgaozqGXJDYRqbHPV4u2F0Dpkb3gjucFIJqp9ApylmByfn3/8TYV3GXrm
w0CMicImh5BNWUTMJHKs6Y61D6v4pFPc8LMwTlZ+j2uPJZy0+3s8D3cINn2Q9ps9HyNZn5838/L4
DBXYQHCDFdI2sYKv+UDnb5swue4IwUPkHEps1oyxi1S4BPcZwFAo7XLmDbluYWy/WtdKiIdcbn09
QVQGPzQWcO399yYBz/ZFCSWPcfv/jSJJR1rDkxoMmzrA8OdqWV43S8sOthGyjJuoIbjA5LAQjVxz
YA7K2ZtcDjT1Jbp/qo4JMvln6SGYovej/zJ+RUjWJO9KZD0g8scHwoNRV5zHWJvE3QN1gv7PsB6V
juFc6yja6tUETF6KHr5xXo89CQx83eR0v5lu3+9FV17ky8EbZ0P3Q5V+nGhzJ6gtf3WZqIZEqQ+0
37CLrahfdGJBxKdJoHD68WVVrxjFoooRcZtSgAszU7jQCp0nTYD5GSOkeFWEfAM87hFkzyRBMKyd
GvTQbirkqw+YiwSrVx2yH8pnEkry7UeT7JAbTfywXuPszWRBBVGyc1k6L0cSDjlA0jAdFq4Gdo9j
Qf6qsjkTgEiIvcJtdZ5DnjFxnGBCp/088xGlMr+Drgy9apHpobLQIf08By+M1KxU0+IaQdXsk2w5
GvU8QNk3I1COJADkLclPooa2mN6R3lKELzwnvDYADzJTgExrsa247lp5yxKWxlSMsLQJnkKUq7JG
TwE90gVxt1a9jRQ9uMH3s2AdPK3nXewLa+R5Oh7fafhzFc+21atPAySSD7eXs9bvz2R7WSL8jcjI
pFRWBd/fxt9S7PJvrwB9LAmEfKymxAOiBpWlyG4F6+fSas0e3NTGq5Ox+sonaZdQte5u/TCnf74m
u3ec7YcEYQcNHfAcSSQwfWy1H0pd6NBZ0QKjxHJYqsYlSEOXktvQJ/WP+p7npyj8/tO/p85I+0xk
zWe2DBpvIgcTlca/49JK2TnT5vBHyx0zr0CurUiQ8Kcx7VvKbr48XvMrOgoux/3/d8nXHbZuQs6W
77/Lggiw3y1FwVZmUVV6hAmE5pNmM+g9nthaOg0ZBGPQdak5rYX7UZWafzYp/ahcd413HHaLrfZg
U2MR3OfUJxp4RCJbJK6Xf2HxjJPtT13o+kID6F7jyNdJYdgb8rqvlyb2025S3utLk342AroI0uYu
Upyov79w4hn2pZDjixEichEQ/K6jm+lSAxcgl4DtD/1Gjf++FsZ0DeoUx4qRBuki7HwXoNuI2zSW
hZqKPrjYZZk7Pw2CsgpYmEG6Con11/kg+z8nS/sl3OHxcFtZkQ/wt+V8PVKz6bTmoBUXMcQfa/Bo
CDAFhxuoeGcxKyzNrHydmF2D2VX6DqlV0nk5PpcE/Qi5onbXuBl47tEnRFEFcXhnn1R9vmy4Bo/G
9j/ivGpCOrji4Lb0yFGJ5f5Gk3OOrSGErsAQswEp2cMFwvE54qTmUzC2XK0pdlwQ9RFeCfAVrfE9
UylOXIKtIkoc/dAsKOPtuNV21HR1xr1NuSUUzG1cC6t5wU8T92fYVxwKRJVfL0yZpwV7+jPfALC4
VFYwNJUY9ynqphKjqcHHH/fujVDzWEVZkGwj3mOVgTrlekQDw+TU0vesbNhTctQvGb8bKHjiS0mP
dB3qgZ7eooJGJI/SozPXw7Fbu0iYnOpygJHKNt4+Jyw2BtkCIvhtxodF9DmsMxQLfg2s6JdKHY29
upR7rhSJCYa3ltyCKTTCAkRz6yYZskm6qFqMH/TBD5WmYvfOYD5hStD4EyzEQo3RKwe+3FfNYAnf
8dlHp8SjplFz0J7zllvDPa0Kv6nVtWXbud5D0LtmZRDtgvqxZVqt7cS3gyKwm4toxsHByu6ms7Jd
eD1fhJ/TmIsuoMCG8XBSN3826fuaSPsGrfyQrNlkmUlKk+CVhCRhjw+76VjRTFIkLm3LAine1TWN
M3ozB6in0SDdnwP1uR3EEaUvWO372Sc/NnO4evQ5WxA2RZq5/dzjR+huRI75WB3zuEkg/dZUr6v+
bVzYu4ZH8XvRg6sdpw9263WoKUrAvCzS9mqWbIjMDzpHIJ9PdTuRjiJn2RE+8FkTWrlkjenDgE5x
HZeMPB0er70B7W3ZK7i6nyKaN0WBRp/WrakVmZx0OvvRW+SJSP10pyaMpswlzRxt4nVe9h7v+BTL
knR1eA1zXzACnt4agIldoF+SmjRM23t0LNAxxQOxQ2q/zAjM9ze9BVeKqU1U3HvfnxL8oFqBVLWD
2z/qMtmfciq8CXV0N7zomuf/2uCx9ilD+eUxCi4TguB/U3z90RUY9brW+oQMY7NDCCEIQADBKWwn
XW1SK3F87Kb9FgM4lAp76fnF4vD8OealAD9UiX0bptjRWS4XyaCtPQysQG0E5mYsC9J9R1uR2CAh
Qmna0OEibWEB0sk37M2qL8AA9wPHnAjLLfkKSYvJepI1L43omWWUugeqGqiOKhfcJiEgeNyXagDH
p0a23P4/DYCnQptIYZ2iWVDMlz84Xc9p0zeFgy+jV/VNDPk6il6fCDenFvIGabUDMOYy5IMaesAl
dnigHRnt2sGS4V01MCg7grzwZBx5fGJ2Phwsw+meOJTTz4eDD8w6nLeWP71aunJkHlAEhnOwrgyO
Ue9m9xhfjndT1dsajINGKoHzkL+fiklbc1H642sqdeWcAN43x6iyWRtjaoNieHwow7P2uLhX9Up+
FYMZabcX0gGWw5d253rRK2YfJBxrGFsVYhHv6ktyM3a/6PqnyhJ9cee28ic4Sg9Y5lZNK2G/XjYD
ta+gO94qkV3Jaee09mtOURnIexBakZyxwpxGm3qoWLGOswNkqObdJeKSJ89UFEe3rKCMMdhgDpkw
q69PDHsBX844phiqrk8hCwg1kCxVEcWjGoNt8HqzRtLJMY6QpJbRcwafBgJziw0X8G8oY34IuVMY
i/QnMY1Nw1RGlfDaYS86MoEmQzj2PYBrTNhPYWguODKrBXd9rNCYbnsx+UbSLsegaxnmBPeg/Yey
zmhpDi9vi1v3dpcFNbR+QNmYJCZrobpjMDbn2AxtLWyaQv3wrYd/vYWExgepPybUVFIubPn4zPay
Bku/PSksIxHbFwGuzJwBxZqPJnQULZo3QCfsf+I8JT3KRa2T7EBGlxdUyI9zoZUjDEISRUDZppG4
0WtVD76ISIMExMOj3vkA0+ZyDaBYKTlMgMj/Zyzt0HhUgWlraG+bPkxzmsOmqEErpW3BdzBwcSrk
bQw5i0l306Oq3GqQFWMiZQYBiCexrFXYX4KeZXFVLQbbGAYByuLjilweX51Yb4f51s7hy27vYr4R
Y56kjMftmCCZT7i5is2DbkQBFzKIbRI6fUjnGeMPRKl0SSxe6WGgZWsVGowintKuZbRvf+CakJ1o
q2YtyJQyKGzpGJivTD+Kd/fgxKb6Sfkqh2t6T4UayNxuD0+CTggRfWAMQl6MVIGqTgm0JEhSoPrS
vfERvP8mz73J5xaaMY3YfnAegS0oYyPIk9vGooo1OfYgzh+BtRlEv751OAf4uB6ITyHdUCw/Chm8
sniiyj3DgG9WrJ6ov+7xGYxD2bVTh+RwdrXtaPDpa5NLtbJ6aiwlolOyVgOMlrDFgjeFHMHJmp2j
tvaO8Vt738E2fYDHRQ3FXTX1UrSIGwlAOaZaPAZhAy75AFZ1iQ7vm7/Dzy2CqQYnYD3c6xnhQV8e
0FyesF60sjg6HMmobrrY3RViYu5+Hb09Hj9zwzmToBERKTx8uJwzBk+igpgsvoCGk2f19j7sYMEr
cf+WVbs7S/A1RvNOxx7GAd7MpZQm29L9h89dPjvehCkhJq4ymmzP0CQJX0IngsXh7hNkTX5sStyZ
p7f5TIb9ZKQ5bbxVuFyJyY1xcWlBwJybiSpTFGPFbAS4O690iyB48P+uyukZxfbhh5HrZGD+SC+9
k0moqjkMbYR8X+/GONLOGc6oyBVko6AiDV1gGwPLVIL6Oo67YENoABOvcHAZ9tsTCJ6aX+38HjF9
J/qnDsHfbNI5HgSV+OXl5/Y1eSOZSiHKRCAyRnpvfoSLb846OrEnXXouaG3ltnHC8bY6HzQH8j/Z
cuh16QAdpEiXPX2VMSbhpkLKl0HmvqkpjqYefABrQNIXI37ho60aGlxo9PrhGBaXjp5gcUjHla2U
DeA3M3DVQPy0YMiPKZ3pwW5p6Y2rdjYoh2OMrmdgP0HsUXXZDrncxjmiOYSPg0GGemqEdRfCX4g6
RjeCm0NtooM75G6z3trK2OsNuBEeBv9vYVPrhe/PJ794FsT5sSz7o9VhjWsqLeEX/j/2FL1DRIuv
LBJDPHyHhjRorYMN5FqIC3D6ibYbAQtu3NExo0hLFEyrWlky7clJ93AzPWk/WrBRm+2Jwr3pbu6t
EnR9WUgAC/qDt904pVy5yfIuCLFvLT0VYTbaXDaScDixhOgSCGFoiC9xhaNhC/15mOXKqrsCxqw3
j0nwZ0HixRYK4cqp4/4mzDFw5apRCS1ujVQSIHE8vc/tgwwQbRraCT+8XIyD69N5J7YiCj6o55gD
OcZZw6K1zvj+7hyiWwN2KIFNxriEMjObG1Z7ySbsl+MwBFBqYqg5SlHx+ZHtuGyFeBE0X8tg/jod
RMAblXu0DSgXkmZE9/r6fY0xfZpXEXvlOv9F8nVbLbD2Ym6RZaJ989mZsOH0uz+4x+2+9TX0s+9O
LaxJSolrpjqmAHf8JNTv0db+hx6S1mXw8q4EASbq6+vysaADCrOyrbPLVsG7+yV6JH70oQGClmKy
XvrrpLtPu4ky9wpD5k3bb/alx9EDM4AEmY6S7vUKNiyl9UBUsApjnv4+QwPNrPPZwdY0MCTeTEFB
xj6aTbkyN5ZVn/NexV5skWsBY/o6oYM3Yo0WdonsEX4lSf28KLkq09Ahj4G+ctFSggL4DEXp6VF/
rRvJaK12v0YgYluVVL4IEvPeydifuE/Yh6NqxHP+uzhRO7WTYjwn8iDQD3tCypwCAS4PCmM0D/OH
PeE9ivESxNG2v0HBOdZdDkmiUpxDSVTxjx1lmwKF8/AH6xs8uCeWq46CnrxjX9MhTDRC68wVdFp0
rIwBdiwhgVlMaFNLwYKSsp18GhMyI9HD7ADDhQEwEA6CggZ9kSOTQrRAGJm6gm2z8Ao8O6ytkKLG
qaoY16GBLGnfNePUnnJdr49hPxRq8vDATVcQ65Da33E3NQ21H7NXFYHcR5Zxm7B+eWIlhtfnptJj
ROW9zFlJk3sBAVE8ytpfmHK83Oa5lhy4QcCpU42I8xylueMpw9QibkK9Ewo7Xa1dGx8oI3EoKoAH
A35veJEk42DpJhDH9JgzwRmDW627BQoJy9fDCISVtAnTkhTBdeJnxe3gUHIceVHAXTkw6MOM7THV
/bqmt79c/D8CSQixCtacK0oRmhB3+9SRnaaluyjpeqPWQjgDmN6VkMDQEfUz/j74wao0rMzTKP/k
YEw662+FjT2jOQtzLsaq4v6haPW9Nwlm2xWzD2f98F1BDxI0zOLMFlas6/3bjY4BbmCSr4vI979Y
ov3nwvPXU8p0BIoVdjlZwO778LxfCxITPkqPm4EMCtXXdl4/HOqG/qhWKPIhjJBZHxGBrMutYavD
AgWfHq4TAYwgDQ5G5nOOyBtSN8fW/ZzNV+IsDDnA9YLJ8W1po9qZEqpG7J20llttjJMHluo90pvz
H4seZtZIBVvpUnlvgNfpGdHTGf3XAXhpqh1i5et21d3Xf6EaNWEjpWAlF2Qt8TL4pVvvwU/sA8qL
9T+LElMCyJoCEC6etCKafrWDPtKm0OvEFAQq6b+Hos0JZ8j9QxPyKewy29C/DNxp1CgDLx7ELqe4
zWQZCQ9cFVQxHL5B346T2kzRNMxzbLmCTmzchpLaOigv5nYUbLG9p00s4IYK4Pw23NjD/euPRzpG
R3twK21VGcV4egOVkLmM3PRShbVI7BxSELQA6Ljg8mPEyWlnSfBhgP7GireelmssHEEVnAz1skWm
5qQeTkECc2yw9VFdYdGCr1/ma5pWCf4q+3Q99REfYenzCT4tVGaTMiWEpMyeTBJr1jF7EMuxbEOk
524IzqO0EOoiC0Jq0jXkje8Tdbq/P5QIHMktI6iunTKK7f9zSBKKtWE7uNwjdFQWIU5i7VVNMFl4
eLiiamUuebq2EEzpqUcimE6NtQ6BaIrObYCLXGDhZQNHeNJ7bHtX3cSnXOh460+/41YYjif5qC6P
kT/pYl8XsaW/mQR61gYndPAaeztP1ws7FWWoSeHjZEflhz2IkLXGX8TLr+nC2bXJUYKlVdpuNLf+
KqSTet4qswIg1/k+PsstEnitvLBqtsJvkXsIeH217BUwiJ3Hvh3U8H8OYu5lgpfKMfkdxCnR5jrW
KJCuRWvkR/NHqSaDjmJn34FcQQevTuqaEDpXoopkzO0bJFwgRE3RQNJEMo4LEZJDYLpNjqVO6Dbb
hj26+h4avnXtYR2xapDBaCUzt/s2jh2HldX4+Txbu8Gx9ZMmGLbF9ggsXlq4H4qTPwosHBiFvlFB
LF61KfMDmo5uJVFbvYmumZi6ddfPU0XQR6kt8cK+QnZupm0rKuBAIdKXuvAdiRdIehrdjbyIcq95
HN4RaBfnBgmqIKFFKp35GIt7Ids1bGb0X4JbaR+/vgPA0raMZHk8w2a6auHW98rjiHYQ9qzpg/cl
ZLnkW401A7kcBAhIL3JpDnr1kIysaaZAB96uqkFjCEtdwWfXJ+XL5O8CyoUAe/Q93dSLpEgpujij
yqKz5HoDQLUsILAheF1Xiy+x71Zcw5dkc0RU5YUBsxb57MztHrv85JILqEEwye+i2VdDn1sBqjJL
qPfhWSVqx15EvlqEGXefCgn9/mz7tCBUkqbU+Dg68Y1gs6KrhKIVcfTlpGjhNm8Ajq5OuOdo8lN1
4fu82uaS8bZy/ydSogBklcG4iMaP9gf/rSzWvFJCAZgH8uAYGYQx+Fp+bVr6TQ/q/K8qiaUDNYkk
J20VyunKuVFM+kXbsIzI0HuafiR2FFSkqgPJEKrPai9TOG8xmxVkxpoGNnkRX+1IgtnuriGrSB9q
1oLnXTlP9zDJ3pKiqiVOYlp0ZVB70gQJnsvFWyBHryCamS5vp7PhjhjMuJb9f9v0pfTIx83WXCbh
uCI1rHaI3MdOEgplwp/7CL9gIQ8cgRxJpj7tBLy3lqY1H5Ssmkhq6sPe1i0zxxdjOu2YYnkS8eB+
Mm5buY3mw84GHDReP3DkgNvAPbfQ5bf3A18/RcV50mkFM4g9pNC+Tw1Mmde9oH1LfMWDAOhOjGji
tf2dWiq/dLVes6kyAoXbvK5h+2ZTVZojIFWyiQsoPyJiXQj83GM/NcRL+mzy9Vua/PRNToNFGeFK
JePjaBUn/CQWspomiHZJret9s06n/gb3cqX2c5SGqXRCT7DJkrqDlztumLTh63jG4iHjZ4EBsdol
SBXFB1QAu8iCAArCESRmvxP0xjBdiH/FjuX6IKMpyV5JExEDtqVVzzKSZFmK7Fuhd4DtUGsPSwKF
PdZI7fsN2o+WXK5YpajTWgNBF1FW7hVZLmL6PWYtTrmrPpy7bJ0gHa6XNfyZgp5k6HzTbUQ/edFL
Lk6Wo6NIjSjtE5VoIX0TtjQZ+IVYmNl19ovBl6i8W1gfuEW0aqYYzCx+vxTlDq5olzl3YE3+w3Lj
fOV/vPpzhkC7AB3y3CkemkRnfxl+GiDDtZmTgxNOMpwcy7yfKgIYmLKBf5aUvqQFZPUNmtP6NM4q
CQSZRpgsb8fhZZDglj1kAi0ZaPlyoLayfivm6goNM4aflC/OviVi6exLlm+8iQQ7qCy9gouamOg1
tC/zb31U4C6yDvoJBkI5gkYdeCm+xTimbbkS4IthflSyY0QUzy2/jPM1NNS6v85DoCZaVALuiMW9
Byzy6cQCgQadPXLL4zwRoE58owDUyR67E4eCfvLlI2P3/f/aepg0L1ZHYHSejB1JUi2HFsiWYVzn
eE18Y9fmeifQffm6Mzdgs17/4SUtLZvy2VvRXsKstZV6a/5N0ldjsV5i4bRf7GWZ2SzxbSihOIhA
hCi902KsKEEYK4pBEKeHn5y2emDsOwheg1E958fHc35lgC0nEYMGl6nAV/b3ywWdO52J4YsxHf7b
gR0drWCi0ZtynF6FP1gkUd8NM5oKIffSpsacMtkiR/WUrUMSRr7oeqBGd1lI1CacJ7B6SUTmeSV7
9qd3ly8BVrHx7vFjWWmX49MZS10gB8o6TpSZ5n20+pC6IdlEp73pn60WiaMAcpXH/AJwqPieWhKN
8lKnWAViS3wlSA48FEBtR1naIQhETqkTlF7NVTe7Pa9uoa1QdFcS0k2CVwQSn+uAiKUJjSAQO5lq
uBXRyc+n2s6/iPa3f/Xmdx/BOPYa3G3xUKcKqdLwjxbC4dhSXv+8dvhvE1IaIIRkb8kMjBfvRMPV
6pgDRbkE+pKG7HrfKBKeV8isXEzM6xhaiFMioeLnHnc/O+2YP/BSyVTrHmNhCly+mCRb4Atu0a4j
AMOuYzg/xjzJHI5P9JI6ArQPrDREb9WwrPmnJP+TQWIYlvETsfdyrMCGvpIfYRuDecdQRo71KMfV
7L2MoofJb4u9rqVv+m+C12vLcgkCA9s5s1PnR7WQGuTUn0y15BNozwVeMDKnpryRzQx7q6AAezBE
LODO8b4Qv0jiWjrvxr6LzbYn0xAKrByhlZMxc6SfKYVxAJmHO2tT+AistnUHVOSFNxF+JOGPp38C
kCegvCjWWDO4KxdyPtJBB+j2RKxU8OsOYfPEB8j3Syudwljf6NNgMq/KAUGli3UtHIfsxZnfQEv+
Bxi3UOSA+V7KdV6PzQ2yeo8zieKdk5Vvj0VyRq6Bt5Z40Gxf9HUSUDV26QRcsWDCmSnx6YLUIG1B
rpZ+FuTO+efj4ZPdEVUMKY1COWMQiMza09nptdKmKQLcrZbQBd9RR1vgvH+NbDkyFOftZECCxIDK
M0rx0M3XjFxVdxb+XZ0hu3vYcEZXoWOqEqz7++rZ37R25UCCAToFE0cKqZXMAQRYDpwYJVXP+NIl
phehu2WsaHcXRiUdxjoa3NnZQZhHedP8xaPheh3GojGk/N+sFGVNq0UseA8NwGMnAijYlKCJUEyK
S/SnRijvu9jHB+9vKvYO38xzqkv+S4gSHFPgh4JivuCPNgyxWlhU5VjuubPB/FePVcLRkvxb0vDl
sVryLVo/skLJsxjSWBYTdnzepKe/FYclaT63DOFwewb7Xso9my1k9PD5PvIUo7fThULb9yZQyegh
rlIwprP3tS9aScSxSKDa7lk6cutyfn6wbui1+DA6r+NFOcCA5m65zMB7Zi2NBLdVP3hAk24lkdj6
KjISqEjo7a2CH17cAtcXlcrIBPlkQnCq77LY3ibU6TmVsu74y8g7DZfSPtPSI35WPmvFUzdz/tKo
wqO8tqPFfwV//L5TRbVMqsGCKlxyJIjU1qMD+eS1Nyy6fCs8JJkHmq8fX5pBWGbqdLsa3g17di1m
HqczOlUOTStBdiaH4kh1QDBfX1e8Af4uqMeic9YSy/1wcNO0OLzVM3rkAMnoPtezrKvj5cVuO2Pq
Sr7GcIL8EisBvdSk+SJL+oJfQ89jpXzLGpvARCkl6B73jWCxVjB5uLhH2vu5gfuv9PKWinKP8jIY
fAEK9O6dlCpMSpNZOjOH/G/yVAvUM1iSfXd8Q/TLX+Dr0L5ZtHZM2Sdkpv7svQwCW1PGTBuFlpc4
5/A1tVH4euXiDnG40e9DV7Rbaxi99XBgmazI8xT38IiebZEi78FtHERb7x7Hrrl6VRfBimn8vizc
xhNUmeAtAUPUMVvQSPRDLREC7AZyTWLKHRa9RxYY7lHKssXm7woLRyhTJAyPFfdCPbs4k+Ec9xPF
nO0JsPk2/+cPQqrAaWGeYiAoDbWylW/OwxGiEduBccbCeUqT6/d8HfsVNPNfIiyN3g9ms034f7M4
vrG5J/6OrSKARGsjd+lF0oI5UHWAGjOY/HC5irzEiDeZm1e/36jb9RNWg0VeZ86Au+WaosZ6uiFg
idClQ0n1hEYaVgVvaDJCy9g3y5ZvW/ZyQM71d25Ny+I67KyrjRvf4x7aUodJwI0HmxM3OQ5mcfD/
gH6lYdRqPXdYWAB1lDohBbqZn0+8S7oflRRoxYZoGovZ5tyaU4f0yaj+Z2AVIqKgIQf4klypwrIT
46Pimvmm332OhgJwTEYtv2f3p2Iz6O7nrmX+v23TrrwZrn+LXud5/Oop7RrxSP99SIJyMQ997JpB
tGxxIyyZkgBBP9zuHsQofX1OdF8U9B06gUE1qh0uzO8P/+M2GN5wi0h8kzikqIMO+WIhH+FotMhA
1C43oTzNuRL10Dtiahp87O2AA+T1RLfp9Ap9opEjuxlWDxZBferVZErq4IaZdHKP9Yd7qDQ2xW5b
PA3u2Iz6XK6OXRV4ybtsTdRTslcwnjpsnM/Rd00t7XbgeCgR9ReQR+BHHJTT9q6/wplDwdLlseBX
PouxUq5pEHOSB9fe3XzD6ux0MSw+ETkZtM04QjihBIFCGHQHikuoz2NCxZdxAh3tZz8rQl6jTHTA
+7uYr3ej79KYgmggD/luDhrAHt7g5gLP7ZWgFWSmlQJEhgQxFiyxzQoYId8xMBQomrNsk2xIlDzB
avS56ZyVHlLBntAYqORimb90iqm9ddZ6YAj4RadhuRQnHAouBidpKJPb/Sx169i3+dsP+PsPO+9E
ptoMTIjGvIEHsHDnB2d27o9K8O0ZO+9MszrAol9Sa34MQuyROAFQNEmaQttG6UjVaEIVFaunNn5K
kR62dSx/EbZq9uluTPY3rAuj2t7e8srRfVQ0X2f5ezDZM4wYWbAdqGvrg3vtObjfgGvnaspjhyxX
EPc0JSCuDyHd49dmmjc7ESo8OAkSnysvJvLDI8VR/eWRWZS2OExbqSSZTurZdagZfJtWIIv6Vfdi
sG/rgWgpri8f0QJPQRkX1VTcjufD8hhZJ5EbWOErPPSQMKEb1WT5fwbx8hHEnyfglHMGLbcL8BAV
VpmypgNIkAEY6jCx+uPx11o3b7JKCQ/t/B5DnmqJygGs5gV2FoJ8WwwwFYVk479OyGmXaMBMUqP7
egn14mh7waxZqDlSUOs52YsozYcnS2y5HtXBjZ5QhLWAi98OFMig5vt5CRviS0HMafEQXqhLoRvb
H2ObERs3NUp0dWD7bcOi+9Wfd6wUpuu3ho3zY7fuGnud9pfclb9Qlk2ZiMT+fKEDuil5JkVUr0AW
oItUVFXOLIqBUb20QlYsYU/WJPOyJibnh6G4viS0mM2/Cn+igV5sx3yo8Ishq7XJNa8mWb8QamGF
gP6GojQqFH6UM2kOTaszRdNo/wf/gOj9w1NrlHHML5hCCocvCawn5zkkf4nvcJAaxz6ouOvAclYr
aCL/T0SLzOPIN0qlJurO53lwwrcR3vtSZCkM1TjIsG2foj0c2SvilVfSw3y6ZAIkiD0RJDsOfvLb
tSl2rCgRbkcEd8MpzmkLmdNmdoZj2Xh4EMb2l7tkk7JAn2US3zI+WWbnFyAbyEU3sMXTNs0bX65U
LQmJ2GCeLgDxTW7vI1vq241/K1+c/wNwuf/lEWifASR5rOMK7gvCI4SeYSHxCp9SfqEjD4JZXlHN
2M2uzH2GrgDJYh+Xd9w/0eTGKXXg4bZzgTIHNafs3xC2ZJMrHRM7ggZ1nkg48Qa6yYlY24INssoA
no6df/g/5GhQ+fe4hlR+LDHzxdXiqSUjmY3g0/wNMA3wqHwY0M8WwKe6ahY5yMyNxscnvR2BI1QZ
JuHmrDcb1zj4NBNyG2ViDjbL01awwvKbuBN4I3awfvpZZwv60wE3inqaqlAxyt2rExhmkciB9MjC
uLivB0/ZrL0mzfdg8Pp5jfxy5hDg2PKwdfjqN0mpMq+4wZxjuLhEv4Pm11pcsVnheVinTOy6/l6+
TNeTxEajIWvR8Rx7TC3Dd9LqXQx3ziI2fBj9BqlabzhxmWHl94/nx53QlC3gXrpV/07BAKxjUCtj
aardmdv/fFHh4fdDi+W5/lQ/AKalRVdJolNz7OMt31trwDP0oTN4EhbUmrlSdn32YuWGGst6RRez
BLC9QEKz89oM5Gpe2sXy88khA1hsQU7LfgA0rU4PJoa6qbEgUJ/AsbRjK+t3iSbkoUxeB0PLOxUx
DiO4kOAWQRcjPa1+UqlQmlZpFEPdjiDDg/2XO0HPEc6qEvwT8P9L+on1GgsKkG3MfmZIGcZyThii
Ult+kE7L0W8c8WQFsPsWwPn8ZPk02FjA9lf9Nnif1sqyQTT58n5I1BqoHWnpkvFY5H+QRK6++9Cw
o6bUDLJZYeYpcsCrT5ZoZmbPPy8KUZG5BG1aT0+TB7eRHH9T18eizY66vbmxj2/8xypVhw7kCJcc
EgvqRcTBWKy84Xonojt//wtBHsFE7N+9/fEO3zMNfv7mr/XEcGVt4s1DTlO7fQrvDHmqfy6pP7wY
tEs8QDv9qDLm/KG8tDUAttUU1TJA1BvS0Qzs0eZT36jVpHAoJ6/UuITFhwmnqHvObnHsELhw/o7T
XXpUNFXj2dxi/DM5mr3RmmoF7xydY9EO/4xEWbTg1ersHJNHVGEQGMRSImRbp8ipXHjXGRBXQ2m5
dEk0+vX2zrq2ocI53e+jBEKc8b8pdO19qlIYqds0jSjKSfnKNTlBk8jftVCRIcnmfR1jrN5afUQQ
LjHgD0WgpfGTyldYSp3KzYjC6vVtCxbyrSNnUzMUvryZUT11QR/m1ueQZ3nY17UJuN7Qch7jOOwx
p7gLZbccsH3V1hjMfg3WE9b9HZi798iph9kEuPsy3BCTsm8WIg24YAishHCQLgir6bMrnbotb0wx
pRqdOIg/I6Ka8U6WlMQl1pK0QIZx6CovaVMhjPN65oaYnUNMxUYT8APfaPzyWYyDGIINQMR16vv8
TIE2cMyyzs4hs/uoJ3hFKh7rmfg7JjRpBZtwb3rQ7bZxMbxUKh4A8ap65DvL+pbI+L7pRpnsOyyc
B8mCLcloTutoksVnobDDyBJjRcnwLBAwJklP5V8beQjURZ4iSx6hy8fDCGxHN6dk4sPDuMvliYBR
jHkJVAMMUZTUf0wYJyvTVD9+01QeHtkBVLo9SEPb3y7nsFy0sr6SZAbHxCT01oSuTZXj8aTo/Ldm
gxzfjcRXScBb8lMxQTCWRLc4fU7MixGCYEERzjiDwCbBJgc4KTTIriYDFMOof9IoZSCGnZkVWmd1
bVp7e1N7nkrsVsAm0PBjn4FgUGyeVBy1z5SpU3cBWB32NZlGr5T/KpgLN+85G9ArT4qOzLb8f5n+
NFzeaE72YbG+fzvCH95gLg7drJ8IvLCbMPTEX2ANGzULqiOynd/JuMbpbgBkL5/qOPYs43JhMQle
QaiR5h69/Hby1bivxFvVgIciYnENezWMrpDb8Dl2FJsg10DQRb2V44dnJCUifbBafebTfp0xT+Eq
4tSV+OYT2ymTiv10Z+mp0BGUcEW8RhA0w3IBCHqumqc/bBShlBIIXK5F+3hZoLhbfemZ60XzdAgP
LrVsrgMi0tdDTVP2zJlybwL7w4UlPoQRwA1jZ6fQHd94WFyBKaV4ItUccl7cNVcTibg8v2eX8AiS
YpEYHVBH1cOrd+iM0ZqNOQOsQSIgMxCZ9PX6Gx/d47JQnmGv5MDazHTPSaPLphnmppaT5SE0GCbq
daTvDBacOw2PRv2ZQpgylP98a8tJx8DqnVIWP95KP029xICHMHRTneNg3UjnXxzcebdBTqL46d8T
60d/seY6mnbHMnGuPiZzeO0nege9CWkrK3YvEzE4qahuWwwDPS2NS+N5YN/ajNbuUIE78XsiGD6L
iO8curToLFvSwhtjzb4terUJIC6oXc3NzJ07ua7HBzVhp/FzsQpWXgROwkev7w9rR8KecohXI3r1
aGQKil+7GKbk8bWxxA621kkCCllAgAmRa9ZWLIXP7RgJHT4E4YTDd19ZdLIcNW98t7IVOsiWU1bq
TDAeeGjjA/04r+W3o1wn7KeuK7cQFerd0jD45enAXvFCQzTwE76UpDHG4x85dU0kCVNO/oDWooq9
Qe2iTc6S0TIPT8Tqj7P7taBZGYK7al1X23ZtMXW58gFYqxEqKCStG7hAFJ4wGoKW63UCl7DlHY9D
2NwJ+PlWrpou+6ChEGXiB2pIXeIA5erTaOQEQuCmOVPIX4f+G0PXsKP6ifrLMnxcBTqixasMryA5
PGXftONwrFkb+tGRjbCUL615bSiayLX2AyqB6XsTaT9GiCjbcEA/hw4rAenuNgTDzgD9zqOB3bR5
6tWqNq7KrxjywF++vKZrwmxaF0hZcDdI8wJRU4PHNtUnBKMhAujbMrAEBJ2iG8V/7+dgp7XqBt2w
NaC93daBQz4EXdfMXzdC9PjhWO1pabjdvg+OpHFzJwsZmZTPsvIEAX/TXwLkh9UjY5i++abpfr8W
n00KgqO9/m1SYjw8zSzNbaSvnuEdMU1g4MePs57OzmyZfwrkXCRmr47Bc+IYd82SpWGKvJiku0NN
mkWp5CVrd+hD1UWHnCaZCoelzwFQ+wZ/y/+E8q7FCIFKtwk3YizONw8mZdfyEPAMKD6GrDnDZXDK
igVtSBPCxPis4gvPmvbM4Fh6E7/NSpqochQcohpTUFXQA4B/eTFeuRekN+1NqvFw0QaS+vn6Qblv
EGYdG0Cf4Hi0oQj4gt7nMcngjXCVjoj1FJYZaaTSH77kLcoTrbZ9rxbh2ULXSg0G3z5Sis/523ym
+SQVRhGhKcvbbRd5ZLvoJLYjMaWsya4RKggeLPozXzwCnNsBqmejzv/s91tEXE/RGlaJQJ/JtifL
iDavu1JuaqaQGZoPpAQn1DsrQtmsxlZTpP1bEXdHgv7UpfeunnBCi2TvFYuC2qDAoVZBNt3CHa0R
VDXA8k6B4OmH+Gak+A8r1Q9HdM9LJkWnFKXfKgRHWhqDffCqQlZp7CM+xWaOHh1+oZp2oVVFKy40
h02X7tXeBOUzhjns4h+OT5pMdpfxmcltTCqMt32Ig7iePos0/BASijmaayvAaD78jAMxB4qndPd8
b9LVWPC4VzPNd7n2Is7Xl3jLYGySpEBiskV4TalekoYS3psWhDYGobJvhWj+FS0bBkC/cjzKOPyM
hnbmseCteJdpIXstGv70xb+8QtRwJX5ZR6aFeTM3PE1dda3QwjCzPPzO+obz5zxxKXJW9h1LCZaS
BUPJQc7vzlwh45xA2TDqI6VzIdgq4N7046m8wNEAbx9krTl96rS1KByL/tFvhgX3d886je6tJhQx
lMtnLYshffN+sUfialCCv+/QzhInwALf9xybhnSsXa44+DoS71k51MwybLR3IkBFF9oeB9jbYUkX
jDtBKQGRJmKhC+QQd+9MTyGLGD7p8Z0Vcy1oynL1ufYjOxfF65Nam4eT6wSJe/g8BJpWmlQGIiQv
EkS3rC7hRpU2D8H5EjPuExyTKvPQHBFOTWKlqg6xX1E2ZM7prSl2B79plAJkXbBMR2sirPiGqukq
oPICORcpOIg2eL+O4eC8hfKe1TE7kQ3/eQbbUl19660YIin+OzARthpeA2vNpE9Y+nvanLJfT8ai
VjPHvK3aVluNNQ1DQu6r2XQWCszltB2yPdVt8EJysiQLPl41cRoBQ8ojX2kGEBKWF6v3wbTaq4M7
PCPOKKhYSbdDryxUgna1imQKJNLB4bsdx8pcBS/Z94Wd1/WsTV01kZpoB4OL9ZhpPnf9cTcjVYDD
1Q5IPLJAOn9EufPe9FAhTPe6lvkKTPtgT/d2zSQQrPhUmOsGv7DkfSGau7sF4Q3E3p5s1saJGZ6G
m8V8xMKUhy7mvF30rP/0x9FwRL0EGf4VMHpc8YMmLa+XKRwKuZ1q3B0bAVmj6xg+rVlmqfY1R7CA
W3jXfccS+dS6Z0OEMjLpx591kYoTeXzJ+98YmOhOvaptfb4rVF+9iLAaVsTVefF/9/ozVPiN3bYI
AN1lH0JjssGV0onh2zkkTFzceKc3Y9ZWOF4WUEWjLNdGuUjyhqi66fNxnmuHUPC1unubdnl3dZBx
u1k7SgBVvhEpLznGjwaoJ36GntWQh1LUoy6PaDdqGrWoqyF981f+NKf4VPLfAYUBUzyK0NQ4DqRQ
XOkDyGkmPlD4B2vEBZPtnYIFa6FTuDriAaW166SprXAstnSYJ3sZECNmNcUa46TOXca/NKADXhYw
YOClT5LRkC1w9De+j7H0raYcU+fg6b1eRV+kYSt1j2o58PrL/0NtnXYLfI+A5DtL/cjBKak0051w
sRBYmdIKgu4KbzuLWE/DfpQrDlCrKyqF5EmsY8MGYfRGFjCH73Ijamhgk79mIOa0T3m28a/ToKXg
J4MeJiEMbW2mqmlualT8lnbSeWAY/+9ULwFq8+PNMNMcS+KjlbHlqHQG4VfhF4Mh1Ml6F1V0QZcP
15b8qKIx1NdcjxV49YnWpWo5QLBmK+BjyLMBPi6IEMPXrX0yriYqshUxgO4I5N1Y1rfI0r9W2jt0
sR1JF3xSzPVibR/K2dvBYp6fbKZiq0mdbzR4ewbqNscyUBjguRYAolZk1mDuhkDPwihWmh6E49ES
LrGHn5Q/zlODo5e1wzeOVQS0bE06N8F6qiHG4XiZWbsuzL7WV4nKEWjqtvXFEvhr0F4B2y1f/rTg
pzGFVfGg7CkFJcDNUgvxUXDqssyVwDVVgFaPvLxlDV39YPIftCi42HhfgPqJZSWdL2BC+25Ocmxe
zNv3VXvo+tkVPQRxGMuRnJ2xbXFeogm+ow+dLDfKRuI+1cjtMy3DfAv7d1z86DAapoA0e5AVJll1
jDvpcKqCHldytpPV3mWwdrgboYOFsHlQj6NVpbVDMwf6CWDOBo5LwTux7164xR9jSpUThM3Ajkpr
w05KnUJczWuDR3ExI+mjP/8yM3et/kXk/FDmHKIG179PVF6LBelG+49HoK4Tn6MUjbsRhxwxFvyj
bDfxP3P9qmchkd6hZeyVZHjBaw8LYFX23x6DaeJ5kRt8R3CSN0y1yKa/gox5qA3OMHjuGr78g//m
JX6hs4vyOivB5RLSLOO5uGBTzY/YgHe+MQkJ/E1p5Rikhou7Mxd1s+ligs5SLrm2Vos4I7Pnr+Lg
AMLF2mv6uwV2yigws1+/yCyqQNcJaZmai8Z1NvSTLZnXtYWCfBJ/7Nkk1+hcROeVEgjsRTTUN+Ac
Dz72kv+wVrj9BdoMK8EpM3Og8PMfL/maP1CXzEibtfdQLsubaluNKlIxKBxXs7jeaeRwKYklL+i2
YvAYe6HF27hdmWwnA8HhWhj+Bb6apGb7Lc3DBorXI0T7II9eiDVJqJdtSaV3jDwHx9DgKnRtfOqy
WazFG4AJp1uj8fZI4aXV4ed6P0xsrSeFfoGct2kgIwJEp1ldXxM7I73Mm4QXU4TplK7X95x/YG9G
iW53qAPItkSMbNbdQfnDzI4B2TYDLCJISaoK3wKLJYPb5ckPLoJ8/Qm9fVvX6+5H3yCf86cLzYmw
7b7Ux6ARCbe5pdtavXs5x0WAi+f8nezPmZTngz9HUv48wkA+AOnXceux5Lnsbhf/7pCU8nuT/0kJ
856Tu1vU/0kBJhb+fPLMYKxyskQ/4u6orcJ885zaTIGoU58Z/103hVm+y6rxWdUGVJVnnU8cKkD0
2UWuqgbbIdyCkpIIe2cr9dveC05zmZ2jbzKXpehRyG1Jytk62xjBjLgSdTO7QoHX+5Xmgid+OWpS
RFkhOFv75n73DJ7m4TeRuAa/ldx2jQ02WDgEIGvUqu7xu2NG75hEU3GehKYOKs5SwZm2LqYARFjq
7pB1I9V8hGAOt1mFhF6B6pkfPiT3IA9KD7wNDdg4+NVPDGUGCVgVN4b17qNTO8bYgYiu/CslbxFT
vRmXSBuOStbxhTnEF5PBdk//uRnczPuauTr8bB4uNdkGCG1SDvWSzGF1zAiSoBFtdKhslg0z7dOS
qjxT62NXi1l9xViq/vNuaE4e094GzsAKdouZ6FSyC4G/hL3NQ5+o3u2FwT1KnHbamASObnCBmpEe
coq8bBDSM0WcO7H7izU3Lh48dYwuYvputTOeI7ny1YlAgYMz8yW8X2HXzdS3XotfxxnLt1k8rCMQ
c/njwCnKOmPNB2KdwYRH1mS8VD8vRKiHefiqNkXATKu6OU+WncjcwZkuJvrY82ySI6vs6c5c0nH0
s3pmELk/IyxtTyvV9YUNr4dYUf8Nqyz8qPqWmkud/rPO5skSEj6NVJdni5wJ1LbbGatk19aIJgXK
YsxYEAUBumFJguK/SI+yzUU8LKRHJdANusRVW1mLCwBPfAi1qbAe4crE4BLZwyPRZIK3FzfdBpZq
eRqmDnpnlnUoPlwVhgmkuT9XEnTJoF+TLO2mq/XzsPaI4eTb+CQwwv3qF4xztkR2Cpt/ZfqAB3cJ
mIxZ1/mNKn5Qzvpp6Q669ah8LzCjiP3tgLAVk/xdtneWvDzWTgZOjQcmifxrmFP5EIGwXhc5a1R1
PtWbFhlUf9mdPxbTLNK1ESdIuv/F0QIY6EKD+0vIXYg1Dr7GEKRm6BuYUPgHnMd9NtktMnIEgmXL
OK7ewUm8DRHrlIRuYcccPdnuAaRwqVvPcTCTamIQ/TPCc6GyCtiG+91p3yEEnI5iVh+qesM6VkcC
J/ZMn5auUGNTglSGSCKGXE58NIgHavoJwzoNSpCsK7PJnEtKRK43QVfrqYrJAhxwWFNqxHEbPDMO
HP/NWgWGDQKhu2gCZEf+iOwGszAQHfHBHo0uNZrLmez5Z48XxivyWWvGOcoGmVfVNE13dovkzVfJ
s6Y5PLbQX97XXHp7jrJqwg1Kg7udBEDdHwDhEI2s8KSI4BU1sDnoSMZiSmPAohlv9x/Qdnsed0R0
R8oL7hivimQPIdk23AJGuu8Wie1fpfst9MNOWJ3ChoQ/Gw2eJ53mMCEF9LagCWUNnxbZ0ivz+avr
TJ+plfFv48f+KYa7MTfpsxZ7NNwcQ9bEETcq+iku6EXLfXsEt5XZToYFoK875MuDfBjmtZfNyAwQ
iTmN7tch/uUZOYkpjFACbF+R4aITq1jBhFgZJvGkwlE/Y8DsfszNZCsgjzA+lTQ/Fs0bJeVczhRG
NVxoE7I1jnjMIVm0vn7mUjGm7Z9hCrNuIWwrA2bamTtGyC8N/7Fi9qq1MaBUY0nlP54T7rqOesoI
nxETotAgxxsvl6cm3NfozVMXTA+7xI5jYbs1UEyEXl0U24SsoQED10bDtcPY35FKvojCorvlJF8N
EyIgSBAGVPC0CAX9Pvk23AUBZSiHf6W2QZVps7SR6fsmJY7kiO2NJ2p9t5Gy7++DvN2MkotOXF/B
bADES6e1ZT/TBh7a/qAh34zgHQysBFTr3mUzZ6UdaH7y+6ZfrF+DlecmicSSb0lv6E/ztvJBzbqs
BUcgJpJxmbr2Q9Jsj5H+YnDAav6Rw93zuiz+oTPF/qBxTR9HfMLCVnxSrulI4agTi3sVJ4cJ2jXJ
jWO/oB3AbvgQCDI3frCLz0Phpe+JElENdJeU8dE1hx215K9Vyl0IJ2ky2aFJd838CxTQGbpLQR/K
D7wNa0/Vj/3MpSUPUxqr1k1jPVBeHtRAXe4YE89km5ASrz1tLBTBIBWtQ+QmAwM2JScltesZQDf+
3s5uHJcFs7Md8pXZeOTdw2r6Qrq4BzxkhhCkTi47ke3sWngpxeI7UT3o/jqt14XhrBHr8iyBF0BZ
id9X99ETrlFak53IKtoayZR+N2ZqlIest+shIuwhZeZO7kbiA28wKUkKv82gTkt66Kr/oVcsu0mf
3vgT6vi0EDweom1FcUMjHZ58ziR4g9yEpzq4S7LA45duX2D+zZaMlV/EXjy/FtuXl8CUqubaScO7
JKBESYD1vuoYUfblB7+sMxhm3yUBVDnEitLKPiaMAGjTn1Tex7QzyRX4MccmZJq0DbIy1r9fvqkO
g7ixcBPv2us/HcE5KJnLOYMpFPgYWtXmCHiEDMt4oea4if88775y4Qv+DnR7inOXXpiVa84MFB3P
tC/edicIergNFLe0ikg9Oz5Tpf4MoEHRij0tqjjVW1MfQ2qef0KLST0HLHRv0Fsku+jlyxUXIwP8
H3PY9/hvmAr66OgutFr+LoHinDnzj2wO/NCjnSyfpUAyDzTgNTBLoJbfX62KFAKDi2zPizw4wLNy
wmFXpLbrNMGiZ4NGmo69am/UkI9Wi7nOyQBRWMO4IeU15ORMiD/WWXfcDrIJbZUY0PfFpe/e+VZ5
Lj4Wr/TwNkqOU6GUxeLVvN5V2qdTOEIYnnW1aOJJJqlTPVgktosWcCygDGMUyOPF8ew5lADMXjKL
KghC5uL95VdJF7DPDqTmv26Du1Y6RGyqHOmVVuGO5zhGwnQZluV5g9W4HBACsPmxPnNIK8EjUCWv
9FEkAoQmF+TJkRxzKMzevt/pFq3gaoeQBTTXBanZfAUYlcAYx3s2TLyRBGcLOrAC/5HmTA/dnopp
KHOCikDYilEq9Wpi1c4R7MjYa3wP8df7zwfAYntTRhpqhZMiqcAhivNkFegSvVk7KfGX5CnkSgmY
+OcmyRvrKrJRHGG4aCznZvTCDbqYH/VCExyboq80KF0in0P5/uGfO++5YuzbzDqOPKQw4K0NEck+
fNc+mqtfiFb7Nb/cjYcFHVA6dGkEx3m+3TT9zPR6ZWIBCYze2WnZVJbs2DNwB9PdK+0nu7A8fqCc
lbeVMBqO8u8ZqDULGVWJ3sEaDEbfs93lLIz2Ig7pjqHFaovl2LoIUF7g5w02fe03o0JMWDYm5bdG
Kt5bS7UOhFeN4X0WOIJfTwm8bRizBpI2cq7aHXukqArYdHqjnwvRa0SIXIWRBUhwF7esMyjoYez7
e1W5FOx9+GXYBY1Wx2IHA7mX937c7a55qHves7Jy92wi00GuyYbXfrx2J6C6HW4G7l4rmS7ATUpm
fJCZVqyBwMMMcM10T+sTaAMKvSI5Mxh5VUfhwD0bea5WrqYrGypussB0/4CuFWcxxb31myAcVj+3
qGGIHXPdxvfHTa4CKBXQh47oMUc+Ef16E+pjNF8orACZILdI5REe9ZltIq+3pQfDZ7VYZvS8I1Qy
n+Nmt93BBzJoehKYHYkTjiyqxwKvYgsfbVH6GgrdcNcSpt/UimXDHFjoDiO4uSp8SZ000dnMBV1d
sAmaB/l6DxfxlvhDjbNeeHbl/uR4PgJ9o0T/Osdj5argfujYb9lkLyZ6wZRivXevInCIwRgIb/GP
ba0mh+rfE/cYNSeIs5zt6WS+vGwrqXkwFkVpu0KoWE1dSIVfLU5XfVs+0XnowhafmtIntmS/zM9M
M2tQNPNqpiI4yZYVtVWl14vpR7r37485Jg7xlN+9bi76WPZaTIv4bF2r4xiDQQNvIY+kUF3Hcfmw
/37mcp33TJ3FVS1U1tcM2E1pZCB9kIN4VwWKeiSdbp51FvmNfRN0aFYJ5NKiSRLYFSEk7JD79G6S
zwGKugd5nCjF6cYQsk+sl2leHV7Ty5IpECg2upkvuM08td8Hq3Su1UFjBDOzHYhDlu0Ad/no7EI7
LRJUXsksxoc8kaYmEsSWiiLiFrHM+T21kbvcHh9LWwZonWs0F+o9tOHkmf5R1MzlzwgY6jCK0vAH
af4eNrw/cmSTJIC7WDYASX5vzsL2VfAd9LoTfV9NCTn62do6g6A00/ZzIa9fYvSDyeBu2QbVHqxC
DoGzFCIyhIEHZRcEGC5pdERODGvq2sv3T/XnnMYJVNYur/9GQWHjOWg7gpNt0Kw6wKyjuk6zH5SR
3KL71ZZ4Ajk3cRQOV4s9NxZRxe/9Rs7GF5Db6MlhMJTX9kjL3yH2klNZJh2dda0Iumb6tVo2D9Gh
mHqCRq62hnB0lmIAqGcrzLsOm+x4FkA55xrxhVhjx9PE3lczPaFbCOE0O1Bchazpr/jCMiKQRJHJ
O92dqgQe+OyOD8hJea3xu8b1hXglqN5B0s5ZBbDDGAGrz8NQUFAviXNvz6Fkl3ei81wDLT+3myPX
To+jqvliJn0xUKWrhL64ha6pySz+1yY7IP+rsVqPzYGWlpaCBvGkX/S+SNOpA6eiXTXbEOToW9hZ
RCnQLFXyHlpNLAeEphI3nqV4wuOLeRYa00tu0iuK/vpfrqPjrDy2WG2zcaxYrJ3okSPxPCdlIsw/
uqHKDugNV5kD8DYmiVepAVJfGMKcPdao3LHZgSzHMhu1p7yIvPcoOXiIJ7ZW+h2DEn8wwacUBiUM
esjZHgi7DOJixZTKTLUjlowzUe9GvME6nqccroYX3z1pEG58+mH4hkW0PJxtlyGhrwe9HLc+48gB
3ujuFrIsEuDK9j5JfFY/SF6l2gcEAifrJ6/KlMCBs7r/6xIDGT2BF8L2wsOTKHOCAIDBjrBLX3i7
MKNXHuSHrmIzCvKvQgzEOQy8GmF7hRTZcaJ1ijeMNuKC8TZjXUWYNIkcqrl3i1KGL/gHjO39vA1o
KF8K2u5Q5IMknUswdjY2vdAErTd06pRQEW5oMhSOWY8w4CAAwmKRjoCqPJ4A6KRtFiC21yN0e4kR
4E0cmYM8zyX8Rfq4pJTW5Sf98CtNww7YyyIodk4vxIPYA/XUND9sQ/AAFu7IOqrL6WPAgLmiQDyu
Giia5o/BqZs301W7ASWlR6oZ03vBgSydVWQzZ6Zq15LQfTZktgtHq2YcY415XCHKza909rtFa0qt
dSDZ6TCrfDamDhh4tJpEsNvwqnCBJlkyK6iew5MgsiSWbAxcWR15gAaWV6B2LV/7/P4fxDGaUz5z
rOifnr3+l30Z1xHjCATqKx4VcO5zvqxHgXECJVS1ERLczqE9+kJkwNF/kEGXOps3ebHkC0Q6y/Lh
crMwhUNZgIn2tKgBjFjOPRAr5FIhESMl1KOuul+XME3HylY+fK6bimaPwX3gd9L5JVwvHLZRlEb6
upeIKGeby9xhVLGPHLLZD7fAucnRvcBMJmNSLjAeFx9M9bujODOR1361Lv0CwEq9H/22vEvw1asM
BhrOfshBxw6RPt9jF3ZXJbqSWIq2eTWV7DSEKNOVaYKlXE0fTdkGcXNGTI0zlbdoDVuosDR0pplh
dAiKVtc1gZfvugbBeMBlrwaLG889Bw9GwBulIedF2SnUuByBzeuN5qsqv6sd2deq/rCW0sadqEmo
jRKu5v9HeWYOTIjGPqRry3HTkL3f7xIPdX0arovZ0L/yyvmjHQPaVAaLQt90O8vvGYNbKNzH9Ns6
UKOXndN+SgPB278iMcdEnG38d+EtSTfBUEjM9EbB+KVvxe1dX9omgz8rbSf0OtiNRZKQs1Qjr6I1
DV1BuplNutQnWrYc/9KkWLY/uVZkv98sL97A46f35HY6cq9G7weCTyDtokyOzEA8NJ5cafwVeHW9
5tGq6gC8xeeOW5ON7GyA4xFIwMSlhjJvl7Mq2RiIvYDfeymARwmcqtUMe3UWpcR+9WC7zEu6F0mG
mk5p3KX/z/iA/8bjCNKMRpX1E6IgAaKZvNyXpKlIZFls3c1zleoMQpPEv6q7TJWsRADIIOLp4lO+
AaXeH8aRVhZUDaI/zjuYAmez7vKKDdnfA3+0bnIc7uFlJlM3EL8/fZBm4Fa8W9HoQqz8jK+Ie/wv
X4Y+fmp2/zskm8qgdvo6roisaF+PC0OztWEVVg3oapaRpyxJG8u4n+buXGhX4vlUuDKkMN99BSBs
qc6vR2RZcWpObCdZNsA8pn7x0RDeaY32n8cHyesypsedjvo9NLEJXhhg9jcl9v8akkciO8yod7nG
II4h3jHuLr/Mbdaq5WK2OWPImWt/C/7QiM+cQc2c/EIgf6yv1H2lw3DMh04M5LKGWIpdTfgTjVM0
qjy9PJxdqDzVb9BUE12+RbBYtP7JCrCLNpay1tWBSRu6IImrc4sfOM15DEil3r2hddtV7RIOVsKL
CBShCQD1fcSx52XEeCuxk3is6eLBJO+lFZ3PcLJ51KEy5blAtuLxsS1GFGozc+iOwadF4+CCKnSh
GPNgZAMUqBT9YFFTPLwbSfntOC/ISs9xyquoawg8atrzPDFUvgjej6PYSmC74dFPdAuWfLnZsX33
4IF0+1GEJdEopHBtuIQpIOQRLTPULs4EDSfoD+SHxNEHGaOBejpcHVBYaEn9MA7tA6D8/bWt3Snx
YIqD89QlZtursPGmUpREDek4b+uMuen50kZBSP5RtCsTm57x7sSOloAxuK3kU8uimwNyQoSJOkvS
335Xwg+za0oul6KqR1c97tvlE3sIAii4WWtYYDG64h/67QmI3iINeLxO+UL7/jJ5xLwo4DjkP+EH
ib2/3s0CilZEb6jVQVzbqNQ9GocSxvFrnO6z8gRcwwyIfYzhGSs4vN1ViRbvyKcTodo4uY0Fh1vM
EU+WvW0pzfFPrUQJzU4iG7riyxMTNXq6OnYK/AfefpRCOWo+oFrtjip9HLBknlV4mPd6JMOeKYvl
gLzqkLkyXdH/6tUolR82H3gOwPmn3nZbQ86yJ5BVIq7mYQRQIThv8N7Ueu76i4h1Qy/4f1Qx5pJ9
TQY8Y2BIkNBChjkVKlYIURASIcUuOkh36+/2Dd6J7j0+4LtAulqAOZeRk5nCuGteBwPLPPTWR5UG
nnHpRSUeRwof2rM/qCu5B6o55IY/YLs1gNo45Ku6h8QNhwBW4zVcRH7N/YXHMyGWhs1KnXvrYtvD
QNZCrbvW66yIgrIwuTSWNPEruhGD6vRO7dM4zlTwFxc9As4viPGsFsPWcQjyGvGjUOfv6qffz2in
SHjoinPCL30gF758EyoWvL0mweqVVWC7f7Cae3Km8tHBpD9DbPMup4O8y/LuIJ6rDDkt20hwSnWi
LE1ozmqYlGaMPnnrrfmM0AHWxJfXmy3gtIfeKJX/eJrpAQnGmFq0DaBHN+U2tUnOowPTR18linxd
SWgnmQipKQCELlLC0nu6JNaP9Qmy9iI8RowhfpPWVbEuFSIqRLlsS6DSjw2ncnWw0SMXchBVVwDv
Ktj10/gQ+piOsBcb48jcRB97kL/5nanUHRZQ3UlY0M7jgqtAJ01gsJRo6TiGVEZYKg9JCcUCfHzT
ZZsf2xV5hZ+qq+JpzL4DO0BbY5h46F7rLWAnnnsxx1QJjJTb9W0h5HJmAvVeMgWagf8OVN77j4Id
SVg8qW6OloEo5prjWapZCFfd3LNTo/HKZX1+qEc68AlVjUaZ6gYn2C38vjvcPTQFesyJbq8Nmnc/
u0M7MHuGjaQ88A5hCRnrJyO259284G6t/o7Zp4ewD8q1Kc9xwlkBfHY2knG+6Jw8ZwxX8uTI9Yx0
NMcmrCR116dW7Mi2pXqc7BXkSpe43rHfrq3YFgipphFdplxvzcMh4IcVsIGapGB5vM4KjniqkdVp
vE6kPqtqEJYrv7jJLG1kp3ForAm5eLRjQ03+xVhZi4TxARjA8hrT8hFsxXutmO3v79m8tRTgyIDh
HSOMWER/lL70vCs03xnsDgo4wvY6go2CYf5/kTyH80d7Kj0vwcKCLHhaIWT0i+8Gqk3YKr29RyiM
BPABdudY1JbJtzpszXSyuUclOWm580OEiERIvdx/rO8c8sDnhAnVVE4+fCB3jIpxZXL/6/Q2SEnG
oXilTmiFbMkDshLiTaQ8oqBoTLhtYsyZt5sD2alNNK0yt99qix4T9fuokAWoZUXzSgbdtz+/mDQs
+mMJ7LbO+QHc5tbi2XGOvFjVi4NEKNUKhpIbfDnrWh1wFVBxZMBtnpCPtLl2s5nOWs4caexduXZH
D6mHYeAlM+MM2RyvRlu18LRAkd0YgdoRCiqt/L+SvEqZS4yh/ZEVYdWTjL5a2ompeiYlFxe06CKO
8KYKymnvUTuSIjlWD2lsanxC/TQoH9yzUsaHXEOwDogn1DbUd6T/ZZmM7p1tytvKS0BRjRRnN8ev
iERdKn8nUmpiB9BmkugketKY3tAY1Yk461nXK4d9nmGn4oo/9r4XvUAN8HyKzqzndIjFeTahSwEz
QrdmQo/rCt8G4Plqmjx/cI9z+mLuEFhyiJF+mKeCQieEvwuada5G7WljtB/uirG8yrz/Z8urlSSJ
ZcCCnUBqgdgJ/v4TkFVmlmpUpPp18sZzyTgZU+q06plAkUIDQWvFLhVaN8Z9hqGn1RUbApTIphQR
7yiz5nlJqJaLHz4JjkCN1+uEZE6jLWqqmCvv6cuKYd4WHD/LxhUnnf/GNam8Ml9LjFhbYsgD8aIc
WVvtcCxrj0LaWaebQRe2edR1fNSFPiTSnF9mFbaIgel/2MTV41RrjbVV8JW9Ugn2n0rwy/SSzvhO
IKbSW66mq4ssKNrHSSEkEeyjDgWStNhr3wmxAS94rBvJf/C1aiz9icAtXBNlsH+nKq3w6b3UlYDW
WYU50UQyI7L/WMX8IbZ+sKVSlHLmJBvF75eZbrf0jFcWjmYxgULnwyIMRfUMSFgJBNRSFd/PNOOy
3XrtHKlPXltOv+DXlCgF2c6CNNRcySSz9VUiNHx/ICOv1CHtL3bWqixUGWO5O4eAVfHePSotf7tO
Ko//kqywAl4xeCVaEtoMZCPYaOav2UmY7kUakntQrv+ujiCmG04nl4j433StETp/N681syn0cUTO
mTUX15rOCeAl2MsHjcSKrvZ1eFO/zCSM1n/y9zerNKYwOecv8HgkZpUxtri8nN2DLZBNA5u6k7d2
k3++wlbXC1Kjc3/8XxFaXVAYOmiuzktDs0VeKeyQVm6sJMqepdEa9l60aIiB8cvszZ+9zjd1SZ+S
1zMK7cL1w2ziwMR3nCYdqfzLHi5nf6lDZ5m/hZkRjfZXgKTVx+W9RZxg3u3JHRmHhlcPRyldU+FX
hizr6P3QYU7gzGR7612UzCn2YZyvKriKOJR4w6ihsGrPTUrNsVocQJDVPXSpVqg/s5VbqNW9LJP5
zsNM7nFywD+MJI2PhgZlF/h4Em1m1q5T098UycJcWeV/tXAwvRkHeYiggEV3omIVQPOzL5TOcH8b
LBKrQWauh6G88yYaR19wLNC8zxdLtMOLBgum1yIQBzDz8Mx+lMZw5x3rzSPVUCQydaX6CoLhsr0j
urbsClNP4y+d7lA+I7cz8o+WpjfHzTL1S9dQwKHSYb6dTEDkmweawcaz3Fdgo3s5CSenUw9Op3SO
7VXvHn2shLqSXcPwdAcoeNrlnlBT3CqYiZwXz6FShkBXeYi2wscgyCkuXsxeyOytUs5sNkSelZLt
DHInkZMSGLmgrC93IOdPTaBqa8MutNDJpEBlQ9M7D4J5E0C1itsL9aS6pm4wgV+WBVhSqx9tj5hS
c5Ge1RlD4GR2tpiSqj+8YMMptuBdo4UHmFyUbT0auhhEHmvCChkxGTFJZceyl/peAGRmbVB1aww2
JL/D6+9m0FVPTsDy93Ljm8ByTJOXg6j20TGYPAZv2gSGM8B6pIPMFVGwO/0UmTbPuFVhZa62sIEH
EHtpkn065N2LIOjuwP5rPGO8Tm+zMGTW8SFalcwLAqZMtXp3voAJ86ZguEWkY0x0pr8crVMO410M
+0Ky2P8SGEnhlmCTrP2x9m2iU67lrKXccJCDNFRxf7MJGkg+jdvk8x/h1lV8Wb2RQPmt9gCFbPVx
M6PqCp5I2HiDuNumXVKCotJaSvQklfATGB2HWv1hrEEbV3z71GkE4BBUi0ZSDoqXZNn7emImmVK7
GKJD5XPdnWbBBMwlK+rUaH4VP6qonmdFcbEZ4Gr9sbsAe75UNDyIggAGqzgHS/FgrZ113FbeVu/8
0DAl0GMhxOjXU64D9Lf1cN23xia5KftOAtdAbW5h3JwV+hnb309OCDJsl1iaTb9KChVQxbtS5/C5
GoaVrueVts7pBlCwBquvM9kDpTj/dxXq4m6gG9xx7O9wFwk7UTqyPQM/ASvKPnDfwDz616jYI9PI
58tPqPEtaY4+Q2LUSuoAKe6MQl7cIu6MQ1J9WRIV4AkAUiDl5VqEms1RvAtK2Rge38Wwgn/g4g/f
/bPg1B8jNHbUc7C3aU6HFRlTcbkk4l40GLlsr/gX8eP6rn8diUJ0A9uxiQqpK+z/R7n0mfhTPW9O
ONmrQahyH5dTsivBD36anM0kQ95mg2k7eBNuqS0M3VNSTqoIAdudB5pDvHeG+E/fMcCRTdqGejJy
wmy8nRmoEFFZ1d8yjOkZgb01BFAPP9ru5pvJ91JR/Iodrq6HnbENXYZiwe9F/qnNkQdRjrnAsHJW
tF1JJTtKc8QP4ns+3GZZs4f/I4pJqfUwO8YMvcvpw2LxikiA9VwDNsInFYSOjYxeFEkktpcqrMkw
WEg5oQBB7Oi1MsUImL3GDsDVElY0xqAuugVL7owYu6dA7TymaUcAgqJj3NT/tv+vm5eHtgpemftk
e8E0uDK39GVpGrDMAcv2ePGyK5ce3UKq+URICrhdcgfmPvR2gH3Hwyx3WddWExGsW14hQ+ktKISY
mI60GxtHJpKeJF8xWaLMlAR6Ehy1QT8jdsOwEIfqgQe1hQ6Dn8L54AdRcki5NPgk7z7dXT80u4Z7
J9gpVZhGIFDIIsrJvskR8XX3efY13TS73yeIWLCIY1gP3c3doFli8n/ayFV2ZPe0l78055Vlsa5y
D5QOvfEbW2PFOWyOl0ahuGIlP2Xpp7dw7J/RUpPH8ZcDnTvFiS6qBjzTN9n+ngka4KIQJ+vKuQqN
HyN2OCwtqDwyb0TmLV6+J4sHKcOVHm54eYRXRRGC0ZAG+44CDMAtxXvwLDvRp3pNKDJyyKmE2uQz
UJ6PSN44qACcI4q3t5wfXoJ7vynJ8MEYiEBY6+S4fEtAmuAJvAvWl5/gDQh0dGwuQd2rZzdoM1+f
zs9bpCWxMUbBYFM4QkVyhsLpLgpY3tvUasjEwkt742q8Ujvr/dPESfrvc4ow5vTRH71VWEOHoUWD
DqUVTNWJ8giaepBnvGXrq4PX1KoTSh5MtYWVCvgMYV0zcvDqLIB5kraza4rPtneqn4nJoooSDWuI
tt8H2gTP1lbFDVp0dx2gYB748FnpU+9T8P0B0aXP4eg1ifuD5W99LHrgakYn6s13qk9Q2EbizWfV
LTDNGkwl4GSDe9hnZg6Lb/at1+8k3Qikmg/7o/rblUUkeQUYHXAO7GnKRCV5Qgf+jvLfjWbTmrlp
PPT/9z87x4jQpVQMCvkic4DU9hiDN9EeUZD5GiA1zdo8VsMe/1Dw/g15mAprKKq3xzSOHoegHg4p
hOPH8J0aZtPEiWu0TTuTQIiV4gzVPievYOrrul+MDPep2wbaPDLumVA+VXOfVIofIz+j7TMk/erG
32Cgwkp0rbX3SHBH8TyW8H3/lg4QlyqXICsZL3F9Rz05wreQNS6uIGtI5akKMDqw8PPLSQbcBDuT
Pzb710UNIpWl5wEZGChJFv6m5C+mF1YXPatO9obQ8jO6Dvi/ZGwvPuUp/XrYGKR1tbUbHkNUO321
TwqjdS+uj1xmOGBPKvvoQnNXXldhfNGCqAA7Pj9qjmaXs8BnxxCpBl7+H2D99MIzqVcBLhEsd8lg
2/55M/4jYVr2JyUQsnRn1SXJOkC/iuaSRo2BtzfrFX8OZCaRq+3lc8OKgWBbQzRthvH79+NmKZA3
KRP56GxrQ79wvb5NDU0EV2V8Q9pPYDO7bC6Myzh3VqgoEX1UaqsUwXJr76D+/JWpqsyBBNp8vjj9
gP8qj52O2kt3gUaQEPUDE/C4imM6Zb1A/qRjU9HhujL0H9tDxJpnBbG1rIVv/hacPVKXQoI+DbuY
cnRkFX9XksOVEM1snxXdpr8dtQQN+0Nm/jxCLAszwA6EupYSVh8bFC0un16FVsLBbw8Gkk8N3l4G
o8oXDmVbXJXFywW1Dgxx0USqQ/1QrA1OMxAU+hqCc6zg3l8D7ktwJJXx0TQTTZFO4U74C86ydukr
ONvglAqIyoZ7jhuC4sEC8V5VQWHfVyLCIctHrD8eN7ogY3g1+7FS/JPppnMb9xsWMiZLmVrNmloT
UuAuB3mp22rWZHWHYUbhW9ya9vivGXpHT3jhHIasp6ndcxlG0efxYfBGdNoXCRcGxprMUc8FzJ9m
PvPVG/N4wPJ9meH8zEuK3kSGF0HkUclslS5ugLpbuvCBsXmlBmZ92doUrWzFGy3qFf2K0R+plHT3
/Q4dozZY+pH7dxUB7U1s97NIT9r2Sbm8RcjmP8HvqpkhovEHsB7NPw969s6RvAWe7U+X0OC4Ah5e
FOFcq8MdmVJME3u7nZ+axSsYnwIcjvcZW1Gd6AtnJY0rtyXbhTaG/ficVwvuDpeWCO1Q0pIfegmZ
5s4WkQtCeQOrmbS32Fwo+5u0rjGu4GhjNf52yUW5xH2duQZhADhhljpvptrQAmK22zDXqwKYpI6R
tO7Il+vPd6DSIiC9czyB5vDF+sn5EpbIl67dHJStXhpPps/pD77uNulz0gytAG6bVYQsfob/kfRl
q+reS8wyZa+595PvUmpUqEC/RmApRRme7z/x40auJdSnyE/yEUQ+KerPR8Y7Ms3/EhD82h4+iZ6O
CUsXb8VyO1nrWVUHyAIOLOtKea3WeBK47w0+JdZpSbCx6moimb36SfwruYcyLQqgbWhyAuG7Y4uU
GjVO7GLFuv/mcgIGPtnkrYGB/7EFxEzkjAda2+NlFkJCUNKMweiNUvH9THtkFWCqgi/uA+QXGyxt
4eaFyWALBxWmaHv6rMMsLEYxKf4xilcJoSrwimoG9y5OlejQL/XkXaDNR8ApU+M3p19GtnYf30Jn
guJiylL71SHkNEaD7IO5tBH2MljppMb1RjKcHxgJK5J8vNiC1bFypj8UNX3sV2VBBZPruFwP//RD
q6UU/Se5N+cpAqfsjNjjhYVtD0M+thU4wKYC9/Ns4bMZh59/6gW7GDAYvFzd97ZYjap7LP8f6qgE
dvX9Bp2thPw2wjqZVRUq9CrgnNQenfWltIJ1em4eosiqKB3xr41DcEplHK9MomIV0XZBjkhGpcgt
ZO/i1NoDEOE9aUeGfs9U74OPK2RfOgtspfOP+rl3HJ7vfI9v4qcCU3bKFpV39MOl37YHXnyoJO/Z
MqZB/5uKvcJGYZxKqo48+RZ4JkiXbIhXR8blwTI+fYylk32XOYXaPaP9X7fyAOT6CGUsxlWki9Ae
INNk71USz2cz4hvmbqAo3tigZiSV0GaxxWElxC5FKYLR86PUfr1j8c4fv6bLO0wK8XTtkN5Bqqp4
xGyrtlgJOwT0FcJTC+BoCLgjymirZ3F6tvJUoAC2n8E+zYlEhnGRSi43yaf1y7j/qbA9OelUlmbC
a/P1UiZLblfmptgJFgvycde4tllsyKrMMIILEnuVDnSI3fVkhlcGAkVIRyk7lFfdVl8slDHEq+Nm
FlYw8c3dFBXv0lZ6SJRp2majJb125TJQzWI0XRzLkQ5hBHEN0egNFZFCBuptR8gwbCQY9bGthUcF
q34soLm6hUizX4DpQw+Vl1CFCowG1p4lteAe1soI1X3OjdcLgpZsL0dqUpV9ixTkAFHaHLNebOg+
mnaJSzGt3S2WQXdVMduJFq5jNjXT54wvzzOwdn+zU4FurnvsTm9LK6Aj9HnZ3cBF3VOM/J3J4vh5
tGt8YO3DnWlKRbsVuSkpiQv/0HHXohIhp7qKZbVy4b6OA2Ru+uu4eZKnGFslJQEopkweRewDzzlP
HOLJf/0LeOX7XO3EJ2XnDy/NFGK1YGKMsUxOjXRj8Ih75ahRZPh2teGFstYCYGD6NRnNcxCF71VR
BIMnXAs4plinjoM90dDWB71SWN1U0rOBpBXwSf1BMcuLMiC+vOUhh4uDrjD6yC3HfeJY+N8ef2Ga
z1g8iOOmJlGqMw1BOlWvvGuM5OGrVgEprYnKq2Tp2ktFMeRAR8GVOANSf6z0kzgdaRwMHFnaREJt
Ut5aEUD1NJHw2mC46U+sFlYWts4BDCe5jxvUt+GKSMKkrnHsROnYJ0rns79+M8xaPDBH5UCT9ESB
2QtQw2Bb24KpNB9wnhL4Ovu5u1B5yfZDPRDqgSZimDByUqd5BYo/q29C5ugLMrcHVON3WL4fskFF
zVzwfwrLpsmD3VZBPMpOxE0XnEc+YQ20DUQKhjoqVhLMcvEfc1F5dAZRHPHIRXTfMwApMMU3O/Yh
eA/vnwTmSHflETHFfpL8phuB95ic0i9PDQTp4pTnznL2k/iV5zLNyy/VuNw/bo06UtchdX+LAtbr
EGXqr/1BRRrTONtuaSxeiHJ1ruJqqPetZSFxMyaV9IJU3Zjh8cPqioP2nwXBmhrTJYlNrsabz0VT
vx4C7w1cukWuE5QbXbgsWvGKtbDXEAkMt/I6NRuk4Ip2rMC05zmlIi5wUuEyktHwvN9o1E+5TSAr
NSwB+lUxs/5hhB0nQ3oB8Ltz4986ZSVctCPGNQZjRJfkLmiwqr+aocoa8bbL5qiYlUnx1jWZ2X1w
FqmVOsAG7RK/2ZnDE5Oi6hecWrCrea0kdshKA5JdhkdG6RLAxjNU+Qwdeal2D6+eSsBE7Q1eB6lT
bj/vE9eEB4CS3BG1T0KCvbZJN2JVg+KoreiUoADyTSQYMoiPNiBJatLg5CFh0gjgISIVhxmy1Elz
S3atwLf+FCAgE6gQJVnHaIuxIaWL+FtRe9fbQBhEeUSeLIGSlUGljRD2ZMH25pqELEwi1ItZwKfd
SZWJcmPxDX0jfE4rvIp4QIqHcp02pSjcbtMO8xncZ128DRT9gi2sT/OTUDUxYbplIngXC8ZMyHNO
/VhfIYTP7tRq9oz2O124eG0Jk9f1FVG14KxoJ8BWByfoIOLY15dkNxrYVqoH1v25Bost9iC+PA09
GE54TaGMe9GxWcRwNHXaKr5ka9R80dOYNSpLEfAcZFVjnQS3/3l204N6/7DrwytcUqX9gBNbuV6/
+u5+0MTTumJ62oxFc155b2hRwe4uflqXMhlamTbteBIGGUgRhatYSnfFdm+qT4fQD3J0WsAsiqsx
rfol5sWTEUhNRMT0EU+RiUCz0EeoI5oKlZoKhgqVkG3/FTdTlL8s2BMs6hSDPIXOt48PJp0JuQ9r
aeNdQcSUzWhRNPTvHk/0ntlZljS7xGvugl61n+IPJ8zP3Kg5S2viw5xZI6U9inOgXxdlMl8CynWh
Rnz6vrAZISkLoeHuNKULOQv4gx3ecNOcftRBMGKnc9NMll0FLmf8Ytn6dudypROueIrlrxqKFA2M
vJtrlxXXX+7QYX07R/SnY9LNT+1+HynRCtTWKk+4jUQYdNL2hcYBzbq5hzRhXPTGaNN7WKMX2ryG
s3BpUO0SVWXrp6zqFcev7tMaYcYC9efE/hhK83LM0gl3/6Z7j9BNfaLYZBJLAdyUQeqbHpJVU5eM
nyITs9+5QW2kOHm0zOEB8kadmXNDBQhikECme2k945qKTkzkBkNhRp0Z6P9kBHvnLRKojsQU5s5H
SqyzyPhuoBpDDJh95j5wx386pSUPyknn8HWoPuhqYB2CgyjqPLum8EdX0KD/NrXAzyVFcyP6/VHE
wNOvS8x5gnswL6PplAI1sXKHRtsqr6sx7asZTbFGnOnm3KlUhuxu8FdFyh3Xemy5uOaWcRx+4brP
AVGH6DxgM/f25v3ppYFAPEQ/RqIz8Ilp3gg4qRVf8kTep22b9lfX5zYJWbwvCsUrrIRZdsqGUjoP
a5SB70QyYW+H9B8MY8dLy1GKB8gAXuTi4FdfzFvHggi9yMcOoD8GfBxUGfmGRACY4+njRK1Ppp+T
9NzSP9qBlmCX9JLvpSRTtFHmsaCIpXRkFbCBfdeg7S0Z5qoXl8/6++5AFnVg1Dy+WoEbxRxkaa9H
FE9MDiPcePc69Rh7mOW7N/5BLRKbQTECJam3EQKFVUnL06LnCtGWeIjq7sGkkKVDMdplx77xTdWt
auxSscpPTMRraHSEfCHqG4epui4TzNg0UvHYWg7IH2mR7rqYyQTiSW27BbiZTbA33HG1f45et97q
zRPUx/03cVhg1y4q9mHGj1CaKomJA5s+jTTH3e2OKR07O+4euHG5sl0LsDUS0tQxGhcQSYmn9BfN
CbjnKQ7Owa+MdIESdFIXlNi264Pwx/upo+ko8LqLKiHLOG8nfgwLbXI6jmp883F4wn3rvGDNXPL2
1d67kcl9q7u0y7RDm20UimU0ExOWasTphzjxe2/J3GGlXXHp7YB0rYJFwEPGEQv4bHREsmqHfUpv
rlcsR5/tplQn7l+y+VOabhpmAz1w2mY7Y0GPM41YBHirPH/j30FJC6TOWhQp7EI/bDDixuapLWTQ
8etO+f8+kn2er1iyC5tLE/2gpjm80gYTop/k6qN+iYncHO1kzQir1j1/uwG4vBjzOwH8GDwjCaeu
eXkThCoJYq7pjT45a9LTGgYKczT4r8PiyCDYaE2J65EP8tY02/Om0qDBwJayi4VoZWVgYuEoZvpc
fh00oAdaFsjVDQUzo+qc31B/ZkfneAZMQNvKLKDy8v5PHF+stP/Pa/MNxQ5tCjnSQDqOuUNNHLwR
YmCpkjwDRIez/trrnXLL0w8AAm4J38FZ5+pG6z/X0cRZR5fir0rZmQNfNrmwU5yO26EhjSiDUmjH
cl6PKDCsx/ZM8FQklMXsnL0i6viSj+Gx83wEku6xGfxIS6TT0EMvnFTL4Pv7/RjQIwzSQCfSzlh1
2eDbUdjZpv1b7+zLAltb0ptPYRqliRSeeKsFg3j/5LJ/qy6U3RXXoYzvh6/I49PA6CHtAA4pjiQ8
Nhgzln60DgzwGogSIBZjngNDmynFOrZzdKMrxOaPdFsBD5CfPsMMevOP5TPP8OkFHXk7zxXLk8uT
Q3HPrzw8GitLRfdd5a3mE7+gJelfdtvpFJEK4r8JNE78jiASOqPh5ubA2bEc2WJNMO4tgojHZ9X2
r/U+ebOCbpFadQtuD900cfGNTNqOudbiq8URS8/Nj3NGNrr5qdvKNVmxXSbKVnxWg3OxO2u1sTce
83Wu/k1Otz1kfHfxvlH5kKeDtCV8pnXFABNA8jdl96Vu0Ai5CWNMZVl2SPHHHn2TmHjehYXpL+Aa
MtlDvPhyy1ZPgaR7jaECcd8zKLqBbra+7IlJ2YU1W+DjR8ZZTP4V6FAYyyW2Sj6uJzHap+9Lj7/P
ORMV9B3JFs5jLm9tsf5VCjYHtl7jJ1Q/Innmm+3UVEcfBJw11q73CdmEMwI7x2xB0HSxJZKkhwdp
Q178EZIE3+dLvRUXpbbnUg7LZYcbrJoPzqZyd3EnXU/ymZdJfzxRq0xZBn6bT9aX7kuo+JLBV7RT
JVCZ+ksPF5E1yWlzwigpBhCnXrGbspKqTxbJwjGEsb+HiPWgOHCK5ph/irO2bvsbz+T4nyYCryJ+
Y7s16UhtphiDMt6xyerV13qT4eMf0kKR3CK2nuFZvq2qN8oGFAw0dWm84KtlHx4lxm9I0iBIE85c
9PsXypaj67NINZSvmWcP3h1U1vHQ5VvNpCSpzdMvIMvUIeLdOBAy9fNeetry6BAwsuBf/lLGfISL
ixjs5W/unUz6B7kS9JRrEe9FbvZywJ/YZ9e0rWakanVOm40f9mzPvT9Te0ZdaeDvU44Yppfsp7Zs
R5y2tHoHQ+E6qyNqSGBxSYGbt7kgSYJo/kp0qpqhYcLBMxtRJdJDifpL/CRzEbFWKPpjTtM/zJAa
GXbFFquIrcLwbOZ8Cz7tFWD3cG+1LFENmWM/V9bHeAUgiYACS9fmOngp/u/GGggU8nFy/Cfc/y9R
0C+DxxHfrLaBanXuXhL3gOIrNUpEQmebZnVWI9hS4bHisZ1srvWPjronyGBdzbVdCUaJBMu5OVZC
zs+SNUDaBw4wIefFZJSa3/RBINoBTlytmh/nZbuzEsIsol4414aBtE//rq+uqycpGtk2S6P8xH8Z
aPmBjYknHkXR1Cq8Jd+u9OfrVshBSOIaayZL20HJeU125bxP8mdPyuaBwA/t/ajEjnQv7XXmvTa+
VRKMKXcWPPTS3mAbuzTfyPE7K5kO84jbHBagmHXxwLsYaISA7e/mDLA7z57H8rGIRZW35cTJs2OG
hofh1NPFB08KvF4vKh0sWkaYzeXTUUEEzyn2YC6C5q9kybHNY+4tG8UDzV7Ik9fhO+yDvxpdYSLi
MpByU1vCC3rSoab4UobrihWZFncl3ic7ywkPrfwSJUJSOXLfHij4JJmnGMMxYYQdzctbEpfBKBmY
gLVQ4a+F9GiWEkimUJkEwA1bo6y1I5k1fs7WpfvlL1L69kiXODpFEw9KR4FRn2enlZiDc75MGUv7
eN+z4D77qBv5YrVWqxgPJhmJL1IcW6BhyaVXOGIWwF0F/j71Mazt0xGVgGrqOmBW3RadRVu+ZB++
o73tyKG8qHeowqYMAYwwNtlhD8dkgAcodYSMANY+d5twKeZWFVUtQCFLzsk6m78bFl5TjYWVfeVC
LD0u2HxeuNgHFjZYd051DaNNM60BqmvcG53d7kxstjQHzs7YxzLY8cPkvXuxhoTRNgidu4k52HXM
NAO4oiy/bgw9g4u2HCpUD9Z9N7Vb/JSrrer/WCFqNRqxEo4wAVqvsNemeBnTh9YgsmjxBqrc3zKh
a1+Bm7peUpLhyHcy85KDO5JN47/JyMuZN9GssppnOE/IBJK5ac2ae7yuHEzc6Th3wXy3DItrQb60
4yQrVtezXHrehlNVr5fBreWOgWWbnetsTR+Z5y1J6vIVuIMjKPzGPbdsJVFjH7eh1X5j47lllALu
MSmqodx1jRp/aNWajQTihqba89J3o8i9bETEyYLXgHC4K5kV+Tglw1+fnHuLRZNIKCcjI1SSagJx
iXsTft4pQoQViWo/n2Xfeqqf74413PVs3HUbx/O7cuCNitmVaw+JPrnGP8EAfmbDK92CgyMIH/La
3Djl60Ua4GrpEv4PMj2M5V/20BLUQNfnx9Qw93bflDUoVl5FGS9F3yFSbMaaYzO2+H34QQPkeiQa
u3kBWfsVYhc9NfuFEhdtWREeUQAeES1psi+gtF39MWhZ4CEnygvCdpCTRZdFe41jORQe7MZro82X
UuNNgEdRVqdIpMu2b0O7gt9cyT1dqABRkGbvmy3HmlrLQ56udXMqiMvWagal2gNeSwTvDqxRIl0D
nP/vrHxIKLWdhCEAAkn9zTH/lWJsoRK3WK7Z10XrtchYTL7g+GDg9i52dNUhF4T1Wm8vBzIUxVks
7BUCICZ4K200d54Etoy24TOE++n2f4Pl4GNe3sPlPcCggR36AZ5YLf7TJlxaomtn2V90/iTt84vR
aRcZnytVW5jsfLz14QUR23zO4UDTunqj3h8lUZUh4NlCiLqV5FwfYbjUlLl4pqObDcFewv/7lYY/
SPICGntf6SadMO7iwSFspzTN1bBzs0PRPgf8x+I1qzjpRo1aK3DZXTJLuFZ09Ao6VblcDowWtL1j
rjpbWj93vMuHm112CcDu/7cDxE3+N20g0aIkl+SaG+OVQNMG0q0Xq2KOr88fiNt3Kk+a3RkzFlQp
OgM0xoLFCqkRkxWjv5JkleHry+eqe/zMxdLJFYuMZ1Pv1mdFL4J0PdGSAgCKGNHK3jfhaskN0n8k
FuIgTo8R9FXwcUDynGW/FwS/tz1YM8/DdFyPIqBSa6wQGhDzAQ1wmzLO483QUcFexBOvmUhQQu1i
XS076ZKCIhqueBFYiVz2ASR12IlD+e/oDExwmDsQFiHROBPw22TCGGJ6bC2YPZd1gcVGV/G60IC7
jTKYJe10QOtVXZAWYIo2oM2FpE5NrpwYwRcxKhcaKuhuhsHM95+xRxfGhDvFen+GaU/02l1SNlju
E0dYW8iLrdbibA1L96eS4ltXf9Bu1SNU+GFIXMBurl7roWiaEHhdTa4SGlp9/Ql0kjWvANOjHCsG
2jheB9mYA+I4g0kTs/4iMAj33rBdWxdeSp1/OhuY5bHe5VuqzB0c8w7TJi5z59w7A1HNoBKJglxP
O+AkfYrcYnfIg4g+6TL1MUjorY/teztFZlxlku2oL3X9Q0bmeIWliqN9Dcwmc8YTwYTAW9XeZ2ZP
r/6ZIvo9nTLK83YXggu3Oobq4FZgXqutt6egTNI3ldMQsKTXCHLwGotOeWSirYwrPeMf/amge34C
LS/1gxpw9pkz73IEdYElviS5rtx1EbQoe5uiZPrSwL2YaDQLInS/hjMzvaUg8QFpZR2AtFTqLEa5
vKPTqG70iKNTJYz3UE3av1/EpYtyPf+laOVMDkZFHmAyqf+GwD77LpfWASp/b2EE2XW09rIVxY4g
e/HCN45qQSxcaGZ4tV/PhYsfmTuujIst5JqIC35XPeNtIozzrq1DKNP2TrS1UO6exstZfG97rUAy
pONMnKYmeW+/0DEPR50dXItrBqVT9BmAR36QmJXBUv27yeJBBIqgxo2PWAsR0XGeCznZpYg3U9Ry
e3NJ+aWmtxEeWOxeQtfZDQIn36QJQA/EEdU3eyYKEjmsaeonJVYbcsVUAcpowhzcicVnvd87g28/
gckdvkn9nmFpTSRtP83uEfiC/BkhnECZiq+YhxfD5v1rpqsKUYOz+i3ctx1e+oKOsNg8rFqydTSd
Y7xxiIPyffJl3siYIDZiALe2tDOtuuTkOZAmQSNC0QwmuPa0Ta7XZEvcS+Jr3jzrqS6HEW4sFxI9
yvYK04nZdzJpDS/YKCk3AlnFaFev8r7dnYCSuLmgb0RrUMLn95kIw4PxSvDUwBZXvBmrjyC2TNAu
y8cbepRi2DQK4XmLXnJGvMyFlcunowJgaeX70cczXUvE/K8KeWs9A+aoqRmDPvfHOkJMoouiHSaM
COkgqHneDKWbqiaTKlxwcoS7Kl+6Osz43gUvXyjknxirKfM2fCY3LPX6U/F6b1voa1HsIo1PBYTs
FQosH3mLu9OiHTiBg1b7Zj6ocV5RL1xAlr1Y8ftuCrgourMW1WBQ+ty92TaAmKRlJ9j0VqOzFFt7
Kbw4cNSz1Vn2ol1wS4773AnDOJiqTiBMQrCpwLNSmxgFdZPRllizTl0Tfnfik0GgQnKFZ4MRAmNE
DiyubPFTupTLlgN1V41xCg4BK4Z74VafvB0rLsYMj4BXqY+AJWkpKyVgxVFdHAN9TOlaffyfwBWe
Lhrf9DX5gajX5Ib1pu0YsIHVkoWjvVE9Hqi1OqD8dD0Bn1kyikdn98v79T7rWOMiEo+SEgVw71Xd
y5jeIqhzjIO8rcIrbgIKbXPcrmmkDrl3Iw24x9ihpZFtlGaLSiiBx6e4MYq+/D5ndaoi0TJW3WdH
j+Q58Ij7oDKEheTi84Sp89bf8YLH17UzpTMi7TEodARIhn1hgfZkVSUa2eHYemGXyrS24t5IEP6n
apSSaQCxRtJADxivNMU7gBve8j8983+DVDp8GwtSo3DvQCNk9AcTeGKRb38GdoeHVmrVR9bzmSjt
XcGlR5UH76A2I7BQkRdvpcDsUCprAgpXPHlYPfF15YLW3QCs0pH4/HakrwLF8jBD9csk7HGULR/n
NyTN69zDVIJM+xiWKHDZ4e4dIFr53KfHKmIW9sL72IE7EWg5BD+/d7WOHX36h3b9HvwGkmfnyfod
RzV4e6L1gTw4U5n+9Bw835wwPvhxaTBAJxarVraCF8Xh4MHZZDBZW3h2gjzHxbXtEA09jjCSKh55
c27CxuXI7EzndWEibfTYz8DdvRxTF47eZEnulHfNWVE1UUjnNS7io0aEgf+j8DeBJ5qJBnxAs6dZ
fx12w0cjNLGLIJYBNkN981rcU/tvxkJ9RRDl/waoFblaF35lwodJM+iFVmv6lKusxmeyTmah/oMG
a6lJYT4/TaaZMeGKfHsUoye2JG3hDh/il9nfT419eHqyq5rFKvQBtY/Y/xK3FWc8kiyCu16EY2wd
2x+t0GwoTqpRIa+u6/kvUFeTQWFb9PEbKnQ7hvYI0aBP+hRUcH6LUtsCoVey6B3zQdiltG77jJj8
ph8x+RUDrTC18a1cEyAgJC5tb6ABMn7wA7Dd4bwz7kpWlcj/bCIN/g4i2m8QJLkIuhwNC+DRKAne
X53mArs7QgDOtMqOldxj82hSJw2e9marc6nbhumEn7TTix0R7jr3qkCMHo15RdOItkRjMtwM9/ED
ePfY2fvUzS3pjPYQZh+LxhOHXfLrzuyBNBIZ5Gk7b9CM+8/0RQgkKtPLxAKqZfFlihcueK/s+Eg9
pbXshSqFgK6YHfuYi3uGZemDzn4JlV/ocz8XgdjWRxCf0i+wOIDIkMo8a9gmXRxQJBfbNBsJVlnp
lr1hF1APD+oCmqRAvbG0B64qsvFoEoInxsnw4WWi0Ez5NhKpJgTac/xavS0Hs5ZDP1a5RO1QZG2q
HPkxWPe3KDY3tvvzdXlvoPhpGLp10LI3ij9M1N99t8uNdd5ImFd1URJzRu+4PlaYE1aDyHxXFmDg
k/MwhXbC2TM3hRPFtEsSDphpkYbhvcsPf9deABGooMktHAa2hAValWDk50ihtRnYZ977j4pO0i31
7qs4CzSGKFco/Zzksmtmk9YgG5xc1ieoOuzYUy7u4wjlYrNpQX39LwK60Rxbs4beVggNSzAjWJGu
Fu/rJ7RFpUcqpjNzNZ9uUlfZv6r1zCIJXXR5jiMdubDZo7VrLdf1K8WPlHVy3D4yvfp7pCLu1dNP
SsSZ8qBiUKKS8wcx8GGUd2Wxhzr2aBRQY/acGfJpsRTUa+x7egVrVc/030P1jgmImA6Vy36MLpI5
XKh1mzfylZjLX92k/ijv2uJnAFdvwrG3LNCO/beTeU/BP8h899baBA1o84zIfEmzj0yBqxctEeHV
ggtGJDh06ID5042kho+rIOjBl7Vgmc1Wl3lSaHznsJW5f/kHHENQ1i+NBpn4fQwnEfQKsCn74DJJ
+zQWOCILy+jsgw0uXsBaRhautFZB2L9RIDN3h9FBcgLgWAE+X43KZtMVQ02yURwSGhGWGYhzF1o6
bRIDBUs5WDM6hOwQG00VTFBw6hHLoyykzu7hRX3faHC1UwEqUIgfKJ4V/JZM9dupOtC0tGvTRju8
zOOwZyhMrGVgY117bbhiGoPEIgSCs2R5rhX6Oe1K5SZo7LaGlcdLip86VdRouNuqJtqC4T0C4eOS
ZR/pu1Gs/HKvCaybxCE/Msb1prAQFG4YBdmnqvfz+7KSf285pxVCFhOO1aTZdFCmqeh7905Sx1ET
mq0TczXWqItCG+S6XzR+c1B3t0CdgBFknhTYZ5cp/8EVa+VjzEqYSkhcl8+wj5KkzZEyFiMNZJgj
9EVKEX6SdLQ+v/ILL+Ol80lbmexf03CA5VrbLDTNeQtxDj8KjPAfz5sqibOt48RwFQ3e2QBoz8Z0
nz8eN4bqh7MqVjkmtz7stuA3usKr8Y6YkNw4l1TSXEg769YpbelJSDS+rGUjqxbqEJIjXj/AtC2n
fqGNmefTSQpTrOiMpvZjR4leuIXRab76FBSf1zys9Mtczzm85Bu/vSEBapwmpKSebvBgLcxIluFc
O1o7JqPuNq1a1ukDywA1n9GYBNB1TGnWAx/nm6ugeac0KIFaIUPnHkQeuf5QL6SeHXaqlSzOOBP0
596eLe4jxtrbh5iqog8B4kAtc2Rab2pS76DvPBqSaLJV2w9isRrQLoLvBOiM3CQ3kw2Z7QYmfvjJ
LwlJklwx0Pn7jGubmx7ufJPAbDKaGE+gfNpdk/e1H4fE/ydMvUxYAoDV66lo7X+cNVQCJsQSmOvN
0MT9Q+beKimznM5ASkEVFi94EnWPqg1My6rN4vT3KhORnSsFLU5FzQEjVgjo76kvyJtpZVSj/L4b
8svkP0dUw9hU51HWYKiJ7e8rIHf5xDyhW7M1jDdOjxFuv6Glg2K0EhPf40PcJnpt9EC/lfrSd5bE
IfxYTYpplNuwZSkQnLcPdgl17t6V3W3VEiYd2Xnqohx2F83nlFfwCjoCuuBdlK3C3nIb7GL90o+q
+lxbUWwjPIsIQJsguyKaR7ndTxhWSakvAQonim4mO5RaY/Z0fx1naiIf3KogM423Vr1CQn2F1mrX
kifSIcoDNgXQjEdKTVT3d1H/Mcd0WOwO+tFUBMDgA8ZL7lmevDZTyLMlO4uMhlYOcTqt7WH7Y9qo
KFRvyG1pltm5sWhga1sZqeufu2T26ZfanfECXU5ADQGv1q5Tl0W/E9zoQpimo8zyHqChVwNRZ7n4
JynasKiqFsk9Hz0sv0Rw6e463KkLNk2zKeCwH76zC4DUCdrKHOrbbTzqMubQzLjWcdh6oj1yP6Nl
LPGs6wjCL2fD6QhbYWEcCAbvy8WgVQd7+IU1NV07CW9Ix/5ROSK/fG3xXmLlbinqtWYs90Z3coul
mRyUYs/ywFMftJF2H55w8B6nH03zWTmiZ8ePBGTwFfy9SWarqDw55wt0pMwm3yr/Bngkia0UxNzJ
AgyDMWrFLCVjprwxC9ut/tebYQXGxWXwGArIE4zhIp6fsBw4fwtYX4LsnVpTnL2kupgo8T0IXjj3
9GLzvMYAViIIeySRNmflkk5u4jO+pA9ZzQiK85nDZpKtW+dtuMW67E79pAD9sfCMe73H4Z3adLMm
bCNkz5VbCbS/R4j+SMVKSwvFVPoLk7zXyui0H7Z0N3Ck5MOcJqH3IBsSXGKODgn/EpxFqP3jchws
GsHMiLAv7SyQ5ZdturFP/nt4SAxNyT1E3N7kcKVM3tuEMzVHL4lOIXgi5gh5cCdJtvV1Hjwh7fMv
w8pTK8KmJxBA8gzWNFHIvxWWLaBMSzv39a5IsCz+nqfoPeM2IJJs3ku6lwZ89X8irAAGlaJR94KT
B+d5TMdDYaCdie07Wmp2B4E2mLtFlprVB+OqKJgaqF9jgw5JICGCBPuduvPx5sIuWSFpaf6TrgYs
YyJ3NGzcpBqZJqTT0Xpg4USL3LxroOchmV2r5XRj418gfi9ZQetByoYcdEH6U84XDW/ENzcjNvPG
LdlWQ1FD8jRD8X8gJI8L1OqYnxTZRGUL03ASx+QOhuR/qRBDNvvt62TaAEXV+xvcRfGsr/lATWAD
g+ib02yOs743GUOKzPG/eEM6DRPo6kI66C+BabqT4bYkOG8cyYTDSNc66OLBjHe8xyG1jpkcvFDr
sFk/ewDyvbOUiQIstnAzEQ2e0GHnkUMfvnpVPFF4JHFnIxwHRpJi6EXCd9+n9fyboccdWJfpj9nF
xoV69QoGTRQKNQ4aDBv12tc1w0R/so89GpgJ44hQxVhLsi8hAvmqp9sjnIm4VaYr+EbB9aGk8G+Y
3tk46P6Oj6IYn35NcdUeEXgWQ3YFFE4EFSci8yFAEkGn2upoD01tye5D2rOEfjF1Kvj3mrRq1CjY
BVJilh4v8BMDgsVwgKVjFGeYPkWUESyHZ/bTn0+i4Lmx2s6jN3gohSs0fyO+hC8R2SPm/dHjguGE
8bFU/Ods6SU2r42cjeZai3yeF17JqtPE4VTz8huP3kaGmsxVd2GdeRo8YebnP4eBhKFuzzD9WeEn
2EsuEI7JP7dZyZsNqvCwHaekBmO8rMZIOIH2Kj7KPsD6IM/PFkK6hZCTTCAv+4XcZroyuFnARBCj
ZMC2D49Y24PnKkEsaWkSBNTgniQJFYJJ+HDsgCUxsGuVZdUVWkE/47tDWmGtqLgzZcyVsfu1J4k5
UEnmtZjnhU43JcnNWLGTW+nTG1Kk1/uXOICd4EZgHtkCh/uB8a2VHh27C4ey0QGwzW70BMUAi7aq
H+Db8F+ATm3bWP7U8oEaT1KJ0dlk9lD59Cr+w4rwPdp/tbnazxS7r6o+iepNQvAvCvvrrqB+hFo2
dr3f+2rGginaeTkYSsoZdDTye+3xyrlbt9xOtcfj5tboFAEuydezv6n+exiJTefkVYjd0arxOP+n
SOI29yTpQBG1Z5fFt1/l1d5NANge3ezuO/r8DQAQGZo0rVME04eCB+CCTTtg/dyAu5uHt19wq9y4
tWyMQxrO0lrAUCfyU3ki8r8Q9Fx++wsukuNbhWMtv9OKYvTVjxfALr8OoF9rbeifg5r4RxIEfRCB
pUvZzD7/BrdF6YbuBkhaLHOgaYIgwWw6602P72eitr/p8q0VXYJS3ksAfBKLCjZ41A7g21cPNTPY
nLYrxTY0/qHxu+xbCWAungE3nox4nEZ7w10ZHQ/KXNBmT9eNR7lAweUKr8DSMOctxG11fXtFeIfn
/6ScqU8ATJI46C5CCN0CK16QxndbztAxQN2vNiq9QLbSfbc4OHxXTsygkUrb9wsQCqAlcIc076dH
mULhFRXXPTfp/G3TR62rjMxr6LFHpllvek5IBeU9lIjOfPGoQmzqWG6Pawl3mmOmRb66+N1/sxxt
Sv6zbdmqyhprjeSR0CVzevj/M/XUJvCZ4mlH7MJE2DVWgX3S+S00ESz084PI08R5NrS/to/9GF0y
bFL+Mqx5sffiXPIy4cXMWAn19x19nZSu4OWKP3HAx42I647rwVopJBnbdKGxTfQmEJrtZXJ+5Gk7
u83bL2BKrkZKU3VC1m9vs0XfcGcQNY68To0e9TdCmJQ5/Bs3OoM/Gt0jtECoInaIM9WDA25zwh6v
9eJoFVNFlGjGtz6DccBYoX6c1XW5KW6AWbWkRXLOcdmhbtsAQ4JDmDqn4oRy3PkPSqmq9yaON5Vo
CWJ+qbAn3URrjTWbEW2fXX3MAIZ9O+e2KWvJ6ikeVKbHZKhH1Wk1dVVlqkkLKa0sjGkftUs5Gv0p
p0OWVvA5puA/vtn+A3o00EfnVqJOojlr6VA95KFYsX9BK2mX7cqKgACLB+s2dwtGDqR1BOcG6OBg
IHnNxpW40YXhL9ZtAwfURtW1IQY7byoVUpEYpWcTKPddb0Fj5qg0wydaHFYN7DCjGdIBOGTMgXaA
phNCehQ9EHBjEZMgj0CVLXqEIl5e3DKLeoLNs/C+ODbq0eVk7NvOlUpPKzQzJNJJMSlZMpYDXe6B
qxY5XL4uOPwjUWudXUz05TaA/aWHc8KOI5tTCbsVoWKEgA/SmWQh6rkkSZiHmhyjPHVH3ysMfLH0
W6NY/WOKgQZ8Dp+WYeGpSngxqgQawT2Kr1BJbn8+0pEzuYU1dmIsQBDj6b5Kt1FxVbU2+0JGJd5f
DevzbGud3uMVD3apazJ+UzqXBYjUzqlsVY173cEpbJGFA/aGkT3AvLVeZ5Mea52lOvs2VSbreDpV
/XOwYWLwZ9R6fIu1tptT06ahj4AVEEs9JyhQ4Eo9eS7Bf4KDXZdGymzOHTW8NOTm6i9+XIwalEEI
uI/kyWIy3uNkk2D2BwiluF13OUdCEHF/y45e+y0aVY4VwGjRshizlDBBi1pykuVJt0tldqFnRorb
RlvxT424xOqcdDrmiKaqcsRPUEdduxMlWpLNHFpcSlceNnYIW51ics0iCTt0bxH5FZF+ZV9okSt/
xErImgeVb7gv/SFity5C392b+O8jTnnSj0FtNXNPp+P1x9J9qsC+IAqrlARHfVFj6jfC4q13HcAn
LoaadHmTCdfvnaiza9nI58ViRKJMUJENDFlAcYthF/OFX8oP6z3pgAaePaR+QqSxJ4+DHa1JopEq
PN0Csd/sot9gK4k+jOQBhEe5g/TU4Lb/rDjmgnUbYAKe8qVnAaRuxpeCxRgJgSEXScJs8rIrs1dT
9PVKeKhFSErx5vPl0czvI4a+KXnK+U4JV8u6jrXCXJL/PKT+GFtWgMg+MIvnRBFusfGEmsKe2PWU
lPRbI31vaOz6JoWxKJ8cRrGNrmGgPK4gS6GkagtGuIrqoPE6a9RqtbRGaaBMjqQjE5iGn5zyCTFU
068Pi1y/8JlbkvijB4n25/Hf4rB+HxgbkEgOYuhHNCf74lj3G0XdXwlpmBkR/N8rQHCMLWk8P3lE
0kqBd4YXnzxUk1OKRYsY3OEvV7R9i4v/yYtB5ej2Fn9aNKLpUuybeQtZyGefhWCceb5+blwi94cj
jf80GIxUpbvqTYimgFctkpC3K1SGHhjvVH/6po9Mbv/ZAGxDCVF/kXtTp6Z1VXTBo7uTjU8xfoS0
gwrWrxfwiU3aSKty6RzJNelCmEB/cnetdItgRbUz26a4mUeZVm1JegmyBPGMAqe9i3GF5eJXI5sj
NBSnXHZOFqw8nTGyWCYQV3OQwIUpOFT1dEFEBMg+6hTfmJQn6hHf+ML9ol5Q0r9lFbf0WTnOs9nz
uj0t6ZGIQpUQ7vZMYgFd2WnOzsGGvMFGLX+s6ddiCfFp48dW0aAyciG6vtlM5IAeW9n2ACvTss2+
riufEgYZz2hQuJtpdR4obV+lE0tQl3MQ51qz9U7etNUAVUj1HU/CNGSifezVbJ8+hHBH5GwdEA75
CeT4gopMI5DOSOva+aHo+iVRAnSbowslzq9yGbiWX17WpvAzluze/MhrbqxuteoORpA1kUjH4QLn
qNcjZm4Yi4vuHsirEiznDu3Ekrav915m22FrNWNs9u3qZQqYwi+g70RCZ0UyANWUYscGOEYkkycJ
GgtwUD9X0gJzjJNAE+GjmOYKsVtXmEd3A3ASo07DZeoHbjR2yxt3LNGgFbNglMa3JrfrGxEgVsxt
t+xih5r0nGxT2hoa+uMGAYnUpJskR8NSGiWGe1rOJyv6i5x6eL5YrN2U7U7k0B9nsdaHniCOJkso
/s141F+utvCmt5rGE2zONl1/Q0AHaDD6763SGK+nYPoPieCC94tKaIllby7IRSfM1vA+QFmI28Fd
hxpc0mVbNBRFZpQPMsVKRtrRvPKmLeQgeFG02vPovTjiRhV1QgL7VOT3qVhAblOsg7pEm+fTdgwK
xeVhX7oDObmrGWXcdmFIXxN4qi87zyT89wB+perMC7Jm2iIIu3vJ87hZLseqoBKna9d51S1etnNV
f6UAQAFWOxQGu+CKzreLmG3IylXcLPchEnEmKxUOLFT8kwt/tWMNVsgMOGGlJ8gnaPcf9bVR7+xj
jDj53asHRjLcIYm9YOSdSbii4X6QaAEjK48TNxLB+cFeE2z4yGsQgXO8YHXOxUb3tX96r0E6kLav
A2SbEKserLpOH5tnYF3dhiKY7elSNiLroI6PpXdYuWGyUti/RFiIku8esPyN6iv6ozLRCNwEw5CG
Tb5jO5HJJRYnwUug/RVEbQvoYiji3Y3Qr38F7bvrKthqc49wyLbUtOoD4rQ18Knxb2VLJRET0ZtF
XBW17NNt0mzHi7LdICARVPEXMozo03yLcJALejevEC2lIsNwT3l0g2JOvB7D3K9m/JmV7kuU3LoT
LE0YseCekWD5lCSznJtJdXS+GKSiI4FXeLIXuQgTF6z64JG4J04apegJlyyKn6wqqzW8DOvGmfOn
Rk4D4xZRJL25gA9nIfMqonH9U1MqKuy7RRVQ4uHiZL2ZJbTcMGAa7b0Ja8rBZNr0g53cjEaO9vft
wvYYFpDtHUlPYij2EOhTWKutEMPnWbx2rjtkPMCqEBcNua2RJMQewXKoNOuF5u0QyjEtIzzhbT1e
PNUlAWNytgWPPVIzK7vkcK+AHNoVffmRki45e6P9Wy8MnZyjjbX0vDg3yUiZTxXWXyOLE9P71N4v
2B+ngn7OvHm1reZPzXjCWE7JTL/4AqBbOOBpmhur1+JiGkBxIRqC0nA6oGs1KYbekVsbsDHB4llA
BI8NzGqby3fB/9pQdHEZmmZHZ+wuehmm/yA6BDAMc02GFlY8yVBSG4a5S2xt88H6OuANt5cDxsIh
QfNgSQP4uoS/K/EMWSaSwfGfyY2rvy20tdCCpVHVTo2/g7O0u8qYWv8WNJvNynON/xcrX42/BqDA
WlS1ThgOvbSxqG7LLE9AnR8Q6mjLE+h8OMvHRp5yyKEw04X9o5uGtFDl1NwOoICfQDyBkCa/q9v+
rAElvJ/Iyz/zC1RaRoxGI+lhgtVgOfI1NxiXJNtw29T1bbP/L4u3Atlw+9/OhfAxBkuxlhw6EoZj
z37faBOrfN5cG/JClRddFSwHbxkiWaX3tdAK8IWBDVDVZeCxn0NhkcVFe6FfkZ4dgulSZ2E8gt8Z
Oe5HyjY8A9xZnyxt+krA3562xB07BE/jMm/L+DpjTmHqUlRBDuZPfRvht3OUx7HOBvu67wdwohG3
iTrskTUVe3YsKch/h0L+JD4jqaKzmQErx110nG5rFWvEUxspRrhX0hOj8lA7/eW5fuBhUC1kMmLD
d9sc9SeEslg3WouKMRdUJe7JgLNxspo7r7Vs4MRKLf7Lg8qurEFn9a9pIRP0n7Oe2wGiUtAP46TK
URn3eqr+JZ1RlKzGl1Pv9AH7/iU6USFGwgZwEByfrv/cmxC2zKTyzVH7Ltnaw1alAY/ZIbD/X3qI
40UvwvnGFjOPPrrZ6cCf3RLPzjCGkMmkSoPt1vGPiygfgDulR0TWGqhjBUuyPE81WInvwXDyPuVY
bWj1v+DOwhr5lmyktrqIcrYAdS2pSjAoMdPlQip6x6G89sdEKoJnqs0Wq/I/v1/UFw5AiQ4VNNa7
IY9xnahMCOfBkE7fOzSPmCNyLdUUhZkXkILXCiZRqn913yZlmRZL4rgrrK4GaasgchxpCEHNlyav
B689Ih49RVLFx9hVvG3Tv6ZWkm5KK4kGtTkxfZJ4HJh+QAcXiMe01wRBdio7J11S5mfSoCxvCx/x
2BpOcpodlab87364JSzgF0WTRTMi/EIXUb9VeVerkIQmYk1IzqltFupLGwZ1i9zR1eBMPLWHB8A2
l9UU+hwVLGLyafPevkO/65jrVqrtIrGrbGw/a22FJeif6tkNHv1TKjZd8pEOWfFBDBrfaQnS784O
GSBeSfEkkc9/ksCPqiZBkJ08T/qrqXhbyveKgqFZz90HYvMsHe+HwshU0MUQIhS3D/oT9TtIZz0U
MQyRff2N8hfbFC6iOc+QRXWLvs3QNl8IjNtPSS6gBPmuzV0Mgz95T7fOrTszpEqz0HYB8t0SGPvb
YRJaStUr2Cu6oJfe4VKwLfmkzp4jOEuc9z4HyudY2DBDSf3PnDHqVnev6T3+ytW6gYvY0Wks00bi
7K7VivBsGJsXL/Dl2fbFHViKFlwQ8sNnTmbrkdAcXuMIBVhCg1mdYPlfcyAwn4r6+k0QhDWpxg4a
wJW0VP1ItaLuzDf3Y1IQn/KgkEbAwpKRgJu6FhaONqrlFGPIIZ3lCpeY1xEgX6n1gKFlZtzN08R0
9dymq5Kg22XsCVLVzZ26JhG5n7SGYJXNWFKCf1cHZ6ARNOWRVpS6B/xyZb8gxAuKRzMiRRr10Cow
U2h0PTHALWtRYGRHScexLgRa3aUhXhHhRRhgLBT24oI8qGU6cNvdJsNMKvytAXjWx7Xlmw3BaxoW
JUROSoI6/E7+WFNyybjiT2XhBZz/7vs+EeFq4SE6iXxvW4o+p+YU3TcGjbtGkAUdvqF1FYaRBA6C
PpDQGLK0kxTSPxJtzBkTY8DAWBv/MeQGou8b/nTsiqvX1zdcUtI+urwYM9vnJqNFWRkdfPZ3dGai
0tvcmDQoj7zWtNph9L6tOdvjOOvOwuQZcWXjzChwXqig3I/pneLUDyBc6QOlKqOTGXaReMfQVkdy
3SX6wOfYUIW25NaUZnLwGnoPMiNY8B6ESwrOUszcE26TDcTuisgN0/693q8aaWnRMQvdqdLogkQM
iRdJqvMZ6hQPc6ZI7s+PeSFitExXn9k59twwYNIQbDWMzzHsY7xUMf3xQ8vRHCavrVG+aGaPq9Y5
oXX1P4voIjyksA3OZ7AsKLU8gGztuNNNbOA4NnEi7Jn1gQNRfUUmGzFkGD0+MWNWn3QyV/YmT2Ff
Qdmb7zMUfYd4fFXiB/9GUFqlcOQdvgdo2GVZhmWDjS58ApDT9mT3JWb/WSrBkr1s8p4wf5q1YFd+
h7tf74LRLEY1TwJMioDPD35JkIbfApPXSxuSeasz0oKcwIon6bmnN2zYOvctdYeL5BZw7lgxQyZ/
5pmv+WNIqHCmmICNkOfhjJLr+B60tiLb34xgFE/njj+ySv4jmfVU21hfDH9lKzspQlGW+sQCt1ug
R2IWdYwUagdFNEPafXV5Rd4TWSba3Qs/dloiH8nUcK4+jlhaa1CZxMO9F1Ddsy3j7BPg/jyvU43g
ix8aTnNswHmfi7fD38/69rqMpmoolMi06g9B9piTQ0lToUlTbhxvDt5wlLXZzvYrmu19C6DU1xJ2
Q5N2M6CvLFnA3ivUWcZBDQRr+X7VcRQ8ie37la9MjsIoZzEKON79dzrrMrQyp1D8lmtGR7dkPsM+
kEaHXoIs66u1NQ+eptAPUq3AGYp6zsWS+0VojD+ZoSnK/NydhW6b5b4q7/tr0f9SZH/UKXsspbNf
O699N78t8xGmA79e0jhUNAlACGlD/B4rMEPalKpnWJ5lc8hW8KAf1v3Ba+z8qFcObgoDrY6qJKhN
tMlZ542ygq/KgHICG0RWVge/ImBElAK5Mhx1uP/GNgIbht/74Y82rMlPvpTExc+wyCOJtoY1hecV
kwVUiOe17aMSbb+ufBgT4rOyEdnkCqfPXCG4ZFs8vmmKaH/c1ylYiAtoJkEkfkvOUxpaWBggMlJV
7wJk3ua8/TPLSVCsZXuniAEOQSOGIl0TE14fq5HHM6yKYMNIoiiKcIJY9LjF8EAiRvzIHvYbukvc
0QqD1YqPuxxrGsV5bAG7iM9fLLxR9i/tfNP/13m0crh2GsKCO6FBMsA8Rl0Mh4Pg+X9iZyV75LOQ
X2KPotLOUYzy7AOUiLLuiXiMxz6EoDfsMQGMC4I6XuZKGtYhkp0Q0hOxgVcGHC5ChNO7x9CMzjYz
h8+G7afDf/j1ro2vv/hpiOAzgyLLd+nud/3I8I2G8GSUx3s0LgqiHWPXnabAycVhSjYTOy9wlMq8
O8V0ZhauDCLLqkBzsY/OKCV1HzjWMOMUl6eeNe8zlYK1Wv1HWbngfJNunt/K1xnggABp+UiJjhWC
ATTyOtH1hek0DOGRwBar/M/Z7nJdIEAulcVZM2djlxHwIJRCnes2/Dxn/cY0yrjyDUdsVcyogZSA
eD/LS9OPsSmSAIXiro56izDSNy5kKbYPpMbPf902B58MZA3tCi0rI89D1vyb+JlWlbK9W/UGqMox
dUJTUrM613eNpA5iT+qtowIXumyhhk4+aCxZhzov37yICRm4Luy1UC3dCNIHpAa+ezP1Z82i7Vga
gxdZ+kC6MOGmm+ffPT6ht8x4SOIx4hJMHaXe0crGaeud3ERM91CPLcGEMy4hqWIfphtQoQQ9+USH
9m4oFer/XihXoQuYbSVGLzWGWKkxiMGaxAURtI1Gd4sECPbMUPf5j+1WCuqgUa/fNl2jLAdQ9E+o
mtjb/uV1eEJBkApwU3zD8AaboNsrI6FFls02iKw15PwZ0fr4rVlfpkKzmF5tbthXJL/177uCOBxJ
qYgz86RxPO7f+GR69TpnO9daV7323achkOm7vYEPUbkBomq5CGQJJ57YXT5zCjYmeVzYPXIPzSe+
yi0CS5uhMD478nem3CAEWBF8lztlbmvaTxB8MIOXsMu7OYjTIfabJElwkHK5S7JTAEMz9miAMwdb
jb/B9VHGbFY/XhhQXFlokS17OfN6RYpFJnXP/lCDh5WSEOi6m+gE1fwMn62SfGxAbNLrDspo78tE
NvDG2hM6bG1z4NTOQYgTotYDSpa8zfWtcN3mGHk48Uiabl5y5jy8wV6Z3901yaK4Q0Iv0a9gl1zR
cM4MN2p5UjnvhZEohtsgUH2g1Xc2t43juwZy9NrYOY+uLCXl5dFDRvbQi8g+vkyDQRiD1OTmfLKT
R+eCurmTvGeM/PfFFzq5e65rULfmotmmW/N+rFWszhBlbRq7zxn6jv2ClmZZBw29hQ79yqKI4rf7
V8vkN4GZ+nG6LdQUYpY2uxyvzFTPM9JHYxTXfPAtQ0m5JiOOlyf0SWCnJ5GgwDt7UYNq3ZFbRElF
vTbLazhoCBiAk/vMAKgYhL1h97kUejtTL+MzceQ0xfPz3zxDM+LY6XKn0ZnsNG3qVtj7WHaV9s/k
6zs2DBfPJ/MZfDJb/ICsdDXEcOQBqByOCTvWa9VPwQVKCITybrid3EZm4A/id2N0M/6ctWBF3Ekq
VwRICwTbxVRKw1j46IP4OUBYrsXiiGLNxw8v5MBUjIRedVXCtXgdHelOD+nYW/WfcqlgSg1ENofz
Ypfvjjb7mruNrcAm4pnyg2gkhiZ7SimQCWydJyuaeqxp4KZRYZ5MdX60L1UNhGxnp55sVLaQVpbC
ob4Mzq/5fazSkb9ljTlGO66RisnZC0sethUtcZ2A6DLfAt66xWMYySzuBcw40TwmHfBlyjZnArQr
nz3x2V68BNsKEW9ODbwNQBcNoBv2Tnp1Y9m4ayBVEM6RF6D6T6GnHW2E8sgDHpPAs7N2Fs31gUge
Uka5l+17ITFuvQM7TtV2y68gEYZmEi4qLu25IGxl5tOtR5BSJDalutHpd1QJNzP/IElwEvWNNbaU
DeMjNj6fdU4p9DPBJ7sPjJ5BkJgYVnx2GbxQy0giJ8SVeP5zQzuX2eR7eOMQg/Kl6s2NZy/LiJQP
R/BZDhJFB6O70oN9Hfqltn13VH2UAWK5K5ozAtibdE9gN61otuoxQpGVrHw+jeLqpZYPigpLRVkz
XCIf5HLa4s5j1kZGILwO+nlcXEZyYuTcVZHXvJMFbinX9Wu1nZoZWDNNyl1HOALbrM2E3Q1ipoEf
CUecrdIUDdceLAX53K6Cf0hGN0oAYGdNGxVxBWnELb6LYgvuBH1kZjVe5HwHFVMvvrS/FcOuXDMq
/1dRo6RMcvIfD2jZfTjk1xxiypya21WBh+m4r38y1SfPfWQV/zRK3Z6w2KYXGFQFJVzFvfdj1itx
4ZaeglLzLOUaS+Muix3lnNI0ZkKRvWEi7GNYqs38TdURKWJkiO2z8RGID9cpxe9UWYbVJxfuIApv
7uFeQr2G/MSqRnfafjMgDO5SZXrE0At1qZN0+aAiA+GQgmXz/uvuNDHeOSqGitZzOqMWBz2fvbjX
Z7C+6HjdFn17VU71MdcSt2DqPRgpJsIV5SRufX/ipEQB8+a8/h1BQfrwFWaz9Ulxc3nOP8P7w/ty
FgCdzEQLMjV25HQ6dM/1Nh8K1IFho1c/trxaF5drr8zrsl+Ckj3nd4JsgmM2NQoXNsccPwYF8QkC
uzfo0GN4S4KuFNf282Zgo7ZJl65L93k5tr/AV6Ami4n4KGptfcbGSooFNfAjq5XooTbOusUxM8hd
EyOw2rBWvDhTWkLmRVVRL/ZvG4jc+wBChdje0KtMcU7rAtOnKyc6Dm2zX5RjnDjv/R6o65GCjdsN
SMPMJh4LUK4Tmgp60GsvhHbBTj8bE8sz39CQT1C/kPaUdjmNDOhXpoYHiG6cy3rgMoVwuRlGrbFj
CiR8u8RdLCF5E0j+nYqsl+/kdBcATGLdw/IgURWSDwO2aZqvoKNn3VqTaxL9DMOijNqsTuSjwibL
GBbkScQMDDkFmV7EBrBFxBvKJa3PVIb190ymxTnYmndodpo3eJkVysYfDXnDzPFUgLT/UvroLY4O
79JsnyVFtv/8M5wjmhQRDAYFCvrPd/6k/WFsflhr0SeydS0xlmNjZARONECWwc5yhhU9M/YmSLBy
oDARa801AAHRH1kde8m077cbo3q+pR9f4pbwAE4rV4e21rsi1mfxrCbp/GNdSWsqjjdcgPCCbHlP
SbNWDgRF90NmKRMKU0dnoON92TnzqsVOhIAB8D52twb3hxZhDIX7rb6J17kXhMmrP+ORANag9vRi
pokF6Qti6O53KPcp0TY48WDdLC9YZA1+8ar0eYcHGO0SXDluEUXMV4gpDW6nVnqiqW6sfduS/BKY
AHzmRT2gOfxYrTC/IWOimpS/8hKWe44zmwOMDubELXneZCZ6BUIeyDFec8ROlqEiU8updHNaSO62
hd4rT504D4Mwgij97tPZEsUYu0rrs8ZyaJ/07egVk7HE9fQGQIYUDAdKf8lCWBfCw6J2xKYgILjk
GzrLS143tgWn1ezXlMhFEe8dxb8IAB7CNi+n5kbT0lK1UNPpdoF8PW6I0o4QE43AjhDzVbdRfmXW
nXjY9BmobhF6OJIvC27P/wZM7fEHnWhCWXYkm5GG5/DVEtbYoaJTcCOAjm3d4+DWCZbkIGmzm2rG
36lOMjfjbwNydyylBs5HAgKni4aaUzNMfbky/YQWj6zvCsQTUPYlRe773yuLbB67HFPJx2LJ8lq5
eLt8mJzd0n7gyFLx32jgZVkl1IdBIBuo2VC4YxAynRp5KuiAV6Y6vyNo6yuIJDvNUmcGO3xrkR55
n9NevHB2wRPm1fztGiSUXdR1cbvPth5PPxra8hMQfljo3hYgONKW3TYVvn97o1BQTHxJa3NcuyBy
aviL/Wz7yUMcUc3Fp+JJdAR8uxS5LpI7Eszn+1FQKQsuClrinWIr7k0SOMrQ2bDAdLOvihsgyNaF
CIpqqYsFb3q/Gvqg5nqERwnqsSB+NOQGC4oW2KGIgYhfcbDkIcxn1S5VCnDHDZPyLzZtMD0H2bFp
yO7rAsbGnZzswKEH0mu4xerD4uR1lNV7Y9pMG0QRSVKKqEdDgHlHmqiioUhVrIuz20w4R2HlID6X
PkVRLN89Z6FcTPGuwPUPwdNRACn6bcViTDXU87S8+YNSv8eRQ3b+ZrcjF7bfEf3MvO27urflZ10r
+qxEdOe0Pr+2TGY7VIA0YMvuHhIKJ/t0QUtWUkM53P7Z5WrsOQ4V50gpafon2FG2Tem2I2lbtnux
7hid31UBeITihCPvn86LXAuawMrwUDtS/kdWRlMVr6iX9yTctT5wxibVVQTxtXZAzi8MBNpVxsHM
fslLLgNrywG5lY9X0NW9tlrrj5jG/X1xCsF1z2OhXqJWiwjh7t/WCqLXwybxdcQapd93Uecv7+ZE
wfOR3SMbZt0u/MrYB/2JUZNGpNUMQAer2EtGxWv3/56RaeEcmeeE9qQCLZWfJCfz+gbX6S3CXvWl
B7fHh5RUjEeWZkHwn0lH1k00E7H+Yv54zoiPzw2gWr+fSVrpknMYDVDiTGb2yiS1tzIYCGAJbA01
/O9syPGHbKQZIpEVuWveEU5ntVRa1PIDK8aYExWueKp6aG2NnqU9xd3w6M8voqRH21CmM7+shMmk
vHe7+dKvbpsfUfkEeJTzSWt8YL2ZLwq2re45Wmpp9dHGgzVGHp39l/tVkF9bro/fY+WtWVBFI8Xc
tKq7R/rPNcGXwDOvzYk7lYrQEYeKTXuLHMDRdaVhL03qdo3IHsPx9GG+X1rAE62kZGl3EEIo1Jd8
AiPKWk2ReIe4dq77A8BcIPONafoF4oSsUOCRFtyiMsbXjV3fSSpVzS8V0JAxj1voGQoLTtW7wmKS
xYIB130lLy5dp1JYMCI5NH6zcoYlsO15/SHETcZ3iNehtmkJndjxMXAIV4Sm0N4abJXGv0IGsVn7
T7yFHDl2VR9q8lqoRb5Uo58pwwREk7p1C18IvDCUTSOvrtF+Ibs5xl5Hgnwv4IjNRnZvokipNiQu
RKoTdAKlm3Qw0EmF9Z6WM8UhYgC6Za/+yOwIKeAE5QgC9ZHbPf5HjASK1rylnoaeNDSdRhF60CcM
TwSPEjAmehJ5cgEDITMjC7DlMpxaB29a3bNpX+Ujsf+orWm68B9SpUxDmFVP2EDW3oAQPzfcjnRF
TYmn/W6Dsar7G/tskspeCWUJ5rmeUmZCsUXn2a0834ty95qfU7ePA3oTExKDw6qr1MNLOehGde8A
J3ByDKiEXnJoAZ2mVMoETfmXWAy60Yfp7fRjjTAubChy4wTv7RT+0nrxC63NX6tkkYg3wVXrkZUo
zy1n/u9fR9CCwAOGhZh1rZvyvBGeub3VFBIComRvesnz4uKvOusSFh2yDfZGrU5qrA9/QqBuqPiM
E5HKotNAkMVt7g3UubZm0ZNZSHCMCWa9XUqhaMd/r8vFRpHAWbhfOVY4HB6wUQK4IU1lMFBZa4fg
v09Qjp4SiDIyr1e6YHS49R59seHL8+DUpSjAw6UbD8g0XbAr970SiaEyfuKvWD9+2b2qxeb6KISo
iM2TpDqF1DZ1lN0TslqmOjbmIhAEiGZ6l/rc0FtRoDWUwVcUPgiAMfWatFgV1fzPAqI2QDvlOCrp
QoHqKp4wKMTMFWgRFQiY2DU0UhR6VQr44xuy63eUg7QWKQVifsaLQcits6nrYIvNFB+bVyPUIDV0
1H02b+egdNybKj8S+Z0uUHvl8SgbKpluloFfQ+EQP2mRvNyyQGuUxo7Oc3Zgb4L5fyC4VrNu4PjD
Up2ADcmUy5cDcC9FY2iXJV6014Bm+0gN78YsZ//V9b+hf20k6xPUZjwCF4znS9HyD8z8iu9Fav9F
no2IHBlyjeNmx4uhix/yjjmgSpk8LMB5Ddj0KR/t+A7l9+uwN+j34ynI46tDxXxc8O8ozAYDHgbL
qBr1KldlldNxBUFyNn40sdbOxBC658qqbj+OInEuPBkg47woJ2cfZYNVMyRn8qwl07m5nUkpGJRt
UM66/jrFN6iZgwRtcEHqFX5nDeFGP3C4HZZ+xSYyOllTPrBlS2EZNau+JWB8ZZwZqiS4DuwThx3E
u11KqjHwXhvhtJGjP5pTscRWnJU1PRM8nqV21jE2zqgEBC/thkij9NfehVJPjTQEIVVgk166XdJ1
2EdXfh2IJ+Gfj/7ZUIPmhAPIGEVAGlEFLvs7+RsXSEA7GF7v6+6uaJojjGZCr6z1Hegje0SNON2I
ARr7hOuIRVEBl32+EvpbWX23hRA27UCD4dIDXbIyxCnZHNePqB4OfDetJwncDLZ4awHrHVIAIb2V
BCz/CArEqf37NVSaiYIqo2Yr8uplGK/rkg6vS8jxrrgdXZUHvBrCVn46sazEQIpZWmuVuXGHyCDQ
YXckMOTKQaRzoUgCFda/FeG2bGH98useUEysecBuIXu68DvfR5ln20aJQAxXdItPrJ/qAbn87Wg9
N9qAqHH9ZlxzuO/LMOcDa5Y76dhaX0t0Msll53TQUq/zRuurppvlqKJsH5H5K0AN32ItQyC7zGSy
y1b6OQp+F59vFsLxWrsARSn+9yN936cwMnfvZqlU8cFskuOBMPfnHpnJgEI1GjPWQ/m2n9yMHbAG
stfqoZCnJ5hrKGAbuAp/xEaMSZbzOR/PoNjHDPi7qABCAfREX7AjO1PDmg5koU8H7XjdANaTRXG0
0NpMx4oPV/Cn8LxHE7bA/joEoi6Ra5r6E7IDGShdTzwPUichZ9C9Hm+Fo8tc1pwVqWIBnKDVi0D1
Ocol0xZRoHLueE7Ar/so3X89o8oI61jJC1wJtzq24c5QUy7aGDliE8/66O3ESCAYCi/cbOwb0Pj7
5wBYslzrXOxtC5CjVMP72wmhGXymy4BI6SX4pECedZ67py0bZYLaEtd0OPxQmHyd4SulnlxyFKg0
lp/L8ihvndx5NdhT8V1h/ByqasQXP+qSwJGWyCXZFCx3TiWLQs9IL/zi5wMeZ3sD1f8Qt+kQvkob
12lvAzQBTNcR3DCOrY5nYBZdiOCoOIp818SF5bdFny7xt+m4RowDvDOO/f7Ycl8D3s0NgssoODxv
DGhqzfimAO1eBZDv8ManeJhQKawVyEKXo8Okr6f5XPHxMSb+g1Wy/gwscbjWa3fnY9FLQeBGOlVt
qqUtk/l27CiLH3JdOxR9iRmFjWlrBun5o+Uxhou+B/R/Mp/89mDIeRbxFoJxHxit2eUwQ3lh51v8
drkNZV2auYCDMRTA3NxXUNo7abIuZEXxAORaTKS2lH5Vgi2X8+c/zIh+CeTT527rZPU4PxnkU1gO
mIVmu2pMPp025YY8LLtsuXgpmygd2edKdeRTukJd6/a7S6fAc8qyhZGW2hB17285D6a5nlLHMVms
mdutLJGvG3a5N44Mos59wS7oFSmuzhj5Di/6Y7l+IEupF5LsGhvwCuW74V3UN9NsmSSV4uOZhmXY
DJ0eadHBGQanDmxsv7juGvVCKImBRzOiPNvSFd+ckAuxvT2/3UnknHLOjM0ATmR9bBCs0KQ8pSBp
9nur1xA7traTRn5RF6CrzBiiogNXCOEvxiRBbDH+7rehmj5T8SgcLZNOzGOFR/pNYT1btU8bj4si
LghZfS0icfgx5NlscGY0VPPeGkn06n4OkG+VZVu5QNoirwj6v5uSwNuUSr3MGwc99pQR/yh7wulr
BO3W5rCj6+TONFdi20+sKTM6+Y9Lv1RUzeCwaKKNAF3iByEma72CiRkzof/LTEfGHVjvAmqKsT68
GPSfeoqXpEMQ0kms0jUSoVwOEJnVaFv5WFEWTECMGSQP+vKQv9VPFbqja9SJLFSXBNsPLB3JrT40
4KAxMUVCnhlZXm4La0WBZ0YyhsUiIhD1SINiv7BSqwPVZsN9k7Z/5wbgMOWTNmDxty5PIs5Yi2hD
Wku8plAUKwxs6iLNif9L40n9NXx7g8Rl0P+KjpvqqAB8/+TV6nlq2mNUN8z8E5lsI+diyIBkTiqN
bP1RZ3Olc0XslRA5jL4TR9Qo1/bwHxrLOBCjmVkbAZLXiOhrsTQvLo7s34//NPK7S3x0nB5GgoWm
RNVTbscK9bVMtD1mvrEQQfT409zuapRPfypSkzGvVPurPVtSVY7CLGlvWnVgwwNq/wDBZ287LiIp
gutCxIz0wM6l+94gsLEgk7d3tEvmAn0holDL8ezqrFOPOGuxv/puY17n2tU2sD3Njm5mTG1kIB87
G5tiaoTp+sgPXKqlil8MESmV2q+x6hGqEUOi+UXLy03HWOSYKsJkPm7tTBf0lCcyznKFrzv78nyZ
amtbAJongv/FW+ndfLQ6zNzO5GcJWH89ocu+EHCYehFOJJHNmGrBWQFqAZbycDLxLS3IUmT6QMiz
dKtmcQbUK7AokM1hEs2bFB51mbT+W5Nqz0Up+n+XM6FLpnTb4PMxCbPP3Jb9wVWKA7I7H51+xa1T
S09JUcRnghFcdbqimJXlissge79OGa+1Itn7SL4zOAU9kVlRKsvjCWEt7F7tEZNFBn78akc08mq+
8TLtcOYUavCC3t0FfuSqoZ88kzWr9EKA/ErnLGr89w5gsaXaouw4Aig/rmHH+CdCIz6+JhPS80t7
NCYmsQcRar8PJoDnTjxrt/y3xF+l+tnXYPlzNDTQjSXOEOX50PLyNR0m6iJispQzx2ENQIrrapWd
B8VpIWhfTfN68QyOiIBSBY5zYa1FUqi41nmBjjvpcUS3PG02evp2vO1jvUI3Zlfxm4BWgvuZNkfE
WxoaJzSMHrAc9XpWgZsHYWzbXFi45skqmym4oCVprkjEtf0YJVSDYNdoq2W885VenWPkWPx+DEyp
fteXYQwaH/g/0+x5WJnM0NNVjgYaC6jKGoa8r6YKHLl5vBTIE6LnzJ+sCZV8qsXOoVoZNZ33HCqJ
yWnzjsYwn4jrDhcpjU+idtl+dYAbvKelW2p3gAigZbu1dS7VPHR2ewE0H29wQFD/oT+BQf0Y0jKb
YwBpjmft/N9UKxoa7ND/nq8hGZABYs0hXbNL13yovuzYlaA88NvhxpeVmMwgOUsHLIAXXBWzm3l4
O6e56tYmg8aq2BekGmLJwVF6hmDcz0VTD0/436Jw7dsiRGbZsGbpaoERSzR9bMImZf3OQ2vuMrcm
IR3OpoA3ulvD91gL6OI0+DlA0fMONz3jgDvIR63+tM7Y7+3hMY4vY5PEXXZB/o2/imdP03VDk1fX
fFghGv/a9K4wnCHG/mWT+4IOVDLycEx4P2ELJXA5a+hWVfsZcSQnZt+sMLmBB8nfvkbKmPoOvFbg
pIOVrOTl/FUjPkTMOrOCsXziSbM+mDpjKpQDu+pm3/jeWGya4XJEYttLooHh4TXiSTHCFiX28mRQ
LoAwfK8SywKlaCIp+2c2pfQyiOEELghN/mXbxYWFbOUZe++opkoFq9YlbmqxI0vfILPBSS69Scu3
ntpbjW+RtqiOVpYQlxa21dKwqtrT0bdQTX1cYYndK1hC96SsY4VSQu8h5/NkYmazbr5kEiJ194uW
aQAZXpH4Rl6sdaoufR6M8q18hCz5Ux+/ytbmKx/JumRmSRZ4Sxm17VW9Raijef4j2xCDh5t5fvGi
WC1USLydPUptd2Ocz1cjJi7LbyE2Sjw76PPphj9hnITDsWGtdi8Y4sY1u/jUI0rxZJBhVh7BrmL5
iThFLbEYPWwDCQnsgpSPpZ6w1l+rnnoXFIyM2tX0tpZ2o1VTYn4ty/+sAZQ24/JJ3HwkkbL14RB4
Eo67Ze1UslLiR1L/GXQSDrqNkJ3hVExlNRs6DCMUKCY/8hJ/cZlNUe4lD9siEOAzdaL8IEnQBiUr
yYJlQk9uoU8YMztPiyVoBFfxnY4u6GCMdaLUDjfrzfEBlzhmh2sP3VlAQdoDoMS9OthAnI7RbOuu
omafKYhoOMPEYSVC0sR1RP2/1yGEivirFMebSdzYgP5iZoIkWHkSwL0fV+DoqOykyLb0nObGieNd
qrmfKXZfsgp4wr9eOKRp3Y/NgFBbWoPlQ7pCKx4d7gok0ycZ+j4fSsoi/oIVBh+4SXT3gBbHnwRk
beeONIwN1IDm6G3flaeEWrZoWRJmEKQmGvl0NELFvnrERa9ZUNatcxHtUPp+2B3DDrUj5p04YA1Y
dxjSLmYoPxucu8asS8TxPCxsat1glaDDeGaWkBy5c7kVoazD3m+1F/qyu/giFKwvellJhl58Nmcv
i3r8Kx61vf7hKeTbpe1D/Ho7aSxeK4x7USV5+9UFYdu+qGcr5nJFfV9R5mXMv/xoGsibP/3J0W6z
2OfCU9/sV2Jsz9vtZdjENVaJPFxcnfZTYdXAo/k+iSQnamCSs7DB9x+Gen+E0jllVS2SioiRXLK9
YJCQxC1pIAczad38FMVX8yh4Bek2sLSvKeFXw+xZj3NKY4Z7eA2JusL8WZKB9TEiAjsDioQZNd/y
YVRzpdl/qHDHYief4Xn0RY/PwBHpnM+zoHDtVZg9S0ema1f0xuTDOEfN3POcLVSMR/+RVNYKLhjI
MF/d3NW4Z2HvJh6EZo0Nbql5r0wJVEQpIrCY+mXomB6Q/gBk2rdVdCu2xel9kxKMa9bsK/6D66Kz
O3rU4zDniQUtsKTKCN8sPP57G0HhqYtvj3tvSx00xC8t8LOKStxehGCNfulTFPRWCJdwRxE1VV8/
Whbd703EP3sMtZAMNcY046VSgt0j8FyoZCMZQxB8z+0B2nIoKKo1lH8J2M5a/Le+sWmURlN0HZEb
gBUwqdCcbmLCVOpELsaZWWW9gJzDr38KipFQo5xnGWlyH6Hiitf9xqvbhZc9VjvNyud88Q0kLT+S
BFWSWXJNa9LYfk4oDgrAjxiUJK5s5OirpzvmhGaQ/G/XUT8Ofg+L5VyTgUdakwOu/L58c6qk9uzD
Cpxs5rBgmqn2WJ72CxXZhpGPAeedLe7Svx2kPphvRhZQApDPVMbs1B4pfOBw7jp4KgQ6trm77wge
ppu2Gu0CpWHLF6fyp1OXcsKkFIXvr3/u+C9SnV7DQZ1wQ6jHP2xfNKJx7W/Y2CdqwjtbLmK2Go+T
S1uwPFEOnWZiaWj3yniGjxFwV9qmrsGS8NVHNnNA/agL7wgf1GvKDKuJyFq1bV9p7VXJ5MOm/D/c
LAO2vZSCoq8MTzlKgoIj6EuvymUpyzshfgtQaKj4fkC0g0NMoyU/WvjK559uHP77kROXs4FE08x1
RGHuS7tBDMpj7C4yTqvEXuOSu2oxVzHyDkI66i8/XZsJNvjrOkTD/XQzHU5Jvu1LdJR9A61z8qYc
lgepPe6fdiKrNa+txFhio2Y0rWT+75q/0ewc6XcqhUftrTdTkONt+LFRspJsKYI9Tw8sGztRw2qN
x4XTmi9z9u+GiFvBadP3zexYavGAUVx7L4+d79sGHKbwxDrO93t8XXV/LmbcZDrwFuGQV25CW7cc
LTsmAfiY4yvGAZ4tZ2ZfiZAS1f9VgnTpTAWWcTQpf/MKym6OeSqLhE9M8g/eXfJ1Ro4BlAGNzQsk
YB1BWL2xDJP/KVu4ctxzXbN1SfNM8lr1ucraq9iHxcrV0/G1vjGLjqFFl0itr9iAw+cy4kSQiSsR
aLwksE31+KYI15psvNkzhEbbm+JL+xEQPfB9UpvfuFaKtVy/9FRtBIdNYJa1LAMhCD2y9LocJBx4
bMhVz26IaQoXfZA3L2YagyCfUT4eA+9zudNCMqSYDHH79FyfOFByPfpz2Pjy/vki0bOUev2ed2P7
Fu6YlZKW0PTkugoWsBO4+zrD8RnpOfBTw+Z4hX7+RNfE3md+c7OTfOqBGcwsuUGqKoHx2jpdf2Rx
PXxD7NBJ/TSLbux3rFPQNKJ/9b5NEgwl45A26+BdcRmOPYtsdSW8xGn/xbVYB6KnA0ABakrF30/x
76/4V5rynyhMW3vIZI0jyOqnpDRMlbVDZP4x00Hewgh/Nk1+vvl2Gg+UI/neiR4xjhv1ypAZJOzm
DZJwyAOiGTVSrnYHGAj22SSHXkcGs3PN7CMNCCrME/xIoHcyOwHqktE8DwLkORbwKNOuTay1fmXF
Epa84OsmI0F+cVqGPq412HFOX4zVuIR/AmKm9pMZlaGkGGAZn/sbKdXEgLnc6gma9XC7cXPFX9j1
E+RyFk4mmJItrODDoMvBdz+NB8QIux2NCm9nMf3ZrflOIuNcdDAUxiZ2EZ4fFRUxcWa7WAiyrC38
eozOGHDXA7aNWBEipWWNUalAMU1OCBNonoPNBLo6sMcNnkK1jks+MKC1eH3qWILfX/qFNu5DxNq/
v/UTS9SuE/wBG52DXEedC1033Hl9fXykuRQLcSUb4YsBbwlnSXoYmdBRzfcJCvE2dJ2VYqTcehuz
HKs4lu9DdY0gwlonWG8akww73QQn48w19g/nYwca97lBnrgN+VD+qOGqlGbOo6mL208Fl4Lh71eq
cLkUwy6z6hqyGvdM7WLfLbA4rFKKq2A/ARiJcDvNsZg11NOT3MMVvJos7mTTVBzlVDP/NkGUnj0I
M/ZWnehR2nRmvFYgNbAfhpcYEigSSUfpYi2VzEuVHw2a0qpN+WM+dFd6SuNZS1i85euUiiKXClao
700vRELulWizCNj197208Xoe8xIH/ECDevxCEuHuWf4+Cvpg5cfp3G2koA+r9dQC4YGPMpkMpjXA
I7pczNXFz/IugmbHNkcy6FyiPgz5gT5q7mhmmcwqPR/aJKQ2U58elyNmbOfUTTatpzU+8pE9UUPH
a40KL4thyK9yr02iXLfQNKLy8mP91OIUGk8Cm2Z8Xv0UNJFd5IKyWMXu/4tvylxJTb3T3as/g0Sy
SJR5GBgfaOLF4KurfGpb4JeKM0LU0lABKDyePrr+EDTswYFe5GssA7qpTx0BoVf5L4tVjtwMDWFB
4qMVect7fQv2gt2UsV3uMdT3cBVhaqAffP9QJx45zKw7vClA3T/uszInPWV7r1DvMWkZrTvAR+aP
YRSaoAcvpM85MPjy5KKZDjie9G5bqvt/WRSXfzFuHrUJkabfHI2+Kd3CBTDOC8U/kAJ75CILwmDp
3ZDVtMtso9ocegdvJFDPlBi5pJZqmxj8mkdX7w9rQFl3JbKE3h9g10L+BOAX4XvOrNoTd1KpZvzr
J98MXER4TN1fLPnwnEOSc7t3MzvAlqJVxWvNyoyo4WgDSZOfxU5tQWBFzT49KgLgitPdlKqjuqhg
ttuZrUaZDVkfHEXItzWgUiihykijsU3nt4fEjuk6DUafI6kmMr8Dv9v2rNOwagBAvPfeq9b8YBBl
PYWQ6sKNDUve8CzxdHKhyWStxFqGhUk7p2qWQKdcPUlxEoNLiyPHaWwSpYvz5425pG8F6P2zNx8+
T4hFaNMPfFHBJLUkWTlA78bHuWM/Nx4Q3ZxoZoEwBxl120HZCWAGSpjMLe8QsYzVAEuH4KNgOe4e
fL+ZdPUuJMQ0JxN0N0E9tmwCjSf+ByTDiaw9Gyedl2VQu0F2IQsqLt2uLanDCr8C4WqdHD7fEoJF
OcMY8+omFpieeW3SbzFAu1s82wjt8+omXGoubOnTjgyc7///PWVc5oFsTougRmpEFd717/Pp3ATN
D0G1B4mmPoQEG3iPQkpgzxt53mfJmpFfvqu+iKvto4hhuFvwxfpPWN246VRirQU7uKenoYTkR16/
qBksZAkThRlICgqVTIINQqs1sXQjA1BNIgK3utb78KYS6ZGTHA7pmRc2Wv1NA0H3F7RgkxNQEmR4
3cekgZ7q71NufgVk2LYo/6EwxKVj16zClX5x060szl7xz7DlMvlpgMrCufEgrPpWZ5u0XgvYUkvU
6TyiO5ORqTCp1i5pcQI6xo5DJ48Xm/oEgE+qKqqanitM78GzURonwHZ2WhWjFSJ19eVBW/tq2zq/
GtbCfKiHLoj+vbpz1syuZEqEH+0FzWcS5NFEIHYTDKPdfg4SlHP1yxX5hqfgsjNXPpbkv+yKXNVE
ZcpH+xQp2KhVa1oMLettLn7pWD58dHMetAdv7APUjptqOhgQJjOAEXDgMF3DOG32vtFZFucI6fPp
oeodYk5KudQLus20h2Ql+Q47QRs0r0UANqPfHKomDZqHG0Fpx0m6U/Iv88fUTmRLdk/1Bqv9FRCU
Ok18JxEpX0Q7+EvZpASYUPAx3pMVhD13ITWRFFvVJK/u3cWY+iGZdxLkOoLW+XNGMKGJ892XA34B
JyB1ajNJk7qMhoX5ZczaXnGeDlDChQUBMXXw/TRYamHjTODpirxB4I7uNJb130ax3bVWuZXy7F9c
Ryf4xx0dreSUgfu04LyfGj74RGJAZwJVv4ydM6hio7FAZ6hjkIedd+ZDgiXWjSxvP9q/SyJ9HqrE
oJoAuuhAx6CRf0kMLJbJbNfZuzpmstLDXN6l399Ke//aA5tUjxpYogyk33wOUbZN2OBU4ESdlMkJ
3L989CIrlWUYwB89ecgcPetskQnHG+KtSzRdK/8LrS9/FUphcJpUho5v6R/xzpQp1x/MlbPt+D9D
truwGKDUc/QF1Xg91XwFFa4lclV1TRFQsVjQaHHOb95duPj16cZ9x5FBgpu9gm4doF8sJsubG+XB
FAMNfM8cdtYTVM3BAVYpGFl6nCqIUOFv0O1WOr1cH7G0FicmZkqBn09W2sQ52RVcI6gL8RkRsqXv
hU6nZcOpUgy9hs9Jprs8dlMjCFDjTuSbZQyIqAcqp3f87Tc9JGPuD8Oh8bu2JuiYUE1LbA5mKx1j
gO9kr/jiFH1Wd+858zaiGlhJ3cqV0XMyd0QtZUgcd0XMk4Oy4U3gZdkwXsmaWcu/GIE2gE2yQowQ
F2FUlMNB6+74wvFnFRnanc08TcsjVRwBRwi6TEBLEsZ9f2fMs/Eug68xQnVERGFD2EcWc9aJdI7r
0UqhT1vplavZ3hVJwgTeSzPsV/GkPcKHkHO5YblP/8qve7W9WuJ0xX8Buh8SzEZr1xy/STeTmyP/
G2s1tIVGnDpCchbPl7wrsj5RSswMUKiT8unPfhjiJzhjAJcLEDIICkiWfvhCvqqkU/r5QxkCWBMb
5Mx1VbkTZBkfQRSaqMARIcHgxmcFk8CQaHqE7ZGnoOD3P/2tEflb6mo1AC8G7nirgDebvwF2+tTS
u+FgfKp8HA9VwMY2zBBZJIUF9jmkfo7XuC8Kf5iLui+BwV2Fm5sRhTD7wjLvvwz21DO5vX/2Yr0P
XpRk2gZGNu94r3SXzSItkbzUuYZC1XjLDrMkS928gUdmV4EoL5ei6Q1SAqyj+ZKm+gIvyGfvmQT6
S86h19syiFyQZUtdWRkF0OBh9j+zJoqwWqS+1XdRAsRlnYB+2SlfF0p9mFl5RKP/UM+CO7t117VC
4rpkeE9to6ASPFEhUY59nqWOjF3iUleHfcNi2qO+lgx3Gmzcph8sruOpkXhoVzNhtTeBrgw4/los
dcSHDRe2nOXl7CvXBoalt5cRAR9d93Hy8QdwEoRyDoifV2g+NAMR/RIDh5ZfvG09X9pQC8zspeus
LOm+fQOynFfoyxhT2yIqOh1oXk2NrpRR8OxIRhBMVSQV0gf1C2JEPcf6GkGrdAKN9BocD5s3ZUfg
N2SWgduxrPYvoyyAdWfWa9Mrn1BEx5iIIu6VgNVkggEl1mVhvMgRBHmbyFqghBCEwN1pfEOak2oO
dk1sKRoqCSOpeJZ0YuF2wFqQRE62k93B0Ssa961zCCOiu94cTYufZ9HCOLEgY9P8PtY6I/EhHAaq
isTlumMU1KBIbnwrewhfLaY4Pi/iiFsfE8gmXNGXyuka7TRv2tnm/ShdYSo64OsT5m5jQN6lZ7Zd
y/uJmTFWo54MQDt8y0tgi3AAoQXgmOhDXDx3Cyef480cUcchS6DJdWGtnJvVmkfw5dHO1Lk5D+Ff
QSg3eFzzdGRfX1r7+XsOy1CiB6akyk4R5sLy+p1bnaiqTEG5ONrugLdzGr2j/lkXsMALXWkGwwVt
s9DKn1UFAZJiF5Vrhkq0qqCVqlHIl+mlIAolhDKHcsygiTbKT9pa9skGzxQAO1REMh/07sW3E7p8
DycX8cb2bFEllGi2yq394+8AetwCL2cA44YEZLqVhZpMGiquZ4Q/iBsgKlzZcLcU0qKZG5/s78Rp
bhzoJiG88UDnrsGCZAjX7DoJcYsY/Pbgywug4CkH4oLhQOXxGHxU6kThiPALMEJQbRCd4zyQ4T9G
eTS0Y5TDv6suh3pguwHoBpc/AVWc1ckh30e1U6gmC0sD4EgHJnpOORcZoZaK2OBjvRlZ6Hk6aBD9
ZC2UZ0j1VTKlHQB00h2pw7hZsE1Odibg1Y521NqSGKEFiCGDXFkUptcMrLMhOOsiPWpN3nGlFKN3
GC+JFo47yLOcNCKXEAeahuMU8YvkysDbUL7eUl68Sk+Jx+UuHImS7tSlYRRdgKsbIXCOI8G4S77V
XpUsMUHgaZGow64vow388BLVF11gbjozyi33/DwPnL18zuNsHcM21xb7V0yxaEkeWbPnnhJGmF9q
VTKQqcYGZ4nQaHAapZBdfnun6/t0IluEnVqQYoIphNTwgc+1mrWFi9Oxb2WIeDoPx/yFGtOrPC1P
QBtYP3XKdp1qqlg3qrt8PXSJVaiIy0O49ax/TKNnE6ykrk0mOTRg6veIWw/hKkrUPjAeADGP/Y1I
bq40iMsdm+Y5aXLo8AEObkJOulIuTEh1t28yorUvpnb//f3rPP4P7y0hCKLLW6WCOhVQcTrl+zhS
W3AgjP/XceOWZ87X6tZYfPvYqPxMTkEkDjsyBBNjivLsl0PNROaIP5j0HVOabcvWEJbyjfZIRjcw
1CEuoRLSCKrua83Bw4UFc/YgjqnUN0he6KdjHd8ZFd1UALD+JX96ilRZTSUhE6CVYnidd5klD5zy
4QCXAu5l0SHuYyLI6LQ/AKQvv4X/plNyFIpEPnNICewaECcWXjGtiTdqTFbSEku7l0xRall1Q6qR
cEs7OfOqEYCNdZvYPTLZpM/TQVT+nxUL2JkMF6G8MC7NyEG1dRutPH6NNfn8tOhSQ/1tlXH3B3Dk
oUYU0x7UAqwWDwvtX4y21HU66y1GpHq22oWp9TDSNxc404dbbLaVOgt8Xzz1qxAbyt5cuoScVW4d
YtZyvslKlDlR9imsIPzNLAHC2UDHMfFFNk6Dz30rs3qrwaiQuEANSZT/AJjP5hLGG6tr1U2qkTaI
Igu/miywN2nas82Mv6Eddr0guOzNbbuBvEpA16iIUYy/xbgwxA7kILTqJRjlFPghe7DxBfGUTojO
Kpm05EF5wtDPSWUQ9GJRN86DUD3/SJrq04DXXdxG9qRdGebIa3S8Mn/vRsuZ5xMgMt1UmX/XSq5Q
Fn4CXrwTPkvB4wPXF1q9hyxCyOdDIKYiEcivEsLFqabZ9IshGBmmnGRr9ITdrqMMgVWtRQZ5VaHS
junvaPRnype5IbjsuFle8Gbri1T51Zcwf4Zvr2knVEy/m+hDCqoCM1Ag1cKLMGV5EDNVmc7F+qpc
nZMxiZVBW8j5Oe6cN3G58mGPGvaaUbqInR6cvJCbYSy/tVVJcY3rqDvrNXKXMZbNGvwkWBnO2bfE
DVq4YhElJ4XbT4Wzv9w5GsGGpvtU6ajRyYVExVKEL8zHwbr3aSSh9F8jqJZIsIRdXTkJxTdkeAEu
EWELZvcXTd/vR7Wkm7O7l6a7tUkbQ4r8aBX+o721JhsOaKdu7iklLR/2953m8L26BvgW+V9VkXi7
DuURwOvC2r/K0lzrVEbqjgqFBXtUFR3EVTdg6mkTgVtSuSO2ofs/bZtYz/8ANXzBTDMcHuHeEYRI
3qNLuNob7fCbla4G8ZJ9BOLduoBJhUgPoQBWlhNn6PcnuvGDDF/Y8uCJcvrvIJKQ9Vl+UwgXQFLH
Vis5lNwzCpCuFTI2qs1qwasPuZWD+8Hx0lf0FFZPf67dVls6h1mOqsGd2WRub5fpb35XiYOVTEJU
CRVicrQQPa+lyOxz33qzyACDJUXIuVUHFj2fMlz1V/OOS1EgHDS8V08O21IklWGPHNw6hRnA+tzn
7c331cNigYryXtAKvQaVnKOnbhstYPlGxyNGvK45jyuW8r3IaQGJvf6mrISRh3TGTPgP5slG0xpm
pE+55pb8vKWD72GyIeEYC6uOroJ+oa1GyHt0qWz6YmK/LQlgRvrKUj7nz40k528hJkzJT2ZfoP0y
4xCTKAsgS2twhsbAPjqaFY1NfLpsqY6bFXfdhYeON5ucWQSjwjoacr9oKk/PratHwcIqZOCRwGfY
qxbQrjwxeHV0AvhceGd063diamYH6zCTeOcCA5XT2mJW1G4FEsgGhjl2MrCtI4V0nlK9Iehsw7wS
AR1qe5dONGwmxax4oyHW1kDSnD8AXOL9L9b+5eh4IWEbp6NgWKN7BW0B1lqumD3BiX+yOYdJKWQD
fbC8hw7ICMnRDY5UVdnCD1JyMfHVIkOsVlSLB6guJ9BrUY+AHX5p5WmTrrW7g9Eo0QI1m1SRGaFC
g2CA50xXRUB9gipQ0Uxnqb0JEiV3R4m1g5VHjyGA1MslUuKUTvTkyzbEAAcK/A/N65NjFBPkO85d
rgXOUcCPqLItm5pW7unGK096U5NmgmIWsPnZn6STEMjyEtfXlfy0pWj9P27NQCRJgZYJCOiezzjk
W3trm0c0AMjgMh4FyOhS/sKfzBvbgG8pOefx8cdxhGHk+YVkLrVYLXD6maBK1Y/4uM1Djo8oluiD
L+QULOmiVRpArWJZOdBViowwFx5wk0aHphzvTMySAX9EQCwb11EVSshDMtG4zHj0aTzG2QRIVpv3
IE8p3GhsvNB9C3RclxidtW4HEc0N2KVezzatvJECYyG6i07sypaGx+DMCLqWrF8fP/gO2GHIlHas
Pr5252ESNrmpujSCZOYZTZ4Wb6C3oqUR9n9QazEmC+tg5fgI21tpBbHJIuSq4QQyKijEoU51d8ie
Q+0A89bfwIaZAlo96Bsc0zl6DO6zvlNHDPiNGXtOJ9jLWsYjaZ0yBJ6jeCSDZ+/Ej7MBNWIStsSo
KWfdGKUOjfimZloFrWOkGFwjU2KDyLL8S53h7UwZVPxNLAzBUEE3gA/NMTHw1Va2yljxHTRYRu1d
h+d4a8b4PtWV0Olh6JntETjJFZWwkKUXGwdFdvyY59KifVVl4VavIgxpN/P7gYLS4i1P3fYOV5fD
loF/MUyIugILcLGDp+AJ04QrET/D7t+GNVN2JLXHHbJ2PLZuomwgW0TanFJgWibwAuj4Veasx5B0
yWnupsrAZ4be+mwTqTRXlKL+cnZJ1TJKQjN4oiysuRudPBZ5aHpoR4TATjvRS40Ew3hvGvq+ZysI
s665zct0C43R9/MiS31FiuvBMaNBb56Wk/dVSG4v1/QonF8+5BAbQYOTUebDM0J38Zx1GVzNmTXM
/+dQzpSlTrnz/DCITV2QQEXoxd7la93EwaZDzGyAeEz+uifm8hNZ269DfJUWv3oC7qp1QJt7qqe1
Y7AMmyfdp9jRfurhVaUz7i5qnC/UCPfzOPvMXDdV7x216VT5NfrAgzUvnbHyLXHDT9GAUh2ZGN4p
dBQWuSICulwNMnHFFG/+dN+0WwjT7bWpe5zhqOVDBfmCmCEz/48FVJNIR4ZqD0GHUqH1v/nRe2hW
RTV9yk9nncokdNLBbAAb9hvJTX8+FxY89gwV4E0qQLGoez3XU1UFt9CIpPr8PaToszOgWTkD1XgL
uL6NFfX12cdb8LJXn8wJ4dk7VkxZwbSPb6AC1ZBrAxyTiuaH7xuFAHcsFFpX3Qg7hXp9izhMDpcH
2XnF9e1DGfLysTevYfpyhcmLQOrQmTLxu/Y9rAs5dVaOQ2IQ7eZakowmHQgniqdUR/YYov/+Qx0s
BSYz3uLWfA8q4DmJsjlgm8/h+1rttY4c465LS8ILjLFF2TcpOAhnu+KW+PHeBcNE2sV9LN8WGCAW
fbCnJhMzzjRQMAA+defsjtsigHsOmvLPdsP0GACokuoMOCu8/0k9ldM8lp8dBH4AUKpNfA1T/jrJ
e+QHJW4IDg7wbqIWXZIMWid+BaPuPg/USzaUH1IEh7iklHj0/g5hCebxTmqkTjYV5c8CkAFBtXJH
lxFaSqYCrO1s2cczcd1TZtUagGyFla/9uhFKuAwcZLCSjt+oQQsafG8i/zaJxFT86eiuMajhqUiQ
VjwjBEDyXsTA6hZdej7wYDotZR73ALTR4c4HnjcsEyEp0g3HyGWYFvhETQqGVbHxzQYatayt9WpM
mPB2ospmxWu5qW4mIkVWZxAhtjL0cloGKUw0w0G1G8V1AovW2wyQc0GaASKCK2k3uSQCtqPhBFrz
kfSkIfAn++pChLPajwhUWQRKtm8MgHmVqhw+acuYHrWynHmfKGlfLv3behicR/c6yv3AWXN+WGYF
jsQONvsGyXymzimbiIhHzqE+3e00tPyIa5H8cwWWwfjVBsvq4sB19W3mAj+DhImCWK0UfsSBySW8
H3NBhfiEvrneDxfpNThupPbRak6bAyzytHf54YxtCi903oG1Kc8AUMIMiCz10ckHuZDk1jplcGMu
RImNtC3Ri/Bkc7NGBsl8nms2wd6YsHD5YqSZcGTa6Y0CyRHxVLShtdoyUnE4OX5UzOsvSNEmBM5s
eeTFxdfrViN8GUQkrfvoirJXAYv/JoTro0DEVTuf24SIHmUA6DGiM2VCZMmTsLWYRSBvDgO+UPZW
OdPZYpLeBtQuj7LUO+RhxmpAA7MgUiX5ka2nN20lsSsxqBW2e2VNXo4mK2lh01gFvEhZ2eLHazy1
atw6HzBoQdVW+PAq3dCZWyxKZldJcaLBDFFIaEVNICDfmEAMQ8QGIBOUrYivzZ37qjSaoGjH4Nlr
TCFqZZh4H64iZ2aH7kRRqZKsbltbllWHNlq974rndAfEO2guVN3QsLwjW73PkdP5fQKEIbkIeoU5
n4C0lFr2KlJdwMRDFLSK37SUff+gKTWcIKbX965XbEkixpws/LiHuKbclfzcFtYA6tjOJp4Gsz7p
WfnLkMVaJIps4zG2nTlPZMKg+HzqXWTZF0PFZRCqn5TufqPmwgwMQlmbgfScCLnankqwp3owAgzd
sjXwqFwymEsieMxH/+QY8CgePrjRclCGCM+N8rO4bTNXoKPiSIWdV6Y0ZhPSWojFbc8FMk/XbVNx
rur26iIrdb+Uz6e71cpFfwxw1WdLVMdrVPrMuE6IWV8BPRhHZq213KJNcJZaTD/6lG8n4/5y8n3d
1dAyC1yK8lbnlshFQLsurJHNFKWlijhArNoS+VA5XBDKcAQsYYZAHrQutIWNVtbKXR+cS+Mx3koO
9IYTrCGdk+5ygU9w8cRjQmlJOj8bWdZ5RNDTF8Bzi9GfkV/H/SYJcccZYVd5aSAsvOxPhUlMHeam
buPe8yeICJczT6CdK94vGAwGm7VbFDs02+Ha7TM4VK84+GiGs0kmL28zKOlvy8U5KOCKKdh1KErG
bIg9egkCnKtwCnJS/Q3tbhjZB0y8CitGV4YXVRt19njAobFJ83GZtN+R9jArEa2AZcFJlgZTCXow
hFRLHolqeTAeXnqs5oRUkg75XKD/zesPY+CESCBDHzYVEbf+y8t/px8dzpJ1JLKGQ30fivUc/VlJ
GY/GDvgoKg6U9RLqKcfYfEB27CdgDc0jwcty6rJf4PZOf4vZXPFymoC2Q+rL4OXVOEu/r4OPHRAF
okYDcKapDcEzt2EW5SBIhHrXmoHlhnWZsLkntmvQxmmaS7B26Y5UuDHMz5VBy4DHcT9P15uQSdQH
RhUm+C0wcofO2jKW/XcJOZiTvW4B0IF84Yhm096SJ/lqS9oc3Zij/wZlvF+B2eLuCYj0A4deAcp4
y2hFZ8Sn0VIQsiZXbuh26/j+b1zSsDmCiKTBCkM0zY/M8jZe9xInk52M1KbC+KYlRlAsHd1YEfYi
o5W5BdqvIz+LthweuRsBDS9pI7samSaHCAo2/KAvhecBtbSLppMMwgOFswFm3XBbTFk95qYlJLuM
53l9zpzuryyS1KaD1jIdoRWqrLaXjHTtNCIO12pMUgcgfwFx0+eTtpdIGVRTBZHyEOs1byepZGzO
FDZ2I4OMY89ihUG9sDZbfl6VOCMlm6hw5MStw7g1e/A4y5iZI4xUV8QVo2lFkCX//bQTIbBSgRNv
O5wTvbPovYVlwuuEwFcabfUjjBGjQ1i8n4DwkVb3UAnbU+2tpA9/lV3Iiid281v5mZJNhAbk+FG4
fTmq+B+V5JcV67D0UiuPY6yqPvVnzHD0Hj/GfOMjBTIoSNNhI9MSvdFBrONuZ5HXq0TOgox/wdH7
3HBR+sFRxzV60xaXyjq4tHaR8yhagxFJ5zX3yleVuPayLL+Du3sIGxENgIvb7AZ3YfBXzuO3LV5l
w5TJN0aGmsL+9/t1dqgF/4f4n/dhGh1Jyj4K0pehIEPcmFLyUTSJfTV+C4domux8Cvl0Xw4UpH80
FQuGAbSPmt42C0XMYPNwFUKLfw2TZPo4WJuuOJBoJ6y3lKPpanc4KAKEQFv0tZx5UpSOoDKUe2Ls
L8Hjsasyx/sXHXzf9BPnkTFswhzZcxs7e6zyfQp57qQxzxah55r5bfiiXuierGvnNKZPgHnV3P+W
MeZtSDk41fjsGHamYFWmUQHxnqSJUQ07V+l6Op9ro8wNa8+609au80u3LP4OwimMg8ygHgqo2Nhf
+wPcDkx6RnQb+PIGQy2VmDC7bhz/qfCN0Iq6gA58fTwkHDi8kQ9POV36GEtFNp9Etstp0xyYWU7E
/HbgO4Gl/p0tXX7a9uYZN9hLXPjkUnB3EeOaUGukL4tvcdue9g1FVF6k+VG3KaABljhnvZZMgrEJ
XrUPjY4yWxVz4TqDUx0dhtBNq0io1nnYuts98DX0zTwQ63yiGdoU79L29H0YkxmAcbgRYYO58yPt
prdJBRZpmrjgzqbk7bsF/ad8jXYucM9pmCvGnDPesBNf5YdKRA6arIMf9d8yJh9+5hih4Pp2m/da
tU4bKJTtExJ2ak2H/zBAFJYc+oAL8tJQFBw2ZLgquDmkW6ykU07uS6KQzBlnCInBo3kTR45jFOG4
fLpiFcRXfHYmIbZBwJNdtMqzi0/X5ghwAh3Udt7Ea6ZuO3JCQpUSl+q2O7v6euXE7uhBPJYZk0FI
xuXuOxV2WBRB6Rsp3c2d+Cu7TVTE5Q6Kz/Pc+lXzAw9adl1nBkWmP8leInVVVDE9fNdI9LQzjuYp
9kNZYLGti0oMQebkfYo5W6Ehx9K9HUeWxnUl7JfRC+alLhQDHo3Eo/z2biI18BfHcMKty16I+RGP
b6CEsIv3WIf0BxqQKKJsDSYLxzJTuGaxnSVMGy9OJRQPem+xK8F9/vtK99/qvRTwHYIeR8H/1yLM
8mj9xBsuK7c1usnW/JYgBVie186fzXjd43O7y/F4tjapICgwdAmV4gTkCJ5C9Q14Rsiy7XJ6llrE
1ffHCVq3Vq5XT93RBDmt7zRBsdGcoNfl1JuOXwTJgB7jMnxDghjIDKynqc0Cm3lGT99WuWXqD1zo
Hb7jiMTNvfdOEniX0dHXNdr85y8DGxK4EkJ2mWFVysGWq3vqB994L1YspuGI5RcckZayWNu58Nnj
ODGKmziWQmA5J/Y7lnGnaT19/MxnX1wh3WH64s3BGBkqcZ7umNd7JiIsxpiESIbfHMRwtG+JSP4v
Vn8b3dv2uuX1KXU2EOs9ZENtRDrk15E2C5kQZdqkTdsc1LLXKZS7DzKvIaPzcm6vx5baoHMYGMpX
1QgNMam+qNEDe5X05f++wDu6Cvy1J0hny+6oyVUY0Zi2OsbmdxQDBJQDu8uqN7Zid1eqyMS7tKIv
c9r+Wp0cyXH2t5XlfoQsAIojuf5LGDEoaKcbzFJoSTXk+OrpV4rVKIMLaqrxXz/Iy6wEh7lbt0HO
2NWumKWnOCjEbWklU/AKoBp8rvhVu3DfQdDQTK5dX3MYRFZZJ6yh+EU2rgloUNrnCieMeB/LPLq1
XCcvlxX5nfsYpa5OCU+iK7N+TeKRSDruTD8cy1dKPY3HX/AnljbcyVhvPypNCD4wGJecfGbbLmr4
JuEOFPaUjtbWD/SHtojQ2R5HcNFcBre+j0QVHhIB53KlwAwrBj7oSIbqCg3YQxQQltxN17BxSDzr
k3cBnaSAtsfkyBjKvMEg0dHTfpCCsrI9VaIl5HHg36mzo0BfXWF/ld9w2vg7589KNMnniVMp0ri9
7SpmVbyvMaj7xYuBGNtAHkENxUNXFRvNFkHa/GyaDdZYMYhGW/rFoHBh1s3nojifk2pL45W5vW5T
Jyn0R/pXAUEVA5XwssIiVuuVyYyhgB4Fap7eiufqQcS/PAQaxWOVMnu3Rt5kCp9Jsu2FCwzkuuH6
THHQPyr2XzKbPXsmhGuH1EGhgrpnXeO1OQyLw6yL52hX0NZgdQNf94T4hP/qgf6AFWCRfWMXzkz/
fuQwzd3B/mzXq8gSEpjUXUBhL0DoLRT4rQoXC/DqNjRi+fT+2mFeXKzRD4VF+Ipy+x+2vqfK7x++
3N98oojMDN1pd0Fn5uWm9GYl7tH/9dGHiI9Pjs2w33YVIBHebCdUU4G0UdDcKgst0N3+aQ5sLP2P
Y6rbTuPSdanAztKHRpA0NfQcTF8xy3cP53ECobEXtNzAV3nsvpj06AsfN+muejRH4vH7WxI5RqRX
QNMXi5g6rrA5dk9tDtMXjUNT3rP3t1w9XfpJCBOoikfiJRzUGopGwDA0gPrWhqgXBSeK8skCR0ih
coonszxCC0fIyE7RUVkMhOa8Y0PdP8xrR26I+BcTDfVl5j3hbmHDkThF3oT0zz+JmthbbDnoPqQH
YoS/IVOLTfaaDxTPiGFdoDbl4AvpsZQ+9aEidojA62CRY88OkYiarojTpuWk+TpZ043LT1xBhWlJ
G4ZXX4jJ8kPs59jWMkA2br/irdvs8KKk1J0dVW3innUpyEsme1A3xb71HrZlpdgJZevbAOvGmlpX
3pO1PHHrmJb7KMDYSJckvc5Xv0g63hDvvVlJwHboHulssCWmpNkVCsjJLlvvvEZSoQJItAITtZJY
JHa++Bt5LaBkiI4As84ut73JuUoag3lFbb1TE+zph4D2tTwPqBkDF+7heAJiSzi9QCFMsW1a8z1z
YISDs7QOV2VOfE42aKe5PtjVuaYHmMlgFzZBmHD9pZeD/r38Pa5C7G/nH5FwJ2iUNN7VyMtYmbzw
1hMnGn0olVbljI1ozZuaoGOg5lbKxiCEtjKw7Q0n5NB0fP4sTkyfRoUK2E8VvsUx1n+fvvBD4Um1
Kk5M/VRM15mRCmc0K28qBEzRQYISi8y4blpbD9i2wOWpbjzBN1/Cun7cFUfVJNyhz/69YmEjnVzT
jtjWX8KcE6laCMDTPkWmNggLG7nqeoUapE1a8HJsAcU56ZUVdVu2qhSbBK/8Zl0o1d5tyWbEFzhP
ED0OIZQsxzw3R1XLQRQWeXjbCYgT/QpHaG4HXvB3h3L352jDvmcqdBlWJh14ZVnoDa02kTG78EEZ
2kdOD3UCfKqylmjSmnckjgB+iXASNf9oz8WRv31bCrAesGPAPveLNjIUmTFM3pQ662KqXenxw/hh
Q/uyZsl3TRFwFFJgSPomsDQERmS/F9Qw/lvt/AotzZ4zJ4k06TFz1wQVMooma8jDl4iD/s6U3kBz
QreUZpJxIOnmNZbyFwG2FaTiAjoIkeOy94a+HlqMMGfpKaCQf6wHoBxqTxsycZRfzumAcHZfH1j0
TCVgX09FuE7Jr/4RFXIJfKfO+isHw2vYfekMMAVhHP334aNS9GEqOgXCixhi6oU9IpYnCsziP5dL
TtiAJTFMZ6eVeiT24TdXTHs8nbPSxUmzpd/t8Hjb38bOAlYOHk+4TmS/GsqJghe/gnLQv9jjC2Bb
+VxqlCKob+x6AzLbbX3QP1Pns/yRHiz1UDaDqMq1RaLFYOHcKxQr1Ix+Oh7dQ36DGstS1l0MSpE6
nMTBnRe0R2wVVKbUxV5cRDHcrIu2pDbvyvNgBury4W+JLFRPB73W/TlMxxxd1Cad2Ew/2x6F/ls8
o6y1qLMb7IgafioOAceMBAyYv2gplGr4NOtAecByOJObpH91mzBDK2BpJs9G2bksNSdkNVj5XJiV
d6sUCMKVxNpDn6imj5tplfkCZrN5Grg+yEI77e11SrpzFBrxf+V+Cq96hkMgQnVVwN5qJqVcsU1L
nGJkAssYGXUVSxbd3mzKKHVLpGrTKEAETfqhUTVb3fDL0h+aOlip8lZGt6rpoCtJJFK54Jr87u3N
eLJU8he+/xp+sL/UFBGIe5l1fGUOwlA5syebRGL8Qn8ToyEQzIYE570EsKZcgbrDGcwrCHAODtqY
lABrbUabVNBjF3ZOz4y4CWNub01BhyqyIChbnx60CcDFfGJFY6/JCJejvTIGDMcHPyy2e8JrDoZu
WM7RNzHtwaccYFqEv0jirlKDVajhS3hg2egef7LjUTEoflsbb1jeuCRYxWrBY1DRCkBPmCV8tTdR
bMMljkzVceDZ8HGH3MF7y4pTewVVlqrbWCbxuj+BON8rbwDQU0iWrNL0yYaq7WnPBiKHlSvJCQF7
8hdwBiBcGx5ZvFKC+N08ZPcena39QNF5xGAWDWCWEMatAdKNplGMquWL973aaCu5TM61ijh066RB
Pp/ciYyikBB6Au3iNbZUlJbI/IqkAu+1reJxfm4K/sRWhkbjiCFzK9DeoCo7CrttLbDBwWkVAX6H
ap6UtxcZkoHABc/k9IKGagBgKHyZOZrRGwCfPLOWDv0kxcx0SN3GEZEZYKkuN2v4JAqK0osL/WYX
ZFyLxUYMWjYQQDWUhI4ppo/wIyK7Ttn/8xC1jh9ilZCUcBF1ZZNeiv5TGzM9D2YWvIYjdiZbQ7Uj
b89gTWqlBY0cx6B5wKU8Afr1SkSweqL5pHtSIpaUSQNorAKZwB4JIVemuc/tLSHxqKo8F9g6edxv
4U1yH4rZsMzMz5YNk8/ne4nlutAI7JiKylAXUy7tRRNNvoEWDSfLhZZKK6zqoXqSfZJbv+YjUkBL
IBkcNpnHSrBOmOgcTNpVJLRR8H3t3rARl5PksWCQ0phL1EBwi4tHuKOt9f6YDV/rl8irYuxb3/n6
5rs1UfRi0adhjlRN0E+hDMxSBOY0Ol5nilD6Q5X4CUXFhAwVzLOdFeN9qaplag9e/SpsdDeI9yyD
BjcKl/rCXLRRrBts1BTbuSLbvaudFKI/OX/3CZN8XJmqpqqsgWz9uqApG9KCxL4mmW6+Gyx2sUu/
5dfgk2oDVD8JwHfBmM9iHTH23TAtWjWjSNqPZFEBQrB7U9xP3thiL8ICOwDMtdJfIUwKsgtSmPI6
U+o+oXqh0ceT9IjTx0uiflY9Qptd1kj6H3Nn2w+EwWKJ8CrKZ24HeDE5FACF9hjypv7XvoGTn7bB
VdRAS9WZCpR2Uf+Hns839KBY6mQ0XeE6+hogZURQeqr+CPtJr9NVqSD+OMuGTKS0H/RbbdVTQWaH
C+/ValZOIYvtgEz8oF1Qg6r+uXrXXyaZ8gcg5cR4DuEBQpp4ttfBTOWJyG5TDYtpeVODgw3PTTOP
tufHfjU1I/PSgpNk5nMZCejJ3SZBYG/kBPyE7Pi08cZLF2TlY506aLmQOJDRk78wgNYxiS8kqwZ2
Yjv6kgAyDCUDO1SVwFmddZz8N7Nwvus9+3pXaBijYHBElNs9NnX8t0IW4HInS+Va1koJIgTJwF7E
Y1A2Bwo9pGWJwLTdZ46oFp3nZ0jxMTO2g/5kpgzFagWCwSp6D1KL9ENu3DQcYM5OPwL5vcFNMBoW
nKYLevJzXNXCuNtr8o0qMCw5Z3PpK2UXIGP8y+2kPQD2yGaE1xef0y63Nam3RtnvNarVwYYrXsdo
AWNPIQ31GIaHiDqo2IuDQiwCbfjFzZvXiqhJRiHFQWADvnhmYb2LNGnFkvn4vtccaQWE8BsUBbkY
G2mn9aVQK9bVhOZ67Ty42RxZTsi9/kGKigM0csiIwry7FDjGXayb7xc9Gj1MVRkXKh41dWV20+7l
LrrSFPU4s6q1lxQdsd54Gw8/Y1LPipxf/f7Py3wYkaYZ7/ugkjOZCRp1yH+AzBPvn15kh7ofyS0B
yAYZKghAxJjoIxDyG0D0j5+cuB4t4BMIA1czGGspapQH/K+hgkesMUU/tu3dPdE5211dtBt+C5ko
1kzg95qxu0Trsv6MI53fYvH3Tg5cSbkvJy5Ax5rlzWP9Alqq3sCZdrZRQ0bhVZkmuUunEjpYmG23
gWzm/GQIi3v/Meo0HYHvaMRUNu6iTN+vXEn02lsn+CrCcDmw2g1gqPTayyieGN/zo0c9HHnR30KJ
lhJxkItVnUROzyJccLDdTuqWRI0uLftSPmIiG9ckl8N6UZmN3As1aLnw4QeYJAl8I+iqbPiKcJdI
3TPYS5CQAPfmc72qzQNNFXzOpdfPFtxa0cH/3e2sOby+SeijXniGqWA6UEakIzOmn/8rhAASGFJT
Dp9RNEmTd/LaycFt5JXHPaDZAVzQ1Fu62lB4kYpgqzlauopg9po1QPxAxU/+PjwiOkktDBr7XGqA
+sUyCTeogeex80NfbzGFxpx4DchtppD0xc6qZwBdBaEVaRPafzVr5htmOi4M1UvUaV1ZFArW5VEI
XVsMd7mfqdbjQ1XLbHPbpdFP9htrMqrM3dzSvFOPxIb+rNb0aXoFQ+PiczncIJL1LV3VEwPWor8w
agaGz5BoBXiDj1JYneXAm0HXQwtSawdecDCxZ41tDIh+pEU146McIwbcjt3e6kZ9oV6Ky0+mQcOF
iu1lgtk6GFi3JX8iER+RijVRb+A8QsfK68cPSUbZ8F6SS1BE0fLu3KZvTypZexXeTbzAZtmv0fe5
qRGSxNoDlpMGDDwXz1D2sk1ZyRoqZnn3BxJmgwm1nOqoPoa3GsN6bI44MqBXE+MAyyzgLGEU74Nd
tg70/VIze6LKQ9rKGZicaaVQSObuvmlM18nkIYVvv95ypQ6p86N1D4j3BG+HviRpJ3Qkbiy2lwe9
2o4poKajxtSXy2IXHPjz5V1VocvWZUUVTqs6QAjEvsY3lQuirqAutkMJ1F4S6EK+uE6R8owu++tC
b/gXDTv6NJL3NgbZELYJQvhEG2+RRPBb8DrnshEywLWWlphH/3cos2B9jCAoWLQ7wiluN3VCJRc4
rzOOMEFzTDfDRBc+gq1Nkns4g0ruP7YQksRFIsdWmx6e6oVWPrw3vNjX29/Q3kXqTJX+eHHNXTGc
a1oQ/bm6qJ/8Vbyh0BH2B+ZZ57m9cLryEBre94rbRdHW3rMJi3cKMK6h01vcjN+SN7eVonbYfstN
bldWMGtGasnj5lE0mFVEUcHYMSpHPe8lvKB153Amwzyp7YHSTH3lv7JYsMsvcm2heTYWzDzYKDSh
nsBc5u9RvbqWI9e/t8rVXDBWF6O/9qP7Z8LKsk/Wi8qx3aIVY+MZLKC/k3hS2Ur5q8n/f9HW996f
Ge3NX4t5kZyxsqtm295q0CPUrVjNoRCkdVWstas4vapPygl686oJ3Whuq26AN/vwRR2Pz9yE8bqd
kcmORh4K3EPT1TYm3wfiVaXzA/exAHPgPuiapaHpAxpdGB5MmxEWGHynCZwwA88D4tx6dHqLV+dd
rUgEX/xvOw/KHsYOgXsMNhhX9+MuJ86ybhfAofU/tfddaJBxLQo8kn+Ar6w8KqxmgJpipDNbvNFv
72zW4xE1bEueL2OY4+w8Mtrw00vZCzkMQOKUx4XYId4oc6KevYUcrcbvMstVwdu51MFRei8pea4T
cs7HkOnW9s5XgWRWh8qq7JL3CGetxgF1vp97BirS5rOgXmu1ep6GKHlbHB1wYwT0adfTug3hzrkS
AkyVarJGBXMVtYrXj9FEQGBqE67fLPid6ArdCmE4FE1a2NoQ2U+ccE/wLbdi3H7d0DbApOy+XXOm
I6ZaFqKeaTN1Itt1Seje+G7un9HLgtyPQpstSwmFFiQz27/rtY065zxNjbXU+kECv9AbWPwceRwF
7SKD/OqtB/qbQ7awr9Wb2+Rs3U/dR9bRSyj+DTd9Kd2yiS+0YX/dXD0RIRRrDqRiPCxyeihvPOv7
HLtmgFbXERNKyyPe3pqdv7jZXIjPS7Boc3cVppG8mfiEvANjEH86KhFt25HkuS6Y+Tm7AwEwecoa
QqeNdb1AAbC88QpgEgAtAfOENabi6dJ8jgGSE/4VzwvpGEOznKS7NLUkiaZx5YixyF4hCECV/tqj
BFmWuv4YL/PCuSz8wfrTrobcWOGuq95pS06onNAI0mcVklR2rVMCL6pKlmPSeqyR7iwqlOOF1Gnz
DZB4JypI/Nq1jmfqwWIhQ+ZPl3yPHi8rzONsbpPb8C4/hW+Eqp+Mr3Gh0XLbfypKj0/oy0btg0V0
Dk3iZbOQJUcPvKz+eHbyBG5zwlfZGuimehKG9vK0IehdZ/vxwTzOdvAcgrDZPJ74a+x1z3g7ZOTx
2KkiMpFwZpE0VsX6Z5myBkuw5rJI2W4W/K6DANuhBAhVxZxYWgvSQQ48MEDPGKTLIPwJZljomAsZ
TGhab5h+GFd4vIs/xUJRYgd/TwYOTtMmHmN8bada3mIQaZTN/nFhDsimWMUy1s+eJfxsIZOWd8x3
xuXLDpjRnXiwtDP3+xeVcwtB/AQXn1Y+0JgKqsv0sFE7FRmG1wB/FqF7ThwehcIfvbJ90qOgfzJH
QajmEkZzC7UN8WaeThDykj8mrj6iPNeh9zvDayxZC3Kn7jZ04UAWgdoSgJYcPHprkfhi+N3kATVW
KDOB2Fv6qPz9b2Dn/0GKRKyzDkto31TD5wvDyWEGm++1QPRvikXU8F+vokslt0nzq/3NN1INvjjn
8y1TFsMrDAi0lnFh+Flfx3ovvCt/psO4c5cmkCO8HP/l5zjIXu3rJPyQ2laXAbqKhVoSnmqvu0L0
3+bzixG96DkBFqCGwJL9Z20oBk/fP58LVTMxVEvlDVCEehRgv8weZNt1670ZLYvtIgDAtjACZPi4
xVr/W2tPV5iDW8ia8J0dThSc3ew2IyM4uZvxoGi2wqiUY0f8dgyn/PZQ5K9JwU+U+VJHTZ8a3cpN
KHtbE5of2/+FrCdB1COGJQM7m1BXi6xa/A5sdpwMA0uDXoaDDNSssVU3nU4qthHkgZP1uW5DReZp
nR1JckGRs4TeGy7/1Fjkha2WaORtTwfBF7a+FYiUU1NQVczGJjdDj2aZeVCsQfsUGzGkdNfn6YIK
16vNVzoWa+PEojaEDQzsgRzt00f1/wkxDiS1gQ/P5fOw/c6pFFedVHGb0rRcGW2P8X1vlAkiYuhf
7KozZlEidCb5x+1p6PBvQSf74bZYvxT2pgi5bt6PhDvuZ9L6lSyIEE77Tx+Kzf6EuzZDYZwK2pNX
pcpyg0A9ucITVvoW5bLnE4h7yQYwuGIZCO9n9Dg/YRIAw38Dv2tFGBYtPnsHbvvBeZD1w5tSByDI
FhvfPBml77hJ5nzHLQ6Kuo3m9OvavMWT+XC9w0JeJGXse/Kp2JB/6vKMHxa+/sB12gWgjhTBS/PU
WmAYAy5uAhuxAkDQH5c9RgeJXwkCG1SnP+4iIqBgYige5uw+PxndGSfeUH6cDR7vPO1GQmo9ZE3E
znwL9nQKpNq32pKbq9lyrEwAo505xDPIOwpf5pmzTRJK/b0Ca6jyKEl7VlRiLRulqw25WmgAW6YV
BrbRLHDXKVWcZLF3pnHrfF+G2/GZ0/OHUitoBnaBENDyjzNaRkvRFIzbxJJPT1tzwRdkqwZ4Hh2o
Ba9w1PiKz438EMoyNk4dTFt8BTRXTt52g/S8NVSLmbiAp4WXs4M7/uEfxqRK3ZHAf811sijkHneL
ZIxGLX0ssjBbx89r78Gc06HS6N0WEUjIbJR4elUJsp7e5iwUCoX60I6CE9wHl0BCdkHyA0V1dMRw
rgpNJpS5Mydv2UxWH5I4zOyHfLI5sxnEe/ilmQKW4ZVWLPqWwfWFqpkHN8dT/3lprMfSb3PBmzkY
BkGRhLJr9vwnZpKN8f1O2oxoQ/tkGuBae+/hJo8H4xgBc6h1+TiQ4CTPupyVHwAeSUgN0jki9K5H
v7nmZnqoPF4MXZgAei5Wjsz9xNn/SkFNpuiSQa5twEYS4g+Vt4r0AiXtTjOrtdsFM5hArg9VqyHt
rfSNHn65J8pff4MlJk4eT+LYjeu+H1VK0S+b7XHi3ZxIIU8oxi/WZHWKcZ3QGFKw9querGuNDKba
IAVJmq3rqhoV1E9bxNT9rBNV0yz1/FqCm4NAwbkhqQFOIZgMXRPg7MUcsp4wYLY12ePU6QW+Bh9q
c+Eq7bNrY0Rw8Fw9LGdqHDbRTLQiY52UMge+3JgAx3WuE0w0/R7UK990Qojp6DcovOOfx6mMqRDT
ZOpKzV88VthxO7+MnbXIGuTiiSizcLEGGqD1X1N4ug8G6Wp9qrIPEsKYl/FkgVvXWX8ukCbEWixx
cSE465wR/elcdn3o0jD/AyzTWdtgBV3g4y+L82Z0uD6ja6K8fNZQowTN+9KyjpPn6zcD253RTRIT
lACy4w2hldtKhvfxJ4MD86gz4apTOPBAk/yYSINCrxsw91SVsf30RgF700sd9U82iCgEGP7u03eu
ND4SGvsLEgugDrU6qYyuZAuu2qg7OOPKkHP7ybK7pq13O9yBOpto6mO89CNRXbrVcJyh3NTzyAmd
jB/P9P4rhIqKmBs7ia0hWM3QOfb3d3gSvYu75N1JWuG9Tykyvk6G3+jhUl62pHMFPsuDH3BHTGE0
D+m9fGQAyiKnggX+ctZLdTTSDrqAJxNetqUojNChPTvVXsltiWV10S3I5T+w163fEe7CCOdIBUgw
wrLmXJOMS/05xxa+kAhEJhTsBL1DLtTn2MAAYWJiQGulR0nS6odIN/x+QsQ3B/07b5Zl5rRx62Tn
ZQNz4DVP6jaVjG7nMNrQuFyohmkhOenX/6kezZkRNQ9MSGbJ89yOvN47ScNRxuVoFe3aiKV9YoPr
4eS/W88uwVBCc/tvCYRaZc09yU66WQznyzdH7MIiiyMMzFtv/oQk1xxiDjV2mNRNv13M/iEWjour
RV8yrWcHUZExF0SZwNThcHUGYtUh1BbbpqeIZ7s3P9NE1pn3qSXMYO3j47GucVAM2PNDKU+zDuGg
NGiMN1T4fbqZuHBPpuZYOM4ytF7UKYRbDrGUs0e9bVjdAJc+szM72Ks2P7s+Ae30d0FRx6fCXvkh
1MxSC62cz/VPSZDdr2c/hEvi4eC7Hs7AsJN8ES2PHUkjbAgVsj73dscOFHa0M6Dfl6OdpFBrB2oM
ny0o6FLFjlC5vOuhpEgMDfOzjVLd+qOd4h2yqTvEm5bgwtxJ33j6reM6SCApI/ZXP+dtmRJgDFNk
a5FBhYnffx5B9hccNFHtkxFZxsIvumUbYO/gb3Zm+THECqJD0P9nNxzq8jh4807lNaoeLGRAKBpx
TohQiH8eTqynGypaCBHac1WX0f/xv6i1G4/+l4p5wOLvh9DelnEjdLCkpoTAx6/kVFfjsapdmlIC
HiJGucgbWghj667v3FfbaLk6RUimevs6oOyt9ZFKaEQtvko2ZC28mcGNNh7eTz5FjfzFHrzS/j/K
vmZKIvryAs8ULEqeQj3LjwtAo6lO34n4bdK3xwXE5gl1lyMF6RsYeylbxebrlJJkXllv2mGjj13/
dAMnqbJCGxAndxBLraT2MXa3fbKcEnAozC3410LknjBmu1Sxt6mFeK7I2xwb/KEadb4aPTHoJDJL
SlC6nq177oFJse7Srgq2CkBC+YCPqjEyojHOm69XzqmTu4auWt+eKDJlL3BC5YP8XjriyZw9UjQD
erGo+bPTQnJZ41fr4PfM7Wd8ZIIZyX0PPq8ZruVcb1Mpo/Olf9HSlQfElrqM+ZZ5MqILlTzVinXB
isJaie961rK3NLPIXWwPPPSxLLLguydNlg61S2zcIX2jCzaGhW86CarsD0gb/Uqx8RyOUHDfuSWG
Uq68SZIfGWpgu/vsqsdL/zZKcDEDrQHCbx1OYdUEehiUdm+HzXF/nUtLHhUEmRWj599/9B2h39fy
S1ZFX5XOhK8Hh4WJ5qmXrqqwiuC20KdKGAaMLSoUwoOmaHMLQ3I5r86+vbdhwyvkXSinCE3b9xx9
A1eTxhaQbZ1ZSKfbjrdsL5mkA8j0KH1fniQjx+ZS+nHQJ8UJO09sy1SE8MxTXzn971GhzDw8xBBH
Pm5L5DIDV06i2mGrEeDWPjoTDG8O45oPSJc/psrng9J+KlOuk69d/UYoGD7Yrp4B6AQ10xkPwdMD
TIAG75WnsVw7vaR1VrkfFIqOpiBLYI0Xe+YQjmp0E+nMrGY5OS8WvxYLG6bgjgf6wYENXiLN8v+V
zI6g+F8eL0rbJeB067G69wLpv2BfsH8+RXtrhIzQImWpAVOIgI2kMf1OciInzZC1tbYxY93ii1zZ
daO259KqjRujNjlKIYMdqD8mGpaQbzNWXLvmcluu2Rfc+0d3pFXc+UFbjYnyUrhW989LYX2Q9Uvy
QeN2yyFCP9xH8B4KVVEZy3fFMKppO7w26qj4yUXjgZHQ/mChzUSsccPT8KDOPOxG7UZHYG7Lgiis
chgNtkUH+4/GFoEv4XWRK91TAF1thjXjjQYTvOWu/DjVFVMGdxM3Hh1dyratjdfJ0F0APp1P43FX
vbbqfLaDY9N95BW7bksXPHU2CweSHJC3AScxuNBV4mS24iJ2foAb1+knY+qALuGDqSmKSVgu9ry+
bre/N2/VmZ3Eozri8OJKszVjSg0SkMhNzkjxsa06aIlci+aNnKp+20PpuemQgfAUhhnxiA9WCC17
uhmg7J/VowyrGgcdTS/HntjV9J2lzU7H2WHLVkToFVXBMEiztP8m3nj1HbopDtc2EK8tVXTRBUIF
5QF4NOg4KfljmzjDCCDnjuR77ccMfqAfxHM+ApRmwH6YEMF4ZEqdBHnO2xowQk9kDghiOKPIJBDm
fUNMfVvFTxizTta/TRzdjvMBC7UQCKRCxwyrtxI89EowYSCCt4dAw7uy2klMYC07gZrWgDev7KGT
MGt3TovoBhpEcaK5b9+zXfijt55l3mtjpSlegWTc1avT6lEO3cc8H5hWS10JJJGVTTcaoseawHUV
ALcjrA4KbmVhHPCM3Qf6gMuCBPWuU1zLSY0gXlEIZJ2benJGZUCADVSr7+RjKR+XRlvRqVT90/Pa
uPIz2fEVL3d4ATiUUqcGNnoqfJJJKpDMvanTlf/5idySurisBd6ie5G6XB9pNz8qN/DEa1lZxk1h
eDsFhHJo97MngZou6nBuNrjnPwDbf98uJ/sFoepfOkojFFfbRB3Nw0thKo+KJ4ZFQS1c117erWZs
15GfnGOOhPKGlD3rBsTE9vUjIxhz4C5yP2kuxxfU03vWDLTl5OVAxPOtwPdQ7oTDqme327St69Mh
ySCe/qaNH9zBYm5VKTVZYG35oZzpYc7TKMe2IPoEua9V1ODWdHoPE22b9q3SwnbxZY/8D8Pd8Ipi
qvV6L02Ta8kvZ3GpXzWTjAML3ZyR33wPDVq5ZwfNZi5jyUYag+psWu4C2HGOH8hqiwKHFfRYFMTG
X+IDJH2F7usf1lJnTxyOqnNIuEoYRoXHou06sn/JoKYeU5ffExBrEdwXAlVtmsTKb5T08bS34HUN
V/d0QK3tnf+S/BMPd/YhosdrZPRbAOeLypgW7+z6sNAOZy9aF23WnOcVQQ0R9ssmPRCJd51awWL1
eTD161QmL/YGx5giVG6xHmViVc4svTjB7FgRaMgzrmpYW6RCc037UE6W7TghZD8s28OAHJfinbPi
l8Jyk55DWXSUzqJi632bpFNSEgO2XQ5iRBJwS8ku1g3negzHZwc3L1FL4SAJL8mKmp0GoKdWL/PG
jKcMy15a6zSYbpi28uci2qx1UGwp8AtMvxGIQdVZIN3FktU26PJNzzHvL1+GJhAJPp39qtYV0W0C
cF71PEJ4xZd7IQv8jGKqj4NwC0sgNTgaj0tH7eiKcL5vtFijEr8wBSs6tvCvWrmFNLkqFJCd9czj
zOZAntDBmyPDC5JgOtn2L0qVOwgxY940f4t2MT/LGr6Xc5vwFhf33bL6sgcVk++YPSXZaB/Z4VB5
tKsyz6leh5ddz/XvkzZHyCBaF44TZqOQvbpwdCkYBdEXqegoXpsbQfvLvsPM9aHc952E6DkSH9a7
3gctCK+FFtuwq8lWY/zQQwyaKjIO87ER8ELsRfVlcLHxlNTPhXIpPO6exFmp9jzPd5j0j76HMrEm
HUt4slMLSWFAaaxA6yN1p5lTtscoA+iM9FSRZzL6mGpQ9EeJ8sHjtuLMTkjhk886kSi/e0eAEzw4
ssMUmzi2TYJCtGKBMQC0y2InqPi/7ESflGcZ0Au6w0voSoDRZSVNcUwxyhxYV5mR4UIA7BFUaHtz
/3gHxtClvm25OB7CHEIKnTPcmkLhdZzJyySzFAOB9qSEhDL8rzaen7igknGxf9rCsS0ggZDTzDk2
PlVGwO17IVLNTm2cQKXDEscFS/ILU5nB4zee8kUyduhmev9o81Tayb6x+wtnZ6q1gTfgnPi21qb1
y7BSH9tsu3vO3E4i6lWzUsN5Yhg1Bkbj4fOifszi8TaBT13exaB79NLp1PxSArRD5P1qShqj4Jnr
RDrcy6ghkOiXX+2Fqn1fSY5O6afMMmtmN2HDDwTPu3H8Is90waaYmuvs9m7Oo6Go3NuOLsZxBBUj
Wbgk5lnrKTexpdlShDOkzJ5BEuzUQ/eVXlLsmxYz/v4RQBEIVSEADWp9aX1sZdVh6gonzR4r4x/L
k+rKMHxVq3AJtIoqhbmMWiiPQ6NxI2SQTRh+S7VqOwvU/UfxiB9fwWYWizJzAUsoymgpNi7UTVbJ
AEFsBVSZuyUeqbML5pZymsjYz72sPOaHpIAjVNCJFbUEzglJuLFwgf6JfTyfIEymsCz8vlxAoSjr
oaa46BNxW0Qysg5ypHdrm/44IPe7w6ZToNBzlnak/gNywUIsk9A4xlLrKxxqm7dOjmhtaNDBRrFc
cP3zre5McfEKbyTCrQ5Q65oN22hNyeyQ8Mey7bbjzyQAmjlPKLq3DUxoJ6onzuN0R4zMMvVGD71Y
BdyCtYIRSMYwObmGZyYlXj82uCxg0fFdjRr2KO5tRvKiDjaAzFGzeLE9czbLeEJwpGNh80ESgZGu
SJZNuxO8cTIGs64Et0ATtwKXA3DzwzS40dN8R8jYijNfKX7uvVY6Y8UESc6AublPOfFRsJ/FM7g4
pw++wrZYGlTqWrlq7IsxfXM2fxgn56NSgLalCch4yu4q5u3YRCO7CfbfaKFp8x9zT7N3dyatveaJ
s+lk9Ey5z1hzZKn4/jiTggZulPBOWS1dQAw+cSUCImrC8BENKg+0aPQIY4kfj+rXR/XLcyXm9dbW
h6E5uWgdi4bL0Jns8WVztOeLh31oUMeXTR8zUqBRMrM6DjOEC+8oDBCTF1p5VHipGCnv/CCEktHU
AtOJzhpIolnGjbbgVTKQtBN8vCxBSNM5X9feCcJ3xqyA4ZS51HPyM/DUJzB2sT3kvgUsmXgRhjFX
p8b63sqpmofC3PV8g9iobCLDnUydvt0f0uD+TGzOnhrC1PhFiV6Y4Sndg3nJlIJfBcpfaXAIc46A
ES5u/T+UBdN1L/4DGIwoRosNT4oiF1BNhKorvTByek8O2f8/fRhrIpHk8Oom4B38pJVM1PiLaTew
03JjHKKmnkgLfT3HXiZZdEjHtydv8fwLhELoyZ4Xn0bmjWVcTr0So2/ASBO+Tucco4/osvIMnRdD
a1gt/J48smsACgxBU5Jp/NMmfTs2hk4nK3bI++5hf6K8VJWd6ZAzQopAql/umfDGi8lo+mx4u2w4
Z78z6hqBferG5ZfBv0k8Lf3EBhl9ctHjUNjzcLaOyBagmJLhGclpcw40Vy0jxHWXZSEXuAPK6ueT
rcAwxSSHxGV4E16agmWmEZOs4XmeuruIsBaL23pZDiiGxmoi488eYWW6vFgEcbEYjV8OZqx9zaey
x7uMCcXHKBHgD4Oa0bchG1HL+4UXQQmm6TJasndNhT33tbcDkAubBXY4fH6Wtpnxn2sRwlKOWfHK
kogoO6z7GdoEd7H+IEpznZDw5b3UIfKYywp0536/rd1rGlJofFmH1geSpqvXMONuNCLVGaTXbrk5
FVVfBMLX2e0A5bmYuGNYh579+Q5FuXMrgQWHKc/5rGFexHhKx6w9fAsI6ss932wqAA2Eoev37uFg
NDmWdaEu7MKbPvznvE3gaK+DdnS41TUnOU5yQ1VVeuSs/hSfZG3YlYTF1gHckIAPPUJ3AsoTmhIJ
U2Mdq7MXGZm+TdbUJkAZklzcWxQi0pO6jeQ7Ttsd6H2xt0iviLufzQghcPoELyO2AGlEtIf5Mg50
EwfoFNNQVVQVTafpZ5qS712+hZnSC9yWJhmxqHdsbuhS3WsnMdGMrpqXAEqOPFMbk8OTj+lo952f
2xIeLG+w0aKom0ORzJtycWfOQnbWeswJ3Ce3Wjjy2bQDixRX6e7bl2dAVPyFvd0howKwnZnGiLPz
1IWSAzXVm6wdzY931lnAAMbpMUfgvtkacWENk/+PL3/u3UK2FhpLTwbANJV3WXLqilaCzAXQLwXm
ImRdJa+R3V+OLR4kE1ApU/sqH4VPPfPSIORUXOC+qIKXuXx6iOJi05xQk2scAc/D2JHfBETcvksK
shQvJwcLUEJC4GMKWhrvIc8WlxVu3jojeGrEGruXndsKR1wLcdNemHoDLImlLwdGUZqWCz6e2GaX
srLXRFq2IfLXGzpFb3MMBlEr8dI1bbzhMJ3Kk2GosY9kPEE4K2jI2C/6nBAY6rnTCOeAjMWwC6AN
Ess3bSSq25W+MHbVaA3oLGp6rAwnTip8c+KJ4abiaUtw6PuodnjziT7EKcVOUiIE5/DHG7iVPgvy
8a7UHbCs37hGpztKlhgVNdWedgeC5qdV/mLqV5V8ww2/ipDLy2lXkjZ0h9n8SP/UTVZSA3IiXP4J
Uy34CWqSBTO157x7p52hveMWBS8pM5RcMD0q87YqJwlHt4mvR915/5pKtV6GTkPHmycMDvP6XEOt
xAUQQgxR39FYE81tFGKeipg+aEbtNd2/hmESke9N+iq66Lp4nH8QJUze3WfX5WC5YEdeTnw2IrDw
3c9G6DolN/FmrwugsiseHS6/7BjgiePIEH54n6qRF/MYD8S9AfbmZIy3Hu8XsNvV2oV4bWB7sJac
BFzgtuJXZ96jRSNcOkstHDR7H2pQRktu69ENT3W2a316xlBoF9BxT5cIpxkXmnMTPjqLXYDgHwgC
Wtf0n9xHDS6GiKfvPTkr2zRs67WxVmZHqkrzCQk/LnoSEVUmv8O7eSXinqWCN0QZhh8KVX1gRnXE
IZHxGXKi9myG5mA/dZwVpTY0N9sBiFrJLPF8xkTkKoHgc77DrzucBBciyTJUC3Rk9NQiePLmFGoc
mv/2n/KBKYq8/LfMYfyB1U9y0s+ZzMT0RD5wpomtFQJPt5UU5F8wj9mSgxrzzUrLyy0vwAaYJZcD
H88W6TbZccRI8cSVyTOdruiA+Ma9nxpnx3M6aq5B5JLIXMZlSDChmnnGsoG/GF+vPt6EeFWm53Ok
a9PjWRad6zq1FgNZPjEYnPilcMUY9sMKrMNoInDs9V80rWIeLiBvfJktQpU1hMThxUAYLOe53k5g
PiJPblSfB323JCEZPckIrvFOonSA2k0Hhovq8dpA9ZyE9pOD4o6jvgT1lZ0WmnAWbJlUPxlGFKWh
2afz/ru8H0uzj+JyMeHibWwS8IOEXlqoNExnbN3p6H0zYrvCGuTJc1RcuNmpojNRDu5oo9KitU1H
8XGUZHeaYfyLzoqL95hcExRWwxKabWd73lrAlSU3xLS3aZMhDuScPKDivyupNA0QrdUxnwh7cMDH
nJisaAGuDGp55eBXtoVIY8vjopiLzFMD8j9Cb010L6dGvk8h22npUKyQaqmm3sIa7fpwCTyjn8Ux
4GW+YKvM2tWkkuagpRbdjw9Bmjb2RulgTHwdc8xOoQDD3TG0+3ls29aTanI51K98vIK6N1QyBcFj
xAi5mnGHnAHfIN2/yV51r+Qz388Uo/mh4mkVq6e082TyhthgaXAn5QaiAg47xrlwwLicVhkolfiq
Wv7lnNOjElzXjAtj/K3NVMtG/FjbaQqktIu4pAZAGF/9v3+vlCtsGWZSCnKQJ+rC4KCLbmoLh4le
2/fovsRFPdtW/lqSO28N2DVZnYVVQl/c32/0VWb2Z7pB8jFQqxD/O4A6XGg1/y6NxUhNMiW08MO9
KePuCQrpsgMPbazjN+bhkIL6Xg1ID+sXBPhEHhTdOm5Z/9NnPPdtLUTrOA7weq5NuC2+IwF2xbNI
i3ewI0224HhSYRdMcGa/t+07vgMwldrKqQecPr9MFQTI8dlgAUqyL6fliZoC9M2Uo0pNFvh6cCDM
d2CrQxI4m6KuFzXXlQCJ0gx+Wvq0jLZ0S9E6cOgcNj7F2tWV3v7wJVtvbsdD/RLARNiaq1sVXVcC
+0g9vpDP6BmtFYBRjeqMAeJav8XLR1PHme12jVCzjjVfk+3RjEawRlIoc+ShzzB4iYujY9+yJ344
SWvANjqFFutoJ/avOjS87h8x0RT6lHGXI7mrWB4Gs/6ol+fgjBEqbUQUBddi65nTCG7VKr17fftN
B/o8GM0BS5icSA1uz67NAvrJT+CWu77NlVMsPnfwIBQauWlil9RzfMHxZyCxF/0GOa/XxhiQzDQU
vnW8fnTNwXnH4naxfZ3s9+N3HEdFHf6NoNpJKF0ULC4gkf5ervAto6+JQMeFa86RrLGKy26HN6JK
Gc4PQ/Gnqnt8R/AyQPZ55u59QHPdS1OP6lA5HiFFKhDQ+q4v8Bj50HVrjN+PoAnuJZHwCua/YHkF
SKcr0s9PvfuhVGIjp/3QGDqSNwCQhT2i+QF/ClWo/RD4Xh3UHaDt6j86MkjhhCKqgM34UKZp8xiS
9BkyegHMefzOlVer51OOdUGyuwf9nJ8TDdffA6r3iHnhQtuLB6FL+humdXnMq/vYdA27VSevU8hU
v0MNoSurBoNKz8Ul+FBw/LC2asQ+l3kvvRsmhQf2QaNBDM44eKAckMp9OkCXrZRX5Dh8azA3iKb+
kAuvLAWpf1xe+46Jc+P36wWXiMq+a/62hT6p5rJSJ99sbTUXXPXlmlEmSxfaOH1Nb4V1iX7YnWRe
2qr7FaANooR+EoHInDhoUsJODNKC/3lWx+tDwH5x5Fls3Z9atofONjagKJ3Z61JojEOmsmx9PYwP
YQPay6vvsrBiNr8RXSF4S8Dz29mK/ZjMsP253s3kHJq15sP0zxHShxHQC5EAGBc+iHikx5WxsWv7
9qPkAbHWh4aIkJOv5jJWKq6XzSbvfVwOZdXyP2ouVgkRvapDAdmACVJFbm+qBWp6v4UiTUvEr6lG
KMNzjzcsziIrQl+DYw30CH/90DEKhTQc3ZoJe7O8gFxl7IgEKu0EZ9Ldi9XMqyzD2gqleoapth5W
+6oDsOsPZeQNuup1qttfiU6gdHPv3mqk+7Ymp4Y0E9gXJhDWpib4MCGqFKWNHMsGbDu8pjpUU7g3
h4vhfBPmyFmeGFDcXICXxoPJO68JQ6vlTpgjsW7dhIsUsQwyqqd4ZV1k4B7MMKIUz+ZXX7DccqJB
CaR2t/zhYKdlWcDokJzmx6N6+8r013P7rlLwFB0wUyo5xLsFMr7hsXL2+7jmJ8VuthedYP2M60bR
ARfzBHoURen7zLoid4XkwNpM4u1kickvY8S8SBgdU09rUo4a/GwGktG4pWhygelcWd7I7Ipl4Y5L
K25DEHyDY5OeAtsLKMaHXvOuogve/dW1QLqg95/YHOi66msNE32QANougJtoB0WtNv3WA0ma1/fb
y/kckjvlTRzieKCxkOjjtTLXDoYFdsRf4a4dVIdp/dGZzzW76IHVHUfTldtX0lX5qDD2lEDm72Ag
oiFTNIbVGrLY00WRfgvvGeT1vvMb5HuzdBULSkxjQJv2nz3kiLPF8b4l5RZDUBsnq66rSJpDpOHi
a6WK4vTTZD93y9A9cGLuHFlDZhNJtmGRboEhKz/eIS2QhoD941RdYlkmbtEYXwe4LHQ29OCdUf5k
WSt9DP6vEk+cfO49CaiftvpYAmCRyE3a+h7p1m3rNSzhckkN5/fW3WcBOY4vLfLg+o7S9QArTai2
1Xo4TYIt2BTicZWrc6AHZASOfDa7xIMy92OyfdrG8gMZvSUQrMh/1RnoXSlL/xfTf/eyRwfKFQh6
S7IyNDW6rd0oMihF/oN/13HmkreiyY0QE3v95EjUUUCapQehV/2LHJDWfLPZsMP8DfwaxxUgVheX
tp41gkOs3/clwQgbxVV0eG/gYg1QHY0mKOYwqYL6LMeyc0Vjqlo9JA67PVxhM6HMqMfdM+4qUlMS
6lFa7F1SzrLuriv9lZ6U5c4A+97b+a4bNUMrF2ZxlJaymyHf3lmk9RH3kftJ4I/wqjGXbuLkJRlb
AAYhdA13Xt6c4GL//XRI/h3UFa6vY0ocDnzl3NcCFQmAqWsH2f2g6lnEQwis2silWUyYfLZhTFYH
2c9X5i2FzK6TiyG7eieaybEiF8Z6ZS2fVvQwwVxVDtlG2/cPzh4l1DdvR2vI+cqeAnvDppXm/XwD
N5OpdVn4UKB2o6ECL/RCaLLnU6gZkNBsmrh//BE9igjYCQx4Eq5+UqNmESAhYRsW/wTo6HMhZvf/
Nug0nebnmQPMXkiYUcEaGsXZWWpaAMtn7BMV2j5ISQE6jcng0J3lZ70kB5x4IM9V5qoj7efOJF2j
BTGed3RHrpsjaQaIWZLvXyOGP4rPvxjuVKKjrqzZZaAr4WcyqUweL2R+K60QSRF022SEhpl6YZpb
ob/nRd9mL9pDEIPXsPtEX+3CXwWEBHN5xy7cj78aE9PS6TIrLNkZCA/H/VRNlUFnrz7mknCdlb7A
V8IW21ij+zCDIccnfRrmQ3ZvAravb8NvCz39GCLlEwCGYSQaVklpzk0buvnfWW7DTyTSg1dRhjKs
4yHNxQCWqz3h3XzbuyvzFFQOAc77LOM0ooa/18B6I2MpXiB7zVbDityNFiTDVH45G5ft0+dd8gAJ
GIb9CEHeTPa2s+XkkbLUALXej0LpzNmdkLmldoCLyxCdgIvkqO0o08TsU2K2HHl+IF+8PSwu7cxC
XSCz8w4Hq/EqPKz4EXpekUPqxdgLlP5QxER1AHg3m9DLNR+bZWOW9jemWU9NBOzE3ihyP81XNAYS
50LzM7bEJa1Pb2dWT8zOeNK3eF8CvH1gOJLVv+r4DTshpdlgoIiPgRFxJUl+95G5q+yfYk+hHCrg
ES7wcK4k0wEFSQQ9VJna/NpxiHE8GqAnYnnIOVC8iz/TJFH849ZzWKJz8k8xJe9zc1Y6A9nSfdDA
vHJjkN1vpJc2IV6EOz0enjbIYZTc8BpF7I4X6UdzG1N0fLqRvT0SyDjoC9McQgJYToyx+w5vg9ZC
QltzYOxl/KjGpThmHoRT1E7GVO0BPnil5VsqaQiA0L8eD1BJqfr4x4dfyrqzFkCkbb5u5NMexjP6
/rHwp/xi4ph7dhvgXdFQGluyXfE0F8B8AlZGggRzOQzjNFzkKpnJmC0TXSGUMGD3FmFBudaTR1UU
hSjq57ObTVG6yGjCGdRJAwyZSR9KqnBDZ2nmgb70rPQGmEe6/oYAsk0WaQCj49uFGxvq5SEURW2w
C7dHjkNea5kumuII7vy5nsNkjg1iGoUryFsyCsmZdzVV0j8zAB+EUsCVO/a1hV8LWPH+mO8KcjaW
tQQ63U8EAURojifQPKtgoee2mSBhnQmE+qaWajcZ7GcbK/ZMCTE8f0M8nXmv76SE5jZN/7M9ikvg
sLR6PQteeRR9YWFDyWQ8Mv3aX4Gw1tDmf5/me046ZThrWS7dMqFXZ3bYy9Fdm/DEiNnQmC1fgHQm
LRw+3SMRacWcmiTRuomUETXI8CBVWjUOnNorcMrWuyuV6uMWT+5WL5Rj/AGDzMQh3kRCMbtsgVsZ
M8EUPrdVLWymBahTJS9bSeXpsUw4LounMRVIzQbZ6JRWmzwx/MV5iTWIuqVmWnbpn+Qrk0O4FBVk
VAiKzgk/fK65Z7z24lejSutUsnEP2AXyKkrdKOjcv9KlT7qzP2VTWBseuGZ4ZxFDNFBOYtRZqZ1A
zQDd0P4iiehHVbIky943gKrwKXmBtjwvZafcNEYxIW0J2u0hH01GOCtcLorB5i9rouih7lYGmozo
G6L8KwdW7iBafXwn7C2lOHZKrzcFZt6ufr2zMHYgES687tqyDJcfu4OrV2KHhtHve8Sm4si1TPRh
0K4LHEWYsqeEew+vuoyMieFwmKu+IEi2bLTjb97JbE+n/a8QBIipFYBALBjw6v+y39ILndCftGAg
cUMNyh123diLO4hwrWLR4VGYr4C9wEkZ8NMaRaEEyPbx6CInOc2sRm6FcA5D/Gdu3vwbz7kpNsHF
oeuhvVFubncFG/gy4sperIHXm1AR2Uc+z3H7HoELnKUTxgnpXa3QMp0+QnlLOBHzgrKYyhW7lXuH
OG47EaEIzuUBcEAVACzENQWrnrt2kvlG7z3ZoeJxaMfNuCEI6c0LaVbMRTsKDZhQsvS/NtfBmhVH
cFoV5SpTER8n6vfSx/Mn18g7jA90kwmKQUEC4jCmXnavDPpdYYpjpGkEcImssXyGaqPb9/eX4Gcq
8d7xtMOoCZlO32kb+2FUJ+WgAXAOomgEuHXBTqc9D4KCQznOkondOlRwgJO1GNP/pp5SodzORHoL
b25syJyxl1mPisL+lv8B1PwUj0/uyiqTc+QLtl/ErjYPhxR3o048F+UJJtFGLdWNUmJzsGP04Cw4
7f7g0kaXOLRgDQl4H1TbgMgUROlL3xYMJPmD+nmNT2awBBvCPSev7nwniXQJG+ov06X8Whhw3vVE
Ws/ts5DGop9xyDiUfjheiRi9K+fcY4TYVXDWiG74Rx8q/g2XjcSO0pIJ6ElCEAO03qEHj26wqK4S
iBqfFenzZ2JQ2Jb09HycXYX34He+v8C3Yzyeo/ozyLsM8PeCO/MQNlfpxb1VrqnUIN+J4+iVpTlq
W7BpDT1aM78auSVA3bnMExW8+YhqZii0ueQJ04ddU5YvBI+mOVhc7IkkI0c2L7tOSaizAgPsKmJU
Wy2d3R31dsZ9EkvlSPjzrL79Zrb1m1dU20QlDLzq1YDMAZCF8EgscXSbSQ1PVArsm8RZuUUjOii5
zBf1+kDtf4mn+kqljQgQNzMPWaDbyXd5clmlpS8cfwHjI9XQOQuiSTkcBsXDDUnjS1sX3vBqcjtS
OUBLkFh3zFfzlbWjdIgzI2tKO2b3iUCsknsfpAbMXQys6QhXgF1iTznXSZXKuC+CHBRaDLuqIf6x
xCiodP/sImNmc2MZE5A+fCyd9v3fir8jfj8SvvGUGjnSKfW89GQ+ADqnKRkNhC2pzJHHkCPOYcBH
96xaUuawD6PZtpIt+7v4baSodXlEw/oaBFVlV5dmjU6lSAhw1Nl8h9XYu0gRgReKSRCX32VTvjqf
eqarMhw0aXNVwh7cE9pG4d7YHEsaAG+d207wkukj5cfuJEeW7S+soCDLhTLiCftOGdQFRtRpSsNe
E9g1WboYzs0Qj9WZ4eMJgkYIOLB2WMydYIjA93fjZXYlcoZUyI48GOquCZtl5MSm2URNkwyhGD5W
o9V33GB3H0g+q7GEOMSWdBe9D+K2fS5HN97ZBl25g6evmcJvV51v8q+bZlJsY8LF2NKX5MG8vQzj
BgHuXwEi8q3o0qlHcHx5Rnl1epxv0Sr29kQmC2KHYKTTHXMApi4CNmPos6oYIegJW5esnDS3+ktc
Rqn261Oxx7Lv1c2rZsozsuNmMqb0ttrxoeFAnmHwnpH/L6smAK0xpogsCjpbgV7h4dk1Q4OhwFRV
vxhJQcL45xbXMSTNqJMU242mteYgsrecJlIsqdf47IEfqK80eTwJSI69BmVVlwWatTA4QlqmY+zt
X/B3aMhNhq/A+nf6F6dxK5FZy6bavYizPBHQ67HCJPp/+vnW37e4MqrKlg/rkpEJSbmOS65E5S8o
Dr1dvsVuJTpgKHLIJXykaU9RiQYhSb6KwlL2+YpUA0rLnuFpBqGoK7BUOJC6k7kylSwacxGV6qny
V7pZS51DiyuJc9gtV01Pw9+jqwftNy3nPvcbVAefUEjFvbvQqTUoM81QAc0bGC5gH6asnVWg8x7p
CsqRTplbDMUNvY89Xz+hxKjKq2mYwDgAd1BSudUcQvr9FQAi0vs6VnOkYvnjiiSMwJ9kuiVD7m/k
V9sSWBSBaoEDU1k3qz0ZzHMzLic0+/9vCBbMFPWAlZnzCWmhz6IIjQ1YFnrbM+6K6YnVRE6RMqbc
FB2KTOSTZD9+Y0CQW3knk+5QUREI6nYXQZeW1rjsOputbgAtEYtkA+jZWiQNYj0TGI9bPp+Flzve
zV1HwAcnhtVrrcaagiWrp68yipvrcq+29RKLKHxg7LrWuDISL5jcaB/AqyiGEiOieyyrp7SjSvWX
1cI8U5q+cJR/62ujoxI1ZSEv9svcGhAGdKRZDTjEN4xKXiubZwtBJIcR8VuVjvVHix8ZfGCf5b9A
tJWY4k/b9oBxqn68YLf7aACHojwIMxIB8h0Xf8Ih7DHwZh8bCy+RUZTwlb+oZFMjzdAwlzc8AMTL
eTvQ4tQEwtYegnn+gozYKZp7kiWsULp02HMcO/ujiguhjvXeXqrkeg9p3o+XnmFDiQeIebEts5YR
aZ4KwhOUtr1uvKk3aGhqSOz6erPaaA/2a1JtAwnpK8egPsxRE/nt6/Mnzagsxj38qAFq9xf+dq8A
nH/z1Xj5230ytTtKneFC1tNrYrQW51vAxNTPU58BsvVYbQ2GbZpUYtWTRK3R0R6UJUZ8IEmnv94p
rejXKblyE6QNT6UQQnO2fIZQ2ywmEQalcpratqVlhSQWFbvsFOFjPYnm5Vra724LbNXWQcycl3+m
dz2oO0iRxZQucrOXX5gyHsbX+4UFxIRjdRwcWq04TLRjh0QYSudBHBo/Dj6ZDq0Ze3iBfaX/GBhA
FY23+iNLb3XmfLl2T4Wg8AUzlD4fg6u0L6szhmd/2XQuxrgSPnKS+i50r7O9nG2fSFGCGDJ1cB3r
ZKdPBZYOEESpmOOcpuzpN6ArMJ+vSn+kk55eTnNdtUpY3tMpwM+ThmUeQdjILlhFim1DUm9TWNvQ
csffUvJGxX7uyudykt7LNMXxxCCEKw5EZSXjLKER+H2ylb7nwy8mwpxl/pNTQ7kW7HwdYl63Cvz1
RBQcC00w6+Hpj+Q/KkY/qH2UamdPDitTjNYtm7f6A1wlv57v5AmA22Rki4KKvF44BhWaaovRwxXv
5qZ4RvQn0rQDf/UTgWg/iRMyqgGMTOgKOFhhNdzZ6ElSFbYwvCHGmudZsvRhp5pZrSAFilM1otqw
OZEQ4LLwNODqCYUaRw+GVrmy/7b5Wp3NuHNv+Zr+v8YlZaBMPY8U0z4DFen80B6c0rrx/CJ1rn5y
X/wWaI0EN512KcJvLhneAMV+6vbiRHqTKwGBHKUtfiRte/5gzRAWitzUT9jptlz2PkwhQdQjherv
JsQH4AXh35EVPQM0iwukR2M5xzmx4WD0+HUcO/yXXYTq7tLkXvGEWasQJJbWa7U5GDP21Zjg9E5p
xdJ6Ado/M0Qnnqoi18wg8ywYfXYo4iASNvQ1p4CMoAlxB69gZJB0n6wvkYsPXckT02ZbYZAHJ6TN
Nf+sbvYprYSS4VS5Ge1wxEg/P/VMw+U+8fmqucLRF64SDTYpemiYO5+WoSq1qbQuZRzg95Tnnd+9
GRGD6drRVqr1NE2t7YDSRLyb/CyZ76Uf9smErpZy4wBfEXuBwTgEBCjElTsywqbsUoC2vKTdqGBB
TW4DL2qPBSwd69NVqv9jnuOn9FKCGwVU53MxgczxBBqFw4e1t320TlaSevTSRPJ7UrCYwHD3Fkrb
z0TxqFCe3esocnM8T28jYPPI1KUgBdpOTL1ePiSwyCPQSgyN6jAj77j31qX0CjILem5fA+5SNa1K
dTF5MgIVR3byD8neOt1ljRZLb0aU63YuRTk5lGMnel6NwOop3fM9/HpFmSH182VFI4x4F0c30qfn
EGkAqgMeKqj0G2ngWpedYOPaCjEqVKgNd8g8/Z0uLc8RfaWUXoiBOMts/fG3lEnoAVfyQDygOLVE
k4s49mtLJPpe2oLhcTEOLGT60LQXXvPyBtt1Izpzebo16dXqGFriFQReu+iRTWEYhZPfbQ8psL50
f78PuKvyP1aEF7u6rv4hn+b+Lx2ad3X/GFXgTCTsW+VASVHArwNcbxNbTvn3gjMpiLRKWKW1lqKF
1mY9v+eiyw3k4Q4cgunj1PXAcxhBQKa3GrE0Icsg2KppjIGtC7o1SKl9LJkVilAg7QC6/Vt8L0zt
G8JXczAi6sldCma1RJLUEonPASB+fX/5gOjdQxQ9ZozaJzLnypNcSaLVs88VNIyWkFyLQ99sU9Ze
ULlvG9QMnMqrv1fLRQEt4mpp9JT1jFkcx0paj2eimVux30C3t7uCH+EDOK3LXvzBIAb1jcmuB4d4
YAaHU1/o5RTsZ2kzBX5e+k4UrxhlNoB3Vfrf2FBU5FNdXnZwv+kYXX/aOR0QA9H+9zeuMDfyuw2K
IC7C64V7fHE4Yck0isZ80olpvtjh5UA9gg/rqjYcx/dlVRFjTcPmXxYThrJm1eMIV8btYcCGV2Z5
vSTcnMNeRB/XVhCSKxMvJHi2yQJcxK98WvkxCEeBWWwgphWCCWZHh+WywaXEQq2onko4VMfbiyKV
8ZenpwnYWLIUMUgQUTu0fl1vLb70pXtEqWgbGwDFLIKp+xqMwQ4CkiuNPN9QJYOK/5Q0oVXZpv+p
M7ssBqBv0wmnDzko6yRSi82Qt8pbtREcK1wVjs0HFmcDNPV7I9RKHmn/zv+OnOLTJJVpiwptpcB0
XcDUZmU+F0xjr8kTkuR2QyW8Th1Qhrw9CpoqAr+M/JTdbU/+iRlElVY/RhkDCmusye9iaV9acBw7
plt9mZsDon6kNVtEiQfLAR4f+/SC+zxpkV97D5kNQza3kwewVMk+mmgOVHCJOJlJEHdjGW+BwxEV
hhUsiOcQuUHpNq1naKZXf5fDQUUSX9KUbzCsa40WWytQygcv2yC3FQhRZlb3U/gEU1/8+gG7v6ov
QVScnH7V6LnGIjaopZvTDCA0+0XU3Ecd5crmHF03QJOwEv+kAJuMUvtIh70suXgrNrffEjrHgduP
Y2spyHhuT7ywprWDFqAQ/Q6JMRBkhBZxiWKuD412s3l9whpU7s5FzdfEK7ioB4beALY67BPT/vkk
ek/VXrP8y7jE2QqTJQRnXsxUA/wWRT46KyI2MvA0j3PURLSj0PwH9OLYA9saJOoVBnsx4+4lqwbZ
GaX2VvPT8pBqgvUOZFP6J/ue/lc8XTQHUodIF/kLneT+TsX28WnJZVF9uQDCqXn8+2cpn1PolHfs
89x0i1JXJlXEwp6fjKTKrMPPp9Q4UPqXrATFHtpFyr1R6BbujKTqMK0B5N5plpqOdFfGY0wiQ7ys
dCoXhFbOn+zlbiy4+u8aUA0dopOLxp/UXnUtj3AnJUNfaCjyo5EuoUDeR57gLRgwVUQL9KUjoB/G
Thsnph5UK8HtbYWY+Xil61Gx5vN+q+W/p0WHKhMI3n+fzNYps7VlKy3DGcbSp2ccPEqyjxiGLQer
RNARlDLsTr0wl1XbOkfjp90EdTNAcl92HgoguqcckV9g3hRvbN4gguWTS9AA9yWHesAyzSysoiPM
H+fsHPVxb+mpX5VuhvPt+NjFp8BmQ+YTOVb+7WFlZUtadv3hVNhWIPMWklEvNQnLLR+QVhBDKs6c
EUneajORSril/3SNNLart7z+MIIFnIVv7rGZ9QDn/w0LbamkGJIizot23MkiUYMEWDCHjEWDL+Wc
yN2l1b0SeckckoOKf9/S02JhHWN7XbHognCEtBKt86sj9f7d/IsNXbSyQ7szt4fjObyu7oeConyd
mR1yj9m6jgA8S9xHi6/1jW8W+nwrKIhMI0+GTxkYvjCDbxpJ0KSMQUKj9nUeQTpvm21R5DZK1Pmr
3OTfV3xqD13F7w2jz+u5T645TjudwfrT2wFz1j97KPD8Ixsp4bQW1a7IyPmAKb1bRPemf8HfnNAP
jsjJGEP/+7ywUo41CDhC1ZzkRgrgPnvqDMdqfuRMvhJM8/+vQbDTkqjxhTC91ILLqmlvFVz9mE9j
l7uQw1hciOzX8w8pXU+0plGPgDLJM+DIPqR94uEwb3UchPD1bSXBkAVpBpIeL43Fq3h5x36kLE/N
tau7sFip6pNvg8qXmg166oZXJWBeB72Z1nEQLMkVUsuOuwBZUAhYr1nrhgPBRNZUjUury+VYSgeA
mIQwMIh115lCD3jzsH65D8nrQoBZskRCYHJFMRN5TEV5Dfn/MU8Yv7cVvbLuhMfTRoUY17cidEh+
7FJLxz71XVJnIHQk5ZE9wM7BNgN9D48c4W8hjJqDn75oSL+O00AFJTyoBrJFT+ZB8fzi33yUNss/
vpUVzLI11WN3Wt2Q6VFJHsdLwnL2UZdu+02vBLSXWfNHwc8ZQlbKfxW/7qM2OembqPt2MFZHpx6Z
nnCoMe4uMf9iMzTIJLOThCpvYQOaMfXtxGYeC+uBaaS/hQoYXWdy/FKp20NC25d9WSmYK9NMvkue
A7pWHD03dpU13YcsBw7BcWKgkvJfOgU2Ejxnu1TnCfXfIbIWxXvrfoU8XWwcym5fP2Q54aznlSF9
5qe+hFmyH9lo0MoCte5ijbivyI4pqRrd/0RH72ywgsX9TANvTx5ue3jY/qMH9XPEviy9MZsyKb+a
Zs/raZN8Eik9Wb0ZrOSgirOB7F31Fdoe08yw9wfPgLsHvXN0ifmG7cBpzvkKu0x7tUz3+54h/+dV
WXeM4SFeY/NEFB8dg/1dAswDcz8C4RiM3oPvYZjX1hCyWjWbbtWvUOlooa7WuxtcrrRF/A/XNlXT
QF43F4WUTFgoBj0ppRwvbxB/aUwvdfenCunsx0bIs1pnQ4lFcomfvsCy4agHpfdealoJ5b/AiXcU
jG0ZO9LxnSCttX7bIPbL2PgNhnmbLE3SzzDV5vZqNTaA0vcEu3meb5RJB1yAh6W93dujPqfDK9+N
/U6RO9ZMveJdJper7EO/6jKE0z6p6GyzqJ82XjAz3Pm2+oCMYdIFrBFr2uqWMrGdpz0/sTlYMwQz
Bt4OKWwqnpzBTdp++u6J9xL+WdIYbWFMtVua9dxo9MAiGSmNb4qkx70J52C4wZh9c6DwIZVMLiAh
tG5XtRIQ6eC5U3D+WJZVqD45mToT8J2AVYQEt8UBZxMVEk1m0Gq9q/iMRZOpxJhXf/Aq71ppcEUV
q7mp26UpxSSIzozp/vITiRrsENG+yuLH3bZo6w8Rcm/jqsk3LhbLBf7ZL+402MRwXenzcnpsok7K
98lrzNcD2fNnN7MGnN+6vf5eMrPMOzlak4l/A7UOn6GCTLiRW9KjBCiDmqPtPcoz0WjuJ32dqQ3V
qh+KzTEbvX7/mSkeBlAqcNni58NYzwgaI3kGc9sx7ivMDLv05KnjGlW7S+3CNXfggirad7vTaug1
++sLwt4r2mOwcVgX8TmPSYStIUGrXKk6Yz+jm/N4StKxgf0XI9yuLNsyySThz/ztm59Yh8geDtMt
IQbIfyCBfKyqF2/3SkhnaMIggON8ZMpLkCjoBX6UpfxYig9A4S0bf1N3Afi0jFE4SXSeJza8qC/G
APAbpM3D1pIXKZ8xJJOf0cipElBznQ5F4ZHsJhXKB0aRWXnX1WuQJJyuRyKmOhYgAq90y3h5K9BB
3dfcAu7ZfMm5RVgjSb7m+vczNCzNI8Iw6nXuR9VReDDrXIdQqk1k0tZIvo/+FMmcXaMyGp4BNmEy
YKYzAz5/k5gW3OtNebmvY0H0Q9WBhAL7x+pVqa+uHLhOLNx35C8A/eSnWjbz+KCgIqG6LmlJbb50
Lvkex1Vorx3Go7PlFLfZlczxcy54ZqTUjxpKYFzAGdgb1NEXPE6tXGV3zJes+Vp24pT6BtbaQj/O
3kZ+SNQjiLl0NffnzW87FIK65Wt0+J7e3GeZa5ypxhC2B0XP/pQ/VaIi6iS12eS9I6O2ErrDEafU
DWU3JyqHMYLqiMwuCWDV+FUxULU0Oh+GcnrY+D34mk4mRMzYV4xUCoThcjT/ImgbvunpjrVdIpG6
YaA6/BYlY6lBdkcdoRB7XBlmLbtqvuG7KgWlBORBE+4gOAHsDHzvbT1FcdNIdNQhFNmJFKjKEAeZ
yHRBrqwCVOS0zjg01NFhv1dAzoedXNqzQnLGxq4AMp3EE0iNb5OiP4Mpt44iBBCwtaFVaRIs5uBS
V6hvEx9H+Ez3Zpa4ARNvqVDEW6LHF//vIcpEuSZjngolMqU+3suTJTox7RKrHS/FqUODnpWFPMKK
zEr1XM6vG4X2YbxCvnX1AiEOaScVlWI9n/bOX+cRc1sAElShN8dgZQRsLkPjkZncYKD8SAdthnR3
V+9bJGG+qRcmt4V9bfgcxX6YYY+7SBRAb1QRGBqMTDfotYiMQPvOhXG7e6jBVMilIBHMiqUgjdCI
WYf+x6YzWh2wA921WsyIIc1i3QeCBNH0zBwSiry/mTs+RwXunrixfxb7p+0LmmSwieqOyCSXe6Re
ovMpWAlBqDupBzff02DOliZAukqkIAdA7ZaG+QxEOyBOsNBdznx/6ER7m6AGzN5VQzi9kyxw9ycT
0q3SPlMXqEP/MF1T+86wVYpaXFUlZNDEqod2DHpzhJcE+28rJBJ1Vep0SerRyI2MfL908tSpMT/g
wv9c9OgI6WNJf+k9r2cctjPynZyNQpBwonUqXexJ+Wn/tjcpNsKYjpMkUM5oY1PqH1CDqR12jeMO
jWFVmaMHb9/REbYd5qEjMxeorTvAXtseUDRg3Bwinzw9ApOIfzmWoutRw/wHE27b0G/IUbKbTuYd
2dL5nkDjlXxYNChAFiOACucaote1o7EQkQJPRIXcKx9+kiCPTHOB+R8fr2I6REyOLdR+/DBZB3Oc
IwndIqatk0nMZ9w6WWhJft3BLN54FQrkb+2hl23VtoMUnuOmy6iiU2/fD+V021Lule3L5IIpXuzb
DS5/U8yKqad3klWy7DaQRsy2Nc8WS5Pa69onHrnLwV8faSzRQcSafpbv8L96dBQX/eG3jVIpF5nV
MKo1Zm/06nGoPpi3XlAl8Cr98CAJ0PeU5npkQs8So/GzChPALeClNiik4bu3q/tshlSq4Y0QGCet
8H1ZYBU8ViEkN+pNtpn/IUCCAcEUPJMt9OLkKLPl+VKvcLkMYGL/m6hXHAZQ2EaooVCNjd1Bbx+U
0updot+EYEYdw/EtEAzDWuTkpGxN42iS1wAVAEgjgAycph85ufk5ZUKFjSv+MgAAiyuO5JaSezeL
DiSGokYv7PMZiUO/Bt+qzWS9jeJFGe5mW0J/0yYUrpsbG6571/sd+JTEknHm8THzq0hm4sWNCBKX
3bXSTrqYlphvu7WmNoi36jJ/AQxMI5chXk/ouPEi7KXF5HIfA0AfN/RgyijxBdlCfeqVPeJ+mKBj
MlRrQjIO5wMXgS9UUp24CrarQvrvQ7Ymj8A0lLwU4RMiOkO/wo/8UazJAL0snBAsfx7SI++8jZtL
RqhgKRrdiq2tHQviWDi0ol8EjE9dEkyl04JXuw6y+rU1dvY43mpv06khjxVMLBgs3xAXxnj6I8Ke
zsb2/7IkOGXLVp9N+XggU6A0s7C0fh9G8hFytt4RaZXKrl4nppW5S12sHNaiQOG/ov+RkBWVM1hB
6DEUuuN6/hX7p/KwkeLPUbdYayvr5K8OuR6o2c4/A8z7kWW4VYuQ2TSogfbbN+xN2etQT5f5SeNA
BHkVGWoqOUEfqMkynWd/SgPlyuNpwmI8IyAKJcIZMSz5iS/skpOrNgDNGD/yY2BA769d8QnFmu3+
i6FnEI/g0nNL+hxcKkn49Dty7XzaScQkUZzK8B+4FuXbS4k3v0XGYrSYlEwZnJYVUzu3u94QqHJd
kyWpkogS00S85z2TpPiJUl6xkE86f6wBqHCoxGBbuWtGs0kgsoo7MrfDDAgfI6k3LAMsgaIr7j7S
uOWVdvvj3RmRoTG2koeKrp11IsMQSX3jQSQno/ohq5ixOmt1awNMnlIGrRcFLXqzMNEEUZUJmXpd
LaZpNKpNQEYIxaiAN1I6i7SkvA9wTXPOF2AgNsh2/sxFFU+/rOW7j+fGY5St0WrCJhy7sLSepshm
6kkzay0N8wCbt+S778mTMpekW/kInJYQ2/Lm3cLznhepaFTcA24GOszQiaPiq9gfqIuZ34TsSNqP
LhbicuuA2FRwzDvlVLsZtAo2CgQmWIaI1FtugspqLtBHbjnyBg9lm3JtPuNJERnkDPhhjhZvL2Hi
0gaQ5VfoLV3neZU27FIOQI//O4whghNIB994dapeHTOerr7KoucnETU0RpP9UkYuqFdQiU22MghC
pjP4amCwaWHcPZnCEkNCRV4xXFB5jKQIBFQb8ny172b0RY3MgKAGqF0tZxPDQzDImVwLeo/l6xz5
hhf6E+6Er6ip8/5JdHjTZCX/Bh8A845WC+LFZsdYk6fUDEfcMJZbceqk3iKo0rrh5O9OoDfZv4iP
yqbF5vj9hahA5myHu0duwUSGsvDoXALZs33x+RZ+Fy82OoMfGXIcFkM6lINcbH+nacl519YeV6tq
eCJoF31ntwtjXwQ9dmOzuyHhDI1FhAncZWiKfvyzUzKFshhhb1xM0Q1yrxVHVShXM3Zfgz66tTSi
SIqRac7WgnK+1Eu/QhOJFk5wxsxuJ30BikUKsJ+/13aWqMgMXBYEUQVdqiUlxBJTLZPMIsbxEIbh
KQkoFsWU5Qf+wXhQUaRc4myAYLLR03J0Vn2dccipnGYs6aYEHQ7ijDlpjMUdC91D3ZJ+elGD61Tw
AX42urU22YfMzjRuRwM9USCell4JdqdnINMjLH0CklFKirp/B/G1yQe2+YVwArGxWLE9g+fmUIDH
7Zx0zpBq4cctBJFPWwdjp7m6JH6boAqg8pj7MtdveIMXx0SJ8oDAEKUVUllW2/Ib4D8BFcjF4t+M
R7p5jtzwB9t52SdFLRg93oMB5xsT8lZXDegGGwyMLd0qx6lWC75w3494nSS9mD67xSa5kBgj7sl+
l1hX6wJq3SuRwddJCTax2BnheGO6DxZdJ56qD7oFKR5rC9s0j/cgy5zMryqHfxX5eSZyPKQSGt+E
Cky26BZOLdqyOB+nCxI2LynfHpNnpK43YsnX1nDtfXob21Ad07gMdBt+O9tqdzFh8zJFfyYdZHiq
Gks+NSKP8kcNWP6Sd00cgHUY/BTXBQghSMM7rEE1TTg3JFkGXGDAYtDjie5k/i7s/27T4LiJWebj
bViMuMktdqW/lemQp9q7T3zjqpmeFaXmTEf2fL/HOJnOcYXO5EutV7E7zZfhkJxDt4pejHpoKtxE
1Bs74xOeLxk4OEcYdRSwrZX0HOeWPrOWFRoCGCq64BOfZJF72xQ7vRPEzRKGqkyXvy6ApVqkzx+T
t7iMYR0xYDaWJkjzbazIhFqKxaRvCaMW0xXxacfYUtk4IqU3QdDTadFe5fXnO6UIaW1xDJHeiMxx
alHDJaJYBuETq4+zjVJYtWUzOfGBKRXhdo5LSpWoI/MnJRpsLQQRLM2nKt9rXB8EnPUf8YOtCLjE
ex4a3XBiYJq05FGXLbrtnO58pm116pO6sn/0h7jM4nspDIh972loI7Ih28GKzQChsaEuQO/eG3PQ
5D8hwjEBl3n6rl2udLXunf2jJwrZCXdsyLYaaFq2TG3ZqjF9VZ3QvQXkTSEvTIfos1knWX6/whWt
438ZhVvPEEpMiEZSmKDQp1Fr12Rn5PJK3wb01gHy3EIXXg8uUZhPsfowVotWWlrYW7I7lUCmu9p5
iV+W+0+YFftRzSkyunJNrLY2jNvW5JOT1uYh34aFEVfPHLUWxEPuCk4kWPQJaM3KcTQWlItpLrX+
CwwOP1lbucvgxu6PnuOJ8rL5Bk1glACYu2pXNxDBXDPE1a0k0N7vJqd7fptPF2Cp3cyHNI96K1Y3
qgRwtiGVK8cTvOp3AO0C0ark71VaGUQhoyErpmCSiXWRPcwqEFkQZGazPd0Gu4mOLJnbKBe2YJAS
PEKEKdDG9f1gF5M0z22tRp+QJ5+ieAq80WRO9f0t5PSIWENuUt/vvt7SJ0y8jf6S3bSX/Mv4V+Uc
corcTWzYSBjUkqxTuSb4wtKfDUyXo627Md8QvgMVwPhJzfZNG9b/LipzlOyzhL5q20szZjPEizqG
Pw7v7/nZZIaaMBJwggimZzCX2JAvnHXeDcfMdB+0tQbVeklwTyew8NlHKqJzxBL4fHkvwL70aQmz
gIw7NbZvyeOpoYC0o3HrbrKj2rEJ2PyUcTx6vmLVZjSf8FT/kc5CGsVSuKf9oEjUE+e4Ljx4g90B
0goT9bGfpAiqDRzvCe/CAYM+dkDYYcnzDvQ/HjqlnI8Y9RNAm0mvPMHzg0i/iArbU8QN8uSjabkx
Ox8wolqVxrfXQdq+lyFH8Ctsxs5QArGi1m3BwDRrlrcl97avxg1Btf4WxCP7RQRfSdbmj9T2yUKr
q6pjxFcKF3QtbvBaRfFBbjuazAsjuEeUTKtHpD0mMD2f21Yb1KSGXbPY674ctEH6C4KP47vd34dp
2Mfd2KkAcQWrqSDm6asK3eiSvv1BOhx+tuWI/VOmhikp4CYpRG3+gQp8J2OrPDizoSS/RuJZG2bJ
F27nzRuHP6pVihgor2ac4AiXObVx/drORnNgyD9N+l2hPwn+MH+jaUk6ftDJmdXMzq5SvUarTF8c
L0Dhoezc7N7kO+cneGKk55FNS1zDvLGLhIJnqwAnG4ZrAEofgdkm2bfXizaUiv0zXmk0KhRCQfL/
qUdg66VCJTE53R65YNPmF5WwhcGFvUE4TpLUd46z+v3aMwYt53efrn2rIT8IcDCQbEqh9RgL5ecR
cOchefB+MwzBwomL0g8fNfWQqriRK2tu/TGcl5AVCGte/GPvVb4tg+j6yI+BvKjeGWSEGufw8NZP
VLLMQNNXfxmNS/9ntdF1aQtQ/ikNeBVEPfOffk2Ewx9UyLStId6fzGsOM2Irv5GNJOgi+ybm5a67
oJsQwVrQVwjgcAPPhXcZuSBIu7K/Eqp5j22suv6P1FX13Ft6A7xR5NIxxwK0NM4806pHRsCYDLn8
pC+rJXGzP9rC+hJMsS1w+ZTw9+NKn6m+5U7LPfzjHejcrRudhxRh4bP/UhxsbZzr/sgvg7WugrMF
JaQRShLyM2bzQR37GjCfRNKXFQdNo3fsjQjQREAd6y448kXR3E6ErRE7tH9GC+H9tLNA5VRciVG7
in296JkxyMOFInqdKWWDqe0cdUOOW5qnyFXrVQcHEmH/aIMhIl+i9jAu0L5wd65c20CY1OoveETe
klM2JsBMO0cjdYaoFI/xy3/qwUebSA6IcbUJBhTHtIFSy5wXQjHPV6vny9Ef2zxu/p6Ip0paiy44
h8Yiz6ZypqiLLsMilOiwNu1PhLzL8LePuU/4FCnRGhZh5SXvzj6YFtw5I2kH9ac1VFxBip/6UqXM
8gW4bZQw90rDnfY5Ss9hfbRcgGnrtXiHWx8P4G1Lm01I5RKL4NC8JVQGehJx1NcJ5PEbHIFlMWYK
G/XXJ3poOrsWr35fuA4vxYyD1mKbjN0ZFbHgfX0JD85NLfrqhjGe/1Up4L53NjmUCIcGN9jOXzFZ
e68EP8PTLUxjGNs5LT2Q3/tDT21hmF0ybgutsktqovKe1wrv/3a3uWrS3A5IMzdrYrXbqpU0uuO5
Hk9AeEqQcmkX/vkXrOs61DF693TH1NzwFUFLr4v4Y4ZVmCQH3jrQvfLG/JePLwx6fs6QTYLAH1rz
84zjP/fl/VfT0C6x4oCsAhw4a1RFoKFAmkD3ITFA+h8GBot/1cnFzwPy/KoF02JIHQbYsLEVAbvQ
mWD2wcusBlLFNkLHbTvfp87+hgVbtmBPDdfweipzBP2CU20UmcPI4o9HLFXRPiIkl2OOW3dSGZ63
8+NPvD5P17NN190qYxbotHUcvQJetaAlNs+hW/rQA330qJ9abQ8ASDikimfYBtaciIKEYT8LAOb5
9Tl8N2pDNfnJpOKPSrPU0cjOAUMCNq1fKxXKlhKiSoSh08POPKaojlFSnRXDrBBkiklXuHQ/wdTn
x4lhU14WVjsvO+89Hkt+PNDELDDR3Qz9TxBUP89Ekgu0p7uuDwhf29JuEGjDiDhCO7MCDww27PRj
bZ+20Y0QUBnMtzX/4h8Fa85aocHCyzgwM7HidNOkTo7+MCG649lc2z8jogUugONThthgW+z+rahy
yOdUwgXkp51hUmHZQgBgCiiAl3KHVyVRs4aoqdhlCWya1bZXsV6hkv/aN3+esf4qV2OFKUL00L4U
/CESNrP5ZSO1ZpBteCM1Mhv4f+F3VOP6Uc8VcDB4+CcfC6kD/RUKDOwuOkbusLp+XsdaQ/6nUrp0
XPmw2vXBkde3ggfXQrAp1TUYrbpN8/CbqzQiV3FgqTF3slG7IWcnTspwKff1oarSWwy+2Tk531vA
hzz7hEpT2q84XSnHUw0VFVOnvjHeLgRCV4myApJsO3xm7RHm9AGVOFerfkC+n9c0scRUJiydlh2M
xRGBwi+Z0ishDWbMeuujTYTwTcVt6vu+8gUG+kSwWL38gNlf4xpuxDiL3zBDkkbMMox7wsSJY6Lk
asXuoRifoBrYnB8fdl/KDliK/WzDn+6sAq3MOtJG4T+lr2VlmBTTvLCk3Kieyo8hMzAFEvRBYye/
q/Go06csoN+y7l+uvRaGeJK4dSTIN5HbVZ+4uJcr6JRMkkeLObjlL93ec8gQBTnbtv6zE6kYv30V
huYZjPsilOryThaiVmfYYHlTEdYxMyEu8i9sVHommElQSyTASOdx87ohdcA1JPz7AHofThxY4vxO
4f93nZzP7kdApnNAGd6sI/scO+mHhfj2iCkAYlqeeo6PF1ZjdUBW8nI3OA64fEsfjEmNxnmvE2Re
vgOFPq6kC5z0n/UwfH2pINpnLCqqMNi4Z8NmSSE5rBG6OPVUQbaM6H9YvTQhH4Jvboc1cncx5Dnj
Kd40G+2wr2wpATUa49YYUQU8gtSPysN8LyqTtCDacVtoO60FeEeAjsmXhdvSHYgisefr1OCbqxoO
SIuXBBkbjnVcsbV8AIIdUUZR31iNABsaSKnI28fA09bZ+L1UlWN2fv1l5rI924mhS90Cw5E0YXSb
198GKju1SXdPuQ/iwD8PZ/GSSFxO7cLm/XCFuFYMiDXfXyuwd5rPLg6noZqNv/pxZZpL82JON+C+
rSFGbAlPqxV88IqktFCYPADSHjiOAHPguc/2/ksxT/gDKZiuQ7DyC+d8r3BMYP4XOdI1mJM2pttP
UhK57ydNDT83K9vzXM7dXRPtBMxATKk8hGjM9ZTP49CDtWTBXAMnjUPRN83tcagBfXFfIrIRWaH/
tvCV/K6jZw6mPS5MtyYKQlJlTq9aIxemp7E4BOwaU1ztpS9pqEQQaN+w49iGyp9RvHFVmuzjGUe0
56ygh1eFNc6qP4Y0EhbFQgp0mwvi9u5QyM21+10QsBuZ+X9qI4kPC3nJybqDtAHJ1sXrJjIooYPd
MlrDtiFGrigFh4Sg2tA8brdYA+2MOdPuUY4M6tC0uXcYzwnjnt7RxGf7N/uQhuM6TTafuaAmYsRQ
0QC1ZLpV0z9RTBb+mnBebVqVGZJFqQdXQXA4IxuJ2ncUDYwgLI4YPrF0BbyZxlF2ddVX25T0AIXq
sy9jbm777N6osRV/T7yeuRoAy+cl5bJlv0OkSZBlzFjDk0tGIp7k2bHUPoTH4tVGPAufHFFjLnvN
4ghj9JQjqrdEfu1k6/QER7qS7Z8TQGbDB6G9aqex1rOTE3A+E4G/cpsnEEhbVgERGjANxx7nS+SX
wz6LZqv8XnG7tzv3nwybR4qhuIToqpG4OnT/qCOMvTKheiZrEqK/LQMvTxAmkRd9FJ1Yy8QTYis8
ApAv/fdSitMkguVivG7/cT5YUNeKBUgsT1ZuHwebGuZMdRHc0FSA2ZrhCIkz5PQCzbiXJ5pTjqE3
LfYvNo4STb6+1FhDAr12gGGpPI6EnY/G3ZBoqrx/Ks3YJ0m3Yam4YN5S0tufruQJhQa49pt+K4mM
+1tw6b3cIOM7u8Kb2Zqy3fiL//O7p0VkAf2gxN62SHj1ZM4VOY5Gy+oc/nlVeRfzwi4DZErZCg2o
nHJhRtFciTkUA5e0gKWf619d+uhIk4jn5MXJzjbGeUXY+BscER7+be2k1c6VTjM3c0aoP1oT8rcP
BtshXY5cNH5TZ/e/o9nrNbFFbW3qCeiVcvk3bEH3emDGYy9ftLYMgA0zdXdshHXkMc9B4n4STdXl
wZ8C6gzfK4KWhRyJCfjCa6Rjo7VaHrzT7E1znb0QjqzfvEcFRthjDez5uLPqhnBlmOCnS2VqVyny
PENaBKkmyn2xqovlIqUnC1KpnTaObNGAs3CrpIDf1rQfahqIh0pLmMQ/nH/c7IjCCrC0eXcHlUq0
8jIB3c9JQU4IVrSmkA1qyPSEfbFm0NpedMEFE2oJuTZ5npeeQNK7Pt7KqWNnFlQxDaeOgBOF5bKf
aYoOjdAnud7kIiWQB6x82ZWHJPUHVOpDt87DPi8YVkGjO1Ue3A7R6X/S9AmwGEBFlMjIQfXnOmNd
tUsGrnI6csat2DqvvCHlL2dsoBtr++5ifx+6JmRyrfm2mYgpzYf+YyMdRq43R4vVrFQCz67oi7RO
zHgjRaPGMJQQtO2NByu7d3b+aZiEqf7YM1rzaeVPrUy1ng1fpPH5mH3oMV+SD2tymAhWtWHzHeUi
plFXlX9xa33vEodRO9XGdjM23a5IYYBKgt50rs3JtYBHjxzGC8XoB5VMxV1Tk+ksS5mU0MJF7OLF
3CJJIT2SgMYxJxSIVPDE0D/I4+3KYmZCA/AzV0vOQdt5wa+UAu7mhk2ULlJCvgur0cfRZq46PWDI
j8tk4UlYE2KG8GDBpcUfAEfLDffdwBlYFGH2VdOtumhx8cFByiF7/lW5XLoc7l7pYgKK846+/Z9A
8zYd1EB6JBXK+6eUNO+bWFgPnB7oxrHGGmhNn19HEiD/KHvgwiCm1nLAiPiCDY8A7mInxcp9HIyM
YhQFnn5Iu2o/3/OmW9XDw1TJ/tpAIFAKc/hVc3/G0D1Mxl07/9DhTUVpnx1nPoXeDNulzle2ADnN
TvC5DuwfZqexwGoRzUiVRk2n6kQhUdZqUm5T3KJTiwGzt+AQRPvbDd16lqqrGZI4H1PTkWVAkACd
ya40DPaeKQrverjbSn/Bl7487dlPDAgAeNsyICuI3eizXatN5qXzKW6CC62V8CdTcOMtWG6iEPy0
poEYJZWIg6plkQrEjOY4Qg7LlT4H2A6mNhk4dxWdJKP8JsRNxBpCokLc/dQdgRAYlL5ULtsrQbq4
TbuJruDyyVTXVbgA8DNls7SzwXl36gzU3qfWFn4euWIft2+wBbd3IRiHx29Z0OJ2oYFXZ6Trhw1c
7IeAcgfhMxclLHxNsBfHM9KkQ7mjgfjgJ6zjjX54EFdF1miw/lRf7z/WMPuemwNyBw3+RC/14zCc
YZuW4R/h1fWVwwtikTGCORzXPGBl/vlXW4E2aImaQ6ti+ee8KTfdIYF+ZrcVwScCElpmtFkUGJJS
wyoeafZ+gnF/1hXCtvbOcvLY8BnTVEJXXbBPvC82T0Y9K7zqPvXznKK2S++C+cWRrqXKWj6WSvgL
5lKpghSvduWGEIN7Bz2sD5zT3h0pi2iE2pg5n3G9ZIf50hcGzY6l8uffjEDNunERH18fnr9qYE/a
wb9vr4YBe9Nr58JoWcKylq3LZbx1WlnAyyxnep7hK/ijLM2l73AePky1G5eYwFJETN+KfZCh1mV3
rtqynPDmXdZEvUlMivrrwGu911xzf0UrSKGL6DdQeosFj0/atbd99zf1k1sygjaoo2ds80AhUV8g
brrkZHWyctgsbRoz7zkzjeTya181N/SHbbt9VSaxMbYRAp2ukdU4d2gOAb6GGib8pD/EKSAhtmZv
k6Pumz1UniUjcgjb0PklWr7o5WWhNKPeZZZamHSdPjyEb3H4qp7LxvgX5yvuhVqy5GwP6Hv1alEP
x7JdbL/fTdmR+mUYePn3ndHtobvIQBCs0Yv6zeK9Xn4jsXfXAQzUEDHJqwV3/wuESRCQ+PsxhWAY
uzxhhGF+x7fqblNx2maFrr5LuFXHXvstzn1SiZZNCWY5fkPW17BG96PKtDV+p9aIiPa9uMS3Ekdo
pm/l1LFPRYfktJmpI2wLzNsAaA5G6NGd3XGvDwZWM00j25T1erAqnvpXQsUa8ZoMecOXan0Z1QTa
/zPPhEjItmoK4ACTMA1SsdeaT2ro/AiMmqd9Al9tlyr6t0fbm/DYsoL2DT0OLLCeebfhHaVMUCH1
3gJSuYn/rhwvO1qOw2wKKbT/x6W3Ybs3gpUV738RZvnTuTxzludUmcVKHgubMiInS4JrowYsatwV
OfSv+tP7N+Y26pQ0hY+0wztt3+MN5433v80gRM6FZpR6ASgGKnloi6aErchu9KcKawMk/NcReKSf
JcCEcgB7YphSdAcw/rx5Zoh6mzsDEG/Ry2JI5c4qkOXC1gSzm09z3nMvo1lAEB2EJ9HJ9uzf6IKK
xpdhftxUb9XVNJUS8yC3MQZa1SovYBEC31CkElpFYwpMIsFQZSgRCOqRWSZBr0WbP+V37YGk+h0w
xmxJ6lLxsthjE5C2LAD07My0FZUzZl+ClKWNkSQgH2HZa6xywQ7SC2fqAzKjyoqAFPURH43B1SIX
hr6hRHdzWNJieNz9NFtHXcbeRGuSY1MgpYTdd5afTaNvYtCW8NSlE/4hcwtPTUzcNAx1CW0xrkrP
TeFaX066H+wTUipMoeDWENnH4vLCnDprUA58gM5cR6B+EUqrzPSfqMMepknatcpBEbASJlMvwAST
HxYlGxyl73UZh/WKe7xWgGNKkeKFAqJYuBIBGw2yIjMRFOchUkDtztLw2SYLy17RihqMx/OtkPhE
vzjnLOL9PSTdIIPQa74Xp9vL0+42U9c+gvgc39nDvPxo2s91z1A982KTJYJhYKY5/NKyIWiR+tMD
jsTprdeGqj9bLKq1t3R2si3GIjJ/MH6Dt92WiXkcEN/ktdW+QFMY/lV1+Q2rREOMnm+ibrPSiD0N
czpFQInA7zx+qyP0MbvrTsz2A+zqIu6BctCzvGI+hT6kIn32A6Fg5ltZnbthiFS29ojhzIV4pM5e
WFARUsGeHSyFIXelUxylsGE6UiXuZdDkv040ouH1KtTAO6TVHOOKCFm7YT1WPr4Kyu9zN6LIQlhm
e6mF7AODkW3k4HoeQ3nvwZpAOVmcu7xVbRIfXG8MaQfKeKGwAFqpku86M0RzwBLGFRBkrUYACCWA
vocNBwZ+OX0dCk6oqfHwcUKpYjTt4MD0n3Ue3XPbetYLeL+65IzBEy1I7eBetpGpQsRKM8xdnOkk
rzTusWhMcDt4tmi3TBKhQ2jHr7v6dwZKH+E+RA4P1AzR9aG64/+yKJ01erPHZLLfFDwjX1RhOqc1
831/N6c/CcEXelQZQZZ9s91WdDbayAFhya1MRw4qmi/hKwdnJy4gf58t74ff42kceskNMjFdXXLr
D7OoM+kJQEgxmYL9LjYiBp4VeteS7+yiiAOXzaXrd4vESL6t76VNex8GNJnbnrjoX4QL8B89N6gA
u+lig2SFRbQHdahhLw+YzTxpeN/tWxRNv6TXFykU+xHUd7P0Rs1QSfT2yifBT6xgJC3Awu3mxbhc
QPS83EPYoVWyZGrmq0CVLEn/0cffcJH8EFl1BVrkMMp5SVaLkgZBEKEvDcZlJv0hLcWyIb0o7elh
5NMe3urG8zIdO5Nc8mUs4sdKwuDhqe93BH8yd1eaXLBiLfPB+ugiMrY8Xg6E91S9g20qnx+H9JXu
syElykgGOGDiFQNDdJBVDdXhrz6D8iZnhyloGi+1FtVfxsnE23Ju4H8AZE7tSeMiBBeBwNFPntT0
CgPrB1ViQuheEic4t09qeDTGcfuO3yDKGCawhMjiqLP3FHlzQygiAvQHNyFDUHl3v0d5+7NxLvwW
PysjeEzbvpsjGwEEcRlx5/tKsEBWqEq9yivfadtRbFwcxF/5I/89urRoamvTQSLsuPb2ZYz4oi3y
ufP9t4x29hW/Ab/20HhXVjQ18Jt3PUCPbi21UybOhhIKwXMeVtKYuefF3lxpm3lV6vqrO65HUMgs
TRYroBPMgSU3PYRSKsgFB5EfMi6foKvNwboHuvbdo1mYbQ0QHgcg8TkUwWBDKvD5oaDk1Y8vDorZ
gsA7x2ZBRfELDf6t8XBDuC+S87AAo0v2JWqrBiVbUy9/6iQeds2K+iPhTQ9KsyKN3U5J+ZM5ywL1
nTXqIutv8M0379HmuYMl+Gu1hDMz0zBRWq1dBj/wVDlzHHTTgoQ36LtB7vJk60yDtXdpUwqDtUGa
JWslKXEyNbniyVdTbIkV+FpSe1h/ItkF/UaDEv9orH19lmtWDdse53BgJMs/PRZ2lU+66n1DuCt5
R3A6elo51I7WDwL0B0llL2eytDnvhpGw3Wu/17EHTtt3DVAQLWedzcQZx7x5iXyI52XmT2DCctT7
4NWzG8znAgpkNvmrk3EQKsjkm4z9OkeXv/eFPPb/nUNHVScJZ3rzRPfR922doOlYwIcJOjRtpYiT
FTeEyf6GzvdlTT3vmyA+9iPudZTPNbWw8EyFXhOUkvK2vfF1f7vpE3Tlt4swdP9xS1zBapdsW3Tu
W0ca5wXrTeANzS3/vqLKRBIKW7pQA9mMjptGrOnAvpPEtCEEJtbVt0OzTC5BiybK7zh/RUF94Uj9
5ZoGZByCNLGy6aHL4aFnpKGgSLllAPXdU3RXZlnsGmQZTWhTHLbJDdElRaB86g2C9FaE6VEcH02a
z8wWMU7gFLCZyGCDm8/VIfPUwNl4d/ELPM6dh4TLUt6bYgf1lWhsY2v+BgbnYC20k6fR+8Rj0tnV
xR5BkVsSB0iPlLOFRVaVpVIfI26nhggJH9mdqSOdjOZ2RtLHOxF8J/xoRjKN+BIQUiNA59IKCAu8
u9gzGpBhJn0E2dnOZkNpYFFaryaNR0QrxjlvN/IjF5bjR8rA/edQvWdLHVyZwPzWuJbk6wuSg/Sy
BYom0zMMh8vfD5aTizLcjGlwlswrxBYKMGI0uQFapQ7xGD5jkmRI65RiJezy/9Ul+bqqMTniDyqc
vQRICtcOI6SDHWrZeDOdevVGUxi+ykthTRRPG7lUcrnOGXSsqS67UPhDieAGcX5AQ5K/D/lYudAU
oxWisyVsXV4pUeNVrUeqdH5PihXSE5P/pgHvgro+7TUSqXczZRl/7SBDoR+pTT3lyTKxYnnETsOB
uTQa5Ta9gQhYIym9Xnz7q8rdZcHRVDq65T0oXyQtPhhYaIw4RRnI5K+FqoZsQBGeU8YwxAA8AZOO
gIVTcRJcSliuZBeOA2cRYF5vFZ26QFIE1z+hs7xh+vRZoaLSWB++5ugiF+ySniz1BxQrh8y/qQ/9
aKQMXZ8As7yPem3XvzpaPPhdDoR96PpWIOHJ/FsxQFmUWV68bWVNbdJOu5qnWALJTbFQT8vx7JOq
Fkxa8q/h+vXy98brFXBm/Etmel6/KbzcV96FLZAlM/Yv/fEpT7p9m3gmCFaGhJqGPNN+lOBQkaC7
5k9VFCgAql6hEfLCfxM8nRieRcF6cVQrUaa9Fw4zZm0Y+yHViiZPsumirKmSmxMCduFuIeWk/LRa
3HPgK+TCvSyRj57FYUwY/d6Rlw+EbGNqtF/ATwlB11ozY6g4Kdb3kKa/vK4Hbv9X+6FA65Ut2C/Y
pWTffHCJx5Vi191o/tc5Az3HA+QL5Q/HCesYl4xsRSK6pX4Wk/fBpA5VOTSQ4ztLVnPJRl2NTCuY
jMPOdOCzvFs3bS9w+794UNU5g/KLS3giuVzYypfexFRM8I32MRGS5a5hABREx+KFTzADfE4nDfrP
k4jM9Q+wYnbzeSXt6Ja+Vt5B3q2WhPPTXqmGVpRq5RscUxpR+Zf75/8gRPRzpNyh1kRRt6s6qQ2+
nUDhvbdyQrpvsK25C8PlCFOx2bdyKS898OHLnIxswmUAoBILo7NLr9t04yO8WZewRgWqFe4i479k
d0WzO/8A0O2purvzZXkzQ6Wv+ylTRWEBtKDcu+FHH7XfFX++5jUeZj/lausqiCsY2WRFeb0sjOOV
XynnJxrcVdoZbFEnOpIT5doxLkK/P+2J7ujl+M3VS6r+TPNrA5QBAM+FcOLG3G9hI/uSCLsWo9Sv
lDihgAlfgRA0f23Lz+JYaJtVaiFPwHLLsP82YkvC4mG91LQx7gXYbjoGJk6H/FBN1P6Q4G5hf6AE
mPyCAgD7rvGbCzLALW5w1OpG7ycS2FTxhsAiMxMjylNLfOvnjJp2/dv27cJykgr+Q2DhNh5GJH+U
x1x9YLoRDbPsLKfkpTtWXlBliMNOHhriB3p2gvEotNhuPV/iSWHmyRwFYBhqnBUg2kBE+hQ2tYNA
LSZAEFotNY8kA1CNOC0oe8JSbwXqc1Pjgjchk4IiIGSa9NYcLqax13NbeeDYSdUvZ2D46RBcY2KY
63dTmiNfDF8yC1b5QBbcVNrhlywKrdpgkUXQLzxPTl9rpJHxUK+NRehWxSyORk/XI4DKaBBAyKGk
BVtQ6thtvz4ECJWZjKcTwkhfxHhIfprYC48Izp2oAf1uF+O8KDTkbBTnAW6ZmkYCiMfPYSTtu0bI
OAXFqcXqa6C9cdLVimdNE8AIFB+2rUkWFtMgP7HAt3eGEwbgybFHnjbyoxkVp8RNkf7um5qghRBR
qrUZCuXpPZIyElYaWP+XZW/XhzxGRMd/S5dqrUX/HEvGicSBk2u3knu4xdqbKHCswyEMFaW5ISWj
kaY54KM/AYTOke7aCvjlVEz6P1K2Z1BBI1sJWGN7y7Ly5SUK0coGDKASMEFsTgVY+GAJ7ITQ/09n
9pTAvbHvC+K7HH+0jzpngvXoyjNVco0sYr/03umNogd+o66Q+Yc15Wbv+ZCRhNylwQmMRW8Cw2pm
xYUYrcs0pkt3Iydrq6hkM+XK8rsaqq65z2vMqEOhjaCBocnVbMlx+5MlL13+nZbDczSv2W9jtAUn
naUUVB0pV8EalPBMeXZwRCVjie1KAAupxjlndFvWs95MdjMvmgM52bUb1dZF8vulEq2HLo4IoQRZ
Gubfm9iZhgb0PobfeYAPpdRw7/QOdxLHseSad55DKjWa1TWHLQjL5QWOsNS2PCJ3gNK2SsYBWN/7
gEamZtIxpehM4KWJWNfkmRAjhrvk3Evi2RMsGg98zpUmhtGKZHLC/C9DCjdHUX6M602FRm6Ywus5
1Z4jYBh39/uNuNKFYDmAEgwQzEfmUkFhoSpz0RVCQGEnYwf/bOi+93Dx2QoOYEiqIABwRtO/ZxG4
wU262oW8BnuF1aUWsVGzQuSAfl/ea9j5nTfBjFsxAaUA00byGSkS/dXx2P9M1KWbvykVEVUPnsy0
dafDG5SVw1KDZUyJcipwhp8auW6x2zwG3v6u+Zzf2ElOMizJibW1IlksbQbN45pA/wQ4HILUR46C
2D4MPsXE2pMxLhQj+YFr3XgURzneH/PWtqCo1rdFYo+MX4XCNdL4+IUi0hJwSXQXK4z9bG8yg4cd
PmRM4hEMlryqNbudGRlP1WO+ezZWETrZKfcvcZ2d0mFd7FbpOvtLfkl/w2vHRJaifWwgaCwX9rr6
9thJrFOpSTmmw3LJDkR4hZikpA4uvPZt4s/svtT7NFCYHaWJUF7sznHwftCmsKSZhWOuADsQk85x
kiYVedqLty/iWCxIhyqqEnSHuV7QMnzg/c4ox94NTecD2isk0rd2U+lBm9fzsyabYfHQwOwc4IO6
zYRsx8hjCQCfKJ9lmsRTmhy2/wgXcSNI86NGamQarq/0adQhCFQJxjANUd0IeViMZm0JHLXT7GLp
PNR18HZy6s+nFA4to7VbmEgsOnqV29D9/Kbi1fIsrpIgbDjqxpv991qE78En8yIQF/gQVmvZUvIe
f5PchDqsygTBpI/DP2tjSxVwFJ+ZTSWLH5nBBn3IjXU83Kh9eo2CYmhLzJD7OGgzN1c+d6fIAQPZ
RDHpTzjCxrGvuH8JLW5n+ALl7radKPenLrGkAIGFA0IzZrYhkpNFWrbv3krYHZCSB0R4q4m+Lroc
iXSffPNbE2eOURY4gFeerFevPEIo0KDJzfSGgeySWQvde22KDf29T9Pq/G68KuxFnIb6kwKhbgUT
bOlX5jIfbvfTlb+dT0N5cQKht0Xkrm/qlT91k/KPZ+hg55rQfkK8Gsjxfo2KgHTuHrsPjRW4rgkX
oem3DIwVWIhA/lnT4CbopcmdiXLQmfJ963p0kbW/jWKnb5Qo35F0bMHgIBrcslc/eZ5U+CvYy/td
Ibzs80OfU0xplS0S0vdNYvLEf9WceJXyR+s/Z0GtEjVqqMrHyBNHGsv32l+XuFjMKxB4M5TXZ7rH
NEEIOx1KcQj1QH3L8rK88Gf4kb+/JjULNmFJjwh4NzkSW6IF/uoUfxj9bZvdOGxr4HwZXYdNn6on
6c7dodnCe/qEtEf3CaFjVoUMgy+01mMU18xiOE6ZVR3rLORFzr55p311CMmI+m2n5Ti0OYOWgRRA
hYaFMXIEHl1nC3soors+X+2kKNp3QeuiYran+qThrXz4lAFpVI26HdNeT7UhEExWIrO8mIKvlKMS
uuMaiAsWg1zC7EANBlOUTR2ufg1Y0QfyoCkG40jvZiMHL3CDYrrq/SzjQNxP/+Wc0pvAEtJD2OWg
GqF+25eXxFu/kWY3Mq+swL7MDxvkiKTs/GmT3s6v9vOCfQyaQMhXsNCbnjGuEShCXDN2nllWu+gu
lXspjaItQEvln0febYTguu4WEgv6s35a3m1ClSvJLt7BqF3i4QLW1x1Zmecwe+4u/qM8OjCV3H/3
26uwbEP9yCd+XgjttLeYrkDTIGHMwcwcIoDvaD8RB4r2y1mAeEwVUbkjgodwiO5FgL+e/NEQAv8E
y0WOfF7m8oSbcPzgaSRWoPuTuq+m2za+ur7UHtQysW3YhOK1SnVOZ4Y0in+TeDbBaewn/COG7EqV
nZ7yoHWuq8S5ztdzreLMliZ36+LwZmNRTvL0QoimQ/iSw573FKEVfk5Bmky5UKBf1F0Ar6O1Ro11
IB0aZFRkiNrvLrqooCEAJZUUvxHJlipi2PSE9lSrk1I2D6uu1kwFc3pl4GBaLNMt1bIF+aKSfj7P
wc4HL/pHJrOCZhdAgbUdJJhkDq9slaThWlLDvpCgOLO0HkbcAAifpWOOM2tdMN+KCohXaZL4Dp/s
lIFZSOB5DSAa59b/UzpI9r0wMQEabmT8AL7vmkOqYFxEGVVaIYQufN8865vdw0xgSOgl2coD/ciY
M5tPnavpyaWkkjmuRsXka7sE4EKExICRGGfHvtWts3qCbkhAmU3efrTrCNSeW8CfT0c66LpJfgN8
jgQ9DhkvAC4bXogI+1UfNHO5NSERc5OXTdFGFpdRLtzBl2WC34aRzPC2toXiMPFlcar4wGsmKTYM
Hszd3bz2iH0ZeHdDP6AWA8MUGgLnkh380jQXWeyGgtiHPsddtOmn22diaw4KguvPGU+8oBjaIf/W
mL/1JCcHveCvX2ZN0TfiSKsx3M9i/ZDdWMdV7HZurD4JIYrjjYAdzefub/Y70V6TlB5DW3NlAJ0w
6tZ11n7wjgoP1K05nnBJeP26cCyUZKTye4UfOvzV315tnaZkf3DEHXXme3G91sw+rnJkY1syVDMh
yaCqEk8HzNs/OgQlL2d8VmmWed05E+KUe8GFXZBRhuWBmLEoDWLkCZqwskp84Fn7oMqR8wCa4Y3Z
ZioI3h0eT2uug95T3ig8IgWfJYHDe28213S2gxl48GJRgD7TwVfxK8metxppewNVzQhY67qOYTOk
IuQDpxsCF289uTm2O9BnNb+pxllC3gy3SLINl1qqrMg1zDFwLaEDSP3JKZzXDn6Q0/GIAppLY9HD
sMmmuGFgxr7h3BUXH45cC9PP4Q4oGWPWdwzsPRFgjw9Cm2lOZto85A7MNahwaG3HPE61ptZF+LEi
4Xr5h1ALZPCZkaDCgTxx9anImgnm0c6lhZvQOa9yFrSwpY3cgYQRediMrgeE75ujwClhYy71DLqt
QVPmaiTTEyvCywrmbT6ABM19tjZAOEMuKyaxgu4jXkZsRW9HOXV4jtFyiwV3/wqCU7tZkvTjSiFV
Fr8GQ14T+MdR/dvn1BnVF+Bgi6maXG2kjNbNubHq59M3MWdPYRex6hCcu3qymPOdipCkM3TDn5KQ
vXbFejvTw8ruLas0Gx2iCznWKakbuxyMoRTZ5pn7E/IrJjHnmrm6Jih2nX+QGPqi9/GSl1qF1wQh
f4R+ewvdg2HdYaMqIZICUHBbEH89xdJ7Gy+naKoDq6wWKuKEHd/5vuvPtHMfkaIs0pLmGOG7JtzK
Ds3rLjoaxwIT6CMqiHZ41fXdsUdEMMC7qi8dN5A8TD4zyFx35yf1zMNBV5iir6kzx2UP1Cc5xwiy
zaSm//2BkUO82KmoSuUDLJcQKnLSCus/G2E/XoZC9oq7U49pkbBwie3h43jPQvNLM1w0R7k3KCHX
vJwEc53FdItjIgfSyIBpLZ/nWBEgsNz8in3uEGfhMwFUZlpTkBEOOaO2TxKQrMRl2oS83aGK2woP
SWP+bmfp+wbL4KFqVbmB2lQynEwDjkAIrDRf7sS94wb6+PIrKX1CrDIiVJKHoDkJ/NPC5kSpKPR3
/9ZEHzi9IMomG331R5wGYz8VKg0v49rULfOL8yiXGWWImlwOEBJkKZwpc25AB5+lS1LHaHeO2zEz
0RT3Y8ZMVobWSN/aSOQhAApjogpzKYtID1yKKMENvh46dY0g2kYb4WC4ns048dRb+sO3LX5/8cGZ
w749xi0knp0bpG+v0o4ZTvbwEVnwDq8Q8A3u+pLRYhdHTmt9AzBIBARXo4Lyjoc/VaQbO5eKAQWc
foND0dxnRvXxfGC4/iMvLY/m1FypfasltifsDmQEigunkReMva2EsX1ox0SFq5TF05hj2xDa5pSR
hYMikeWlBdtiFQlrP8czJYDlJ3fuPnYsM4rsrPHSnAgDKSoryZWPpOqwdQ9UguBNl8zBQXpvvFLm
uAZibgSpI4h2caX8xemPK6ZXMXgcadMGqlF4W5lPDChQLaOnR9FYJnmTmF3k+L+XpKJXIniFeTOX
eTDBvfvrdISKGymJyNk+t14pdJM1jvqdy3VtnTT6K/RwU1mmmvBR2E3IxgstMzRVsaLNMp1pi03C
K4Ey85876g7aSX/CBhpDEkqzK5VMmW8iDxEv0X/E+Wv42DtPgPXz1VaiDgqdEPrZUXH7ABuj9maF
7M6M2LT8Cx/XeN5J3FU8R9qoMU4daPWmnJBvkc99iy2Du08U29oQ+JUaXDdwHCB1VkcD1JjaNQHV
KmbSOOtVFVVhVnCV8W9oreV62VDIwAzdi9n/1BBLQVw2JPjaCBgv4DYktPWCtb4xwukPs38krMR3
5rXG7PXiaVfAFmD3SHG8qOKS+vBXHZwWuleDHp4dWLn7f/eNPNtDA6EiYh0XP+bz2qwOwIfzbiGw
SGQvXPmT6PCPTvxvcANLu6GNPw1Hkq8KfIik1WenbPUUAMiVuQD+V6jw7snYyTH0TsDL/UYZ09VS
EuTtVsPPxfalEGKrNwZpBa1yGUNII1/XRrjwxwmjd9AtMwm5jKFVqlKKsUBjRBm3hv4oojObKw60
6lmlboJAqWCj34MzGPeB6X5Ihdjn/LGMLQnbDfWosx8TLxgetZsq+94FbrIemgoNKYvAaBlJmrg9
lItnKWUVUwre3873PgBWH6kKnULRimb/xJwue8RWYcs7VJ+AyUd85XssWQpOkMcmfwK6Gk2hqu8g
6ZRg/rssGiJWc3dO6ukWsdO6UH3OCEKaPJXenLD0AlqL+ffPSt3neaaDP3NHZ8rfi3Ly/MDlxMrt
eZHU7VrFAFus+4N++y2bMBlYViK+rACz3dmVChIEggiyXoUvZ9UUnHv4IcIgcQcL52QUl/zjWNPq
SKjaKvv1LxlN59TAYbZnCxplBjn4GOpqnsEL8mLwgEiB4KK5tA4wzX8MYIeNVdSBxlbMEJuO5k66
ZOr2Egb9XHG5L08Ta2AW5UOHJX+Y2VKDZktwZhkJmIHJRJ0+EhP8c5fdjMb4TmlJwq5aXhCKW8SS
N2KipWldwX62mlpD4CADyGSk1O9/DecCQ4l4E7LuGjNObhroWrcVSEkFK02ZQDPMRiHWZ8V89nM2
l40ACi53+4jEEzNwS7S2h/bUCSGQM/5ck+hSa3dgjbhTdAQkMhKFGSLPgZYhimM5ivDLgsfeJBRI
lp0ZW88DkVcSKJfe0saYJ3QYJDeH9X7SsfxPKWEEaM2NY0AI8I73TxwL09gnLzqhJwWnMedkcMtO
sNE2mNDf4dSLeBtA59lXcz5T9gwSNYU2QINRkY12crjM2aLk2oaOkyX5pgmG6OUXbJ2DzVuFwopl
UHrCh3Qb9JFRLJZ8uDfs9PhM7yVnvZ5KjoHLxjSSHMbaT7+TA5yIROOQHXJUV2LTs2IeS+QSax+2
lV1n3TF1mDLJJuUuwEFennJViaDwTPpKY2h6Xw360dwhpgZDvKy1C7T5XMi473Zbf+aAzXbv8IVf
gVKFS5AJX8qu688FYdu9eimsameMwepGxL31j9bgNYgQ0A8SG4N8agQTOtOulU981vZfvWmHeViK
iN6VyXt1gtSj925yhiu8HvbUoQ0HVUF8rL07W2IIlW/rvzrHitMl0PCH1COpU9/78z5h1m8EGzSz
sgiF8pfIiKDSq5a7HG95POO905vveFrpBm8hdc3gQiUdycNbDBKcaH4koqJ/VfLe1ti6rWKau3oc
vNjqTIQAcBZNivy2DV0leZG3oTduLQV621IvNq9J0PET2zNguRLcN59ABSK17VsQ5VThMIvsAV80
i+1kor3AlsCReFvGxoFyzuX9arTl8zlPlFPM220jU1kcnfr23+8NfwyPd+YHPyp8c35lRV0otSy4
SXBpiKI1rzVWhbxcrI65j3Et7wlo8Zf0aRqO3G3WfHUm3hHWguAHmfq4HziTkgoGdsNdcFPOjjYs
oiap7GpjAEu8ZCgWOnLP8i+VCbLS7Lg4xkxKdC6hgfdTV67X+pnYclz+MSLWlhk8MrShL/lrigf2
JZZhGZ89UVzpI10843VoznbnOIF79ymPpG1C3Yo30iXVmDLotJeDvvadY8uT7HZi2skEOlOEjYBl
6oAQnL82huJ+JyJV8jJvRbfEvEnOe+Sbex5i7kJL85PkCeIYda5FBjj+TJmXC3QvPMLcBK188XaF
0gBT+b7bh3D1kiusiIqGJVUsMFL3zHS96+FeJj2i6tBM2sO3tzs5ak3YBa5CbsaG+Yj71uf73z6D
8MuXkIElO6gn/DoWrv6nE0+J0z+zUbMJJ3/QhEh4q3+l4nVI1AzA+8QOLgwd0grVgSZKX4BIHHI8
GSmLKuYoC7SsE+4XfJPTPKviBdcQYNGXe9cOae1mV+drvkDJT0kBsZofkTRIiqt1A9ddf1ICLjuy
zIDWHbyPG+7q99BxtpX+j4v4fX+fThZXWwnLzde09NMVvWmYyFKLydSwoY7/mm1Omekfu91mzhWY
uM/UjvvQj3SiDpm512LhRcQPnkxKRMRTIY9kiSgoUkv9r92Ra21E2WGxvvXOMebjwoWR6W+VEil7
smb8rGBxJhT8Cz8BCjnHuRgd6qTeom3aquY2aPjHxEPMU0nCh11VPWuzquZQ0JT0/z3zbTkFgkg4
JZBugJvwP2Oz/gi7VT9YPBx8UdkwQHDHv6ZGqPWf8/6y+JgX9ZDvBKB7qKwgRDTU8SSz0zsAipVx
c6v6c8Aax0NkJXmZhjcqKlJJ5/l9mQnY9NiOMzfnp5gvXxgIxxna8+2uFSK6bEn92ofghA9ny+VO
7xpTQkb+QLGu9lWnKz3TUmKVJ8lcx7FvgSQAJO84YT9ftEDswDCVfB4rZafg65euP2d0kboZWYcW
/UZKtZ8Buf5bvmHDyf3W7ojt46FLs1dUNdnwoG4MS4bSvsSE8KRpOoMbpjEFDTEXDbm2UY7JwrAe
WfeQXWeCqutOoYRxDqp9C5pLzGRPA3PcicwjyYT+KY/JXciFDWYYsidbq2Dggd2b4AZ1I+NEEFm+
wtZ9maBXKs2xXjL5UO+Mze2ZwBxSN50msfC6CjgFSHyFeEYwjjVb8QoBZ158+f8iWnlXdznMHAZR
IXx+ZuLH/R5KPdtXiEjGbdJcREr85YOrisHGi6WZvrzqi3ieSU6fE6dH/lDnYWGFX+vEcjvE3iaq
vi22jRAHKnhBlfal9qMm/uF2kjrw1MyZx6Y90kE9IyEHKYmXsaOpsFxetD8EXm7jawNWJqR4nIVR
1ufx2KXirxnAwBdSvCu0Bme3hYbO+w5zy43GiRKWTBnNZFOyhH/eGFckz5yvBKNamvhvpBWA+BAb
9THRDyRZy8OF34TIMV5LnuTYKGywajNikJcPhHHYfuYIG1QWqB0RGf5DdwxZ41lScGgIfjZn2J3p
NSMJTa3EtSHXhYXreGv7thk39LaCCgenbsVUeCfkF/WBN3VyxqpOszhnYCkH6qfmk2Pi3DbqD//K
wptzCdcScDdVsYe/I6nE2aU8lbPjLtWy3RGGjH+YyyA3+phRuUtL7b1BBD+0ApikOL5bHN7ofc5N
hmXC0MsSomJhgZleobaXmAJrMkTftoXsrLgRoxf/W39tjg7IR3j5RfOJ4c03+kQ3UiUy9fMR7C7y
Jendu0/zHXWqxw1scodlhJFDC7mKMPn5EHaXPYT4slCN816wa94LwQ6HZJkXffIUsBOT8tASMjNv
B9jKBqgPMlMYDxDdftnrRCzjwRNkcm2vh9588+0aKQ9wDRGn3Xcg/27Rs7cFIyDidxZSo8B96Hsb
OOBr6AvY/pcW4wyHoQ7C795SxXMH2xrOtH7z1rj6vnFZly06y7F8t/pS2asEBtES2aMt9yOTOpMx
WyKDd5+9dC3VGjZtHnLVwAbv7Ss7zQ89qr6iF7Cg8E/8aZ75DPljQB+Tg+xz4HmpZr8sfXVIb3Gr
qQRlnDZPqMQzgFvGHNxr2/01u+HS/V7EN9btEBJL8ESt4fR9ud8ePYi/slnmtGydjIYZl/wlP3E4
CDDD3YVxZqVd51Ln2ub1WGLKDWROptDUNHb/PSHo6puZJIB7UGOmNqrh2v9OeiE5iq5wpLg5aw2L
+5jjVkP/Q2Yy2M6qMkeesi3tfcKPEeIcxkCVxIOufqe/xMKs09RRWwO0daYFT75EEJYcsWhNZUTB
Z3RKXkmuEDF+aTLeMQyJSMUZEmjtDiWsQl6mfvmwoWkazGl3qGuzFOkgAWtB4YMHG1UyJSlBqSAL
p3Pqq9h5YQT6ZWt2oW0iXVrO+d9nGtEK45EdLqhcnN7G/bCHN1Ok/qn+U5RzNGA1diA4Ko6PBVDS
MAqdhiikGTIsa9hK1WH0gKjD1LESGsD4uTSkGHIuujT1vqpKBrIuy/yQg5x4axcyqgkYkkXpMYpY
+v12EBV/aRw5DLOu4Ktb/fNNd1hl0nbbgzPJLDDxdlOmPns5HYD8qk2y/UrdzfU9zZO5nFFJ33SO
fzcY/VRKsuu923y9M1nnwlH/UcYYkzEQh5xX0MVkrX84yphqqwZjqVNxgQclUso6bPbEctNYAfGH
4s4S2vwJjGuwZLgS3JwrQTSR4Szxkm7FJiltMBMjDkPKONLkOkyDwUFjc5+icEyTwIdbsPUnj7eB
xhqn/h69CdxZKJD+XfbmBSVnpr3BG9tHxLUh50SjMgRNqZGChC5Dixe00shWjFpWcOXZWNWnJlG/
urra84A1E0RCDqvTcMsIN6ZwlLzhSSK73REDYg0b1lpOy0f4YKCapgISmSNT+4dtZC5mBmb+lR7k
TLko21RNphSPRTxzAn3b67LaM5FjwI5jlIJXxGUcPQRHkdOdkZXPNvNEKB2gySFd1aOKaR2ADZKW
iIeTKYyzS3Fi4IAFO2rAfWTj7QYpTH/Ws9dpwEMrdzKTmIwpNVdOL1GtMIy8KtGpJOKJ4lvUOVxZ
fLsa9EakHh2AnBiSTFJzWoYp0Wzboq1o2XTlunlaAOglsNSMG3HLbqgw5gW/gXFA8UifHB7VuqJF
JBr4lkvqNAtzdqVlKL3L/a+rHSpeL8/PQnFPtVktWCC6ZKrCpXoLiCkMcMF9noJzK8hR6kXLSBiK
agdVgLBqGpgF6C7Trr1CWauNf81WZ8jjccbp7ZzRl6HP/bBcsW2+aSYpz9xaTDPx/m5hT5qzCtQ2
AJInexQFJjG881SzwY47orWvKmzOxHsdstdnvzs7gYSwyK2PgEBXxyeQ4Xy3NAITZ9fE2OQDV/Lk
s8ECd/IBZQ54/lhG/GdaKhtz81h+NSxIAI89hs8AwvMjnNWO2ezhpBAuQCPhvwlfRhvSGhnkSlvx
HRMOezg3tli7qR23embQtBafXO700MOfOdUXy/lkIubbY7NmkLVrmIw82I60kGyNAL5ob+v52Mzq
NUu4S05uEhETPeP5JkH5pQ7QqDcdxGsz9DHp5MPJoXC60gQNba22+OHNnSA6bsvJlBdeG0dN3Et0
IpChpwZ1NHLqRjSWpZCFJVHfbQGoLTVB6zzpa3kF/co5iDHgPtTxVx5DAVx3bQbzreKpQ58JzXe0
RymyAMVgABSERbcTfxyoJHjsmlkwAi+UH0SxqSog494tmFr1ngHEKAyBuE8mdzH0l0CT18qAGEBg
4fWO6twCQHNMQnTa9lUHdzmvjGp0hgQ47foAUJbTYJOmd/dv+5JxQuhwimzugxnl0veA/CAJKfVk
kjeHC1tfWGuk7owFiqBKo+EDfsVpvxP+ovFRsyB4fK4pCu+s0JpBrhpKKOsSAQdiPjjF+b1O0qVb
CRyJ70C5BXhpoccuqKd+l0yiEluPeNXI/UBhRzbs+DiHH1vf/QkKApuXr0SDGtRF13puogTiT1FS
nkEg/h7cyvBmiM/Php3gD+ELu79wfmJipcNuctk0ruB8r/lCOtgTExI9s8hLr0FEfJaGcLwNDbte
2cTGuiPAI5T8a2rsiIShiy1d3ll34J6Yup5ixyxoqeiLNOeJzUMnT+br/xPQVcBF2q5SsAQG1aRU
Kc8rFZO09SqdhmUUk2p5N7JpTDuqiGCIKHsJGM0XSQt6A2BwuVfNP/BHnl8cjSvmc1dSwhionU36
weYZeAJi/eTeGEZqMpY3Kd1aGwj5hqwsBoV3zH8CoVNuBwZzFeMWTwQWn28uZLfAh75x/Tryud9o
l7Ju9VM3ZGfdyPH2n6pL2Nlh59OOXnwsrXx3gvZZD7UhH522AxiSysM3AFrpc7lZn8TVc9Xsqh6E
lOOx3UhPOTbcWUaOlk4HAFTUoQXnK7mU3MgecA5uMJpQOLwQrYcv3zNTkEjLkL7TUk0DjUghiUAM
jeVr23WCvPgONZ33iw3AC06i6z/XlenJ63vkUWKxO17SacgAldDuB+krKK/2NrY0MpCA/Z5t/mBj
MkgM2IZQ28bSzXJ8U/DJmpmlBqxKfUFKgvTz0zlGd2C7Ei8d1QmwmP5mVngKVu3CBKhzvbPJS5GO
+WuEXi5OkwAWI3x42HczW4k3RhsrUcUGA61SyY/lc3zZOsg70n57WQcz5lSWwfosqNzxFx9xqHNy
33plJFtQn1+a7aMZ3LuI5hfaXwSV8Pd1AJF3Fg29bIXcPvd2yhKGwuWp/6sf2FpuTobPKDx2+NMw
uQiRPZK2Kxr2wkfRa5E+cOhNtDEVIbjGV8SteVmd3I+XlcqQSod2X0w3WIj0i7THEWqfyOJ6F0G1
ZkiTVXucGICmzCEKQzt4B/16+RIpOMjBDuaOyiaHAL1bAqhf/wHxdEXTccVd74BePzCVLwQ+ec2E
NrIyuC9fQPOc1h8W+raXp56YhNIQPXEsfSt93n88vCa5SRWevFj/Bh1fTq5omC3obY+ic48LFhly
VyM5KQ/hiDUt1XHSKn9BLPHqzgD4YAhtndYw+PQavp1IoUEga38tYTxbdCxMhqo7iPy6rn3TybtR
tKAJ+FNSR3kkIVJiL/n281tYH06z5kyyH60pgwnpe44/Elty4m0DTkUiv+L2YEKAl8yTTsfVP2AH
NRtlKT7pW08Xj6wmFewWS9tYRG6pffEOTqKM5SYpEzOyevL0u/hTn1TDZJTBE2Ea5DD1TA33U1P6
PRm8ArBB+M89NKCDBRscCBjFBgcDltAfFg3pntC1boYp/9WW9I47bc0GoD5Jxch5i4TEmSZVGTKi
cZBXh7sQ1iberRF5taaAo+u4KjCqp1EIqlFqI4PelLNaUYibp0WyznGvvHoTredGM4H2OzouQWL/
LaBIqfESKbiysUBT4XvYZBqUvLHt9TDrmXiXGS9ilGothLU+UnMKj2c4IInY53cdccnbDZrAt86q
DOw/ostQPf7khi1Q+D7abDOPQ3NeCFGpUoIyYEmt9C3vD/b3Ak93YlHMIgBfSCDugK+8HH0IPJtw
L5GY/Wuzjgl6CZJ+t5HvCx4G8EaX/Hlgc1svt1doMd7b6XhpmG//x9B8wCCnnjgK0x7nz1ztVOZV
KoaUG9Qa+JUYuWy7q+awe6VdGM4fdDatwHEpiyC2QBTTbgbapNbEsKZcx6iVLrQvZbHoAeBtv6Yz
2kZngZmq3IXN2iIzOdQ85ohq/KVbzBwiwRaqQ68WGQWvXr6aFdxF5nlxC7WWMvd3Nh95eDLe5jmK
VC5JrIx3zfoutBWGmBGdloSo6bkaACdLPEVZRiMmwKHiOAcxkxjL+E6f0pOP9/zUHK4/Lfpsllfe
19+Ob9XwJIqVGoc2uUEjrQ0Zx+9qGbdENEXKNgngpsyFPzra66oZBbTma1dtUo5VulA2lx/7RiLE
z+v+eeCYXADOyYTRAstvX8DoXzYbXmY1gOePUpQ3eqSucW0VbMFZUgmJgqhh0/URDwMMJzSdNRMQ
wVmTPJobZ+PqFmiu+l3SL9/l/QVM6Kh0NWe/VT3Hq1mzEHX0Pb0fdWVGl8yaJsrzwLR2NoGOXc/u
7/EoZaLMpuJ4U2gPyYuqI48e24HDJZJerfhz+1CUU5XiTRTgBYmkePIFquG3tni4uF8iQXZUtZDK
uKB18c/A1qt92+lMMBPH9NqgIBt3wFgiv77ujkp7KhkP/rJtpciJsdVqSPC+/H9fEq7CJZBCSl0T
i7nSDV2DNEhTXdHGve8EZbyeHadxq8WoyOdLX6EmSyWh+MShV/KVe54COsjW+IgPQZc38KB6UBUK
KrLHny2b9CnynAsAjE8AjVngb+5pZjXDH8gsHF0UihXuC8uVC8lawZXnaI3Q+phqYY8gyxCf95aI
sRg/89pffdPHQKZfw02fJlQzFj23yDMKfh93f7o8aCJXfBEMZ4tLsTJ2DzlbMo74cEXJhpuivBIz
UOnC226jRVW1tOiV54ClQIcweIRpXoXa2J71evjQE1iw0HtLmRcIasO1a1v4zTOZwhcd7XDvorIq
pd8waDBXcWWGQE9k/IvhEi8L5pVnyKffXGBY4JUPtW2J33faCEtorifO+DK2dvZXAZDnd04YHP/8
048NMhDOmhPlohYPrBpjHqSJ97E+cBD4j01ky3GYh5X6A4LZfmgO+ALySBmutnzS3C8+D8VjN0Fe
BX7X/wJhM1wxxoZe2qe/jH3TCIWa2b8QYnPGjkgaokqGIMbxGJC3Z3zQ80OIfIDd94WSMu47ZdE1
fubi3bn3clK3NVCJYpuUGzn+UhgwOXVlRGMzWt1P6zGcOmXY1HoXjGCOYE6IZvba0+xtKjqn36g/
T+Kiw8F3x31uyOdRmPK1A16422XSBKuSnYr5+F/iSP0OoC1NsvmSpCnxTBK7Sr+oSItm+6fbbyJk
fCitVyV+/Pv/50Ujt6l0gKQrx2YeIQJOO7HF9Rxc5jD8UxOv7tX9ecG1K7uX3254w5hpLQ++w9xy
Ot9H0wosCCRzsJbOdr3FVr28mSjvqO8Q1iSpnXpHZPq55oCkeUrLoUzIRGh+aP9H5gPLchD2LVyj
uZIq/iz3o8lYRBeT0L1I5RnL4S6UV5a90jgpm0+F4M5YkoFM6FKQLzNDvrzBmKos8ewyu57fy+ij
WbYSTbxRxHLD+XvexqOCwagrrlFjGcLXGbNNrjNE9OzJVGDLSeuawTpu/IINI9kG93Wi5AFd4O5L
j3WTL4UmI5Sg+/AT08W/dw1nyqAHnoi4FXwRCmSBi5+GUhSpgItkVBWOcKeCoTICucKjdUyat2b5
mAYk4UtrMrX1gVVBXxzsUzZZNUQ27VhNUz6Ngr4hEagJKv5gPUURkrW4ja6B65RhLnjL0vTsNEQT
KpL0ARIUywOpvMWBTzHdfvKXQK/KsK6ZZt/i5FqWSSWKN+T1dexsdu+QzfSOCXzWnXZBfQmzE8mG
xd/TAgRXRRuAmRBG5LmIqZmi03n5dKHfOv2X4j0i1cjKe/75ZkuuWxU3m11Ko9m9a2BHko95BXA8
hxC0d6QANk/5vewsCYWZg16/xFJu+psbaTTUS3Q98Br9OT/ZZdy1Md8QG6Vsb0/zBcKBjpcqwHrS
0Ed0fOFDWhIXB+MvY1JvxI0DpdHpohOEpcZ8TEdGWYCCEKrI4uwWK6ncMR0JtvBGeY13fKWet00D
wlDmbKDWg5pNIsdkBBMHSRum2co7USYP40Y+q19iUTJmrOfMBzvp/RYy1l9OCxyx3sczGb9OYnPq
D+yF9BWXIRLvRrh5jttBH5QSsx14Qcf4kiVp8QggI0wWfwECRH01SfGZVKPzo8LBuEZp4l/DMNJc
+YVZJZ3GPsqpkBGH5aNqU0HyR6rAkYbmeUvEd8g7sXfHjTUDJ5shhU1wzmHb7nkpmB8fj0UyHAcs
qubobtFcNJz9efd+ZYy7jckCGdEk+2P3FzJT6OyofF0fmJnjzZ2z7DcnV44jkEWzqinBlsOpLWXK
aHbCVrp4qK666U6t4nR6lGYJMWC4MscGYDsg9xUvn9Ji4jSeQ0GlKTVHCLFKkS0Jmb5YsVZXMn9X
aGq1rVMAZOr1ZcehgtzILDCmqopjjiPg9wXXxucU2lbFNxu3QjOtbVq1L/Qd3aP4qyo1c+yRaS54
v9TAOsmKd62w3/V1Ac9b9mIc95YW4yriL7AdbOt83/tk/nlXqTQTvy/39vl8qRMe3MVV8TVsLVbO
JOqQM7tCbxmBFmbaW7Aqq9Y65y/XfsAlNqGh8EkXvBK22iomILD6VDXhOsN2L/fFf5IeHSP0LslJ
gHBl1wVkygy0H0xvIYhnOivIsklqvMDLh4iz5katbXMDE7ktgY8NQxEoZ7N4k3x6DWJYCOjy1eY4
v2PBWy8YEgETYOL6v50e0DwWqlcxj+YSpdfK9ewv+wXinTsEH69zXz0IkDh7oM68DeCsdVy0a6lJ
zmFs03qpDPkhDxRnNEDsMd2qrFfDmVfzlIx1TAWfdzBm2Au4/tErCtsmmS8I4+h5Bm3ED5r8B369
sdkVpR7g2MBQor5v3OPXWyKWti/YQ+dyy7xx1wP2LzH2dn1MqEuZA2+zItYrbcORklXtRbPf509K
0vCTR0fhhsonMHXIVNvX8o/OPXJvNjzlqcK/OPIhDNZXY2S3XhBrzkvQ9amo5+VVOdWs2lT1Mqro
N67TT7hI1/qcT7feVWUedZGjlN0g2w3N+UCI2QKF09YLSrY/TQLyvb5V5U4wtV8NRMCZhQN58dYi
JWYARQwgpurqADxvoHWoWQl/7+wF4puc4Q8SQ6HX8ewP1F17gKS9miIUnRV6aA4aDr19FLw063J5
saGbv+lXtGo45NLBcC/s636SaHwUDce+4edGs0qrunHSL0bW7OujuG7bJX7pc1R6NWE2+8QLDlP8
X1WQJ3lchnIu14EDrJl46Oh09n2broTGtzPVYk9amHIB0Pw0tPpLJMHWfUygXJSIA+1hyDEhsnQF
HaQq0K4Y7tdy6JIaR+kbS4RoG7gWjy3obgs4Wr3g3OhcT+4buIZrmxK87WZG5M8/guDkhoTffCEl
acTjI3AoQHgZva5hkySaZBufNBOsDBXxCwBu4ft5Bz/0MQGt0NmxeNwQeTqk1YHdWmDK4WLeVOCE
CNOn4ken8ENN7DmocLOcs/m9nW/uoMor6KNwHaIvtYH51pQNIv+XpDtKS58+tWjhc8IPu2nFbwg5
DQYSEo8VJEk1n+PM/C7wXhrKSmCjtZApDcBfwLmAoHoiT0gkNtXKSnRucIKYGlbhUmwzXIlenGV/
2js4T/1LmkQZyF9vsq8lmgxghNeOnCoPa/1wbiyK9vNiOwHMEvEyhKe4nxkOzWZ6dWJ5dDHwTkX7
LmezdOe1+1SephvGYIp6vJNevHKFNJRguHSWUGokX8WnTXtPMwBNx48MLaAtWkLADcQf8L8PK2kn
Hwb1TPuIja7Io6mdBB6T4Avm4Cj+7CybdhkfXBuj4674NZTOVt7tpCkQjoBYuWNDbpjmahvMTNXZ
JZPB7ThgRUgsXkriG3ty0YAr40fEFYKLT9N5fQmkp2WB5OXvKRV/wkj4Jq7GmZ9JmRazbRUWw9C2
T1j0q1FgglZ7T8n5bFyOVyFpcGvOrGAZYXIxMrx0EsEupSX6gE1tFKjgm+W/zCvlvLzBRokUqNcX
Reem+7AL2yROT0ACUrUT4GYXQxUUySMBaE0t4SSnMeOnzLlIgXVErXsBoWp3oBVJWHWJy+3lnmp2
lFnFRIpVJAazPft7MWkuZb7Jn2NP4mQQBIzBma+glgwuw13+zzdJ6/FcEo4oCMiuJglwHoPoHH37
eukyY1DFHmZPl4XjujUbY+GrfdRANDR0B1DOoxxhoKVFTMT1T1/7pRehl57LHI8QeMtMlmWVwnfn
Z2W2b5oR0D4TPQb4jUGLil+7B1rlJMf+iaVRqic/6nGZ7hcQtsuiypFotfvEje/t+dGFA0MrzA0I
XG39xDGcayE80227t6fufwg0det+mSNKWJvZ2T63bDZpUgVBwHGLwOAKdkYfNIrK7q4QeGbMyUhT
eQhFfx+3PfZFSAKEWrdivbUzF7V3GiUPcOfd9lrshqs98sv1/EpCxIoVLCxVTHbjuj6KKct96zfY
wKcOmSO41/TK7EoZn0KPqxGKerXuYuY0xVGT48qDvXGuihfgW0rcKrxylnKHsqhF98re1vOSs6cl
xp3uLMp2fvsDLBlZlNE+PVIDbUQZLZGP9AALSZEnVYt6zE5nPeaeXEdVnXXqd2dqaF7T9Ldo9yPB
Qn6SjnPy238kytkchSF7y1thiCW/PDQndO2A2ZrV3C/H5rmGmXwtuju6DLj8R2sD1SKqtscg5gCg
3+NmJK9XTLZYTjkKhSCzp8BGqnz3TAFvItVBT7Ll5z2DUyh8toc/i1/xfKsWPHNytJJzKEHQhajU
W8knmhUKp7PR2ibqpXipoHCQcmMajUXQNrSKij8RBB6piBzY/yvLmFCDcqiSYAo4etrEBW9Q4b03
sRBED7SJOytbXMD6UYNaw2mzWdn3UdmJrBNi6q75sYLCj85CPjcR9VvOBTAesZqhi6GdRdVAinCr
SggyyT7LBt+Py28qZvn3Z0axv7iRIdxUP20n4gxJGuA2OL+APoTFsetbCKb8jl4B9RGFPq2QpHTE
CCkUBsjrhXt23YkbVTlVIgv8rs2llGTG5sP8I5z+iq2QJGOEzAjWvONHE32soRGJZSnPh1cA7sI6
rnvStOktUOXuWT3c9pqZtHZhiyY2lEEXqQgvOFHcOhpgnTFNY+F57YXSj1T4W2OTeLzGYT4ekXdT
lumffxAivk76uknAOTN1zhmyqRV9ezHb7KK/rQOU4PQS4F/XX5lhvN35ePBqgx39XPmvsRPfgzdy
767/saUoFDOXRJsUsP0fkHpHC3w6zjKlqZP7HCS/uRiDZKeAA4CehIiD0g4YPs1JClNWn5fdGnSy
wKY9dyb+SR09vMh21v1/h9pOHfq+/F3cjUrTGxYL8i6mn5lvLa+5KCZZPxnCUOID+ZTID0jj9WGy
E2UnI0C16BjTQ6VBKcm7hkiTBxCys1Ha7iA75h0etRvhKI1sQ3FLtPtfPTOFacYYH7p60zKJbUk7
vKWXfiPPGspg4U+PdjAmYNxyWi5LyIEI2XVS0DoYjiT6+707c+rRhsj7SS5qiz4ZfVkxiuYvln/s
anHZaDSACS3nX3W+ArEJNzn2elv3pZ5Fmq1QUnvDnOQKjemiW5+vKYCHRWTv9QZHlycgJIBuGQEK
hKfGwVMs91ziukkMAJMxftAYBZZCwnBQKHES1mPI2dcyzkubWvKdbUR8ivfnYXOaorSz5resuz6n
iHp4f/pau0AW/Lb+GJSuvICewcf0f33uSyK9/cg1v7s8h6j1XBT8aKcWYNTKpmeysoJdi4OeVpJ1
AeoJ1vvarZuwEYhf7vvIPRxunBOzbTPpdoKthGh++2vfQpc+zn4TfFlgksekOVBPy0flPw2UcO01
u1Rwtimmid3R0AGI4BihmXp67n8ulQPGh1W/GXc8hg2TSB103if+pqRn9lkURmk4lIdjiwjomZ7u
3RTiUXmNoHo9+VV55IaezBBGlowIwx+bwlVFqK9rtixQ09o4DbszrlPicFIRHsMdH120juLComdv
jDbAgDmckFes9YpdEMElC/r89Q1FxoIqt16tF5ZbX+lvCtKjqQdoo0v/xFwWJR3e57QBgHeLdZC8
YpN4JQVKcafw8mQCjJMOQ0zd1Z0hmL1gFD7oLLwcx6aIjnRfOfzVETgajoAaAvlIgXZfJ6io8ZPY
D+zKokkzLhZn/fIlFyb1yBXmweKD1TVMdHITGv+R7+BCQOYaVk96T+xxiW8KbVSEKwkF0cSITFOB
Py62px7eiZtkL5hF0yqUTTvYtSgomu1W7SdzcsPGv9OXElLGPGDxgbktOYTCCTsFAUiSx1mVSdZF
S79RhAnJaC0gWtcfglYSMiXhXsx9AP2JaiylmUgmx7ajDLZREam8u96ArbZ985NC5Ntk5UAO38HI
VrXm1UTTf/VQ+CYu/iFYfnjISZb0LZ7xLZjhSBN+0sS6R4SRs1Db6YtHc4O2INHZ+EhneRpSvlIf
Ev7rF1usOJWvyWoQQcYhrCnuIyfv9HkeIzuBHzf2YeoFhhGf7OdCJ+xQEB0dMA5wx08iJqkXkZlM
fXd9K+9mWeSHux/LANu1xaDLjCsDO2SJFP4hHvDoS3nJ3e2fWg/dzcryCB+KiapLuqxsjBb4zRLF
QR4J1xnmChTvZ/554Gjxu5nijqZfDXk9QKRCwYulJ56Ae1iFbRqt1/tSuI5WX+xsz7wR9MWDQqUP
kTJC4BiRD+0pawBjUwuBmTsN8U8OzjurC3dh24ihmrquZTFNy9h7h7756zUVEa8Rqe0Dpo+uNSuy
NP2OO5nHym3Z0ZEVUwse8XfxbJuwarLXiRDBnUJhGjLZBf+CHgqB+56i+NWyzeLVaFHxdsH97grr
Rz2QyXYGsnE+QwilD+wXMSRxlAota85TDGqKA38nKa1z919xosln2YftPIbU+T+Gvn0thI+FkOaB
jXf8KpTEBzopBApEMh+sLg/GfpVZxZ+pYxWsxvnNwwpx1iOt0e104osW7MQviI/ANQZ8oxnwWeKQ
vKrxSvr5QK7V77tQ138tJCkC+5JC2yBIiXk6SjndK2VZiC1gUZ0an7ZBx5thY+iAtMERtWrGTijp
m0guZHTJVWtQZ3dxv+lqTzWsScdkn4KdeRKAokDhRGum6H+kYEcCpOcVeXA51p71K9gfIomVGtWz
4HJrH2z9cgMS6CBi/NqiuoGTlwC9HXSBkJHGWLukEM5YJd+PI65up2ZqW7uNGhVpJA/TeMQj7bA+
ySlIqb2wjFX5V8GnUFmsILqCqIwtCsx33GXPG8iQ10i/ICsNKyeWh7kYuCOhx9jHCIFtk0kMQUyd
F+agTdNwCOwh7yVI0OGPyCDHeP2lgItkn/gNSUeBocKsT3i67dSbfZgFeR94b9rsF6fxZ9C/+wOb
/jjsnQUQAVZfEQI/hUIeyUrFcfSIIpXop7R1KQhlU2uS67nXqbfYOPVqS/zF8wVk98tD09EZmSOa
ZGALAFvScdbKEQe/gKqhyqG8Pz4neE3Gf/0oAjAEocwPSeQ63Xr7L4rgHv6qUzkbxslS7VS3Pl0z
ePmolA9Vd7BoPwXEY2UrA/OIRxHRAa5gonvDHX6P0GR+3Wnh9YqNNf7B7lJ18YBBJR9hiZBh7BxD
MMTe4MYi325yU7928qgDBuxPVmNBORQmxTG9T4v8L5hvlbY1gRol+P1tcqZJnY/EdgQFuac4Llyt
lyHezzBF3n/5mHhOV7JVGJP8tV2dKOamE+m5so7IsmuNIbysR1tJLMXt+jBmJ4gS7ZBfTBNXUmig
kUG8mNd6SCYiBI1EpocRLLqiqn/mbyGcYNJk0NO2zJnFtXRrN8UqlS5epPimOY8bm/r8EhjSHaaC
3ZL2rByRTiZY5vMDxt6kbQuV4sEvcPE/6xzM+i/hprITjOHYrxm1QVVXzhMRmLsr7Qvz6SGqUCCj
xQRwy9A5lbs9FUuG7MioqCPTj/tOMxojZLC8/g51sNQ84YUh7Q7HPFQMk2lQSbF+4EyDNo3Plh6M
foBE9pLsqg6bZgSkTCqArSxpthGdHYGL6NmxGEkOxZi0jadfdIsQKvqExkSnWKVXBscNJ+QX2sPn
7OiGEmUgxs/OLq92m41RLUo6VX77+gPTvxjeIJ3by2jfBqFLgtchmij9pupV37ZSaaTGTTQPbki1
NM9dKaq9FC1+4EvqnrYSqcMfffJWXIRzZg/kDYc2QNCt5qvyUqSZCuPpbOMci2cjjACTZVa93eDs
NNliSFtESAW1VvJsjAXCAIo/2wJkq/ZI0P2sPgKbOnmESwxpPueGH4st3E5wkpKJPC3ItKYfpX9K
+Mta5a6rozXUDmJkAxgpGbBLeoQdgUCrVvG3+8ORaZ4de7L1Yf5hSXW9bQNKcfvbX5Gy85j/wGrx
0MIHCY7e1Q4+aSx0vfWnxS9yYyy4eWlAG+Hsv5kq8kXU7oJARZqCQUrtVsyR9p7+5O+J5NQf9XL1
1sftWg2cC75EkhQNHpiL0himbcU+tIkNrBYuj5KvK6jRc8homMfw5HqDEJkMOiUOBILT1/igcjKN
PYmUNprQFXb2VhBZntBOkokrig89gx461OB7J68HQc9peSIPgduySZmzJjutg11LHTD/1kv64RlT
1qx7OvgR0sB+qgU5m+m3GUKKnLj3a68fCesKN2o0TAliejj9dY8bvZDnk9Q1iTGseawOVboWOZOA
TbMydAKM9fS0J+tzUvnCLl8fTISYyUtdrNf/qXcK6Hp4KVEtR0UbUUPoUoZgEduy5EuXzseGp4Qz
VXsMclAuNlzjDqUVBQ5FjqqUs8JEVQb17mSnFke9P6Ep7Le/mVROWWQ4Iir4v3BZOCTSA2MIaN2E
2QgHbFEOubSMyhpUJouPG7yl09C5LHsBX+inxBf3ogQgzcD4iJjMemanaCM65Fvj4yS6zKfJZWs+
VxzY/MwlP4opuLDv81BgGmRhatQuQ+x84fiWyFJT1z32yUrFSEC7EM2zih0ao4ksVz6swNysZFhy
g4Ma6rUG/6GcykWow637oOpI9vzS4XUhms9h7UM/lLRSazEDcSU2dIU6BofxxlbOTcZEuSfXFnQH
jOqBpMoDnKm8gwDiAZwxKd6vnqsdC0ZP2efAq/lQjEe+wz2YUi5h2VM5YJDn1zu1+6szML0DWzfF
HRvpXzsKlg/sRrLuXDnSzkreBwc0mWzLeml5P9ZzdvaM4FIEtEqMfAXjNgDU/B+Ahih6FSEoc0qF
fjlfmMHE6YyEKZDQP7+CXag+/xcVug5aTcs5jj8/0ulwKphHGiy16LotNE/FP5KLzygqdCxx8vjg
lRUG2xUGEi3eg2+J90K2M99nUbYU+Lu44516JfQu89LXtDfKNs1/5Qf6hFjLx/VD+JIBm/x9A5S6
bU9wC1/0wdKmVucvinApVJeAPt8Lqqt+2IADMzI4IfYeneEr1eqQFddqQOahr0lgkKyaifOlAN+1
it/Yaf0vQMvmWZ5ctISxU2s71bR0zCVeUG/X95mMx+egJTZAWZl/fv7WKPKH+argMRg7hdLn88OD
0xiEpx1N5MGyby4Lu9UpDpk88utDFMziSA3q95oY3u16pR5cwGexKpQheDpMp2OXUR4V7X5WjcTz
ddokTLxnzFMVxu2Vur40GBTQH+XxCb/hicrxjxAPfEE645WqwRj2twCYLXvSvTNDkeEZy9Iu+m3i
ZTvVAt/6YHcrjx2D+r0qa3AIX9HPQ3gQGa8MASa0Ym7ti9BeZ0+Y9mWKh1Fw5i2yAqsws2e3rQPA
ZRM67KRdPM+gNx1Km+l9jDfNLxxm14whQeuqSCLtEURHhhnbx/FQJ76T/H5Ct5PWHMN5+L2wvCdd
oIwRUy/Ru0koCCqLXRU/L5TRD2fWhWPvkpslhTNrLgN3XOAnsXos1Sf6HJrpXFgETTZDuxIamhvn
fb2CaPjbALSXf/GiOgtAY1/gCcn50EbviXhcy6ZJ4MNH2JDB4uyRZhykXfHBJTE3XTgXkCbp+4tR
BvDpSsVuTcS/o3xtblZzQdEjSKJ5zTgN0wDJwGfF+7a5qNp++HbzZ5/04LFU5hIDSET2j+pPLG1C
MYCBbxBvm/ldJj8RXjOzfkVR7Jr+y9x0cBe93APd5P5QVV3lXwIRkCJm0PODQo23ejbiizdnamlO
GmeQlNQ0yWH/U5KcCEGUlPoPcmSLdT1SOTGAUMnBRZOXJOJLlmIwsEJLizLPR8gVZN+5E3TAFNlM
R+Tv2eJTXSd8oM1y62xk43P0+fs+wW9NWWHNW8aGSESpsM2FW5HNDJd3W9ruOgUuQQl2ReUCwhIg
SJJgjgPgcdI472PIwGSaSC6o/7yCsfwX2z1Ywm78sQU98MPJW/Ww5k16cL7/+y4pyOfJoHsyacQU
x+MmWd2c+PIm46G/6rj5XU6DGYn5iEGIrNGLSO9tKlNhqyLvyhHsoM5o/FXa3wfNzg9JG+0jo7Ix
rr96JSVOeLqNYklYNRsoOy+1pf41GjvaiZODRQpNiwuz7vVxflJ1eUCBQeHvyUohbUt4IzKA799Z
koXsslyvEqhhMRh6cM331xM0A6Ua/truz0eu43GexBK6nLs5Fu/6eD01TnjmKi1BXC5bl4OwJXdX
8n68khfkXtJNUKcmPnwNCXBXBj82rNmUYapZ+7kTaNFaB8SlugF0qxGXhR6U8376HHh13lTG0bvL
JbGvTF5Pt5BA47Uf4dHgXMHiamZnvBNetFbWcZbYm2+o9C0mdMA6lkVqZ6Ks3Og3Mn+IELuWjdOU
VBsSXN1yB1rVyBAxMjPVeEnV7L6G6/+MZKwIC+7MfHk+EIlCesnylfeEF2NIcVwsm6jH7UEJxtl0
Kxq6ZVzsvd4O/JfxsNWvpkfqetQoqcZH+dDHdvzqwzGWQdkJElNSKChd6nJv0D6yOvXHmyUPePlH
kY0Ew1fF0FMS8zfEU/t8A8scHdSeUQPgIkgte3R5Va4jkihiSIgxwkE3EIG/0PJBvbCuZH8EmEae
vORUhqPsI7j1U4BLTBG+e3M+qEfCSbXfD6RTbitkivDmzp6anaI37Tz+eUtVbPJYYmrelcaS/ZM1
DuZxcwI/W/K5OvnjRynfAuz7paD5d4IKE4NhFta2AP0XaBZaq3JOE3DbGu66Sae2PlThDIsTfdvb
aQiHplSkQcxd6ETGUbbVfw5CZuxLdWVwWNQQmVHcTMpdBN7+RPICF+yx89N8cSJ7KgmyiQTyAUJJ
rbkEA4XHPl0lJ5C3zyBsRku0TeULXcXX0knohPJ0TOJBibw5PO/rXhAHXiBnFSJnJXnJlzpccYjO
j4gkGxll1Cf1y6fK0ybm/Li467502MebUYYWxAFOSrjdEoLtjUSwedDXewh+OYpY+QukSQa7l5f9
R8H18f3RMsa+tAQvh8mx5atp/zgVXB5HgrIk0aQ0WEiwaZBXjVksX401+BryUC/jHB+cIC2cC33v
Wcj0C+aqR2NawsU8RWJO6DAj4ENydIgUKFfpgmeOElWzVwojPCH8Wb+yAgVl0N+Xcb8W5vFXf7hj
Xlu7wPzOuJcSJNHubcVJv/w3T02obFeEpYg6hqktj/rKamhO5MFFp3xuNwpFp8Do/OKpW18zIG+2
KeN5M6uZ7+I2L/SUpgDwmgEZ1WhmliYXSY6fW/m0q9uC30YbnOPUbwuuACZjhHrMH80LDqMgqW7i
cjiJkk2XZOTPVkHjryOTuTgTqrVStsnJXuTHENMp3jPSqF9S5i1L2TuG811+HUSVNmQ21NUvRH1Q
3yrX4sn8N7aj6nagDdseXIoMrDECr5M/7paYHB18FqXITBj4Hq+nrlzDb6eXDvGy+bs3P4p6sEDW
l8MJryCI9LjLHHzuPfM6Ef4vHQIM1pSR2MbqRBXSq2y8jdYTzW8JLSwyQdxJD+0hN30ue5bwu3fk
yMizz1AQSrdl+iNUqICxuKAousUBDVjQMpn/rilQFqhyfAuVTfR4VZEOVXnZ9iFbAPXLZBm4+LVL
2eFCdB3yKUEFgIOanQWxURxD44ZPaAHh16wPNOKwWO77x1VOndfnmtwh2kllgCWCrxtzI+1qvHXU
IFfvAtBeypCeruuOhdb+IQodMsq/dPBnAXiLcKz/rqoutv2QmudvQjGSHYxqZ9VYxeNFuqrDbWlo
xLzDZPKhKjBwMuMQrExIwvNh2j2/njH4luyeCyaAbqqTq1RZHLpoewoBBKQn/0qt8Xxnbdbbi6Rg
MDaHTvcSR3O10m0agUqgl0auV0gzfKnrsQx7MLjeXfLF1r+8bQ3Wi6IzrHzTUzLhPmVmMw/+VQkX
TXTWFza6/42iA0DPiV00r9HZa5UjW+U6MfXtOVBP2YOMvbf+0aT6DciXDiNPinbQWUAJV78GTTqh
xLlmTrKKoXZ5GKZc3N4HpOlOpR8neZow8v+2/p33J/o23v4m/8x8+VkcSlEW+zNHHLHyscwBz+x6
RR4M9dXtCOckehqSHUlWGH5UsFkTaW8AfDZVAu3ADYPqBXR9EvlkNz6un9O+wFbyf6IEbhR1m3Sr
3YtoBELOqU61cYfUAb8lN+4x0sJiVx7IeA1+FLm5g7O4zv2NChycx7v9Bj3Jn1Y7BaHMRxxcjyxr
LDeIQpbH0A2eIgMGsxRZfPgzrBcuO9nW1J64o2USyHnxp7wZMDNm0Kpp+CwazrFrbV2elyF9+UyG
tt5kJokDebPhAvmEQt9jX4+Gh8QIv4UriOvDliqQ3YRw2rSRpfG02Vn164drExge6kvh9aZTRqQz
n/Z0brvEkQf0qkJDqkxtNvKOwdw3Z9gMM97x3Kakdm0fKCvIbwmUQMRy3juCEYrKEkltUL9FUThI
9LKfp7/VpdtGvgWU9gPbSKxgBNw/gtpw5ec+NB1ynYyRuQvZp+J9y+uUlRlO9Xzd2HlU0JmUccnx
PFlG5Q1/tkU7tvRIX+E/fxEbaTNtUkNvgmEshKruwpDN3sosv1TAOn7XdBBc9uqvj5E+YxLnNpi2
XUlnSJzPpqu27cEi2grVhNhmfuNIDKjQYtqi7XEUk+O6XEucnHnLQ2nYB/3VkS+DjO8bk9vTsgTL
fVrzGMs5dpNPO2/5VVPfdlG3fEIhc4G37VMSfhsZVUCfAJnXmQTmOUXm9AE4ZgH46U8bEZynQKKQ
psEZonOKze17EzUHAq6tC39lbyTx9c56Cpe87VmKocKN2ufdapyUKvekq1GiWq2U+JFWOOpvHnb4
UqsAr8xvrutrAd3+/rtwWI/tR9KuqgCAoFq0f9Uu1ZGIryFiz/66Kl+7ukFV8ujzU8I00PWgRzmH
WBJxEF3dT9mzyDANQ6mdWIqDWd3/BrFh4X8M+UJxFYLV7Ax2ZLzvIGKEc17kGtdTxmib6cxCcarP
mAygRwyy/TNrcSW9xeXW3QD7eexF0EyuERw0vub5JKfoiWLRWKAByef/RmB4fqJQMnCit4OwoKsl
IwQr3qlKLBPLLkmZvBkFdZGD98PgfjuRnF3hw+0rHItX60pefpNIGdht0t/2ClB05vuMKcRXZD7d
VuFwKM+3JvvCL4o12oLbJmcWA9JfDCiZm6k7JzZeetYC9LPY6PuoFvNzxDQtCgHNL0mcdEgQiep/
H7oGOBFpsaxwFoWxua++uNYdtCIZ3wrpfWYlBUgaUpvRhV3pZlzLgorgx4oOvSDTEmlJtYPcfWUo
Q2ZCQzV2xpRciph8yWmXKRB8N78N+dtOuyAcHWOUnn88+g+H6S8DCf070WmV0s72N+cAoAYUv0og
bUvLAkqhdeIFBlclv3NIlXv52aL3hnLI7EDwFc6teHka+NTNFx++Ng9xs2qncyYeikQAfJrak4u0
W95gz3jn79wPQYFD41rJFDzbCgPBPIZphSM32QpLoJgCRT0FWVlyzefNKXv1o0lEiMeAqb+0Lzzg
OUi4dwiiJBxo6M4AOrPLE2FM6GRoLRRWAUA95EiV6y94O3DJhlpzMWNP/xF18cyKzYn+Srk+hYHK
EAX02OfJo/PNzfIzPIm2yqTL1t8nQxWF0oDetGNpoKHnJv2Jl3h69DznnW5euyyqDIjtcVS4WT+b
nIGS7XdONlXdpexll6RvTDG6QX0TDhnCmGyBgRIK26GHw3j/HYd61L90940yOQLwqqdIwHfxvk8L
pvxt1bkSQSSFrasuWeA/rJ74e3l/s9GUMQ0ssOa1fye1Es44QLJqCzLTP14q9ISOrQJaNCD116+/
ytW747iXkHYEfLHUohut4S8IahqGRwrU3mRfbh7YaqmZjOJuZxmzWUngZjW3iwdWlLwQ+1aiDmcP
ehyccKhSPKfkp6xwLp0MMz/1Ur/RDC9qcibERpkOBZfVZn2cvH07BWlcVMz70fWWylqvBSib2MTl
vF8RHdwEeF+qhgPIlo6Bi3/0YDF5zhUxrj/2sg6xj30uGqfLXI45e+3Lksw5TMrWKh/A6dw3coiZ
7rOtEqK45GKWrEc4OJPpTRbq72EVlZs8SR/kZ6hKiB0ziSpDIzOLyuyQ7ahH4P2hbUTur+D4jO0G
dzGEknE3GFgvus+snnhtHUatbxMbzI4x/CZh4hPjdm1Z5/NLvVt2BfHDvO4jliV4UlXMBlnakMg0
chs+ftOVaCJ04K4cWkqpOTZeOaoEVOKRaSCtNAJ8NHGoQOQrJZoBDERB3CkVxLprpjiI/JYvVPdS
oVn3Vw2oLS0rY0Q9wnyihZ6f9Z1Ic1eLuZO9b+jh/iofuK1mxsRZea1YrggroN2grwKHwMvXCIXk
HSxHL/i1lx925RNLxvGfHOBzbKebLS7LVIXPO15dbZKE+2clinkgzNsGLjTjuirQZNrYSttij8XR
bNxidSIObydC9lAACuvo53CCFk2xgHgvvtxr5El/7G0bvFh1ojtLT28Ujg9HDMMh/cJU824FPAM4
G+Y3VbkVjBUi4Nw3UFNY2B6mXNl/tOKxWAPYDnpx7Ic3K2TjqtxGwivUQvxeCvwtiw3m47ZR2NsS
mfU2BPjE7iirQXjn855MQHYTHPmOidHC0ZQxeTKw2ttZlcOnhN25+LQDppRhXt63a+B7TPQxikr3
bh1R02DX8/RKS0j4RJ9JixeTGAMobbcxgI31SIJKLQSd/cSsR6KohXemyjIHdxAZRZKEoOMUwYpw
zkI52YM54si31ElosVJ8UTz56twc9eLTku+MIE5vw3jl2VSDlVRsbtL1iRfWLU5oF2N5nUhspl8k
fLrVzvX5BUlHoz3XRjnts+xcD0OXtlm+9w/KV41tPVhIUDsbv37ujdceAmRNAD3cthRm8gy3mBEJ
URlFqHyu/FL/FURN/2I7EVMR+2jyUsiojj8EHNqCM7wtO4ZS5OTwNY59f9xTZIY3a33IAefDYqqC
o6p+Xa7q8ddFaNnzRrq9tDqU3Oy3tRNJAoEv1VXXyVv9cGjajf7sLuBL3Bpsn3MCOEP4gZaeHyIh
/WQRab1d7K1/PznlHY2029bAOxpppwjGfBLkE8Mv+tP/r0k5Ns7/aZ8cVpLCNj1jSCKomW3UseTo
ySPJJsymsanalRdEejWucOc6Mz5d6zLDVnhsTdD5A8Egx6JJjz1hc6lSlUgRS7wrROFAczs+j5GI
VAm2vhb8FOLFZeBH4hpu3OAJrHidooot6WQIEhgN0cXpv+Re16pedp4/yPzpsgnca58nlVVmH+Fd
8W9s2NAK8mdvLhvewMLKAzH9qzQXfQX7Ps2I6cvnYmhQlGmUXGRSf/uz8voFhED69A9sZNb0/Rg/
gP4mpc8fI0VsLX6rLXncI8HAL9amLFWpYNngzkcgPIWGqjEBL4SzgKjR8fma4Au79pZpDHDYlldb
RE33Bd7EFS+sQzLmxA6lHOyrO7Bd1QCZdQ+UBmy5D6weh7JbJv+fiXEs0YIfbx4ShEScEKaVtD/V
6OoZc19k5I4nAODY96otYrwDNmqDknXlxtHe2DhxfvU92uffelIDqtLYCv45UJnoda6Pfm1B+qzH
UOdedSvuoy3YxOoL+J6XB9hZzSedb5SfweODVrnqlyc2M2LnzLSPTuiOypmveFjri2rzirZAdHDW
UQPWvng9immKN31bK/cD5ASqSMya94mPxbMWK6sEL42el0r86BWV1r2+xuXSp0jus/ben1FTJXxg
F7Nv0aqmSj7ELzTZscOgILqEewUbQ+SdZLUnXiamTpx3ryuvfC6omNec4I6Xcnr3HtHjDdd08c+8
5swvxi4TXI9b1vSdXib+owTg0ZUt+Cw0XD8rtPAk6Q17qsFRZO7/erINzPH87FpeVDBsfXjG4x/E
wEBO/5Ju2cceTR1h8LRG2tZq5+nVlS+HoApZx0z3GS6ICiGqSJNjnASpQSF4QHW6PptHI9pZKvLt
2x+AO97ML13MgmSv/EnTvafz8Nqkimhr6JauD8Xw3D1587C9kRy2hNDD7MXLKI8a8QsBdl9RyyTS
L+6nW2lOjRKbz64j99ygZmncOd48c3Q+ofnI6CrwyBkP4mfpcsL2S+LDeZgjDNT+vEUOdQ8uisK0
15WKqW/sku9UbBc0SFgXzL3Z2xFzCMzCOyb/Bz8lMSfcwKQSMGt8571BuSPvz7S6W5YPyuZaheiw
Ofyvq9hjFdTy9+guWpVM1o0Vi28gf3jyejZVMnoMSKkKyN6sri7A4YSUFjiJL+mmWXMmcuw1sSlW
TLai4bUhkQXrrVfEMjQpwtJd0fWXl0IgBldPsTQeWdVeVHu18PshWA0tHccmYfB/3m8J4iead+Vl
AhSzFe27OzVPT6EByssnMksuDDzR3Ar3uTfpMKbt8+6hL7o9hXOnSUrbTSEBMSWHPr2BTP+WKe1q
exzLYHjcE6Pr1+1Er1sKbSD2ref8Mdsw7XokuKHOi76WZzuOMpZPx0WsfE9aHPpOOXpspzwzGHTW
rhQKHbWhY/RNv0QEP5XXI1s+WQI7QxVaYYu3OmjQRwnSa5RjMtsbmZsEnHmmoTjtrwW0efxElvC2
CH5ppzTLG1hM4wLdlQZNyv+jJzi1+gxSpGQVzHcOxFzKETYkQmg6ak2ZQIrUf5XBBUOsKXp1zVuK
Y9ndbCE7KN2x7POP4R2qhP1IP9V2y/COnYfuPZn5mEnQLWqWY6bI+ag5ceRvYR6wYlOMLDXaPPPN
K2zEhPDT8GeDu9MDYnQap6giTXPEbkMdfgJGSAVFNlEiCMuk56qZXbc/WhuOuOpx9zRkcDkxdWuJ
UznVstUj0epDNYe+M1Dr1Gy+WCPcepefmwoEJQnbw8oR69YArvu+lalKSbzQJspNXKdhX9jFRtGS
lfQ4a5rsTB/Y+ZRGNT0VeMHcKITtD5sR2VSDeDY4jHyWiVhrUlBmqbCDLKJpMpLs7MDMfnJ4T0U/
S8rwLNGB/v7r+3vMVEA8b7RH93tfwfh4CSnWMLJBc+OG0lbuquRLsZjcH7mFhofyK8z7vc5CTKL2
Eot90gjX2Ee2V8+3d/FRx11lyq7Z8gdy1jxU4A7mZl6BwKsiWhMW1ev4C7DDN+K6OcK4rviWAMqJ
zbemLT4tOOjctc5QPcXXZ4OlWQtu0IudUeTq83vHzeHG2ASHd9i5RPQvjpgbrJj8BfOtc/KWPELw
9O/0lolcjTSarcbebvynBlf5D8YFZRtiKNIwpcbkrkzR8dyRozjMSME/soqlDZrOI3BACc+/6AMt
reNkOoTUqoLjPxwi8Q3OOyltebIoScx/nk0OOjjkAkuXylbGgWn4KdUEkPzYyv3Q4YB/KlYouMCm
Hz6pJlU8w4c34R5Apt5Zcal69ssykQ39qUSCi3B+jkDAeyAiJ/ZEEpHCfx6uf3dUxIE27eZ9fhEZ
m0QLFYXfti52ZncNiFWwpdqjh8dhKMc/9aSyHmoD0hC9u1ulIAT+bkzXJdbRVetbfp6CRmuOdaU6
jwMtpJ5xC8TanAtwTcS2RMAMlyJexpfGQM+1y6sxci+L4hNNmgrYSfvM0qSTkv3nIzwiBXKuIgdr
r4CCsIyAdYmnALsjvMDwHdV10uOdIix72Brb/2tzSPtThIa4qDQWP+bqcj51+/8BBMrYspt8Xz6n
1TF72TWss0pI7GVHUQs9cTq/F8EEh6errQh8DBFXIcKssLiTYZTGj/HutA/3f09/w9QLBSvpXKn4
atGuV6ak89S0WR7Zj8wnwgaflKwUSN2NW0tLLWMtsoIDcKkmwOBxzgjzPpCFa/vyHhAn+CWbMJPk
NRMxJqpSovsaYJnm4qZFljn9HMXxz8GPFCulWNYqq51bIjaRgg7WVma016CMvHN2RDvFPgvPIotq
YwYVxawnHl1TdMH7e4rqcgo2H9oFRN0KNCrCQPhWWpqHI1IrkS32WkaWEFMa5ueuc9adnAkEeFh8
DomCN3bAC1K38MV99DtZs5AWXN7ths6nG5tF52+Aj1h5n4aYErMvWtbehhl6RChqlpsnJ2IpgSo3
dXAXEseN2dRgibHhZPIFb/c8EnF2fbtng6KDhDoHy/NOGjBDSV3poKktd7enlyYT/qpcnA/8vcui
x/Op7s6F/GbViVWdXfkXt6apckjTb2cRl321y1ESXscxGAgEBakPQmaG0H1qrgqQY18cREUXPNPH
5/rRHqXoA1qooOrZpw6YnEfOFb8c1aywzsIBBa6RSQS4+b3vvmZd0mIKjc56dDQW9xciPI7AE5WQ
I0iaj93fx+9xuIjc8kNhIFzULUPr0O+WqIENLgm1gKQ2aAaRNpIKJVEMMG9DfjDvdGHt5tSXkSz1
TjQzTZVy5imrbE3dm5JIyeAitFEERM4Me5lJukRpuGcN2j+ft7WQt5Jfi6FXVF9k/DigyUcDnfbM
NS2yeBQMUhMFY4Liie1wwTQJ2vP3slzqQv8EGB+EPodgE9LipdzLXNuSQlWD4AB4SAAkZ5kT4uGe
Q1pVWvMeemCTEZ0iNu7i86tPwwUBmKhoUCPkVL7FhIBA1VmiD8jIc5lJ5BGik+PB8FdBvWhwVzp0
4ZpNxyH0mOJT/y66PdkHgcabxXwIFI/5Qr0e6V1kg+78jjn+gkPqBG5OcJKvwV5vdCHTD9k/qr+P
yAUtlt8/aWoQGd6vIpFsmcU9bROIpWVzkRc+fJuGYARW1rTZSQTdrLi82ehmC/CvCxRxNBpVJvyJ
k9l6uBjAwaX7+d3amJFaijx1Ob/SUs6Rv3pDh+roK1m/zc8RsLjBvswAzK7I4S4/4GePqC+7/w6p
+3uAczS1RsCA14KmfM5HNER/6hi+AsExAeDLn4+Foq1SMiX/hsWKRJzlsvZpxxEshHjgfa3COLuL
Di6yGm8Vdrx2CS992M6K3OFKkapZwUy+jLCQBeevR1LcLowyhkYU9uqASFi9lXYL/RLbrsRPloyq
/wulabls3D6bGQG/nnA1wU/5R2Hj5nUZk9a6o6UH4lKf+Nuxuw3qr7/pdWmYEL6cfXh03SOzckQw
BjVnK1O8ZGGUKamt/bP/wn2gWbqiVs6sRhhNq7QnE38SuUyv2fL21/eGFhFtKTb5uiJBejiOeg4H
MgHj4iJBeChZAYljDEbZ/dH1PZP8/cRvb0EQ0UbJOjwBIZCJgNt76xh6sPeNPo27Wo2QQgkyrjQY
ljRVeCOJKXx1I9jQniLeU8UTPxjjLvvuA2eNUjmWH+nfvpmgmEk1vFtnoQ7qnmFmeSr9IZRqT6+0
Q4S7viBO2h0aybJ02TjlfwuQf/hzGi/Qg+nGaedHF3DLTi9fcApdQRhIcMvrBVqGblSugINp/IbU
SYlMYazlhG2A5Pf7LDCoyM02s9rjUYteyKgE6o+kEyTAyCAYF8fWF3f07Ky21NdZE3V0/dBUdnDJ
Sh8s2A81N8/Awi76YPDn0POsRBv6tVQhyPawdE+H5MAk001FfFgfnGwuHagnPwpxNtjOYJr/DXpF
7HZiEoEUmEOhA+Ba7g7E+sxYL+SQlNr+GAG3pmeWtqxlsoZX2yiIk+V9DCMVvZsDuzIyn3V8RSIw
lX4hUhIKN9CGwAU1vVDLSXWgVliRTXLM+1CSi/xUvcHFyBIuiVN4m9dFhDs8HS6WBrDBHQ89JYDR
1ltujP6bp2ggaO/++gPWWZXZY6qyRYFmREwCefOLBNKYx7pFy5zA0+knpllN6Qe2PS9zM8q5Re+b
VEjhrAV6lnl20IPd5admSggA6ixn6S/ZSb0wv+i6GZx/0SnSgc9QyikM81AaCJB6sO9GNRzMmhfv
h7hWZ4j2AqTi3IvLuolcINOBuy3tHK71GJM6FXk9LV5fq+lpQx/H84RswRWhQv8SADjjMq/ZESnu
UqeA2SSFEsl9DPiJCjI+eWbqjDkwfdY0N+Na73nWIw68cS3m3H7AKAMtUfSulLSgHz9Zl/HUMp05
/KbgOKqfmto4LLioaNwbig7uHD64ApHlwxQ0eV//vCO/4j48i3rSbTbT6KhVSsLELfGLYpr5wlU7
RO9K3MMeOY86z82JRcOGQ8fGnQEDD6MtEvPMftRy/M58DYSG/XHSk5ah7xFxrtdHcPjB68x8XriR
4KLgeIsTK2H+vVK3eXZ63rqN6/R0CvszfLu6551d1+CKdtwkBCAGsRNiwVzDdweJBGwpCmgCjL2E
OlJQGYhiFa48oIdRtd+TrkIFJCoPsF0xDBnaTd4PHyHzxib5G55QKu3upahn0Xv0hQWdeXoS/WGH
L9vtBvRglGCZz5ggMeBWhG62cDg4ud5D0QQ1JuQOZbxnZ9u0gyK4oQCVz6g8RcARcwtkAmW8Jrug
iul4pFm7Ocw1a+kdLMaLpGWu7EKyQplT52+aHMICxG08hio2LIYyx5aHlC26s3Pr29quRh+qBwT8
lVGwiauZJ+Xll0eatOSTjFsDTPo6wf0BYC9M8vZ5RXzkbVlu05TOC/e8lMHp00h3IRiSakJjhWbT
tYCTwUBZ5VgdmXdzcNQeOIyMD/WYPWEKMTfz44flayNnxP35+jOFBm0frMdlxxMqU8483Vt9PO9l
56riISfGtOL/0d0GRIebfkiFxxEVOGH7L4TH2jN8UsqwOxNUx7TE4OQMlfP/7IAKgP4zy7AdsBil
FgPYNwAiIRqAE+Mq3YrTLCrs9gXxNb35nN+Lnzppx3ON6QAZMNSnYcAQl0pQMJ87llJTAHTd5SoQ
IWRvQh0teTz7UoKiRno2sgLLDBuC989ynQCuq18l9QrViexvSGL6nhD+HAOf/0O+OTTFK/Cqb8eG
ZWDH3axT2/XQ20kYJDgD8Vi+VhJ67n5Y1z6Gwk+jo4uuN1qnEaUEa7bgzt6NPs4GgF+Z2yHHZLPH
RJ4bXa96td53unwSLtBFVh2pewJqiXOVkZHPlFKwZKU/CyUx7QTy8wYHOxWnFbg4BsETYxwy/8+v
p0X/0vtkwLJX/ZVf4gS+R7QRM/byXKwmJswDI6MnTlg4hj2Xd/JfsFBJfQZUSqOM9aCAiz3NO//e
WPJ56gmTdaU5EWdX4pX8anoGeexJPNH7bFu0xsVUhl5HN/M6iK618TvklYh632BF6jtvkgFFer3g
mjj2rzpej/SFsOVAFkVPQzxkbonf4/PWUiSrcAwRIC4ifwFyKH+MvVTZN+cQ3TdLiVnRjDwxEL0h
90f0JiRmFDNhV6nuZ0JxBeiPG8wHMbGd9s1NMwtSTkOqGNK04wHvpbfqyJoXpofdktLn0U3Tax+N
KBniTwA7CTGOw8NEvmtftZl8HVRh0nnY3jB/kk1Q+pcQn6C22UstErOcT0lsXvgRXTbP6O8WKR2e
eZWU5/+JuORDSk0vkDAHUWfTQamRAJvD24U64BQyOISxYsl/gDv13fZvBHU/rjTyQdRtjcWbfFms
5qURyiJx9SKasHEFoilWDPefciB0WvstutacbT7zwSYhMB9lhdKYyApDF4qroCI/CMbB2PXQZvIg
qkLkPr4/4NWsSSTvCRsM63ROrYzsaAA3Ah6Fg7sbmBKasvQKOOz7IWk7rRaJtjl/aBvGoQBeadsx
wNc6ZYLqJVg8AlTeFMouui5F6qh0CFmLt+icWB9TlUC593x0ywjdNHkOYcEJsCH5CqOqCHfwxDus
XX6Z40GLSC38qdi86TApxYpCpOBkPS2BTL+DDy+7iIkaGM8a2huXz4l99wsAsdF8hsle/ie6ixPf
B7xk1kNs/hF6qdi1k7Lk03ZzeJKaYracJ9840qAgac1AQwzYMlYKmYy6s+PIG4WxXQ/OpsW9Koup
OLbHIJ4erOeM3ECWRV4FpVPQLO5vsA9zJwH6KCghVMeq4mtGbMspegHNYWtcr+gTW5nrQlSv29wg
tHb2213+r+nyRILmpSA1aFjyeK9a6lSTpaUps1Of9eSQ60ETfMSqTqqIQKbsM71PGA2e25xHn0gb
KeGHnPlCTyCG8GfGTUciDYP/Mgm0nTPCIZaO+ciKEHHs3/VQC84BanK0PJyfmStFU5uL/VFeG/ko
r1qK1htrb5xewV7/RLGUaFcym9B3Xa4j1waYPjDDn3jMn0xYot7mWhDQC6thJxno7tNAzWqXpqQB
azibz+JT/9MpP5urZAxqByW70Apk6iVZffgO5g0Os1baI7ipQs9yxyWcw4NawvNiKmBhyFUGpVP1
hrpCUnWnJ5fEjPCWaLRYAT8SI1JBDyx9NQhzX6SFA9rCVi3FEVtjQOuLwXoqHYw0ADzu6d5arY/O
ZAWwdqM0dzVNrpBNAbyYRLehgcftfYXVUR1HlPeDKqdt2Uo4q9OX76MLxiOU1HmTE6tOC+PzFQw1
tNKfGorHROl1NXBjQlb0QpVIFGy0XiC08ai3MC5tqYZJAaWS7Fzm8KThljm0UeGLPk3QYAAm6kFP
KJ5Eb1RFNIZHTCXTqP8d2kjt3y5PcAiKcLZgVvpfsi2WVrZ7X7j0KyQBPNQi+rbR+qokcKBUeME4
gg37dl2gknfpKnfIIB96G147B+YbmttXAPckio2l08K64PDXZ5HvN9888XNv5QCvP3YZinQKdScv
MZIkclsQC8qc7VPpNAQEiUtlapzI20njwcZYarGURNnNviDl6Or6yoOfqDFjSStysi9yMu0I06ss
LXpKyeXqxL423jVZNVwc14IwY2Y5EF7u/pbXBLir4dNg4DXnfFAlt0P2/8Dop+wlita6eIUZI6cX
ay1KGkVVK2d+Yo3EOGSpTiAP8g9cdm+riJhG7NtzOb5z+IqbWhvZ/kORnII1fwBGlqNZqFiEwRga
UEuBRZUbI1rL/67OSJ3Fb0FGRbT1nvP385S2TaGp2sMoDezLJc7WwyneAOWXpQ42EyJt+NSUbqOK
e2upiKke6qEhQZzvuhSZDF0RI64Yo90aqUs2NdnMokKkzhXDprg8QkTbjWOLORT9zEyREouSWkBB
VtWC9KktNaTwHPkbTGTzdY3UphdsJDbtRLRaVvqc5SYMZv7vzz6uuprwP1i9B2PFtib9CCedDGz2
lFAEc0J+sgkQqCVSG4ndT8gc/t9grEz/7blVxjmCZPlAiJ8iQLkfADZ7tXe1k5zhOxFFb3MkBiKl
+UzPkniFQCk4T7J981qkZCZb1LxxVLbdwG7kbIduE/2WoKRi72XTgG/tO67/W/LDei7tuqdW47xq
rpTgPyKevlESKlEd4EzFILLmdBF2uDST01Lph5Qmg5eP6pzWHt1V6MQF4flUasDE36i98eg6ljuj
xjaFtoh7nP9usNDCKGtiJjNoekkAD13lUrcf5je4cSrqPJDw1Ji6Rmh2fel7zFZPWv1J0BQ5OAAV
+TTekp5Su9+NzgP0bety7Azxiv+wNa+pY2ZFsLUrQM+6Vtt4ThZRinmAP8Pywk6Gmbz1yNZDgjrV
EM2c5BDtd5xknMqhjTWU4ARyRgyxHt/kckzwiyzZUhQ3iXxoRZ0dbzPaa9TwhQF9r7sE5A4UhNz4
DRy+qOfk7FKBEnyu8d+VVJHu5fFxlXUIspCT8wa2XMRtP3wvU9rGy9x+mPiVXup6Kf5PDfuZX+Wc
Wvc/BfyZOLoiTSw7W/Jti+VFHs4ZURpHa3sEV0z57Rz3kVfpVtPEtxJm5uT+zwMw9UVR4q2Uf1rR
H13bv9dgb2ZbVNXgmWVt5eBnCrFnn4UUfkK+EbfuIjfqJfTxAUUyz5qT8y7iLMjmT6Q9Z5TU8UKw
ODyPrz4wDc47oEa3MsDiklkD9GoSV7/bwYbrMhvGZNEb5Q/GhGaJ6gT9/njjntqbqPlbjGconZN3
GBwpPScEBJPBIVsMSf2t4GQ8n2AQGjXNdX+HcFHwg3R6qQVK72CX4b5s8pz12wyxweIQtWt8yA1q
4cRehMUdSQxuekqXXcyUIai2bd9PpGq9VIVkKn9+JRuZkX9KVxcfJk59kG3Tjo6SC3ExYE5+ChCG
2s+F71+fBhExl+h5786L6yiGYMXO0I3TdTAmQFNVg9y+Egdm/Cs46aU26KUmex5MWzwWT+lhC9UQ
JSoCrbfXXBNGMKozoGVu1YbKCihR+/emYrjK1Jw/pLskZEAolKsZ02tl4qCJbcnKlNFvR610MwlF
6PgZML4lv7hEK6Z0LMloz3usjBP83nJyMsFkZd6c4+3eSyWeBs5J5/R4mMfnSsEUClyy9psLAa89
XaptpMLuRlEX7ne4wS55cCNBbzLmsPUCSGDOt6AlO7g99iXH38AGPDcdnDidBEJoIWOC4/eznTpO
3/rrfCoyeOniRePuIDeDCIMQBg9CfhTNK9VknV8hebMtUJzPEfBNRKfZThBPFbrbE5wXYEP0EJxC
5lx/9zVp5BoSzpxiCxAsUwjpWxUfCf6qBeZJsDRq23+4wErob549E/Vp3zBtsYotXkzcU0A3ev80
a3Pi1mxIGcrgLcPpMRJQmJOx4ydNlNSDOk/7vtYJ0F/4uMqbrcyarh7+2VQD4ihNX+rgTqLLRHlg
Gdlv1tsFyrEoe+Ui6QfcTyavZmvzQYss3UxFBaaGeQ12mrR/0ew6PoxBJRNztSFcdhMhadCmpH/n
XiPlKNX8hgQsRvId55dPZMxk5xmCs9JZcMY/gDr4ZUGBeGCyjb02HaagvU9TuKtWX5uh0CXtxoi4
cgAcXqdyzjKTS9EEjs4HPPm8IKSQPr1AUTRjePGsGTW+I6AIZCfHg7RxChVQgEZIox9TOlJhhglG
HoyRBBIvTcIqD2z+mqxdAOS9i6kwXPnVNeh5ZjxjVmtGb6RRMDlNn6sn3/Mf79yiPX7kqMNap2oy
5Bm7sdd+1ihAauOnsZmSuO4yOdAd4xIZSBw7sPkfCbEuA823nYWPH6u1eDosU5uLNt+Aawkxf1wh
UzeIxIz8KnoQ36JzOmxuoQfrxDh/j5wiJVltPeHj6uFRBRRU6D9tnPjyTC/oT48iL3ucxRz4xX8q
cMIo9fqg2uD6n1LPg3z6Pm6iSxP1yk6kGGY3Yj/8kkr7Ka+VBA3NxbaJFbPcVh2tfqSxA/cLLWfg
BuliabRFEFbb0UECdnkV3fvw0CAmxEoilSXUb9KIHkQG2XrKN3dspIA5e9Uh1HUbNRqcLTti/NNF
QnDvZCXaWvWdtTnP6sXiFKYN+HnmmP4aKIfaUturm6sjffxIrpC9vl7oZvCsp87+LeKIJYvESNeu
UVI9+3MnWGrOokyB0bAKNAxh/C7SXVrkScFqHU5v3zmrEMHcuwE+P1WmzUZHlsE0xQJrkx5fbPuw
b7ujpaEQfc9UHOijAt5xYmyhQ/1dr78+2MjhxK7+jfeK1lIlMYVqpzFkClZTVo8FrgnzfRomN17C
ZpSG3M/aAnRRI96n5tguP7/MwadfyfxNp5rFxmZaCk5HrU1D2QAosynhlutFwo4WKyiSS/fy19/D
/U6SZyiZ7BRDxGuvQ+gEqZNgrJAY6QPru9S/uryv8WURs9tPjbm/AQFUuR9KBWOtsRKN9CteyyuL
P1tH70hphtb9C/1IfR0llUcBjQo9oVPd4yQD3Jq5Pp8+gBJM8t13Qxfxfjqcz5AZ8GlhsSRW7Nuo
j5v8fxrpmJKna+wWumm7NPpnS+1w2X2AXqoxQlLtPZni+A1LMdOr/o8CLsFv0SC+AAzqz2CNm0cd
idh/jaNMglrEMxnEZI2sK/MJYA3cqtVvaR4o2moIWWqClSSzGSwwVbE2ZjuGWCCwW+vvxPiEz2u3
CNXKBcfwkww07tYkEcHxKg49KjZUj4nTZ4DKO56zhmNLQHxHZ5lPbBiYxdJJN//uFX2HLEJrsfFW
GpNPj++hA3PV8pSxFxqW+pQuINDdKac2VGDclPlydnwxdggHAScVRH5cb11SZfTHvtRfB10YAABi
k61fCyGO2iI0805Tj3qtp/9dqJuGz/E2kKTmL4/J/rcV85Ds+ejSMylKv1/SHL2idGnEZhPsKf9V
yQSl1Cu0jntgdsG3kMU7YA+ehnQJTSDiHqjwg6mPwxH4plu3+KvalN0Ofp2qFxFjbfvRCoiwwYRo
xsEsOSKKXbRXdaY0QASGoSVAIsFFXu/G2F0fQl383DZezUaKCgyuuTShGGZ3LP53pdM7C4T2UltI
V68d9VbXo1tdBosHA+3NwsP2JurcQlk1XUVaqKG82xIfV2RORKtnna1VPQhYAbfLUm8zyjHXGOu1
HusiFHM9+CT1NkrvJLNziIqjoTcLEEqK5WMJ3yMBeIe8cDjavElROTRcD6JGoQPfDFPpQivNpG5x
FWEBdyauwt6dgM/1in/wRb4iO8n/9SVrZdNBN6CTlNdvekVX9GqwuTi1Xff1JmNjs1UY+/MKs7wT
DUPEEMkouuzwd7NGGll+rsvdQLk+sshDewCXgrZKLf00uNzaBqhkU9odpQ/Gy7eX4wK7cxvK3nPL
MKH2EnP4OsN5AsC9Wv1OoeNuni2yoAsKl8GgTxrRX7/Rkoi6tqlcXD36XWIF3biC4YtbmXymq4Ui
ogRRdfEpSeQtf58r0cp31cgw+8Nxklrlp4V+epV0XMMrvGu9slYkx94PXSHHo8r3kxSwJnssEht9
4mF7RH7ZFEUa1IrqFhhj4qhtdj1JP3A96Bj1B/vjMUX+SG7P695ajIRT9KWTlHVUckceobW6Pmvd
gTj1PUnEzYNGNVwPYi17qS9eIkVe+ib/V/wJpsqcr3UKD5gl4p0Gxid9DfcT98jT2ti1M3+oITmI
kky/63NbUqc8xDfMnQjZREjfu4tIvZzzFPe+ZVjP7fVRY3UGPiCd7+t+YPjbNuZdCbQkdLq4IUwc
efYMXfPAyd7KzLzaKqgpdYStFOwHOokXgkcnkZ15DM+mIAatAhzv13HBW35NNSQB3lx/2YrWmdzf
aS+hHGLZuw+5rS0CyN4Fx6jG/auKni4cqpMxhTrm3uY69RuRYtUZssfKv/eQhYnX4xG1tVIqVRhv
1PfZaOG0my4S/ziJi+UweXEcmipXltZNgTA2wUoygw6o6ZoGrxDeCbRpHL5nYatxGc8aIAMRi+BY
CHyZWQo8nnT9V+8lIi4ubSQSlBgyV8uAQ8avtV80Q/VbjLxSJPzHlrzV2jrUBczf0x42IqCCSfIj
63AHP30qCxsX8KISwKqnVy69WmBMPYT6xVq5DuqCj1YNYvZrtZxUCjSC5eW9+jp2UcF7s2OxCaf2
9uzv/LSaqFnsRKQ503vuCXfzh4dEBd1+tCGiBG9TfPlAkYHkFH7XAn91vmesHGLohWevu0lBxiie
gY72zCE32RQ9I4qmnMHyXH+gN1nuRx7QXyu2ZvNw7c8eOfEjJzCArUm/nR6XxIvXP/zknnzxPxyo
4/AyZZnao59v8y9st42seCEoEDpX5tj8Aic+tUxlI74Lpk9famyu6dM0XNXMtFWH6KL05W1JICN/
HilDt2g9ZGZenngp3mg9esPFCGFnFx9E2vxVQAO+RK1vmLHOikZHS5dNqGY8F7xjnFbeDJrsQ5qf
bZRevbh8tby+FINZEw8YPC+DcVCqPnQv/GMBMpa8IBnvYKrlCARc21LuTVJ/GSkYv3gV48frDDef
K4D7YN/pARQC/3ZH4leSBAggGD3huy9H4JAbHGxhA5nEz2ZAlHsldZutoWdEmKZTNIzGn0yKCyxP
UJ9pPVAxSzOaafqf37lM/jFvi5voIIzB8e8vkdwevkiIpzMBKbQHZEQitC8yVlSPlcpZRa4mxu2c
dNgHrWzEZUoXy2joJvuLq8YboAi4L4fwJNvmCjxvD1Rh0XldD8OSJwkFmo6dl9EYUjhCCoNQnlkC
l6Rohj8prN1hUICeHyC32eGtbaXpWBMkDVtuokS3gsoF/kz3UxhQ/huj4dQRqTlxD8BJfYNNSEtL
gw0OgYu1HT90FFKeinx/TiJ3uUoDBG0kd0b8z3hhRYPaFRQV6ABKb6ywGnW8JXopMVFK0L4q3NaE
8OQoz0vvLgh+KFA+kE6sH8kU9hw/B422NbF6/X5vXkRirnVguNEWCrDukXTRW6nttf7TIwvshp/O
sQDQPMestPWZX3A2DuQ18Eqh04Hv74kqWNE6b50IVhM0kR6HN3P2Pqr/7Bp097DSwlIw6CE09F5a
B/0FR+5uMNOdvVPRaN+91GNCt7DMeV2Uv7P2otHaQNWqG2eEr35/du+QaYnD41MM9UY7dl/p058k
i4GG1KxPmVopfXXY1xF4zMZi6Awzt/toXptNvvmY0w/TW5fF+eikyEXs6uzn1iJTG0Z96P55Xq46
0k+sFTJuILdZMekI8wo5DMGwyOG7EYaz9EMczrQbo0vTTlGMT1AR/HXRv1/Xw6qU/30JEdVhF2lL
esomoqkelIJgtrkHrWxmAWI5OdT3TSv1Sd4jyAeudewrdR/mm7kOLDsAc1NOxzbzq/PZwBzMxG81
o6S7+/KkD+tcS28YGmsCZUX9AtAdLCli1KarLiLl5dYpTGef3FvosPv7FS46jDdp1W7jsgvprjkf
tzm2E6I4OkHBzvYhlXfohXiIx7XH6JNA+tXpAGIDVv5uy5CaXCqcdA5gGsWxZ0k2ZAJO3grUwvR9
Ey2HqHeIoGScMGXNtjQqvSpZJDgJnE7ISXdXCM4yb3WU6hMe7y43gMBAPlR5c+8QBnDFwCKrtWaJ
ew+Pxd470qpxpLDpKHAlhNtxnltYnpSPo4fgoSb1IZRlCc6w2635Y5+mcXjHgHV94aBhEpRvXB3o
40rm+YLPS7mPMWs1mbSb44mQ89Dzq1mBexwwwbpYwcr2h5X+RZP6peXg9YPSltTlk3TXoDa8h8G7
MW1rHpgJh1HyffbB8gJ7SLCEyJDLNM9BYKIxT+SZk00uYZFS8c18IPCDMRLYHZ14K/EML5CrdtAv
A8wCQXl/QlJg5Hoq8o4HRtTVG+4z+2aGKOP+eOjlaA/DnlS+6T0tqCpRfbjiP+CR+CHnqEb2PGYw
A/Pap3y6MPhOUmQUGhff08LzZg7tut+YszsQTkEjFp2FwFNAC8m9QUOnqPt+MTBJ0HgFTVGOjD9i
6RVzZsAm0RxJJ4DDAG3RS2wU7Iy22VCadbluHBArFZm6SDLxR8zrSJCCgmO2xE3APPn1/T+UV8VK
K6XRQQeyJ4EguDWg2CTwQlwMldAK3LCR+fopvVEANLZdnLFtrP2/y2lUSm2YXb3zMNFNTKdEG+KK
s/sE7jUZYQ2YoFoH3EDHQXGj02rwV2JfxQeJ7jXA33WGaOG6Pd+3QQZT6vyXN1QAc7jtXv1BKIAd
ABTMf8KJr/hxCtFXQZON7fPzw4CwAgTbCWnZBHGPVn8a0rgW2DAQw7HOSQTDr/ikISd7Z5/BuO9t
GpIponJoucCy2X2ZhFluXlJpYuH695O/+x7FD8nLPMTLOJcOBCWgO2CsAGqqoE4Lc/YOSnCzDvI9
JTknlau2rn/jksSmkYBeOqbNo29SMjNXZOyqsXkkMBwvs1Ydg2XQF56vSFuMhUEYBORI0CJ7kV2j
HIZimK7MiDriKmE+XF/HOMPoP+s/hcOzEm6mVsyo0DHuY/xrRT12nFzNbqI7RjzMyUA+2JrQOzDG
Z1LN2ClWPREEcA59w03ySkKPIHU30FnIFCQaJ/BZCZI4dQdWxPhuMan+5ax4zMFZix3qJgaR/H1W
/Lp9IuwfjtIXJQsYWr1NZZhTSwVP8VHneh4mjCNw5/GESI+x8ZdhPnwSGdv3D6G105qU/4P7sbXu
nJ/9u3V/jqV3IQvOeN/Lv1Q82vRONDc8OnmJkSr+AmntOrIQ80KVOlrIa5WKndoMthT94JjvYfdX
eaGS8e5iUEaNe8rTmPEDFVqAq/n8uvTrKaidyi3cvCar0ntaN2X8hh2wRnz3O6rwLaKTgze1H+LJ
HzhfJ5DwttpaAVrIPz5X7sGA7EZyxI3aIEu09KR+caoyCdsoH8VQOHZEb4zwBmovCpWsLWunMbPI
FrMVtmaiPRki8YmHENUZQD4Qu20cq1N7f/DMSYvIe9EyoF9Po8cn2bYV2I/x8m+mLBOhQzF1Yesi
ez3VUo6WTTQrPORmtcpMP+l2Jh4uKOHdhEAdhPrcNuwVXImdJxM7jQrDEJX0Fi3qs7MrVIMYbfm2
XsXig32GUaVbcDAI4Qt2viM906HJyHihwPdqlETkAoZzUrDs5zYm7O3hVheHC0cuQua+1P5WAIVQ
n2GY02FnwYj2ztW3KGOQ2po4rW0KaW+Ue40e4QnXow9IkHCQG9XIw2IHS/M2Rz1DZENJRviZsK4I
QIBFAP92CiDDZLfJYYKr8NuS94bA2CNGGQ+CKKY0WR5usVqBLbKiF+bDbTECpX+tfzFqXtBqBI9E
QLEYHPomDADmS7NEacSwQLn7vlDZ0aE7OulPb8saeeVCFX73d9fMja+BNnck8UHphZwq7/VHprUs
oXBhJ/qeXAC1dXhrdK2B/kXPZvNJV/J28fuUDNsrL0U/jEG8iBus2wxNGBArsrlKhS4ZwAI5L44+
FDPIpAz2DlJh9DzW1i18tAn+KVxI66XHjzOsuK0rfUs3bDNbC4atp3rOzVgN50UPEKAm90EvuIzs
GyY7Q8cRcIH8LNelwi0totOoiZl/0z/qri8F4VflrsYg40LtXRwv2luP35UyTUwag8pmIRVkdao3
7yJ7Tts7gPntiOWQrfecgmL7jkJIfibuQ8A8Ko8u/WeG4s6u2OQYqJvbdUN6lfdlRZkLj5i1aFTo
JyymlOZw9LzQ68ixb5Z10KxNqT/WA31mxrruY35RVn9erEdwyuHzDEH/oB1uhih2rlttUHliFoEm
Kis7BQzxFp1w757IZ97BJQIHekpIZRBneAftVtua+DPB0VwMImU/p1zcqJQAZLyxMK0RWCfOnhZI
Q6csTDp+rN+WP5vc29bceMA0A8umjjkuk+MihGQv963I2so79e9A52jrOrHnkeavhfZqTN+6ZgFQ
mHQhFsxPVy3s6e7ex+ci4bgYIiONy+j2motVq2MQJasNsxbHyE1T2+3R9c6TEagPDqNkAQzUDJ77
4Gnfkhc/EoCGtAC7uZ8xVgyqGjm4JySwmooMWgNnGYxsr71iN7id9vm54NuCi9JVznlp9r2SQILu
hwSAOL2DDo39pa3xBjTSAX9wNKXtpF6CpBlelbsk1UPAoTqLHIAJeN4Tpk3gaaqx1Or0MeqFrpAg
QfPTPbGsOCXDzpshIoOWCJSQv73aZHt7WuqJD1lIXPXiTUvOVRCSj+NbAgRp/SDoCxkTcN3QKI5A
6YsJapqjv3O0lCubidONCuOO/4jn+f86qphwS++K39wc/RxTxwFA4gq2dEvqJeQTFovo4LfEf7XW
YP+y+UEMjvBMC3xA7OPocR+94kd4GK4skNADUumW4SrfB1FS1HN1QxO0WPP6r+QqIH5TfAJDWxYY
Cm8x9iYKu4p/j6g1co4jqrxL9jKOyA8hg498NFddgk7KyxFmDc1S54Cohsb5GnUkrnfCQJBKw2xV
+VeBrrwjZUXdWfOSagV7T/lcQi8Mu2zw/1R/PgUf/DTWCp4AXbgxMeER7zSZeSpZkql98pJDUFjL
SlyRc/GSPN4mlRwLONF5D6EcwQbQ8wkbLzaxLfXPWM76ejX6ld+09lpVlSPPfEOeA6D7vo05KScn
CzoCV86uvJ41XwgKkmYNTV584y9ELe6k7R3TjYEC4F2hROo8+W/ztBq7mjqwC5yakG/+ykvZGk4x
yBL+8CjOk0nSR/hpUXhXVJIfJgqJU/qDP3OyadNI6GvVzH0qfS9w+nvZ1RjtyPf5buNcHltEQAFP
n1AxZ4eEipcLG2kkCOCgQ0IdbQnWms3TaanxaXyiLsRIEPnnHYarag1QTwwAHU36p/CszF849A7T
UzOvlVTgd9hjsC05BIXhIhcMdE/s2FBCfKujizVCWu3SFgUTVUF0cZts6vH7pFnVzbrweqsWweP+
HHQmb9J2cs7AYjQt56KSgfXBUB+s33qZIpnRS4hUYLpiTP0u1aH0VF9zV2thcwrJwuJVgStmIXf0
FKT08VZhunSIuJ31erYUVB4zWGOl3v0zADiahY7bdUifkJgbOPAZ/T2Qe27o2oomzxKRrXW6QXAw
Vd5TbkWOOiekyCNvvWeRi07XzVAXIBc8Zs3PLOj+EuIMrfy7LG+nuH7gcB9VPPPL3sK8kM+R2O1H
5ts90CQJ9wS8pQvERHMpBnlJ8Ug7WrQ+4XsdqIuwpIDJcYHQcfuk55busxGMIYjaayaA9JFAAS/h
z73GyIs1qvg7alCVzyelOQeggL55iaMPcWVvz37hd9YWaXA1nxrBpkzQDalWypxOo0eMX5N6A/BV
SXVIqQ5NIVpYHvfrFHGKLTRQrMpf6E8bpZylMI0YIb4soJfGwjjc3tBGTHIIOVMUCAakZdKlJlW2
WC4847RmeUXh5QN90dSLrvIt4RssG8xBQj39SNNtezGFfAg2LYbglUH/61QL7FN0Q7aaNY05ikdc
7SSxhh5I5byD0SN53vS925k6i36gMIFa7GkYYLPXkgpOzOudseppjhMLk8hKxQN99rYDtv06u9gD
DcDwAAG9X0yJLf/oFkYKTdkKeN7aJdsNWAb5ePCuQH3MDiD+ufwA/cQC62lgW+ltbJVLAqVQCtmM
Kd78CeaiZbLwMlGxkvGk3U/bASX4d8kD+xh6+B9gMew17P/6Mx+2FSYCbOwbgbd71juqbogGoPVy
9cqu6fJBFFx84cOO7CjBV89Fu7APiMJzh/Bwgh+X3fvPIEMaJgkijaodMAo15BXUXzn+lUuupStg
ktqHsUxKM1DKt8uf1ATzE/iBk26Q2EZXCNEQpuDajeY9HkXdZzDQ5ZVVB2CiqEQ7VaI+yHsrE0E5
D0jjYNdy2Ltdf8tIIVUGK/k23HwxojEzq9fVw6Zld2uNsRkzCZfxK+nUj4c+2ztqTEa/EdP1z9zi
RoI5vxI+LxN5UmlFcvR/6tnJh2Fv8rYysymxThs1Yau4/MqpVYS+1tTTRiDe01q8OhXIKBPO8t1y
U04sOmX7/FGQilmH9RL98mrHjVynJcBmN6HA7vhgaIwnwP3pFunW1U4tRqZY6mrjivQbaD6ZKLWN
D4L3kNsiu2t2R1ODvMhRF7aZMQ6d3+/kgN3dIre3OGLO+6LX9siHmeY8g4IZfIYg0s783Q6a4IvU
DRnJEd+62Djk+kMeGRNl3rRKKVsIDKvRZk0rdD+55E0oE7uIH+WufdS0a/4rvHNKfj9FLtgDti7j
t4Ut+jWMI4ZG9YDuyqCF6rwQSj7V9YoYrTE1dEj33lFjgpmzvz6fPn7WMJXEQ+wv2WBnYpVz5IdY
GJqp47dAivtmfOPGAsLQcVFk4PaeNSGPl+eoNd9U/ZC2Pt2wLjgk5JZSQOMk/Hw+1iZopM2i/y1K
RDd8V9mxYl+36ap+YtAdig1zRbsxQ+4bEGRixhgk4zeO8TC4VaTBuDKeJUy06wd/ytHoiLiyaQAY
UrmnRBvmfY/mGqsz7HMsJa51kOXmUh2/x2ws9CJAB9PW9BdWYft/7CljvKqe8j9Qa6FmqAx1HDQk
zojpvPPpswakdBe0Qc0CZwgTlxYdG6WnmtguffUItzicLN7EZaHwjrRoxRmHWc5KHrCksIsWDmJn
D+xx+vSIdD5cWa+J3HMbhcyub4vLo4D81YU9LGbavu6w2xEK4mXqSQKUndpxnaGw+RfJQWnb4395
MxRwxMznKuy1GDurrCSiM1u/wFSqlGsjC8NZY/9t0FMlSU+VukvWjbMYDC5MCEA6ojcmex6loPR9
07ByVKuCRWfdZ1UXatjO20sslQGboWpSXIDkXmxUbFH+TtjnCBHCz+1Rh/3w/cUqxf/YSGIAyw5y
Fi4h+JTPvR+E9Kf9XDqUTS6mEi5N3BXFqiSLEzVnG2797TjblZy4udXmcQUM0b1NjjGbEDpfPtQo
1nYPD5z9ahz6hXw7+RuiAtO4bW0VEtbDqnRBgMMifInV5W67sSZs/cnTNBvMyLe1d3+Zvuv0FVak
0VYLLoehFN1Mc8/dED77WardSAJvqkPUFC1Wa0Jtw3Pd0nvddOpWxx/l9SpPOxGNGq+kzc0HIeub
md8OxMFbDSvhhXRsMroVvNWtUHmwu2uB+svccjcoLJixviSlfdGi2D/xuy6pHgbuVacIbxtBVDna
fItHwvyNldtUtHXTKHY6YOcsGagw/WPu8UDC4eAFVpxLd62mBoLdjX5OtB7BiNePtvMe8DZFC7V6
AKNlh/oLjcD4JLH4oX/H6a2Q90QrETBDADs9Y0wC22b9IQHQkm+eC+fTrYUF7McwrG+3wSDM6PNb
NWC0J82sE+4jZad+Ts8Hv+s4H0Xs5Ywkcid+G744aC6TXoCg1dRbzrxc8QK8zg8GmHwTXLsDC8JT
9dUx0ElHUq2VjzK4wDCDIoMd+yGt5iZxhg8PWEuwkH9ppXQDzByxFV9RkONd+a12u9oGH6b2L0Qi
LiSi2//iskElEm7e1vozc2+STWVzlsXH4Jl5H3KGLfwsdAeAoPIlTt4DgA81HN/UCdwyNtM6NW/c
H5rl5MXnn56ssrAY/bxk8nOYSuXGx/S0Pqv6GRdnk/9lT4z/Ei8s+jtwQRzu4/NXtvZKaJ4g1YGT
Qhb1zkBEEa8N2P13ziwV6ltLLSJCDVx5zVqVNuI1gjHpG2pNe28Lqp6M/lUDW1/C5lqrb5zxf5UW
44e+vMkKvcaHNDDqSznkok3dW6m0bMtZHCc2zUyJag6PSy8/vGepZgq6SRteRaeffdr3+YlPunXT
ksWzHrpsOAFHQgAcLIDX8K8ReDxQammeGv3jp2QXSlmeCPyYNV00Lbawtee71P3k84lK5ci2DQN9
lnP4J20tlJ78u2qd+p5xhIbjTK6t5FWPicJYMf/ehnyo52EIx+kxvgcu+sUubWO5xDC2xF6Pj2nu
HwFODmvF2x7Yab2g5pQG7XDDphKt9xWwzs+ipI35urbEWXAFwEJCUi24DK81Det3Ge4c/WFOgOYt
eti9eLHXFfgud2XsB/gCVP8LKfiJrfDmvNksRVidsUVH2IRlQU6KQVejdE2jynEDEeO3n/Vg1tQQ
j2coO6Mb6wmgY30m+sWPUnbfpOvMYK6s4gHHCxI1uC/JeVwMU2yfZtJAtqC4y0HZ7gxVe2Hk5H4K
BX2eG/xEI+Wpkj2+uPnSflg6qF4CBN2W+QSCfY/7T0QaCOeBXWJ0+t7JOvG3+kpGbnm+vCJ/VRvt
nCtgBLWrPgFv5NOCrdTnKXsJ2X2yuvuMih+TlZi9e34dg0hJK/F5IzOA/pMe5LlKDniVtsb5Q+j/
tPZNdvzFbV5FhLnzVkPV2utwXUCgUvlChymoTWKwr/ypZnTKGl9k6a82vxjuMIhF3dUr5fcr2ZE2
kETOQKAx+NzIigVotao+29EtspoNlY9ylV++02Yz7Tk4sKn3zbULyecBXsMezj6p0Mv5EOgth798
yZie0GpwxDYwIX2ezeuoigM3TV0wsoX+COTssQqlAIETb7/Z8YXNg+lXg9E9xDbjUTeuX4EWafjv
SZJ1MYmsocZqfJYR66nuHEYWHIkfMe2BO0q2ztXdfktJJH3yXCxu+PzFWfI3bJXP0Ska8Sh9d4bB
qbLbYAHD9poJLzYsLI6Z2blsmUiPB42S4kJn+05uSkGaxipBZZnFEe1Nze7zBWKVPIxE9qB5H13x
Iblr/gJA1KIEZKwo0IihWCdczeRoOCr8hTmKLd727bJmBOSu6yLlZ3YpmGzacmA6d394t9tY4pWX
j9SZM9qGQg97MTvUJQb2BXFpZEtj6welAfIH+qqhC5pAYWwUAP1IRflhypRcWmc7PzA9OQsfhqO8
MBdPfEbGhjNizm7tbSFtvk7lgpAdGtYMmNfFvxHaGasOpFjUpKjSz3rW37OaFHgB7+DFjUgHKMYi
i2QZ4uk2Fze74xaK3SbSbtd5S/sEGjv2Xr3G2oC5m/3a1v+hVEGt46PQ9QQoAReh8dzQg/AYAfFs
0Yw/DX6L+wS34azNYqZmZWXNsQuEDPKrV7PNJysn4GI/VdG1vtMQApCawFOSIJN2LNKG7L4LdZxn
yxkls8+7QpGUCT9MGCw3N9EeFm3MaezDjmZ1qfmunE/GtkZshKP+QT7mNVpgYp2iIVXWhQ0Ntvuq
/AlcYFwl+cpLWIc/Ew9AEsDdJogkV1/SdyC7ZA5d4Uibw+XDWL36N+kEz3eGF4XoOoUAt8jSeyoQ
cOveZJ9uM0ziV2zpiwQcLO0PtMqulJ8m7P+2EJuggShWP4As+dWp4IQMPZgCmKVgXkUGXK4ghTk2
eDCn6rHuMEaPhUF1wZVq94TfU4R9nrZvklM1DCKR8Q38yMF0dtfuzzwXinuGMjyupIY13F6p4gDg
TBAjpxQ2jQYGYkixHFn8s8ZSuUpt+H2PWQp+0zgi4dFtpvIrwGtYW97XSR8xlXlRRwIOf2xY85dz
TTVNHFruRUoGQnPDAweOOSQ/cr1mP2vmcwdayG6gtWMtLhPWBFEuYmlaF6N0Ikk6C+Kk38l+YN5a
r/oyIUY91cfgGU/DEbfVUd9Jv4Y6FbbT4gNZ2+N55ZTwCiPUwf5d/hDjEcwSBIm2OC2mCItDIV6B
CY7mUg3+lRqFsZq6eHmJTR4VOAHyKtwGqIhQfhmRiIZBXZ1zLTvnOw7dHRmRc+PCEWFZ/3XzG1uO
T1Cch4ZIvBLVbPrYhqPTt5eAPBnUh2gL4qthVoZ6E1ReIymSNWE2wiwrYBbQYJ3OmaP1TaFNt2Qt
uhW35fKqzt4SpSAwX08ahFvrv4ShyS5VqI28BEuO8L8nmVhwGukoXCVPVS3GB6Ga3+D8Mv0pFreu
wIFXaoxzY8OfCIDHJsOX1S4x0PcW03rjc6W82XgZ6K2msm9sOmHDjJJj8zpw+ry56j0xzdCR5CuQ
kEIAoUy7amgnVAXHzFu5yeUXYFd0r2ZIGqBkHZ6Ngasf2QpzzjM3bGo9zt3uLJyvjsE93rLA/MkI
tjdHpARBD+Cm96NqdjV4+5+aTa7FAI9XT4p1IOuuewCJQN0QzwlC3zJQpr4BWrbFUDhNih8dZ3/T
anTwtgTscWp3mHL4b6nY2a8onWEzUJhh1u5mHWt9MtOYs7dDaN3MjlHpktYom2LVteDGq91K3XhG
EZEBHL1SREGIU51woDPe7neIUOTVNZ7RTPlfWjUaoyJ6HyhZLN+hDGCJQ9jCSKeJtYvfawxraaQs
yUOYa8P+THhJjWX+y07JflSiwmrd+TbxpzLqHcbZGl9ZdaLk9SKVHqz0z5up9iR0T0/mpt86G755
bW8vYVOF9K3S8BvXSNqMCtK08zsqkXYIBnIza7MkMPJ6MvBvYUKdJ66D3/2HvqrFN/9LoFfIFtGx
qu7MEAG68f2CLAh2sU1Z8TXJp70O337uhJ1CY42OFBI4hK7CdSDHZVhr4cAJhhi2lsITsD4lPMZq
KrbMlYYvbcx9m6xsJS9Rl5ZUIlfUgrMGnQL3HVJ6gf570ffWc/zJ5ZOzWbdk2oGE+nQ0qrSO1Avb
AeOc3QzP+/ZeE1rud7Uc6fxCR7YEdAxZAiPLFZe57++538wrXe5Bfvg97UMiNxYGUTKBFZ9di4eZ
r8+lzsT9uucPpiUbX5ClU6r3fA2cTwnK8N/ZuA96Twa4QMKnPhPGV8Fa1xejTR7waDPM9zi9y2Bm
39TJ69mzPbjOUVlYvnmUuHfSF/avtRrGoR2Wz+SroJ0l2/rXRVjShqNWkENBWFcUtNCYiajq9CTs
0DoGG6isEjP4kVQkHJL5pnpqnSgGtqm5+qvq5h95EmYqEUTLtgVtHpN0eBwGJfYlv99VKzeBIWfv
SPHxkkP6czu5fXswkResvZFc0HeP07ZinGm3QgZ95eH6hR2gSY+SGX2kdGh3A+5t8nN+UVpptUTl
83SJCTry+GsW9LW/tQTVn4MAXnPMxSPB62tFmN3C6J2nHBGBHoyedZbb0Vabx5P0GGRbzSJRyjtG
B50ph95fRAQA2OLOqPJMvuHPyEMnuSXGVNtag90ijoMtU7p4mWVyw1BHBUfk15LAh0DZsfFnxlUM
fvdKhEj2yqzMO0kaOYMfWEf8/Mqmjfe85F5w0d4TmigDTD53TgLabGjWo7b6pyHPplupin0WTCVC
a/inICdBjBS4bvkEcayMMDFszuwXgULLVObVaB+uFIv9M83imnMGXCDUtpmcNhhtgzhhuKleBvbR
nAtM9Tt2Ksno6mN3KibzlS33yo93QitHPsEIcGagqtlp6McEJsa4gyensLomk8T0CqeC7rxSMw7D
95Sw0XcTXv4egT4jPieO66QY6FEJho0OM4scNu36s5boWWC0I0sEi+6sClXymaUpRk9jDtqhByRE
w6JA/0+7YL4nTnlAnIe6pnSeeaiHrUJxX8KBPJUeIHfnR1UTcJV/dmKa769k56CKBIozrCaMF8G8
eDQxALj+BLc6Bbj2gGLv5VGM6sMFv5Ii1fpWUrsHYmuonFWmABJiEOLHX2cwUdynM5AxPHmPQEGW
IsHAgAOou9V7H7uDgS+eqHiMjN2trJkwNX/3Z8uwN6xz1qtpYZGSv9f/xge13JZD9ZvYUwDz5d4Y
otG2kdnRfPkAHBJoPETSI0QHkX31yvMev73Y/hD848OKthvbSGEO9KV3sSSdS+5ime4TluSJBVoc
JbN+OO34+Ey49avD2OPe7R+31FJQ7x0cbOgWv2DWhdgJzLYWSH7HH6Qu5EyMI8DsfR+4VHqFDzgO
bDEPiolr3xiRHIDSZuQgQxyz1s5+/5Eih0C/xIfni3KZau6ejkUEkSg6YkF3AgkydcWmkzTfMoQi
RsqISA/8KPTdlQUkAzr6cxVxooqus34wV0uWgrHNhlfabk/cr2I/HeKTvLHnOXDl+c11A+kbKKqL
b9HAZ68CFMdegQwtMBJ2yDO6srSWA0llL/cZZcHrmWJ9sbt8vzNQ0LqHX7TlywAM14Z0PdJbKpeM
/v1QGD++LLa42w4kU/qvA+9G9jc++Xi7YyyhZhWLrBQACJAyCnfHl8nI4ggw/gUrKuSjpVfRTNB7
SPCHJPKervPwjtGDSE3SuZ3qSnYKEdNEm4bdnfyjyeVj14ZdJppNJdJHPbGKvfJVgqtqVfvrit1c
VRfcD71u49XyyhVZkYipPqMCCcVsycaKsQHATpJKWY0+BDIaqDY97O6jn51ZNV+sdyZmlKnKAyuW
KhO9R12cnFTU+PxfGoUmWfAaFFQrmZmgykUvvL8nGMIbzLzf00X4qgoDQzfPlhCHCuzbeSeqCRX0
aa1SjvGdk5kgZ2gabFJcByrpmhCR5L4fWdrnUV4THTN13pam6jcL6K1DFulGEr0xh0yDtKI+UHPk
Jb2tRdsmtC1wMeR+k1SUaAroAfugehVyxSswVIe9++ml8KtDi5lRkRwLxmiDaraU/6C/ab2xD4XE
jOB0PhDlIw6nBpOYhz0caPyiNGnza/+LYFGxqNEgNl0epOWf9+pDSfb1Sw9kWohuaMOoldFZbCD4
tK4LryEJLQKawefoOPgD0RC0CbSnsOjMdzXbM1/vCv4nIaWx+aeXzXKqBaIUI83sczZHY8biXY3l
Ubn5oOcw7GNX4bOQgIY0dXgpdcEwNVYxaGZ8RVjzGzeuKk8+wIKKN6/W8asbJU/LMCHVyU5Iv7Wf
9SFVSiBD9Zp3b0MBqoLhixsneVR/j4uQ3tTvWREJwEn9p109ckT979coJndd2lo5b9aMZNvfHMAD
3uUg3BiKSdJpKcXp5A2G03JLPo15Fro7O7zijwWUwkdyJrdhWSX5MkEFzEJSRVdpQY/25zko37Ue
2rRBXEkMqUtWEQwm3QdbSXOQkGtwxgSFTJmA/yvzup8niaLZ6IDT/YEdy/nONJI0rxhBrB15dIkn
pq0WpPgzGdCiXW0Fm1+HVte4yVmLSrCXOvmx6RRkHNtfHXr125K2WA9NCG1f0m3Of4CTgNW2Q7Wr
CyRE/r/HiLD3z0rl3AxCIwdrRIDIptU29Djde/uj58MA0V5W8MEoqOR97oxz5KzsneEq0PbnVZK4
uOp5HOBLE3qsTAOcurj6DNcyKqWmITL0k9/LYJvDuydPbwrGcNLAQoklk2aHpqxnb8NwutjxpXdH
PTUfmp0OOJLoVdZd72Fvwybztljb9mCMftvyOXfcVmwiTu7TyXk9xMRSqxEkp9uaNFQ+irgkxT2e
d5PVVm9r5fuKBR1IUBz5mcTK7Htm96lRZaFNtVMFBHPJpyUN0gxnDIyOM8RyHctEIn0yEpZovrcO
5FmDTlD2Lp3vr0i27B3hGV0KgU54IydHbRuAu3rGKCuB5CzLCr+Kp+YGE2tgej+gSx8jY7OklZuC
40jsO9loSg9K4WRrAebNHTIRSVRtzeTEN85jfYPlOimaQjfP2t9ngwSeUfNckkVhIQZ3sWXTDqeX
q7ZkTVzRK42YVOq/t+4i3A1gq0KLt1S0Vks1K2kddWqcIPELzwXLF78NRLf4VSvRp6nwF425E5mR
kTOS5cIrFpdpcH37wzS2MZs7ZzOXukhqFB0cZphxoGgDPtmLuQ61CuzZNpJkOefKIdYz71DGtBPE
DIQ14KIpuXjHmi0X4prBxvBGCt2lnI1sr+mFs4gJYB1BNDecWEQnge1G86wSXX2RkXT9s9IdL1Lq
6NlQ+ZSh9XmmVPCRAX+pwvz6LGP00jlzoUJXWHg7gL9RJ6wkG9GL5zhdYXgOhv31RA9eLrWZLxIA
cZyWpvPCxoVIW2Lbq5GCo672kDTW0qCFdIIIPyk0VRk75G+dworGZVrO0piOXZTEGg3Po24v3Cbp
FKeCtB9Vn8kWMXSb89PlCkqIS/f6cq/CF8YyR+ZlMY3N7b+fJ8hSlgsbrPH3nP68MQgy3U+k9Pf7
WNY8FFlCdfrrw2oH0JYs7x9oCRRFngEUFnIaUCVMkvYVUFS9yb396kze5HvndyMTXo1x0RF7xciz
2dB3lbY4cu3jioqRBIjlZfsFzEr7/Wbgzt76zIi6M5vqxXH0pHaAafhyVlWAwnkw+hQ8yA0XrQ/z
464uacMLWIJ7L+ZybK0aiHi+9Q93UAalBxQayh/79kykWR7xRljzvk+3DLfWJrIOVgyma8yUBF1u
LRRH9k98gECBc3k2JX+p9WkLwkYmJ7RBxbaGn6K+OTCMv7ABOxXvZMNzQo6wdUAmXJHYZ5cLqGfr
dBmXkBV0xbm4YZXS7K6Eqd/Ok3JRZKBYRxDWBp5EXM9awTlzlZhmNSPFBSh65FEQfnzO7p0n6ys6
jNOA4pzqpId4ITPtKRRK5Q7B6oaffUSxAn5O4UAN1tXZiXMPchRbdWYI/mArsOF2RMl3VHK40JA1
pwyBHKPKLlBAPzjs4wa7Zwo+A1TthxZRt8B08kKjfnS5dltyIRzItOc1+ApEBoE0Nbq0g9B8otsp
3BcAIYVZKTEF/rX/i9M+Il2+VG+S6zvsYsSpSRsFgJS2MMq2fU0jm1OIwyv9xSsN6Z7mzE0TS9iy
z2q+FyUYhcnOnicl5oY0ZZZFLAsTUdZO8wtY0q4PsPNulsvkFg8nGyFSyLldYXJePa6w2Pa05rR9
r6ZOTgnKpUj0G7RKVzR4m/o3nasie1Om7Fb2gu7DCvItoPkUK/AS92aOg/CfX6helGis7tZav9Ie
/uQUfEUoe+TLWp1HBgpQq6pxC0Ql4Wzv6IlEhSrGTdCKxjTXmNE2NJv2ejvahdFoSAlHpwCAFywO
odujtfZkXPtc3VVlOcLZpGQFa9AOBjY7WPIizQB5pSSex/muup38751mYYerF49J1GUlA/SQYrps
gcYYsL4xdg9A0vYRSm8keJMJ7q3l+ZzX+QfMOsSHpQKbCLt5V9/IIRtvVTosQ7SmL1r/Flp2wEv9
oeCRXz3mad2Sjq1R/Qux0Mo2CtkyKLJvibSN9pIMoM9mKKFWtiOvLLzdtgHXJVYGzShfDbh9dqTF
zyv/oEn9HysMjNLdXjnFOzE6SyYY8bmByuOv6aFxw6MkId9kxCKQ2Onm9XJqAJhiu0XwzmfguFFX
5/qSOuaVo2alFnm9dMjO+vK15dyvh7FG7xqCVBwliE1K5QEjZCNBi0XqIDcVfP6C2kI+5fM7jpiO
zpERAaBNqdVOBt+rbOJvODuWJfBre20hly8IDG3u1NDRt1EibvG+FP42gEPTOaBppPRHmNTxgC9O
nSnM1QnzKVBNglH2D0PO0pqhuXCkhrbklj7brovFAJ6FcXamG/OucIS90m3898bF+52fyLGUg4cJ
/7m5MJ/09zCUW1RToAkCYo0yh66EOsYg+I6eo6Xve5EBvXFv01jdX1MKDjFyADa2oaIgGSF18TnN
/mALZj3DW2j5xbyyqJaEcWos4a0iAQNh2fDhmyrgfGYYk1vu6kWkg2R+/4GPDHM2wO/KMUEQv7+f
tZenevJheA62cUQbrhcpytC1KM71jBHIE/AEYwi7SuuJTkvp+96J5TW2RgRN1pP4mdnHYDAA33Mc
esFKqkEAN/u/a9gFFhYe94ybeOTSg7c+QzsI/DcmQse/3jF2on+ROSdlusjh94fIAffVwI5AIcux
lDtYPTzUnX+1gdxALR1Fp/ENqn0Jr+GPU2A9DxBoKQe3fsXhkWfUE3UvTwgFMYjBb48aBtKJt+4r
EnObk3LJ+i33QnYp3fhVfEK75IqUOyHkINVpkDTGim+9qEFXOtlbrmxqrp9v3EEugIwIV2x2svXw
BCaiItWbjX69vC5DFJfkajGOkG5qfBQtb0+kB25dOyVii6yApA8/6jocQahj9HcDcwSV1hU1mTuQ
VTqEaCBVoK2eDMNHzJoZewfr24cNjR739NVDM1Wa4IWelfs71jwmv8d8k99mysWf1SOIcVSsd1ko
5/ss+Fu1rTJdznVOOQNr1Xej20OqfI81T5LmODgizv9fIMSsB0zoZEvK4i2J359gyrj3jsZ2tLZ5
QXguhqoUbETtDoTozGvTX2Jxr5+HDbRC/J6Y645gmdhfsxZyvA+Mv8E3tiCaP21MrOuIx7D2JTAe
y4Cebb534ulvNa1iae1JOWanmU4mrY2emjNanO2ysN7pYX1kFEtQ3tF5j63dxTHs+uHPycAivBi1
Uf8X7W6QJsXZ8w7qvqXNHgPE01wWoATvay4JkssYBrNLeNdwO/eNCRpsot7XPc3ZsEMdqmx81WeH
HzvPkJTKOn6NV5VBpQx/KwnDVJe+M1WtkFGRsTbUa4sxmfgVHg4WSmMct2APTsj2SzcOpkAvbuCz
b84MdL7dV37mr96pbJt7cbarNrxw5G3etmI1RqA5jGfHkavxiv/+r970N88sxji8HIq0vEiw3nUF
KYDT/IlTKXVgInE2n0g+/9WXS0ABRxDvBzIfGDJ6i2a4swb8+bx4Bdh8lIQt18ngjKJtKvSlqYoa
IXULxgm+srZAZfVXgg/grrXmPa7E9MPqMci7o3dW+zQ19HC7TJhG1l/MidTGkSpV4BZykQoPmO9k
GNdacyn1gm6/AEdC2x3ZhCJiygoAoRkIbKi0RxShVwj2CNyGWbV2+bQDmVasPtPDhTh93Fw8rlCs
cxkrWZT1Kbedof5quLRfwQo7U6orY65/CHi6EhGBGiVuQ4aXDOcr4fPAOI1VXvVbSPVmkPLTpYx1
PTEpI7+LShps3ye0/jNnenkuKFx2lylxN5DHCdsRG8mlA8j986w65DRh+ip5DDpl3WtZTo230X5g
haHMQ/l+uSaioWagP3X6YWyGESKDUjW9Mv2BhirTrJy3XO56j1SJP0/peMNhXiNjRJhrDKt0rEjA
CIBOkjFVntK9DmNWk8IMigJIwn2L78vSQJQehmMa1B9+FNty8uA+w2n4zllR9HVhAVlMYz7ukWDy
28dfTYTD+no/VHeBZStVmCykZtyLUb4mT2nttf3VHm3vre+q2Ij34Rtm3x5kU8wxaormbmBr3syP
TruUIEKjTsVN5KLjwMJ3buDjPfvOcCbr5IDRvotpfUXRFQebGX+q/+4mcF+nZw0K7kExHOSZbbzz
aQV7Hc04dcRGzrWuIXSXsC9GjHREDz7T4ShRDrbjdRpAwU/YrzJV4X95iBGUiQQ3djtGGIoG+ga8
6l1JYwdtyAKakjIrWif7CTPiG6pOQHYDVx9TIJC7PCy2j4HYuamAiTOpZZMOu4pYYTllxQn6NAlY
0UFIJZsNYGTrMh8GCkckevIRvkeZLJ6Sub/V8VmPINx0JOQ+oHvJLtVxx7IvtuXs19I57zK5YyqP
aJjXDoLJbistGULcNK/iM/u5ciLHMksttp4ppjzgCdHlirYcfYfyAUiNBooLkPlCW4yPyq1ZQZ5a
uaY+wHyqm7a3bq5OEESnOnoR8CzvW+zRXuV66cjhNC7ByGb+2Lr5uMHRKZMXhga9dNTWV6tYJIng
o334DxNCGVdmG/hXn2ptq9Q9HUsYTsta+EI438PN/WGPknjRqeDyu1OB7ai6ULNYKN8FiyW2zFsT
z4wkhpn+sLdAAOOnXgCRxPU5V+TtwDJrng+syrZO93Nw02MqsTuSb3WrKJ/mKGaE7azfm8GYjtcp
hmOd8rnEtyp/V/Jgin+J80jl1YehUB5L0E+g4M8O7lvKTslsxkkz9HLxd7MUN0tEo3NZWvclowHd
2Qt2sx5zYtzS+fLt0w6+GyXiCYcha2PCSGmGFTw+tWHdomn5+MfBjzqKXwmBeT2TjRVbTN1SgvPG
FD/f/1L/aYmOMedqg20P0CZRpfZzfs0Z8L0vxIoVsRLviBsp9A+WkJM1CHcMykUoe8qZ3h1k30Zb
FputhMaOXQfmkmo5k25FHs/6XodzRtqBnlCwTUXo/2Ojbj2oDf2hUuSph6XQUlqNYcdFP5ZF76V4
K4z8pQKz75vWo3Tmc+peXuLI7Aws1eTDsLCW8iZXtZvYXU5aelpXvgKcf808nFdHXGIAarU5z7qJ
w5fSmY3aemTPHyWVgp1PsaN8/X2pj/0Y7FxHqCuw1LnhaB7ABLMxW5YsQ45LkFf7z88GUjun2Tt4
cdDBCWs4gBEJRPG3l7oC7KYkJnwnQ8m8Ia0Znyfvza0DM/zxZgqTSB2NpJDwwsfMjv/b6PACyc7r
yS+XpaPkSuBuoEoEKm33uNuh1dMK+MTa8Z87xKwiYNn2RuihG+sbRvrrssn3e8TnqEKv0iHbIo3j
ZXJCUysGdWxHcG6BYBaOdmqCMzttqPsqWi+qtd6gxxCsOlpSSuBAplYgfE2Q9ZKAbp2HvIwOjVFc
9qmLSR4P8ZPS9bDnMLi1JIRVgsD8uHK+Q2v9pRnbX8MaTxK+3A33JLy9UJJ2njZhOljl2W8HwH/c
h+fCSTf18+YKMmeCjduilQ/1GwrrKA7ztUSEBCmNli8zwji1f+qCdRUZDlKreK7zBTjX6haA0Yo3
FBaHDY+TlO/+HnPZfu87v0A5b01zrHVQqU1uk2InvCtz0dPaI0mSlEEcXMjdahShP7Qaeuk+maO8
Itoc4RoSyB5Af1rKIA3Ch457Mz1xRoOJfZuw29q/DnPfXVLYCtUVCKRxJGXV35aGYHSxGrbKqPWs
z9WTi4II7uvv5PVMMLeneE/RIwBXWPH9Awvw8n3Uol1ygQiec64n/0mSJmVpUC+y1w7iNFfK9se8
8HjMPrRgIrH4VIUhmT42EqVxbttjE3+/G/F7j2XAHeW6p3H4DfHN4sb6pZm0xGyW4XVc2Euzb8Q+
O8KGx6eY5C/0N4hvnL6SXloCwmchUPG3pb/gwITWKm/HP9zcL3MYbYV6PtgDo98zjK+2zRAyyng3
CHbAf+TmzOSGNOA6kBnQpjKDnHUDzGjaeXMqejx8kKwKQOfodJkdHgpRaGCKuSUlsqPMVTbCrQIx
mojcbCQXL/ZCNXSW7dt2RsZXNsZubenbPNeGNTl/HzSmnC3kN57oK0DNY8q8UxllqYUnjhYo7J3E
bTepMk/keBxWENCMY/YH36Cug+eY+PYsjY8zoMeN4ed3sE+yNiDLkhJdRdJqP+vF+S33cYB9EudJ
ASFzZvvP9ADBCYQTvDNHpaKEd/lvfFTH4U3dVj498vBSjLCpn0989E1Rm/1yRqJiYm4clKFpbvQw
moIAEHbAKb4VVhnANpfbo5g2X8i5TZp+MhUyVAKlY0iT3e+9/C4Tc1DMgsz9FzGrlSbDX7TYhQ3q
t5gmb//pvge4p6DO9YkhzwpkVEabJ6q1TOO01Ghb91kk9xbqi878+2Q3aFe8BMMTsLmPJAc0yXfW
3GGQ9Fu7HAsUv3GyQT+mo1LKylf18Cpn5BdDY7anKnaUDCYsju2M0mTzgDxNGWziNc9ZFVRx94av
7emhUbvn/7tuib4rLmlBQtXTcPFOP4Zv5Dk8LzYhvvWqin5AeALrV6b8EvGcx4yuWtGeUAUOHILs
2VK6I/YX/GDRFdpiQ9LTqiQZ4QWXg6MKVPWOM13tBsbs4pzYbE81JB/U0WG92zagkmtKJ+ghVze9
iyshGPrMRXDES3rugxusqEsHSWf0ab35yf/4fH39NVDTn4K8GLUNbRA6oRQ5o49fBCKCJ+8/yJrs
7lQebWgJy+T1S241/fHD+7FlphzOe2eNanVCRzm4NMZriJIVv4nQx3WYYN37kG/39VyxAsHGKV8f
q+iiGO6lppRFRgC2+UIKxcXK3gnth+Bh++4kq4O+q9LYiB2sSBjL+hRwHhnjvo1VV9jmVtTS9FRn
yfLGGMj7/8+ASotgdDsP2YMn9+S858R+wcFK4BvNrPwGWeScEjIBOiqpU5Nw+RStwE5ub+3HM62O
X+/QGwKFCi2Pc9FumEr3F15xPSKyFmnUCq9DF30HpDfayZkraX9663FxmJGWUfA2/K1nNhnFASL/
rTKpLqRM2xlrtsuzmh4VcqxAzQOEDLMNGUPSeQH3TLJMwTHKOfrQkDb9ZpBBVy0BZrNilCajfiYH
IU3MGv8NtAWI51DrDiNXyaOBoMrbNkkxHvTEmUQvPK1OliOjfaSbT0s9Dj5q0qOZrDBmVVahYito
Pf/a0qq/00mi9lBhwlX3+eyqrwimFgI5getCTcH1bw2kauef5tn4dGxB0KN35WHg+ulvPhV1Yq3f
Fs9SiNzTpHheMxfoJ1M5Guoc1EimuPBd6WdeebPF7wKXGzO1D6AeWHh3REsjUmlDTWcVzfZbW1aO
wlMtFI23kqHHAvElUPHoHDvPDV2dFgy6OrkGAoLeMR0olwmSX9iK0SrI4t1IlqVenTh2hILyL9nL
D2H2CGT12t7nGerlqsDst3Qenaji3NXTJmWCXkKDKFRgRXZ0R1yby9C5JgTpz6/TzKNBjfaRfgxS
nmq46rtwE6MDeRzQbs/8qLPKkTnVrtc+Q2zwEflAyy7hUuvWz1PIfITkc2SktOjqsb5fNn+2LdL3
L9KPdcT6SUbhEvLjjWEReXJAdjhKkReQT1P0jY5ekQ6Mi4M+J3BDzuCGiQIi64R1PuXvhW9NWDoM
WkScbY0SD2zmFQ5XZ86Dfs1hlMm8CQhPq1WHTykP5bpswq5br2pgm4Yq357oITJfuFcHmnLiKtMp
FmeGia8u6MpSz23SflTzxSuzl/hcQ8ZnxfucZNLOBEs5NoiqGupT3j6byMh+TML/azj5muhI8cAw
8ZI/NmgyrGoXJPD0CUPHGL0oEZQn1CievjAWeaAY5Zoab0DHmNIbwLMfYduqblMosk0AdTOLC1r4
Xlj091yw9psy5p2U4Ls7a8lmYKMgUiL68eODRby64H14koOjfhuwhxBVCD3cjNOgXN5P521/RB9P
iXmVR/fd4WZ8IV4hg9s0sB+/ckVYDcgPn+TrMa3S6rsDcbk9jGcK79gTBbB4KP23yc6EriGJfTSt
+Q5cTol66GkbcJm8NF1/7E3x17caBpUOypcMt1GnNNizcrgV4dezLCljnKv5m7GgqvEggCCHLiwJ
U6eGVSyYEqriklCKt2HBzXG/rfn7Qu6vy28gbnh5PGxhmEOmzu0608DUexIP3pOhHq25CTSnCOiu
j9IzGKvxX2Z+2jw+6+paAv66NCgXTVkkdgPexF7vqmr1/WcALcx6lO+5CoeQo2MmUkJFCwgd7D78
qYbQW0rJuP3kiCSEpXr3hpvmJO1FyuvHeC/rcNN8h4aIKD6POyJdRDBm/hTtHejxF3WKBGbdr4+1
pX0a8ZazMq5KMHJfDQezdjijXCs6KNHDFV/6UypC4kAg7PwvaBaMezxixNA+IHSp29c6dQm3i3TZ
bCk61t5S6whg9A2lHlzF8fAlDi7yZ+Kupd1N0cvLKmJyEfwOAwL3KTa59VwD6P1vl4X4wPtQS0hC
50wNUDa71VL7mP0jFS7xfMa3Da/DrWeKUU+xn7krV4RTDUd8FB0fdy8blLsndHyq57+RofZb4/rR
teRBeKXb23fKVftKJKRHSvLdfgNuETQAY6rLP0ZnaF54PzH98DomOvPXD/AZRuXkSxAYLMZH/rFU
tUiUnJR+LbcrHWrGXLphv68tIie0WCqpK0wvkurNLZ749CGBzEBXHrx0tKgfWSMGRLF6bVgnonJK
qGuLoU1y42bsGOvd6qOo/Af5NKKNXxAx0wsmRiOo5euQ/CzctV2zcoBdiRXGRvwb65hfaxBpRgiV
kUWRPFG0Xuh3dMXdPxTKO2rgjbI0/noFwADQTzotPNnGzRYx/aKzbodNGYU0tXax9IidOgmaHgVB
EckptwM52hnGQAbFa72FihvVZ15V591MwJAXDOUXvmfxqSqqIKN/fA2QRgl/aYtEh3mgilSZ8Xpu
9YhoP7qQD+X0O8BLmIJd9iIa5e+j0FoSfUyWU2mq5YwxHd0AMFvaaXUK74J5J4VFVZ3OVZcj3Aq6
FVn3efAN3PsvSaQjDXJjR+u6ShowEjFf+DWeFvmVIOxjAfqV9EgSwj67nHQ4fhmPVKPp+E1ND8+5
Xbd3n7bHAF5Ab8hiz1CR5nBgmgTFkKFWQ2S63j0USMYHpzk+PDneD2yhSr0XRT4XOQfQhFFcTuAt
tsRXilgWZfnlfClpajTALZ+K2PsAfeDhcD+PZ5WS4CudV/6O3gYq59pPsCRBte1st436x8MXygvL
l4Lt4x/nYIEcnoMyr2x+g7S30FtTsY7kjEVInOciDhy0d+J5edWpdvMRD8JGmMttycHxyc3glA2C
PGzZZPLkri8yMALGsO69pGJm5O6HyvIRX2ENzJnrz4fk43qkhpotg2M1MdLl40EKeSA9x7vlFqGW
6h3gzUwdzYuZkRpb/PpbMMaYWbDUnQznsJCioSL6881VUisJwpuCgdMYrq9a9kiEGkn02xLSpnE5
c1e3NaO3lAo+kQT1qwK/mSCThHOLDl2h5UphBVgbXYoJg96isFq88urzJBfwyiH5YrYaVw27vnpm
ctBOW6iHHu9AkHspoVPdIFAh4ouz6IJTlZ6WpY2qsduvTThZAZMSBNZZR/XUUEFuSvMgyKozwPgs
JH1P1K/ZqmH1tHNf4DyGUkNf3dvs5vLMr+K4lnPFG7UW0Twm7/qjTMQzGb1x9X7o9bDO8vur3dK3
FDm0oimebeq0i9ZYLpHcdOkhdd+6Sm4xhe3b3nbLoxxJGF15FNt/LzqE3+F5xa4JJb3EVnm4Bzpa
ZhumVPC3Fq6GwrYeQ6qyRIg9OtuukBQdPsnUxU7S3av+f5LrLP8GOYPDfpaWxaie+u/fPtfTD8WX
+dBvBSSXAGx7frzLu0VYZl2gb5S7ege61M4et1chpRQg5bS/oEGafDqVTJaxpP0Ui9YN1Sd/Ezwe
6Dq/Gh2WUISApTL1g46EpE/5tBZvNe49AJiSsb3M6HHh5yZc9nCIbMG3FWkRUhSySHDTvLQYXiIX
lPmnImpPXxmLEoin7YSrTrn+BXr1b5FEf6QJRS3RlihaBgUCf8WJRh1WNrDHQubIGrWt6dLoEGLa
nh5Pml+l5l+gBvFyL6/q/2BE5dKUWspeULacTeSFwxqxHSXq34Lg1BGjoDly6dkyGA3wjye0v6Cq
c4zh23tRefyCKC51Tl1MfyqbfPPOL62Ax3K4Fv/k2TMCMHdSdurgcPVJMATdJzvya+9Hz1agRrJz
/3oW8TW4WVxknOqcvJzj2GRPxNExa6nRemDlGxQp5rkMJ8otrmSGL/bI8C02a1pmCfVUfqwVgg4q
WYImH9hup4P/hB3aOVq95VHTPFk94zfuOgQHFU3ER98Pw9NwtJraAMVSYvVk3ZjXduQdEwtno5RX
qFDv6rU8HLf0i1/cKkdpvzvXHGPhY08B2UbfDXEPj7I9rjBGENIYnyeTuEhIhsXl/djKlJlboN0+
DPQjG6A+MwBgcPjDW0jdgHGsMvROCeVZfJiLIr22fM0r+X+ahWcv3yz+W+DqrEEtaPCy1qByL1qG
zOjVNfcEu1bxoVsA4+2UhKFARcxWzCd3DlDHEDq7fQz1pDva0RkvxaM1OP4AD1DI/2nPRdlsuzaa
i1INQqfcAJHcXLdwzfYVfidvtR7bMJdQc6OuKuPhKD5CoVCepgnfS746e5lOuiXPqeKVJAnIDJ//
bboIKRut1gaiTjpKjhS9LS8+rr7QdG8rFtNpFpLbl8a3eHvDXZNFJf1xLwJ3E9oYDJdVbMoPU7XT
UiB6wzZaiqTA9PiALSck+yRJlmoEjmeMDcS6f8UiHcZophIFRwk8xaLlURIqCkOc3ll0NHoKQe6h
AIGxzeRQe04e6mJAamC8qYXCA+LRJQi38+zcCCTKd3VIcMdltLxNNSvFfPlq0uwruHElF4usinkT
x+fQbUAf2WXdSlirApEBsMVWaMXgbNJ6AEk2QUfMfm2tl/4KdFTVChuh4y/VkbCp9t1MTqQwfL5h
ZU/cMJgBNxI/qHUqAnmarPlXNyI9VSnNUiiCZv0XhZkbxKdFXdUaiR9jVEmS1eoK1735N6MLj7U1
x7QYFo/XBHajp2jbIGHXBGqHPfSwzPWR1Bt/lXcUZYjUptS8ycXC9Tof8BvkadFGpJoFNZAZBZoT
9PCHj0B8dksOkDmvZ03+oNo3l0r3f7reAQEA2NSIjvvmmIS99opQLKev82AJOHEi9DaVU8Ye1op1
YHLU1r+yjBDG/EcasFMWdd59kUWaubW4GdMyYnP362Fa/wBlbblUXhRAfE8iIL4t24DLxbi8OaA9
lD9gRtbBqVZnYDrIKgYdewdkjy48JMQb7ys7raTyLIjlo4tQDqRCLITy4njMOwckDHWJkzs1xJNw
Mnz1iVpRJv/bgvYzG9uiiAqaaKbhUh0Oo8PP3XrpSBJawGLsPVk4Gf4uLlOxigozCu90j9BbLhLh
NHD2DY3B6Qv1MPARQxhwfDzt2vwzDz8rKphD4kzw8KCJbFkDqaEIMCrd+a4NX4vNRqIlpKX7oZui
Atyk9yid2CrHMwFg7iOdEt/Nff30e3eaCeJFFFuIe9xwVN81PS+7ilAyJxcv655gOPVc6U0PalJG
8Okn1IN4rCMMxhLco1D7E5XtE38qe7+Nivcj6cEoIg87RVYzAijIohYcarZiB5BMiPz1f/Ig/YGz
fh3jkPnWz4I2QUrvF7yOMJbCAOufEXszXQozX1UCfMLuuxbWkpQ6qqwR38UBoSZ7YWGXGUt4j1Vu
rJ5gys81Aqq1ZYdmgJaZKQaOYTkA0h7Z7CSv3AEQJQPTgtMV1GAol8EKxQO7l8hueDyjGoB/7q68
AhicuEOS3rn4ZO/6JSfX7u5XZDQKslT83k/7I9sZKTb4auAcyyqbUX5q2TEcMbco9RNp3linHcpr
rehJ/7bEziaN6UI1F/AzAFYSWjebG7dI61Aa4BfQGxU+z3c13CXm1XvKbmJUw5LKIAFHYiaprNqi
XbEQ1Rn9kJv+Zweg2+Ecs+2ZnJdVS+g1vWvMNxFwRdxGA6VX7Vk21WjvuT+tu1uYcpHftScsyTfA
5u+mBOYIJAVft2+yeDU4jiYB6JjHs7PaB8qz3BCe/QnsfkPW7P4IuKKyv+0DsDWOB1RHwGIICsRj
eVeroFNNHa1v95vBa4QFzZNbonK1bYhzDAqMglh09kZxeoXkdNlF7OYVspiAJlT6X1YjZ9tSUFeg
8xPZAwnDUPiUBhaN+X6/2gcGIVTTXKCHRD+FQrfydgxwWDBWptS4gOAYpEsQ80Lj4936oS6K8ao9
vcbzNzAREqJFYrXJGDp6doo+4uCDPoMTtMZU+hqH4g0r2hQRyFV6/Mqqk4btkVp25OAAuzgMCD/k
4qcfSAEeJmGGGCKooTYHJ0HCIjfQW41L3gzGeIxR+kFav4jO0wA59IND836Fc4QLHAVZcvCdffYi
cckz8YLY3YwGd0Ab1MU/ka7GqLGzztWYkZJj98E3yP4Y7+w6cNOzjGyCHBa4U2U4igmKQjOaBMPp
0fEKqjU5XE5R4yqUPj3OMnlIZPCzqCCwda39KOV4jpUn/xUaimOG8d0jB0Pw7e2RNjWpxQaqPzAg
DR7zU1TwF6PlUeJuSYrkOZrXy4uIm8wMnfJx6h2HcJtFH+ufH2JM1dA7Pe5YT9JSEMt3ZVAt4yTv
CYQCPCosVcCEF5W5/28O+B6/c8MNeSrOUOf31YnWZHWAm2gA8+Ifj1Sa92kAVFzAj2XuXnvZTulp
0TUgPcKypnCkkYgV8o8otvMnRCx0hjlGXu9xNC8TgIw4Vs9WL48zA87H/a8RHKYJpHoWyKsSd2Vd
f5n5QMfl+PcXVcTmjY1HZgJHeQNiCtiGZ64b8GpPYjCBbI4R4gbEOWlJfUBlwGNrmZISOM11gZ85
v8HrPUlOlRcFZrueXHX2Fnn/8gPfvs4U9GjlBK8a/8eFs0nBcIQGbDoaz79LZGOMIM5O1al1aCOI
CcfyhC+72GLA9wvyoHAICDa0+7VL+4yT8lv/p7eq5l9/y3JvG2OXg7LdfskP2s9fp581x9L15mmj
msEXzVCpT2bEDnP/0Le9lfjkn+Xr8OX9xgJ+XNQzGsL4+tfVMqS6Vk9l9Lksfrl9ptWLJvJD6LQN
RZZbN7C0FYPLFpIrsxGlraVgjWCSI2dkJXaige9GBsM7p1agKbfJeUGVtUbvJ0axW7AlglkKNfiP
GYuthpCk/sClMM5ujU4LenxPwpCerOCMTkUxMuBsTsmmRZVqVms0NhkUuMQR+grHovb9p5qQtM+x
GNdOJ51pVx+naJ8SA+fV/wcrqV1mCoS14yqY5FyXBkV+y/6j+9wdruZ165AhDmaAT/XAvpQ7+Mem
/qiqdLbPAVHN3KZUpYbTbYeUc4f114KmMpg6rm7hs1nKZxQHohoCjqPEs4VPIsCKs/AwS5mMhP0x
xZz9Qjq4o6SKvdonEr3G2Swv+Cx7w5G9qcafdO3eCqaHCL7cQ7jprDNQ8r31KKznPRCXSCE1Xq8o
l4hjxOIMD6/8qJ6OfHSWpzPGp5ML58GhbUEOdEhJEwCX1rIlDusW1nTk9DtaPaw+X74dRCLYw9Rb
vB2R/ZgZibD27s88DdxlRmHnUpK8FiVfBX+R2znoJVEDNuNHNRIiw74d5i8AnkeV1Tf64hh/JRwM
pymKLp+j2cOTY4Fokt9J+glRVlYcOFKM9G0ncmuijbEEiQlZEdmzoA9NZ/hv1WCzzbpXy1hbMYsC
1udqn0Ox43w+NJ47CbggVwBsDfyqjB8f667ssMC9imdJ4AXeiQvydgsWz6zH5hnDSju4jlFejebk
XzK+4XZNeVCqXIe0zmpqi2lDm6IzE/voWlWqcEvK7yGyxWVTH8uByfbCuwvQ5kCC6xtJNT22ZdMT
TmU2zz/gPSx3wCTFAJJRaGr1/5ssB4YSJ4RICHe5kPBiJ05E4w4VfyubJ+HNTZKhT1/hepfBnVs7
NwZkvwv8hF5670kGvs0GOU9xP7WIY8StO6W06knGKLD35XsCfJbTL3DWOjacCqnT12dqSc29soOw
uNNhtmYRoNpN3C/yrBwKBiSmrw238YU2qw16gp7K+BIbdwk9eAWi9n+/xHYVx+9/KiZsU4Q2PI2T
R7OGWkgl5VDgO9PIWlPbBgNtLCgdC6NEB7+IHVx1DmyGsCdgI1XVNoLRJV7F+mGKL7FRqIRAzxFo
R22teT2/uEHRIxg/KrNWDwwCNRVmkQCUFZCGYb+vd00l/Wny0B4qWqsMDpAQHWnElOKKKbej32In
+hVdxhaz+xdcXXn/FlV03pqhKXHHiCvAhhOLR0olb27m31FVTFkT2k+cdKgrdOBge7Js5r3SUUfL
O3LqYAYZX4BsfOel4fEjfSKjLGZOC4afaYnEx/9KLu3l7CM61+cSIhcKRD3QAU2GtCrTDZW5wuv5
PO9RftizzyCrQoB61I/b/LNMRlHRLeXwWNLPq8YDeidA0f7JfK4W9n5xPWYFcB2fWzieJRaokeWo
UHhGHIpCGrDf9OCnFde7KLNXt3Eouex4QY+NCgt4LJ9iqSwxLucmuGQkmt4r9l8bGBHIIro1aiWL
dUl+gKstLZGL5C19ftw5Z5fTTF+EqNLQXKEw4Ul1DRe4gDwWXePOPa5rhmpscL76UjV54+NAagVn
DD8g2JSSLB/MFneTfhkL2arSwz7Wdqk1f7ohCFxu8fd0hzlLkCfV39COvognbsSs5dLQkVZcsRbl
JMWTBQBY3f1oEqzNBtL4pWwR/pmdTpqfEB9bZ/yUZDRs+AjEqkTo1Zduzwz9LChLLnS97Ecxc9ek
rc3FGXFnuCxbsrZsZZSii9kt5aKMjZUs4KFK0BOZgELvZcLCgnepUF3Inzb321RATH/ACLGK8bGl
WS9p+qx523+M7dyb/NoOXyPwhcgU9Nn3pLiQWsqJD6hMSn+wp2De1DjndgejlCEVhwhgiL/1awok
sh0RsY4th/OQzlf6mGAcAXL7aWSsduc9e6DcHDtBaLMfZdd85he3K4Z8ElxoPhpgE10XbvUFB87p
Sn2ONnmS0Uvhj52iKeD0W9xxyfmSlS2HoKwKsiSl1b6j+zCizfyp2QRQr7az7hZRgHc4/8fWvatY
3hBmtlAqjDat1xQbazCa7X4likamYBa+ihBs7B3MfWjJb9YmWW2jokQ7yA1yTTZxU8/dG+M4eFXr
4Kgon6iyN/6dYMWSqv1hyjcpVkmoqEmdwmJVwQAqIVd27eyP+6cfoYJoUWR4E2MczC6yvdccTL6C
xWyBIqS5PQemsb4tRZWZrAROi7sJLc+zuWHNR4oSxUxJNO6bgsbnuPM6SExQ9uBtS++BIXLeNr/s
8AcRVN8gEA4SBweCnWWDGjnSVCKobvyjPmK6ymVkcN9BI77eKHj9PRYa5VQBexsKyOTEEMQDgokh
fXnKN/3cEf9O7hnhTuKkmU9cbctXZeudOafs0765vEk+nmPEPFvtVC38E1W3gONu2no+Kj1RO3fr
vXhpW3tyqji8X7Ch4xSKkUoHBTRgS6tH0gstcmHh3HddHowZcLUwHd3FNq84drQjUYPZz4grPk5j
WLaXjwvVo0/qIWNgzC4bt9zaB2R9HmE/QHZbsRI8plYnEXogDdktBp36NJ6yDZA22KcDLaO/OKjE
NRi9B6mv7qjuoK58WQFEr6DKQrBXOTFtfkmqW2/xAFYIucPklGBd5Pcpussi7GhfRq8QAxAq41p2
tqdURVEDr9tsTAUbSadH5e7/BVHrigM4l3A3LWYjenyby2l0heZKmpJ+IYqScnkblgtMUqMDIB4c
pP4UPwq87UPGmiN0DdAt+Ui69pTjxXfXegY9k4/+e+Ix+btjBPrQfYIawI65mkN6Fh/UwnXbcp0g
UIBGyRgQ+pBGA0/MKTw8dnw/k0extDh9A7TC5DIbNjquarFu4CMLQUk87jb20/0EXQNr7lhTFdy/
7VP9Qzt26TdBib7UwYwkubahWgbadZ4uxNprGXrFlu3ppVNYYlXdrjHF+SepSgYQLDD6MlKlGs/O
MYGrRUZiH8zyAsAJB68uAo4KVsOKZbqBLdueufflEnRy/0eiiisrm0Gn4jZPrgAPe/UhthuvI3F/
lTJQj1LeW13eEr6zExkG9WJPsdCQMpWxLGWcKM1KV5RIpexqpQj+05VNZpZZcKkECPmAzLsCGOmF
m3clNPnijIJuw/GIwWcpfx6SjRbw5lvhnqsgb9WwBzjOTBK2RESeENjviP2juLz1nsNS3f7OYZDc
z8JjcAPfWn3iYx/aACwAUQLU0uvADmmpDbSnFlNhg52lIKtuMtZi67y8Pa3xjUm6zkooagwdlHmt
pUoVczFBb8+suUzbAvMQZnxXGnu6+mGYiMLkRpG0jkm+tXTz72H8FcSRCW9nDnb2yAD7Wgeue/1L
EIS4ODhVtRxcq/2NZvuP5gni+mLJaNDghcZ0XVnmGMbAkM5Cfzhl0dLkgFtqfdlu0M2ASO7yra/q
kQ2/M2gHvz3qy3wY8156K+V9WgMtA47PG3H8K9RXZ37qao1aZ0PTxYEfw0dmiURnmdgoFe//FfpV
ocDCpCGaf12PaLf/+zdfZYcure2djBb2oJ6FcQtrqgHHvcyVgi4SnqnQUmjglOSbcFMgzoZ49H5Q
QEhp8rPSCQ68HsX1Z5GmOcxyA8yFbJVjJbHRgAeMIPaTQFwpGIQa4hGJ9yYWYFK4YLRtgr8+go9x
/J+FSZ8/QPPyxzKlI4RK2f6zNLUiLdWtkYiJ1JH7Zjj9feZhnku+Zb7P9E5UCGakgZ6fF1L22FOb
2GN8wP2MEm43Orc8mHfjt2+w7Bmwwxoo6gZnaANfFPF8GgfndGLDaZEGlbX/wzO95/slMMft57vR
mxB83wL9c6WyELwR3NX8YRXoGocVE41tEng0dsr6LsM3K+sjb0AmYpiD+yUHwzsv9CWbpJRf2Tov
u37/dG1vXh4+kwQCluptHhsxjNTWAxvyHZW2wq4TA1PpG6oFYEqpe4o96aKOEfLd4m72qzplhZLn
G3PiNDjkpst0I2MV0wUoQWdh+LW9+kh7NfVLuV0jP6JsrnK1YQEIRReUDzDtQyroNDFLIcmQDr8q
EyXZUmjYY/JtNuZw1hXWIYDj9wanPviV9nTGtumNYIWLGHnHPaiMwF4hJ1HXsuAIeEVHJsP+m116
CzrUhBjMssuhaD9kWYSYY+txUtISjDKNbpbVjfihbushjIAF1y63WH53X2hDqFAZiYbddQhxBWHS
Dt3HDYU+h59fAvT21ONCJLfXYTBSkjvWTnBhyP6A77xtWqcGv60NggkqmIOttMGu+s6KS2+vY1F5
iFYdQyqHxE5guO+21mrWKfZ4dVw1HoEMUZ8SEP1S5zbmjXWVELSkJjsG6NzwuwrgYqzsG2IY454M
0DHlJtbnBaHsDa6sAMMy1SAMCWWGOFat1R6nVzXqECgxWoSp0NOQL26YyLXlTnOzbBKRasf4xvp2
5PYDZ57vBzqdWhJ5EqK2dP0RaptlZ3EdMGbZwJJMgxhdBMsyCS2NyJG+SzS7Xg2chMnyhQDnfrbz
m7G5po4gSvNGlbTzE1H2kvykJBxDYVQReWv3Gq7x7/1ABuWMLf8WCDUro7J2tGPvQ1tLZ3yXXpg8
xF+Gr1PpUUFtR/6agAo2MzlECb+jIfTN+9k8CM9ip2JrT8VFaw6wwS7R+DpmcgP5/bOmYdTiaSEi
hYcwCfDZwXwy6FVf1XEf3GB7E6Plu/mE3YMa87ARWOJGhUMSCYitiqbAfhkjT/055hTehgMM+QR9
BL7q1mhnGDD1JAPXosXTt+VWRbPW6TU+l5fthjEWqueFleZKQKIZVfVJc/FHRzmXrHkIOZcDrJJ2
hNxLdsFTQ5QJg1VVpmwgeDDCpVKclSEniekX7yuq+dE1XkMeRqsLNj6bJ/8Xee9IE2RQtGwcoa89
7RsejyRtbTREKJzbK0VIwSgLw8YEtZvhH/3jMlv2OY/SdtaIrWqhr8ViPBk8gtLroalM31EuMZdK
sVwvdyTicWWJ9ayeUAe5HnOSkyi3dOfqMcOm6bHxg2UgKscOmFvVYLiRErZ2q+JTOhVFOFgoJ111
s8Y8Z4JfH1mNL+fcDUmirwQYR76esXmGMBfF9l167tJG1lWd4CAd77Ve/L+2fa3DLpQQvMoUdxQO
94XS/F4FTcnDOEFXG65NKpCfwtxNSfXefgI+MvoAx+iSgosKy7hkQrZFOxZqali80kgFhOhR7htl
IZuhPQC0kYZfLhO+PWIfHz4aabWOQQxZBseT7iSYxfKkj0SzLKxdKjcfb/DUusqRcCjtcbSGJDBy
/8rd19ixZHHH5CBCwAOQyH7J75ZqccBqbztVwHqERVE9Te9Vx4UCQeBSZigDOcF4QrMOEfmb2YX6
gpaw1seKfK0pz9aK8ADf0m7f36Wx2DM2/R/bM/25Q17rCtvbga/sAA4tNX/AAbIxwQxJbJHRVyl3
0UUB68fsHcO26pgfYcuOlD65u0hnWxE+Lytyhey+qKjJMh52VfJxAFuQXaYf7kDeL1kzJKeCOy4z
Vmz1PGeAJLemP/iCvh6vaOfWvzDfeq9ZB5k+/5/nNuBfvsaqKi+T1MF3HtlYU1dA7wbApamw4k83
8387cDqJpPJp/5EohB6bMgQr4gPt8ivxyFgv8mxhIaDJohn3YqxDJyY6iR9mfRTQjvLni1mv66WK
enLWPSJxLSsyoZ2iRSItmd0Ic44KFPVpwfzI4LELgeWQOCi4QD8EZhoO4MtoWJXW6ExE6zPSJ0qk
+vd7wTYFwbKl+U3PkV1rS0hkP4wkra/2/4QS+LxeLLoiU1HItx6IO7gf9FdtmlIfCS+/MRU+amas
+NJ16LOu5lqKAd5WxNJY1s7iIbWBfL0zns12TdDy/i/Yp/nT2qI8fa2zyRaVldtS5DrK2Rac4TwX
2q8ADYKwITAsWt9IR+220euQtdtVc5MPSSAHmmTnh+rhXvn6mV/3kgTpW0l6QS84xj598l47S+Ed
6lC3tKk8No96bhj843eVz5/Yt3UBHwhex+z0lkNSz7X3tSfK5Czcfsf6l94A0Wt/SH623fWqzuap
/abky3Phr0lnFz/jVAF32++kFKGkCRwd07nrEu6My1TBRxEMPCk1ZJfNUwW42LDBagJvJHi+ZpK5
KRsA2eJIY/Vop+l1wPYnO1ComCGRVejLgDx16AZ6HN5XGyUNCvIypQvUr1ssQDOZ3geV7TfXNnJ2
PanHsiq9DzvjXPus46zpHTJTfYs3HSyQW3UgcudnA/lCh2RHbjE79xlQvrL3kInEWymkhRrdU5kI
uZIOBn4Z/gV4D+XJLg7j95ZPMJylMmTNTWaDXqSwX4EE3mjgRpD4NzEtQKpdv8NB6Q+hvME35pIb
BfecsJEAqxf9S2/SgdTCvIeo275cGOZHo+jaeArrZYJJGatedcxNwHS+/R/tcVDxW1Y2uCbiOioU
+KqVjQGb4HIBRr65n1ZVsJikbObG00JWY2xssKR73rolXCatuS2hbhxAOo64Pzu1tTfMVacSzgt0
zgkBNF/2JfjN1ZLSBQoolSGvLA/nv5mn6Lkz76rEqKhwwMzrif9RKziV8hD9HQMfl0A6HrwgIyW2
MsD03YkrgYCbyf+GngOWBojNPVpn2UtNQmrx/tpKAE9wRkd/Hg220uwXBNfOCfYBUW3Fxzn2SAx7
frNwHEFBwfyX0GjoT2H6qfZkeU7QwNyg/PxiycJUHwRG40W1MkmLBD+3XZt2at47UFRBBk8iS3cJ
1nchItjPxtDmIMymWgDZ93iqEPKiuiHEbxiCPbW6oZlbxXLdJYqAGHW2P+JvjY4qbWPyL7IvNGl2
fQZ44YTy3w6FclkzVThkRswdGWHv1wBtI2H5Bibf/E0ovsyUstNKu6a4i6Q6KcI1kIDPZnf0zjx+
s+rvPanohzMIBOxBqe8dEB10Kv1yenZONLDWnHb9EsVvBzjv3DZrXwxCd3/zT/R4VDTtccUIAvPP
Ssw+22tBrf1X1aVZCDb2FmTYDU8kuBkbCKSvNwgOwYHl3yJOWe1HZvxQp/+pyrnsSWXF526K4TQc
260UPWOlxpAZlbRM7KzkSBMNCY4PlVrjYugSW5vNzDrGHK7Sdom362/0kghrjs6nMMeHf3Dn5fdP
c08hvnCXqqQCXN2pFbWvu2kM0HrWBg0DQo0OgAlf/UQ9uFk4YRzvVDcs1JlYawcato9VrHeZiyRU
oY/woO8LpbG8hZX3FUl/ZH4fsvavyi3sfGn1BSdqhS8QlucNWlOyZiVTM81ubtur9l3SBFl5xrTN
/y2AmFth5f/UPUKAk6OLBkZV3NapET6na/LC90g+Su1mrI8BKBLATI5GtTiwidY6/zr1M69DC5e/
tZ2pBAx/tHEFzlPFE7WQQ2607DEyvITM+VMNIKq7awvjuwTuVCLzkjU3x3tja4AuD7i1Ap0e0EkE
1rpN4R0QUs65AnpFKEPX4vJRNlxGIQj+08G6M7b8SJpuquM2yUMwC2Uc2ipHoIoIrmScbYvmQmPP
bFR4CpULuqFqT9nIn9g6aSk+Sc1aIbGLg8YDtd3gZj7VneWZR4q2s0qo0ccMp100bd5jo5Qx+HSc
4rS51Oya/SAO4sL+KW4kfqcvomz6l019qcJHocAyLwaV73LcXs+lGxtTK62PaK3t6HmEj2T4Z7kJ
QPIhVIuUJ1AhIQcUnSn+fJ6vgZs9RFjJJeZt008Q5vpFwXEEXdYZHpyw9Dpa6M/KEo7KPn+/MRqs
6c/V8FR4rDkegbHRYcud8G6pHN31ik3tLZd6BQ8+HjEMmtBWCaWVU57y9lUnPZw3U8zHNV0NFKxx
B1etFoQWMvQeIO/BkbSP+/qzpH/dEbBackIf2e/YM2MHQZ9Hh0iIGEP5yDPgiPOM5zgtJ5iEE7Sa
fb4rF3Pby82u7VrUc45RypudFwHllFnym4oBDMYT+bA5jGsiYSx8AG7ghH7Z+K5bwx6JDfv5tTYI
eb3eBP7ALSh3WmlT6fsY8nJfKCkILayJQNEjaPEWm0EXppmGR0OHiLmaSbksFb8PolfJnPRkfMag
Kaq6YqMx7r6M4JXP6dS4bQ4FMnnILeDh3w/CyT0WlHMNTMJH5KPJXV46DSV/ovXS0fW3vQFV0anH
WFuD6wD3zoae4eLihKBNEJtndBoNhYMX5T+//Zglsn/96KI29hatoZfFCToAzTrEFgxsl96LQFgU
9JDwXVaR2cjVIHyxzy9BU6bZSXan4+Czh8497Q9Jf+H4IcDWIDGpoHu+sDHfC+q4UdkaJfzqwYtJ
TJf8zSJoUjCEpY9EVetpGLtXq+ADGXqLIwSdKef89DdYVxFWpjs4nUGZWU8hOFPVQuBYF1R2tcDr
GffEC4cvBLPhhNjFmAEyQ6lV3dX9tumXDmbnPCLP80PTAX+MTsnNbsApzchx/XTdSSGUpL3LKxsy
cKwAMHLb48wgUXZL94rH7WxHzYlAs5Dy7JwDaX7gkMKH2t4jnA8MUyPNnWDXsVXgnXumTgADQLiK
4HtoiBqnFtZdligQd1ZLjrXUclj3tWnwewNIMt8iHk+st0SWrMp0s0SGFu4XbBUpIQw6ouW7aq98
VQke/so4vzuYWAiXX4XIHhRc2Lk5c2AmprrZnj2s/6b4dlTc7NgvIN/8PfT5myZzQ5yRjTaSJJiZ
pEVqaf9huTJ1CNe3RH3M6g1vIfMfIUXkeph/REgB9vQTYIBEakJ1zNs54bl8BAzYTB560U+X4L5E
jg8Ie394BLor9+LVQwpUvi7dsUbSuJf2WXZOABenVM95YFRbKhcROzHNXICDEe/htv5KAyCyw95A
Ywv3pqTCFyPJ5IUbVf0tQQ4QxV9EFHImPL90J7RkFJyyvqIMtMUCmRfEGmV0cxZT51s1sdO5m+rn
VOrQ41rqkdbnAaw28u7NSrgbdl2XxTZDVBiJ944xf1eTdzOdJaIxl3z8DNejwjP0eL2UF61Cr6DR
bUbqIS60mEc+jHOX6XsW6dsonwx9C1iozuJIzOrHtQHw33JV45Dfo/5B7eK2efVAQqJFbb5qa8BB
0YVK5UWzR08RTlefhIYZBuKaOoUGml3yhgot652PUnb+Yn8Q5vZKN7NbAbv61bc4yNp4Lf4q1R6T
1NhYqi9y5+1rrSetFvRSA+fo4eBehNjwGfbRqLLcr3ZymC6V/QBVSHKnQRXROv6no/0U9IWMzYBP
3iIPiOiIAH3CLYhJD7SRMSKn+4/ae8O/KevJFw6sYIy5zXdECepGhbdw8aVAU48DORCDz/G7ZukG
ea1smiQ9s1haDhoLM0/4Rlmc8b1DquephKolADDzCRXR4k3/5y3or/ODQuB0OYqIl5VWCrpEMIF6
2C1VvJtLN+n5b7RoynwPzyfu2iC7j8A3jz+w7oLwYzUF2mU/wXt4vbdGHiSrpFA3cIFVvLKQcyDF
D5mL9tojM/L+MVIervqq/nkij5ZRDOVL2700toMleigyrJ8Bbrn4n4yxjSg1JPdj9l3PnAHR9Ze1
eNpppQfTORR9g8z/Jxo+kTvgW71GvU0YztRSfFWko3xijEQOi2fKTJ/AfHNsHF42mxVKx9enFRZh
4D6+xnDgxQImQegVfEmzaKb/rP3n3PoRhgiM8NLrU0fZeMOfqkXdkyVw4ShTefCs1hQ+b7Cw7/Wl
zeeEAol+dw/07TpiE1tyX6GuoHKT086TDxbURr5y/rRX8OelGJz1qFANL0805dbb/myP7GMLWWo+
RNsBkS7ZDjFoEfRJBUsW9HgbYqlSqkQftJcfm3bpPfE+poTLweSpOPIe7clcw33DsDeAEasrOtBT
4cPaN8e0kpZIZ+naZyOurfIsUk/G+16/Nw6djNou6yB7ptbdw1eDyaoBcu10OM9rUl/eBkj/TRIJ
TMwMLtkDRae66hm2fe7p2fvZ/hC66Xv6DXDHnv2qjHkJQA51wFX5b5SNesdQgnbSUqnhp3rxoFPF
792zqrTL8AUSBiQYlkYgB5a+FNiToHuX3eOZQ/BAHVHY2AmnUuM2uEwmB+B0Y3bmHneDXy6zTTmx
1R9cmAXKLY2xcsIc1EhCCn7YSb9bfvV+SLwoaXNcAD2M1kSMDYroth567o6yocSJM1nBVaR1HLMz
4hiNRYSsFDKiih7yHqQcaEMYyPv6ZdzjCy/NOoyvSz/pjQf5pQ+TS7bQ2B8fx3DNo/FMSc9UJO9k
Un53ImeLHszVl4JQ0JRurw0ycyxxPGTaQ+emRGaCqEH+WnVjQzOq6HFsMXv8tp9IjHfQ/j5ZAYRw
jC2oay64xEdYgrrHNmOykkjMATuHx+MGgLKHEk/iimKKM1J0xPjN8jXYUx3B9AetP9JLUpz+pq0L
r1vLiym1Y53jYKNOzB55vV5Xg9UgT0qLT01x4o92J1A8TwpkDYd9LA0pT8h0vuBNZp+bLLDMZuyq
/9I0r5wQCy8EGMDwAvb2tx1q0xqKt1hF8UEWcMXPsEGUFhdNd9peNsHwQwbO1cYusUHjKVgMX5et
OU87IX3XfcvunB5lXWSDC9CjkOHQVeb8zVmNcfjy8IX45+C+GWuNNpkgiEtY/4w2K051xi+xMqQa
YlzNd1quvnXvynLJOdyq6jy7/H2JZ7u4weqK1nzLeBG/2uOaJY2f1u7FIGmWC8rZ4fpieL2TIHeB
p5wLuuL7TrjBnXPRUDTX5np0givHsMICGexRIZ7EXHWJtnq+RjhE+6xdNHGgglzaGUvqSkiHL4ib
6f5s8hhvvaHRHZf1nRc086bmVro+opw2CCtfI8s4lzC4Wgwnu6JakQ5voT/lP+fE5x+NipFErD39
x8U1ZUd8+rSuMyT+FOawHKch7MJ7QwdOZeRbFkuthQXELe4TStzs4z0pr+E/CcgSIO23OnNrFRZx
T8unpDVme0X8Xp9Y81XqO5WOYBlVdBNY+eWpGfC4O3PPArp8aWT7oVSnoNrA/BnaP7BZlVH5d18M
h+f9aRrhwAouzzzUsELbkHGSSf9JqQKTBVfuDeo5AAYLU5wxQjwP6rAfcdzZ+6NT5Thf+FuQVBdW
k1LY2FCgj3dBXF4EtqTBu3ZP5MuMEBkKGrAGKVQvct6KMUojpQCaSpW73fJAVNM+Cs2E4gzPXcyF
OfqF09XeqACoka4U176jwPn5IUiijUWW80ZKUjl7IPdsDjkmGzPFVtG3TY5ghcB65RGz1SB/RhNs
ipadw42QlkdoMyRreXH3vaeQ4EsIG+Y34OPFw309DlFk1HpFLL2hV+YjRLLdq+wYTAYZgTCFXyXY
32+EP4LYAcTfGlYPSHOzryGKnw+ItoaQa/JuqK04AFlZv1djQcT3gVSjQBRQ2t31gbjsljFfllwJ
R5PAd1oQ8hpBs6i9uX7D0+a0mqOandx/7cSUqM/SR53oCWkpDESBfPmSlCAfAOS2fmlu97k6HtQF
AoO+DqhV4iOykQcmFbrggudq3Z8+oJGJYPpe227ROGW/kpJL2l1v81r38S09pX9JV40mZ1mSkOpQ
jM8Dg129f+V2skwRNaSwg09KJx2OYHhhgOHjhR4Gu10KPocih/Bra4vLiwnPWSLRoLA5HqhHZpts
BMUX8geS0B7Rg5LCi6urLIvjGrhjeJwopg8YH7DY5hAjJDJGXitcPu68xOhFXeDwZrXU0O0ce8GJ
voyFnCY/CnLehOuUxdLB7PLh9zBu6dTchvAffqnsYkHcuBbd1sdnJH33jM/iJ2AOEqNACmDPMmRW
BSWfMZsWQny65HmmD6cq/G2H2Q2WRobt3ynDxaYMZDmV3dl2JtKYSvXSs0JAHv1low1DZVtgzZOs
G5lX/ox280CN1ms7H+5+TLBR4fvMQbTBOOv2z06cNmAZn3gQ9m4DezwkiVnulE+3sarlBWZGb2o5
BnuEhM4HF4mhW8CB7iXoHab5XO9PBOjrcfia5p8RmmvdmmXgs/cdNBUGitt6senxDG9kmh7pkWrn
wrSUqrePq2gvbXEdZyN5hsrrkxlziNr/mtxsg9+Kwks5JjuRATe8fE3I1S8iddOtFHaaCpPmu9tE
DF1vO1AQAq1EQDi5QZZ/ij2LJISKsyu8wCm/3Jwvl52VWbp//uTyUizC2JuKiC4mMqZ1yMxfel8x
i1bgMJKjA+bvGgsIDPI+8chm4pW6mqy9xCmILfcEW5zRmifrC497DB85US53UptpcN0xhMYt6pVV
CzD84ACTisLYlpcplG3fkccQ1rt6l/paDzW+cWkuMj1YaJjRtXoDeC38PiJ86B0BcQ15mS/XUYxy
A8acAxs3TMraMCO5PcjN5J3RmCVy9WNT5kJBAgDknBkhIkg82Xdj33cwUjsoLXYYhFUCFMznUp67
t5Rm+19pebyLlBQi2rHxDGUlawaWL3us6m6Z7XJtPNQmiCvpdtvVSC2pQ14nXfM0UYbN+LnY5VEw
5drMyUmf0tulLkUb+VuawqpGuyIF/kEIJmY1Phj7Qx3itBiP9T9LuC/7sKydUbtwZ1bvvP+0SPAf
V0yPMKI1VM9hN6UvPkhVRCSK70LJnhIT2wf0RlXBIKtS+xqntue/rUfhMCtdDxsvhC1f2nXhNj2m
XmqLIjOYWqsb0fRB8p7bPJROs4dVVVjCoWXIXsZp2G05Sw3zx18dVl+c692+9/VSljtiOe0RdBnS
gHFT8nF1nop/xBo1xNwK9DJdSJYJtJCp4c2M9BOqRQ/wdqyMHCJ3ENL2+cwwyOKQJ9rroxJDzu02
ktGYEPHKFUV6JhWAdYXXtOfTykEKGHGM8IoQ2gcEXTxg196Uv87Cr+9HcDt/He6XwRmv/6NO+XOu
0+CxYUM/l57wgyBlUXWIoDhGkHLWyTrd0+579PdVCzXHThzGaAqyCCF8mliMlAgMA6cSf5z3xsXW
BuxVd8Z4s+kmZNVoQdvTBVMdmPPGZeA+W1t6ESG/Ti/ZlEwznKGQs8c5iExUayOtQxKea/Xfo8mz
n7/mEKeA/Y93rjXqvhTl7MsvUhvkL+2ZRcsgZFK2vgFPSjcTjCyrv998IpE4Ip3LL6MfLJpf1GBO
zIG966jIy0vc4eQWD+lOv16KXtRGjSqv4DSVw6Rm+a/6fPr/sSY2LhEMXdMG/DqZUMpbtnxIVwsA
Ar9xJQuMVY+yM8IbRH+DSSKY4ww+SbPbng/caJmHrYVvNJCJcuURjKUKS+KkLj55hlPuVKCAPo2+
YoWz6lYCipgfHC8hXmlBtM52o5lDrsX9LAyxZwFCt8unOMPbLvyRRHylwXJZ6lqeKN9LEZjBhJn2
bxtD73f7FYo/yBEl7Dm9DWtkg/tpN8FG8V404QOQzM5lVIdVxaQKlLzKf5SzRL9xZ2xDQ8dsBLiR
3OxAA0UZcw7KAUMWE2ZcW4zj4fsSm8gEwxc4os9se7YKatNqfZDC2TUkzOzyENuhVBNggW7IDqxN
eEiSvSwRfQn0737zOkDc7HRf7jpZGe0JtA/h5SsQi3s0INmIsSoOZeimf4/5vY0UZND2iEHzF5LI
bjBTC5ZniWbK7Vcbvg/Ky9XjHfea87uzKS88FneUFl+Hm2XyvUPJqf24652AvsQFCwkNODjR27mL
KaKKKF+AkFBd816PCwQ3jjAL43mm6OUy9pSS+UMKxZVjWCbHSd0GGb7yldnvCTflO8XLdnKv+cnW
94BnsSMTgXs6URw9Jq574pvRf6hAqOUXssQkKOcnJD9+agq+/rerXdQRZK8GnCBxIYxwvUQHGrS9
bnyxb7wDkiCXAEcnnsJQlOTzuwj7mtKpV/NClsFTm8hyxXaHx8lfbldbBkWWPBzGyxcOY3WnM+J6
8Q4kEWbcu+YK4u73SJ9MkfHX3w5JDVPf8mJfFIyjruyHHJdV1cnpKYPrjdTzmj4+1lJJ4DIQ/ZOB
tL3bscak3CXDoz4gJFS+Nmb18+wmytjewDSyZO3+Tt1DWX0KWwCLCe9vZH/atMjxag++d5haNSv6
xq93q43dEK9P7DFllbpUZJ8BWirHsTQzpNJnDzeSvPhmH3eteHaatPdc02SpTfy8mxGt46axiIzZ
ID2HwXilwFm7AYWECtguUEtDRrr8VpsRQ3RyJXyYp52G3QWU5liDFDMFvCGs77k5yugB4+cW1mL0
vr+9t3owSYbMxjtBZRJtI9XT/1dYZ6rZ9xcSrsh4S5DtncB+1Rz8+qv+P2Q1/r/0QQYorO6LPSRQ
c82XpOpN4n2ED2js9uMXXd4FkwngNvf61392XC6qkKDJaec9F0Gkv9hyA6rYZLiZEVgBdbf8/Qc9
5QyGaLzaB4StpzvflTpvSKeRxmtfZcVoN71K6SLco8kokWlWWtly5T3Pj75YniG6vCDtUk2ikDzF
+oCoOhIdBCeqnGOUFhCDXQnf7imrULG6YYwo1DtOpUPlkDjlfQW5bLQran3GWhAuMPcKnFRDSTIk
SViZobHSc73GmXLyh/LEdpbMhW5RTZO5MYD14CEzK6c3HTQLituBBt8TTS3cbbv7BE+2rM0O85BQ
0HBQTIAmkBe29BJ9opq4WV/TlM2yLmz9qN6Oj5ZWgEiwO7r73gUlUaiD1tdThD72DZH25p9XopeO
F/lVs87lHpG47FUGS9drRHBPNDOiBTmpkban4oGGEDbCaO3ZAYWz8Ie1dm7qavL/e2vWNVQDTMy6
si/eC0rMaKMaSn2KkfKP8ao9HVBKq2mHCaPjrkkU6Xh+BOFupQ4V+ID1GsVOvKmvho7FxRRgH7Of
sbc2Ttfzl39w4k1dL7y13PXBWcD0eFXr6IOneliTmEhYVzo/ZK3Swxrht7bwIp1T15f+DQYUV1o7
QCs6PToLr0gAUs2Qm0OhANzm/opgnoNsuSBwKYl+oyTaZojbpSwT5WsezxVfhYGlteRFYWWSHGNK
RsHBFEfc/2oSkw/reV345/fQpH1ACS4eg+ri1xHdq+/rBafm6yI1hO5OXdPbqkxqbsIJaKdzjcoV
rpS4wVk10EBQ761x5Hb4BunuTL7gGOOiZqqXJNk6s7gS9aZRdY1V4Q8pfi2iBgXg591XqOIbwnym
Ygw6Pj3R/arH/0P8EUe9vwwc4MQg5SE6dl7bueTzfj9Sq2uBCpnOJhyCzL7YavfsQNYZSlzFEXSt
e40FsyzwFluW0lJUokXcFpTD+4Wmu4aQQXGLvFy8caJQJUz6gR6LyK0N7QqbxnrJGxN41a1uaNED
zaYukjerEuIY2qqg0SMPm+iWvZpEmzI+5MUqOUkRE6glvP4eDUM4reWGA/hzRJnJgv4KkSZfmgAi
b8Fi2rgmC8CrfwZH9HA1yTyE6lOGHJ3jaqS2J9LIuVZSC0xZ7nC86XScO9J3LfPKSym8w6Ac1JzJ
GvwucbZJ1Qjke4wcvMLE+WnahzZgY6m7EzK+UsPnHWN/aOSvduMmN0UjT732VgdsPE9SHgNZAMdL
JYAsZmnkKqm09gEjQlE4x1eE69PsOnjURB5yMZEJfEyudoQBy/PuIH5FLWiO5wdOt1r08jLOu8ql
D7s3IZr41OQ2QmdDRjGUAHcO950jRLQIOqboz5+wbOqes49G7uzTmkpO8TkKH7xbdWFOH7Dn8iOR
rxF0/XCasNsLLhuBP7yZtcGWbKitaISeRHPgtnF4QT6e+RFml3dZ04soBvPbeROyf7drKVuUAFqj
JaXAet1fBrL1ZYEfnjAOkSH+h4mNysbezArqFn1XAe+IelQkSaf9ME4m28ocTwrF1g7z8Icv3+9Y
lRqCJNB6tLjkbIy33olXhuM8zTT8LXD/JK8LNLVHnezwepSr/VHKiRFVXBxWJCUSQpTRgjA2+C2M
fXFJqhaj/qDbXJgg/qEwh1At44UCcauOxUAuogsRtJyN1BvBW8BlP6x6kJhQvbuoJHdJIuTYyNRj
OKyEcEPEQq0FGTG0fXQZd9wm47j2hu2pcv4Ksn7SDNPiiBINt7yBlb+tgz//ypkG9aqS3I13sqOM
4CLjTzAKntAQYvyT4+Ts3mtAkk0lETBjkcibh0jWSYeetvw9I2V/DQwgVR9VtMGcViiZ/XhWyz0o
eHPW65ayyc1EsdDVLkznIDjpQYevhsRzXKc5C/kirVIwAmfBNxgQMTjN6dO9+wR9CGa9e+o5ywcl
/Wk9s2DmXvFtbHuo9fgCZBTJnj+gskWz+Qn2AmudyH0cp0n0KZvuQ0aamSqVyANmBjqS/BexlGsd
mek1tJtXhQrPKV1/DexUOIwuGPB/zOuyos8ISqS2uQvfKVUuhGsMfYlBik2yGkcpn2X/7zRP4AiP
+0hhwl+VLBOrm0H8qf3vSjgsQ6+bmKEdLwu9TY3aywZkpS+Qd7oM1oTmsxVngCsHDN7fNMEIMhDM
Zvq6jBXrI9dK7/NCnqOIcXpGNwtwFeouOFqubpQ1QIhIDPHvH59+3vQwR5/hAQdRmMgjXv4AnZ/d
gq78Up1QEU2sxEWMx1zWe15IWnUEtowwHhC4+cv6gPQfDD3UCenTyLQKViuMDFZX1JylNTWolIVw
YzmCa2GPQ6l11p8PipnO58aX1TWcFch8RxnhEA/BilKN/otll0TnQVKCgHbw38uPCvISebCdpF/b
PD5HyCMdh4plvRSviADsemWSiwvMnJs641vfx/1+PsV8Q1ES/Wrez0qtMMMwx2I9WyBUIlQWMhQi
FXGv5iDzXz1zrRZzwkQf6Pi430ZiZFrbK5s7DqN3VCk1WpX8ATdzFyDXmp9RJxG57OMgoZQfMRWT
785GfHpEuR/W4Q8O9O+ni5/tEbeALdWLIyKcpMbuHgBYGRdgr2i+e7ZZoMaOU8u7uUuvwrarIRxs
ImpRekaRLQdBCHafllNK/dQIKWHFb/h1pknbO6GCc91+yavWsT0uY6g/4R5e9iczBsMnAERuLhyj
hd+0QPi8Ej/CcML8rG8HxRftwPcLzC+kt8wCDsvkYlgiAFoAkCoue80siBWCIwuOJGnXSptlTa5u
MhKNMwMsw6SOmfbcpssf2i5LBMJUt4w/6eymjSOiXg+iIyCWl+J/BeVpulKOTglP+2nfA4w1DF0u
7/+UjzxoPthE23Z7kAOpPjQsvalYWm/QMqtSF4dffC9y9XEOW9x+EOo5KVOkN/Jdl28xrBt8cUHv
sgjxegtBHU2Anjf+qJ9x81zdZ5DPlQWDKxdjM7bveBhH7aRbUQaptyfyBLfLy45tzd5P1CKCE9dF
M74v9c8BfWvg6fVwzJFjDBfYlyZA4eZF70fS5yfFtc2bLgRH6tGwdLsvYJejyHUxnKpLXGuekRJa
er7VpSibg/KJ565ahlVpIMQiqNVnhg9+dspgeoU2WPgT/q/gl2be0ayj6H0qGzs7k9l7U6BR9mhA
8Floz/CgXhie8FE0w1LVC2jkPFR1Npf8CCqFW2v3fwKCOxOUk36mbfjymgWhH+jinKovWe8KUiAE
3ZYCsBFGDFZB9CtK7izlyY8RJ3z7CRhhgj3aDz/+Thdk5PZdzn3YMCYDAiDw5C/kMD0+EICxc0WN
UFAy7IEmSfeVK2nBPqjoDgpyYQzG2wpB8fDbJCWJ11gkfGce3+LZFTkyOZcavhIuSWceXq7xhkV3
HaEpXigeMCJPTCVcG7LcEGzi76DnVzw91fPJE7XrFNGXsll003tTyacBgF/TjKrOjjasmpsycU4D
zGAsB4oZQYqO0U5js6+KqcrhFUz9lSCXdtWXKcqomK/KSycLQFBWtma94ap2q/AJC/kwQobjr5Y8
msqAVR+5xZnGExoWrsw3tDskZXuCG21Ev0cY6/JLxqDKg9A4XF3L/5w50lQB8fUvzmdZE7YouRXn
TFdSo7/KoRWNjmU0/VC5kt/Shn1fJsWsg8/LOwMeww+JkFpijUFIY6mXr3cKo9QlLppjLJhW3pOb
mkqmpD6I4mXiJU/tQRCLBLVGe0mq5y+iwswU0uhdbO+w2o1X4SPK35zb3XMBm4nd2o45zGlqz/Rg
bY5PFZhlguwwfslkHhOQTaxqIYvFRfWpyL9EHbNNSiOoVSEWeLkwTUAwuEDLjck3zzCfMdomHDJV
8EONNUs+NSUsQHdJmVZdNJ/Isu4Mzxc3XRVXKgM4GDy2eRFwVPL7OJds6TzWAXTlnvoL6iyT0DWP
gYNxod08AsWsVTHKf28vmNXZiGPEODg+TjEHASxYjvEOFq7u/ypESDhhUsh0KtuPc/nc9AKs3/Pj
VCWCE9rOd4eRgGryyA6b/piB9/ocx+OI5P1IsCTDfYhiY0AINlXUkE7/1GXcMdN3hLoHe62AqLst
DTF1m0h9lC6Hen5ppZE+JLUokwQiZjaCrWSMBcackSJ26H8BMF8raANyikoZD8GTFjeaMVe1B8dM
bE5CjVSUj+BKpk/XnWEN5hNYjwZcPCh28pHmNiCbkuyvTAwJTz+EbIwdBML60G3IXuqP/4g8gcLK
7RmVkJ90BGE5+NpZeSfnztl9/I7B1hGLmUYKrUdkeAA1u9JcioLlED0wYNFrJKRVXeeTqbfphFsA
CftqVwhcKEzQTHiMYnda4B9PFkTqH2KXsG2g8G1qx1VGC6FNzl79hyPLvXya1c+Ks/YFc1mfz6NN
9O0pICN+MycYUhAYa/C9UM+0mDRng49Y2w3kUvsI9nidcupsX9E0K6/UnQDMWx3LzzSgHJ9sFJN1
TR1PA7jQxKVedwpIgpNi0OUvT4kuaAi9hnsFB4tU9PtxUK6vg/Pp/I/3dTDGcQ+tqQZ3UI+IT9dg
vUGhrpg6BerEj7Vn9RwlYj2zgbNhjoRtRY1GbryWeAKG4fOxjfHn+5wK4tjj7Du6hsmWYSRVUPWq
7p1QxYsULImY6fm9POhQY6rGeTXzg9bVVBB2wo1CHZc8eAUzHmBqvWH+VyVOUd/mZhbuEo/7PF00
M+wBz7Rf6CXDwxzS8xI8Qn8Q6ACl+qitV/bJhCThBdtwIebLtS4kUVSx3Obr5MMdzHJ1aPLPrV5N
T0onKyVvt4nJ7c4ZGB0I8ma5r5xVFWB3N+De6a2jBBy0BDgc6W3fH9lSBXyheqTK8kbElvtcp4aY
s42wzJ48wmB+xOrg0tz2USaNqvBVikGRq02SDVOF624rTZhZEhhF2CHJyccyC0nctQnxfGtTD73y
QZNCRJHaUOycVJFPeuQzdlyrQbCkpn65tDGrsRDZ1+9wrXMdD0AefLHWvH/dnOuhD2oAMpDfcJId
NF2ayb0qEvE/PHCNDlzD8D72FqDTdsT/kDk54HoeqdMsj6Waa/TN89TDOdaeO6rjrRMExqBQozQp
D38kQ2PCVeUMTmt2qEd1D9tXPj+dTlIkjYdUDYF508ZLgVs9bwHI0r8lrtfghqz2q+khfo9YFgyX
IRCXteczNZKw6HAlLAXCVw2AKicD3yz1aA7Lcz3IcEa7VE1kmH6BhXCyrvS/lXdJGwsnr5xnBreA
h0Ws3qOpuy0wZaRPWOhduATmlig0XWfLs64LurwF4XjZKOPf7p9bqI88w2crO0NRMfQmj8qlr0hR
KsuEyzrcfc9F6eq+1ZvGyZ7Q8QqniIUT2Ij3JqimEQVjDufQCG9FCXNQrR3LAcvN9ofQ8fzk+ysv
VEjto+3M6hTJMlqZC8IH4oCZ5z5g8xdqKsJhYCOlg0fzEcceXTy8HKhJPDgF37rUDjjOq2l6AvXU
DMO+KvT2x6I1/3cd+BEErKI1/NbMDyI5aelLEfx8tE4Yyha337Ql/IrpxMyF8kLe52JNCcxnBZe1
uirOri28g6Kdo2cGvKaOW4xtLXgSOu2qO8klX8axrXm0/ZVLS5XcIsA9XX6FZm7nzTs/QF6Diqjo
UkCem59nlFvrMCNs3mIBH2O58jF4nW02kUJURj9zZtOWjTYm1jV4jNCw4doWPoSBXbk8PI9AnJaP
OyndGfdMC6cp9eRsi8SnLhsxSJLAbiF83UANhaP7vF35IUlqvXgtqocHRSBefrMh8deQ4wAETnnz
ocsE2TNJwdRKsQtsEBv6CqHAZaclRlbSowayS0KysUAeFc3mFasT2pJTsLuPD8oKsne8LQZKAhjt
1FQANWHg7ERpE9Rxme8V6wn6F6rQUjXNfmfhdHlnLfGjPtdlqp6rb/KO6fmLQxccwPu8Yg9peymZ
Ls9wiYYspI1bELL0Z7ac4uYi212XGrpNKqQj9SI3ZoU/rt1guy8yrNlvcevYA/nhB9VxBrkrS47a
hg2o6EC4IvIKCyZszkulhOt5PkWPg4mkWwxuKl6Fad7LWMNRiXZAEaJ1fucRHYzQCTWrBwgKPjMy
hHJiRn6nNprvZ6IOtrxm0lWy5hJXT1nANIK1emu+aetbTfjtEOIStfrjB69Q+022XWIrK5fyPWx/
rBN99agogiW2/aLl4KuXSndC0zsz4pgCIGYzMtyDD+z4ZhKNiqrPTc9o2qSP3MdNvPdrSWFimJla
ONx1bzx7TBegVRqtj5QPYKetn0r+0hD/GBm2jdL3b6ctK0xEeFxXFPTQPsWRFHEP8kITornRNHsW
7/nWjjpBwmiwxpuGL67XOtX2dsl5vhAXGtaAdvaNLGfNmHm/cv52MT0gxlGMwEMG4P/v5XHZp4Ed
YAKhXYzgn4a7+7byFpSyoWS3dCK5tLObd1qwiD4HaGJDNVd6SBENJMgmmRrDXtCXMCrHSjp3+QVN
9P+KW7Ncd8gAUdgYhTtk1Y3Gk1oZEOcHR2EoDS45L5JYqR6PlfAqHIdVRo9SR93lshF+fVANzi+A
C9bk+W19d3wG7HZhoMR4pbN1wWkGGDPEef3lEDXfpYh6/SycpB9rRHay5hEWhd3TNq47vr9VYOWE
46WZIQdc0s0FHqleDhp+S8UgB6r8hLXiAMuYubhIcFlhV2bJGJfoIuklvxI7n4erIt1jI+VKx7eo
r2FraFMMxPGk2Af+b5iOaYzAw0qgN8E8XpsqhMOfbLxYvbtQnO+UIepqL6TCzPbGXp9SP3x5zQHF
wvvDBgaQw833SeSz4Ks0XGBhjeezRLa3Cd3/eiNNtCz1SswJZDbrpfXPuUoz3oHcjjvJH4BoE+BZ
akW9/P1zEGS5JeCNM2Yz5+VNjJdwIuPaSIe3thv65teqxD6Cf29qimd56wgtzKQhaYZEPimmsMRK
RNoM/07+UxkmQfozhi5dcvoS/JVsPEO/92TBWqktsax4Up8szQDqMPMQznfZrev3RVCLrBYmksvE
u62OgZi/SwVo6vsoL7CfUx6y5iyBxvVtn7j4HEoB8qaafOKXGvpxeEdF2fjL2/frSohuCHumV2bf
jUAE2RYRotQwNQPkkqS+eB9JowG9nusc2CPjWfOHmVoBbY7P0KZAD+iV12CVqQtty0KbWIEOrRts
O5J62kV/H7a+6ocgdAhH1hHxR+QW/pL1YCHQUgfOVTC0I6wMhnMVZmWBHqKgiRZsCGuGlX6/z7+w
5A7woaEsNDZGI7cXAWQ6ho1jYuJ67lL90Ntea/ccxYRS1/3g1jPT3/DNcTRV/GoKi1MUqzohO6od
oO95ifRZzLND5APOe4pFJOfArZRygB2J7akXen5gi8pHXy0SIcPU+TkJWZ4Qdghv4lLyOoYU1W+5
xfQ3XDy8tFMElwH5J9OOQ+wa2VVFZ2elZrZ4uPhgNK7MWz000WcGEcVjkkGYZBcWxOkZhPrbhACB
lMlj+JCpb0kHeFS6OtJV53M8fhCRmIPKrRI5AxLFsBHCFfhZ48MY7JU/IySfMnUnuuXqf5AKQKJd
YuT/hrmP8auTAPGB3ENQyYrAo/BAAalZjn6oJKAuDo84xO2kbBhm/wPyoz2STiUhWPc2LExnZN58
oWxIgABHphyn0LOM4pMKIzuaPklBYdfLZJbVQDvVxfYaFIMT0kbaPyyxvFHEvVVzHbimaKuXEX5N
T+/30FHYwBxKhiUaYRsrBU50nTMVUkcQaHxvq7RxgvK471NNM1m3Io/KeiF6LFaODrfHtX+RUDDH
tvYDKy7szvsi2wDJrA72Fvm+Jw+iuc7/bZJoDa83eQmiCZseNFzvbKFD+KPj5vON1eLa1BUprNz8
G6Sd+SEtnde7ST7XOPa3tztL4+JFtoD/qkjLYJrHarT1bYcRsqam1OnBZ2RlN+ylQyOfd75C90IS
MNakEJYoyRexWziwYjGu3otYf3/t9SJp+JsEoif8t3WSxYtTmDakLhmd6MtsAiLBtoVRQkVU/e7l
EpNM80aYL6J+ydmXSY150nzU7Se43jSHvgIkvio/x2tzszlr7nuYDqgOhqmzR+dQqpfxRI3X+VFC
1iq3OxLwUYWIIY2s7Ft4y5fBcXwq/mg6nuXovtJ+6VZ8uGOYEtDf0AwTwayKc1LKfagqwjnge1hi
fybLThI9yk6WcqtXCENzBcyh3ydo8KLpE7KJaHyzIY3Cwh3HkiYEydIy52lXGcTA3eFy3T4U+ucT
zaRxsBiYFkbcRX5F060rQKvzoG/7DZIWxnw04A820j35Gj5zPl2sGJkkUGe6l74g3FqwtQn4PpFt
y1U64brx1vLtkWFETb5TCB8VOtIVquhyXIdPe7KmtLDbKzF3ui/lagONGTzr5vhvtSHXQ3YUzVUi
jWahUCDBNAMiD/iROsPMTriDdkmgafVPlRY6TnJsAYkxV3w23k5zckkgdsXO3oU76TWLOyDshVEu
gmZn55bby4qslYoZpBxhtyExlFJlb1Rrdb2nGJSZr32CuHW7MKWQ1soPkVGc+haTllJuPHokAL9w
/20qLu15zpLSqWw90nTXLuIIqqs5XQOOlSujjlqzN+6k8saFMM1lTpNpia+qeSqZ8x6dzybHqfv2
Yxslu+ncX+R8XyC2ALl2mykrDc3SeAH7XxmAzIHaoSCxg6QI5f5WVKSyh76qzhNMWUdpnthHXIBP
dcZxjgVn4LWeq2+LPNgJtT7bj0tVBP0tHLf3Ajthp/40LD6Z/cBSC8UHFwOzFy37OOOxVTFeRx8k
m12b+Ks85zRyGTYxaOH2tQ0Z0TdKUroS9dHCs1nwDdSwKQjBdbcwErwoaLHY64HRf9veBQdg8w+l
2ykEBu4L/IUtVUTKMErrjib8n3Z0XNK//nQag1eULtQE3YLXiKncjgELeDwBCK/ji80gh4SL10VB
28bknw7VTaqcIqrZ4bBW0C0ddmvQ7et8FTO1sJjJHUoxkUVnpa6Qt5sFbfB001kikCg9tZOSeuF3
/bflPbnLDU4UhGAabfLiLcvo09eq+zsCp1dNCjPO3j4farhyF2Jtnh6G2vL/GBlcrhkkeemWHrra
Utpudvrf/kcDi0JQymH+PyVbTV5RXKtGEeno5HuiZOP0gI8McDzxM6EZPI1Hkfmwwe1Y5R74QTCR
2amaCsv5TV3l6cC3LaQvUQJeafZUxru2f3Q/mlKGypdiz3lRN2+RETTuoyg8Crmc87PxdIn76aKm
WukXti35Cb9BK1KuUUFUrMSqMWzhciQ+yUzoK4OoBuMW71+aFWPuM52+BjTwx2N8of6v5Yc/T/KJ
uHNkbYCseKU9OgxNQWRCzqtD9vxZ9k5fli4M7s0eVfiDAMc+blOmuAXUUmvlU3Hlv6rHuciA6zol
CzTESs75hbtFvkAenNaPQSZyrrSha2b2mVygAf6GG0anKD9qjBFFukguq8nwh9n/xTKP6LG+jJ0X
1c74mNaIOeyPKV2ZMyhiUgnHOr3ycqG4u5qL2qRyRReSp+uTasonIBMsGZNnkZBlGM7PUPLBzBKW
CvA2478CHqWjlloaNbzML4sUwRCCjD6aR3+xMuWiPKglkj1oPa8J7SvIahKsGn+xZCNPpKd1yHp9
SkQE0iSbQhmm8q20CiviurUUoAxMMTLO4HLntpde+ZX9prLHBmzay58+YR6MAfYSu+zuGoClDMh6
OyjaiWFiwgeenHd7mp4UDDkvZTWB5iRQCVnR1jNpEQasyuaKgHGKbeSfrD+00ALdw2lxB0aeagsZ
7cMUAUYwAmqAL5v6hQUttSCk0iH+DbTcH0x3634W5Z3oRqy0qahE4X+SvxPe57x7rY3ThJXdoPuo
t4Yxrn9LiJlJ1q/wWD3SQ2aF32LwNjSnK21pf4Nyha37o1cAKoWG3pZ6eonTP/MxhpK0NQWigy6P
0078im2Nd01HiF6LYxFlyjH+cvCnfFw1P9YxYGyql/MFwExm1wAOQ6bxHQrkJFrMsITiE068Gpl/
uJcGPlpHlg5BXrsflgeobMV52fagWK7GPqeuKt225UOAXtBiMKxt1XDqZ5TF58uWyILHl6JSMmP1
GGf0ao8Qcfkt4Bwbf0oDzyN1NQZxn3AV8cxcOTuRTFf/m1ghUceciGmUGRT+a6z/cKutbf/GH8n/
s7c8uArH0+QITfs3YtbWW1WunvvIXvkYtzHNSxrJ4B2Q+qEZh+9dUYld984z4xEsPiYlwgZp0C3O
0o0Xz40DUyNkxZZ5sl4Ja6pYpuSdfvGRDsr1DMl8cTErFS++cXOd1uXRElLrA6uFfUKn2Mm8gll8
7Cd/5aVAEvgjrFUsFuY7krqrSwztQ5C7JVjPsJdCQtG7sFOM4JDm6IGI5yJzLdZH441YHx2a9RoH
XnjavXl+YXTLkHF4Hfr4ruIftbX5eCCCY1gWFkFpVLySO6NtcunAlJS4AcxaweRYQmPS2FUJwSXF
j++odG30LWIezX4RPJ17N00SLTbU2kotNcAeNKoiZaOSrikh94QNSdmq0NAOTDbicrigHPopMujb
GOiS1r7IxN2ev/vlOCdC1RgGXxLF5NBhmiw5pZAl7Ka2n+pJYp/7xovgFMvou52JJPSEvIogo51P
IK9BcEfbKgRmT2zUYiFxfWB9srGhisAXXfGCqDb88UAEjrqdjyXNZXpQRY2HoHhoecNWYpRfKcTp
3HNEA7xA5+5q1Pr69JvwBRKsJiEUl/qfYQHmMkOCArkLtuAc5UkynRb0A3VqzN7GgIcRKj4sQWPc
e1s2IYg9plrHUAiG7i9YqVDjGBp673nRusmjHzGW7Zm7UUzbN6lbr67Ritg/oH684fjXvvcqVE4P
qSv3eQSJkQTt1KvqT1TO1AVGoviuyYmownE0kJkz3bMEr9fCWOtPCswBRgexN99q3JXJOuq0Oqgj
OGfxCLfQiChHyJ/zZGnXim0ZY/TTFlWt5dZscdJB/MmRs+l5vmjanxHANewDGnl2wPuhD03HmD8e
jegxT5jYLrZTt63IxWLNI7brkxavDX/hKTwUN6jjxq/HyZ8T+ipTRUZ0mIkIqDfp+SsR6qqk3w/7
ParF6zAVDBeUGxIRHa4hftMXaSILCMypRJrNHMKMYRL4v4AfDeRKykB1RmL0HqaOH/bgwLt+vKss
aZyE+7fvd4Uul6PSjqbU0eqOUsjzPojALb22cv9k7fN1dTmmkqFVzhApcntMBfB2Ly3QzyZqhzI+
iGNthCO9UYHUlugtHUJxoD7rsuFD14B/hhfNuy3tvWJI1VxJpRN+6O5MnFcosgHToSB/HfNRZNlK
D2+wQgK/WhaNcPUqzYHGpqhk61QFL1raV1DgD3CYJx309yGvuCRm5XBDv9v1OLcQcwbTJFyAW2KK
uFDteQNgUEC3HXrzcT0qVxY3D3hvkOR5sOxP/E4aTNXZaIDNQJFJDpQLkUPGetbCzHSzW+gkDmBI
9jIqMHbgJbzTu4t/wVkDlRlxHjudOggciozn5QYM7TU58iv04GQiiT794hlm1VRYzfgXM1iBZLLu
XcHioFTWpwEnh/DNo9vF//kECBJEsxX8YIVwILWwqqVinlM1+UavvdG9xuuRcexPeo3LJZzAVA34
nkzWIJrU37Jst/Nh0ZgRPX+RFYHjCwWz6XpdyH8lurhN9rZY1A2L0WNr4eoJHmwT8L8tAIACAKoK
H2D+A6h9U7MKeK2pxfXRFkkydAu9/uo+fkyDKoB+bCq1lsXdkxqHhBdedebi1ukRox7ZobZ54Hta
svEiWcyiDAdpETCEM68mloJZwMpBb2ShcIXbozPN/OYFE4W276197Z1uvWhSZcPQpElN002ZmWUS
VKYmZtMKjp6uJryD3kV4PaFNvfT3vl8NiAaF+emjpFkr+lN5HdH4ZXR+K8M6yfeSK0LcQycb/TYd
2h4bTVNAYFudEz9Ht2d4L7Sggg7hXAuT4/IN3qs53n1Hq1RqRJR48GewpKTjcutkODiimXBtBBf7
ci4qDrtuQOqKh0DHqaaVsZTK4Gv3uF+N8DosVckX+5Kqqd5e+pd0ggB3k7wAMbRSEw+F+SU5upDk
Pqg2Ahnq0yLxZFn9BWNEdBJZ7e1SFqEoausGigoQWdnH/gfd3o687Ex0k9RwT+wnZgYMbVEKoY1K
Y5PkoSn5ZDfVoYvCM+INN9vrzdyCRJrmdy3LU/zXTETwLkTTAV3TmRTBfjyrUYMb4b/A2L5FCWAJ
HI+M+DdQQhg6+2cH5Fc9KVkL/++18TobXKw/QgZEKaAdE4Xr+mlBJxuWFq9U7Mbet3XVNflblBWe
4KFfSST6Zkybi/EB5I6IlTghwmrnp0UG6DbM41AWAA3+t350uU2BHM5LSsQTMSmkmi9xDnA4fDro
Ddxj43IBo5Jxr+PtFAAijP+C7OCf/DB62+cdlmTanKOXhQXL6HHEz/PBP0TiSu5GaGWCgbJfVIuv
1wnTnRWyQZgfZMLgID/qTruVNuMbYFiJTg0ZK+9ogPN0hwMA3OYhO3J5SjOBPFnCukhiMaXf+2iy
1GMI/54IvUD759lU4hABqrYvs8PqVX35egEmj8Sh3H29dXIIxwwIAG226xE+eDaLARlomVi/tyhF
XePjrfLSvyEd5TAOrmb4AwFz45Qw2m5PGkxvEc1aB3JXWu2ILH3NB5KNSaKDebY5k/I9NADFQ+aA
r4Q4EbeeVMPl9zkl8dztYXAopmdWbotkw7dIYldnCvREkdTVpiAlPLOE6FkVmLUMWldZvEpES6FP
XMw9hlsPTILiarL0aNH5Af1hhyROqLvfgyG3kj9AQrmh0WlXdPbduI2xbg2ALYPZorNYhiCDHFOn
GydcI6laRWKNwo8VTLJgwz71yQAYQJncHfa9VdJ0ipmOTWtm9Zy0bZy4b/tzuEj9a6y6/rT2UU3z
+M9+DfJaNKzzRK8YA3qW+BE9CtT/uC6vw7xCIlOQpA978TtV+blqCC/Ux5Upek9AUW/gZT9vnLZq
rJ2dn48IKhG7iKn2F14p+NHpzw8kAZpsC+kIJRS+onV8Kr0QQoInZibnFz+EUXLFvkn1p+EJar4I
QLsyEkf/tc2GOkP0q9I126RpPpABd4ss0ori1P8+rglhs4oJWaLLVA8rFCAar29RBAIZfTiFwI1G
Q+Z4FCZb5j9crBnYoeH+hjOKGxTATTnRLeMd9lJaGoGz0DINEYaj0/jS1Cof6Pcgq88KXrZdzkv1
8IE23LDa61lvA2VnjOA2PqZ5tVwjx1RC7Qip/ZHxej+QEjsBnMQnaL16dgmjX+RODv5QBfVOWHi4
AfkfYYKmLWCJZAGjZFtP+v7uk5EPTRawL2sSyC59oyXlYC7hkyScsviCMsz7ULbMS2aeKw2k3HZb
eCgEr2o8q5fbGjTAXSCE2ZRmKdCp1CsGIDqYKTcEmEWWn2iLWY5Ooa2a0b5ZDIA3y2hoYMugV6zR
n1wAw63rxTEKWvYJJwANoxFGNE6hDJcqyFZCGMhdmiA6m5IUuCx9rHrXBLoOOtMRbcjOAWstFNri
6sJX156zGWq1fI3JDK2jTxYvNe0PHebyLJUdBJLiQmRE2r8s6kpVzLSnJV1OdfhuBBQRe0J3qW/B
RMZzvwF0INEDFn+oaHfo1Q6x/8D1Ed+eNJmtinILtZOKQ4xdUtRHSN9O4Ca9NRC537alqH63qZH4
wmrh51xDuuRtITZvgFH9wZ/jNQIowbqfCFryhcOGz6TvDtuYK2xBXUf751RqLtiX+Wa9A1HTHuv8
SJ05fnM8XcdV6GxsLqF0hodkEyBEBuvJqgHfbc80Cuu9m1s/mxtCKx/DBHqxtvTRahBTY2EhVAHY
+yB+wvIChhiJqZEZrXTOIoPNbe8l6he/0uQn3I6cBq07ikUyTwwXFJriMP0Aprq+1qDtot+Pyv2w
Zj4uEvlpsvTfkmZQTvSzlcNIojuPIAU8UWku1L4i8GR1Ou1QUFJcifJgtvEvzvn53aObfye0wM02
rLfWleEyIpgxWaYR5pcNnY3TE4rCnqnFcEZVj1SFRKXMd+c6jwE109xdF6hWLUeL6ZvyeYxcZycD
ixYzgIIre5DH4oSMkBHKT93UXX+oPeZBRdZIiNshDvZJxBxOmPru2Khm9KtvP8V8VJCyFFmnUBp1
JWYaRnQtVOaBMC2n5lelaM/gYhfeQ/OX1yxDJ+Gux4lbm1lvzVJFUyi6L6BCbXy6c6vwvr6DPaum
8d9ToUFAD3bzqsrSB522QzaV8UyZrpKI5o/5TjoEITMXa++JwQqhwRplBRDn5l/AD7BmncqJJHdW
5OFKcomuZM2hiqQ0ETnOJ/n9iprrWkcMD7VQ4MgdqlhlFACBWMkKZYzCQT28oP74ajC60VkesuyP
BP8yC5s5ItI4UhYfo6rAZlX6CxzvcV6b852poPsz4kJBpMKaoDKv9FO2D7HSDfZWrwGI4JTh180p
pIgYXI3w4xdqT/pN2/R+e1XQTdHRjFCIGNl7/7k81zdFI7RYuAPxe8piYtFDoYmoPcbCZChaAas4
drvz13TqQBeTNVnQEp9zmXZr8/AQ1tM8/r17w4VmS+zOFDkgACRPdWMRsfk8hNE92BUSv53+lqyX
0FyI3Oex2+kYAIlcDTa7vKAaeb16SDsnFvrxocQ+UOIPUPKwgUX027r3OfXoCJrgsr4NZf7Gi610
wlTZiEI6jUPDEDhn8bCl58hhfkkuF2g8YZZyEYcWHptkBZwGmmbsMrMQdB3Z6ja1SquHnMPJC2UV
pwOf6+AsDVthdF1yJnjAc1f8JORedbigyOJVQpeRyF4bNNXfkryGd1uJyauntW7X09kGiuOAHk5e
X/jEwtUE4dqlVOKEcfP/g/pEcjlwzzS6jD9yGdUT+H+FUs/xmM62VrZz4ko2QG5nr8hfaKWOZjyA
QyhEGzMydlYI5bRrzQM9yed30MB138BUdctvsC7F+oIoGP2/+M3If++zsgvNc+Tt7zu5fTy3AOPM
GgHb1bLE4pWnMRYg08PB6EO+Ij1x1qGTfQ6HdfEWqDrbXQ/iTsx8CgD1paLgbKlQnWzqE6z65Eqg
BQ+XOnzPrhmIJDmPbHbwmVfEYuQbDNPok6hFW8VKeKPKRLmgyzmpL1R6qb6mwiURWTsEdJtYRtAX
QO7PydFRiKTimVX4dzoZQtry8YvwWVjx0lWTtQZhI70Sa/N1lmkGBV0LIC51TySO/IJh7NSummk0
V+6E8FQHLDT36wiHpOGRS2VfwL81o+ZGKqCcQgkZwlyCOTMRhZd3C0Y6CAgocWyBmOFVrlYAdZMK
xBO4Bs3XsI67DPqyCRXu/miRpHni/XBD6qkbwcDSBQgXGacNny+01f2bQA8rU/nATXo3KXqCmo7I
zxLhn3Wd4m0CsWXzr2d8Px3R41xjqA7Yj/hyDFYr2C4H+6aPDllK9isJ7NO6QsqFjcm82AmOK9US
UMbCSFzD1DzAvSSfCrQBIjuqp0xePMJZZ0sz+ZWD3+DlcE42xp8ut02oglkPEWQwUIu/Tmx8bwXH
A7pIx0Fg3qWKfW62+oakqDmA4m2Y9fUoZQw071cNbJn8UQKQD37RMmpjQFRoHNZ0yIWBIJMQruZC
doVt+u13vLrJ1MTD5l3vTsKy/s7uNOBvFLWan7Yq9CRYU9pXl0CBAHh9aMW4HyxjFdsRDc+VwxKj
YO7Pu037IFp294hZn6Mqqf0SoUbxtu1ttdOpjKQXShoff3pU93bscnV/fdvglpy6qeBT6W1/3L99
ytnvhVinwhZwnhPTqolP6IWMERF5PA8eP0ANw49XyURqiV6rtLfDCL6PYW2MwGk9wBq6UQKwaSCE
x10F9ZxMeeCUtm6aZtJyBGOY4Fa4afhrVFD8BQf/m/DDc8P7HA2lZdAuL2WrD1wfGOelv+m4Nc2x
dlp0RxsjBMHyr3ESbMSAobecyNog5HYQg+aEH6Hx64sO3RCzRmJ/ybEAGywLFddZ5bRxyezCDEqm
fqsSUDR+MtztZBExG96oCTkHVnX8+Q6eBNw/8Vb4OsP/Q8kaIhaXDJSsaO6VWwinQ9RM0+0j2Qjv
jTz7uaR4RD60zrCJWaMY9m1k/qS89B/9glx249/k4BRUno5yOcDdjiYQHUp1d9yIhSNcvjvR8U9M
N3n5lr8VQhRi4Oxn9dPG8I7M6xiJFOrC//s+/i5+6Ew8RyyS9tNAVKuLGeoN2Q9Ve5v5Ri+PccMK
7AJM7Rp6TaY1wvMpovVLMVrDz0ppFgXq1aaIJkEZJUn4Y696wpSC86EB7VldamG+GoQuVlN3yakR
aWDMghyR7KE6ETh4RMt7kNrqtPcx1QdFCdzMFuFErwWRsGxA/f40hs9PPcziDibMtRbuYWGF9acD
oG6KkvH7yKBzJ88KfSNo0XwkHBgy5t0HDi5H9Y+gMz1rCao7HvSsQqj0sPjvgIbcSJKIfi1/Gf/f
Q5kI3zpahcD3Ek9GK26mUBi5qO9SCfBSCs3ogOlE75U8leUKrq+ErCyrNSobOghWZT7/DLq4oNct
B3ZhNLn1uUyJaEkF+68Qk4k++CTKzn0XXeQvQbMPBaWQ8e6H+E/aLT9Aw5rtREI0HmXuQySDnDqd
vfC0JfTT6fTnAZmS4x02lPev7oSCyJ01HlIzy2q5EZQRwvZt4Jm3Lx4I1SjQwl9K7Ijaem3oQxww
KVEXCHagvG+ey6KHoAWAhthXiSWKlRbSAcPhzJ25C0ib8+0sb10meI8wWOOydOwgOAkioBwu+7bG
ng+7yYPX3Ugh7zBRoWgr6UiXBukz50BY7M2v87QWjlI0N0jiopLFAUQjY9dQZfMfoV3jF7+u0klC
UzcW1pYMYsb2X/wrjNQvAedbCNN2RHBmVlHsXU9GFylFYCRT7+ZN+QbyYyki3Nqs2rPqT6HILZkb
WbeaPt0lID9nf4Mz0GmNSJ29VYIgHOrdoI8JEcsxReFqLYd+Ha+ibhSjH2e7QIECmy3lgZWfK5Jb
Y2F7zMKQpIBusgu+tUj+HBViAZjUYOsXCK3q2izeWEmmdzMvdtF3zhicuyOpmuOatPIK7G5qGASP
oX5fjorMmFPboOxpK8sAg8ZkA2LMfJ+ea+6rcAFQgzimOa9gJp639geBIilHB8Kp1RKyBerISoao
qCOEQrz1zV1h/gixIVdgQxTOjFigWCV5JUQeIQ7+OfsdFVaoOB9R5nFZVUmBreABDLlXTzZMc/GN
jRgZQAbKBIpqoewHmHMwUa94rGGhW9X5BVBP3n+PARLJCXrltsmzocJ/V1j/T0MMrUgb3RriZHPI
MZUY+oE8m434tuFrrE7bjw17f4HoyfXvxKtqElDFCjV4BWFqOOswIb4T+vNMUglogntH8qXHzp5h
uL4GmM+HPTZZLPhMim29Xg4DOyr5lbijGVSr47Vw3Yc602ZCO49wMFqviwZcl54b7PB+Ogu9XIKp
TLFuaWiMGJ+iwXz7wwVEDlRPZPb+eOuxNtDyKca1qEYHzug22v5Ct9egqsMApHEm1/8wZl5idoYk
28Jb6Zd9w1fhIMcaO04Ut1v05VyU89SInXvpKcxLS9XFuqCvbnN41oGVhfPldWcjRLN6I5tFtq0x
d6uLx+WGKaaG2e4Cgfj5YjLLtI8c7tMsPJZsHKuFFCRkQuIu+qNZe598375NTT38kPVjjscGTgGv
4FeHE02IrmhIAfaQvvi8qQx3UsVzw1aFx8Xp/oYCk8R4nInHhyuqhxjBTKgxlYqtafHoMEj4OApR
yQQZD9FOmpQz0TB8mU9O0dty8NsyZx1JsQIu3BFpXCPcCAyKBnmLiFRyb+OZO1EqeQw0d05mtFdW
J62YN01sX7639QWNa7ccMolUJxBNp/byFtFvFDY30MamEwFAiDMwQXHdhObDbwTjoAL9ePD7i3w7
0qmHUu9lwrggWH9n2aopCU9bBi3RJa463Nlt1n9cVogMdOiJVn2lxyebPWI/cpvPYLdp2I5lGivm
uFUb+xRiq91fEdFxt5Z9q9sVzEB15aFH3y6sOB8jauv7EbVMEesC4xLwxdNLKf02IPfEaz6sTtNU
vTFuj6ziGOnjj1mmqRcS8iGMNCS7mtRgcgRcAwBbJms1gMpjhETXSUMZwVaZD/j4HidR4aKHi8KP
7E0FZjQrVPj+KFvyRwNwgcNkPULZzomHdZGv56AmXlSBobEGpHqI+kd6X0G6Je4tE26/TYZEeZ4I
xHNTou8cF5W+Um0nV6ojF6V7fLY56bVIcO/2/JSahlRPf/igEuieK9zT+TxhSQNlvGWVwViLymks
16ASjOqyyqd8eyNReLsrLNnXXzNR7fnVBdwwY1VZNB8RBaG6HZMS5Idie3qt8b+FfvhlcSjiUzf5
VjJeOt8Ex10x5bT6sfL1bOCkSXI3LxtsqA5KsYosES/oZoixXrhvyGVrOSyGHQM6Px8MpdQ3HK42
eimMXA0DPZPY9iUtxFCXin75fRD8c+hIW5dfriYEqaWbx4QNQ7xniiBSGDr85muVFml/ySU34Hbo
yZ0jaRj+VVIUWN+YV2hdXvZ9YxOBmt7gaJiBrFWpFvEeAsMFVwVL42zR42UHOxf2t0xFuSoawii1
T2iUgVvX2Fwyo4n6EPrZExghZCKTzq3n5s6PzlLvS1lVPeRb5dkasSAV/yL2klmGUt8Pg+UtUQcs
iGwz/QK/ZimGFrj5qyVvgr8CUQFUQbLyYBqA4K/9JzV3SAU2Dt8DMsTd8Pi1DjEbInQoR6JXLsjv
YjWc/3lWafvf9XoSpoGadFjO5amxajo5PkCTHYlINOHpdACCATujp2RmWntb2SggsJxjRPJDfJat
/8xgtp3q9tUflKy3N90WfTSiapxJQkpBg203Veq9jCZToQ9FhXY1w7vxtnjn3Pp9jHeFz9IXTiPK
usi9PbcEpdAiSpGObQsSSlh5+CAUKW7OjDE/4n8Ai/YEj5jdhIVYViBtfiL/65HlRnVpyBqQlLzP
WMh2IPRBPC0BheMeStSwBd1CHEOaLnSZQ4DLgeEq5S1qQZ4ey0ZbsFaXTcawt81aK7MkJexNuUcQ
ph6pAKYtfNxG01d9LaF9QekCoX+WpH3TABQEdAerUGqqhjkfDbodS45gR405gbyMoia+j+6DBjP9
pVKXnmkAh8CNukFrBY8ODfcquWmu7/t5gzBqiRYLfZbN8kWE9qxX2UfPtACddBx/X3tl8671qG1h
zxReNaQrBdfWEze9xjX8vE4IvPEI+vQOwadsDDOvy3O70bzWO1g1BXnLAJPHJGjhbo1GFhaXt9FM
l3xueNZ6EQKg8YXfnf+egDKVtFTsD+zah2StLspBFAgHzKV2SDq4HcCT2wwliAq5dfxer/aJx3qv
k9Flni6xRfyts+Jzh5ki3P4d5sKyBez5yOTuKG7+nnsscUaa8ejDj5MCk+T0V5vPOkWJ0p6GE8nG
iejspF4Oa4JZ0C1CxxrO0dm05iWvMUyiXkAmLYWgaGtO5AHiTg3rEzUBa09GFR01jPrVYaFVxVS8
dRp0uNJJX4mzztRn3iN7g8dnUW9Kv9GB/PNGQptr/2w4JKqEZFNw50CvvW5mi3/0PCHQzvK9vg8W
Nkx0g1/yFkYbWHCXrp2dBkSalCUopEUtaYgtYV1rmEANAvzLsilIfMmH6vup6bEFW6dxncU/6yXm
v1KCRTmtOsGxMULW7Vcuo0MkFUZmNAwuycKKIjbH/roxf88MPtFzth9VhaMebaKGyTwcVFjLuUNu
w/J1rCoOyvR5ud9JX3+kRM1tzFWmuM2uMUrrolPBi3+kLMZ+yVOdjCRvfaJLc2XPap8t/JQmXxAC
sNutt23thqIJVjTiO/kAbG0vsU3LQ3vvtWgBqvqm/h2kchZTrBeupja1PScDqgv8NkCmkTFZ2q9a
QNJSuLSLabqv7Pbx9s+eyTqKy5E2VRJPHNv81EWxFJGjGrKik8ocIBkHNmgo2l4h3OByYxFgaH8a
nVLEpH+0500xkSxE7xFXb7CBcNYQeT5r6Z9xuIlypPHA6VpPt3bzb7SXh6gpvHn3TDW6V5t7CUsN
5wzq/dXNgI7JhHIA41x8gpa7rpCiLKQ6X5z+ZiUrOtYlvFfExSqXkAN33vbp4vM3IH5Jml7/XzXu
IBWYvZbUVWd11sNkhRk+0bqF7kmsAZhyHoUZ3a624WX6bW9arBJEfxmqcUUjPyBmEvoWpVNoA1S8
NZ21EZbr6Ht7uMvJhmmbwhEbyaxFQAF4cf54jhE9wGXVbhx8EkkR7mRMByZhrDq+C9stMi6EHjzB
uRebrLEAcMRkE4cPoENlMJVIBaBQxpZrIwCN7mFOVt4TLIyErt1MfrTNBZVNarPnHk5IVOjFiUYC
1Tt0otdoDxyZhh8I0MdHtqCFjB9JkoxvKXV7qohTdx5HFFIkV4KeB7aXUl5dF2m7AAvpAW/PY7OP
r8CwxBwjjym9sTDvIaL/mkOAHbtsGsNO7jR97Xx2ljxZu/yMTb65Be3fzcSCVEYEnwdmtCW6PctY
6CikRpLh3c3aO7wiRY6DT1OcmED9PtFhLfxVKBb5U1FkPGnZkYLTnMg1B5X8SR8oq0tqtbbyZtEE
MF+2LpegADDYuWaeggJloJKpq0prkNGh22R3KIq2U0XOdZh15OygMrlsr8Ak/A4wRCKgmpV4w/D1
kiaovxOzMxiYfgTxtnfgRWwz5XdMB8INJ8pEJC2ILv5ETJQojxLk6JZEudh7fftq/DfRHv6u2z+5
0DpZ+13j/O8vid0BR0UGPtTski9SjzuyfFtHoXPHGrfwlqP9XZ138cAnJ1YqAUA1yOddKfwnuEXZ
bmGc2MP7otNWSS4VM2+Lin5IXbEs3G70jNM5GOiun5/9W1+ideAja4T5bIWN3fpfZnX+HMCBBlG8
GiogxlxXkDUKVNTFyhMe6C4VA3fwHMwOaXzXA+yUTr8Gev1KWTfhrmWet4vlxmar2IhCKvpI3+Pq
uXZz0pPyNnX0uOMIwAnL7yW3emUN0NqmTcdmnxLcrWXP1w33QuRRMeF8TOyjHVdaPju9UlUO7/Eh
LO2QHMoLHvNornSwc39YkQhMPFe7MaFlb16C0IUIHNOKc6W0CUpv6yMMKwZtZ+TgHF39ydNF1H1q
obaosB3Vx2E2LXy2hbFw4KYlxOd9cI3Q4Dhff9E1RIkQ7ZsJPFSKpHPAzw22MlhnJX70yADeyb+P
7jiwxjYlpRTPtXaW34yhC0HgAv2QIa3ijT5+ehaSv7w/9pGjBy1S/VnKj9wOZt+uZ8SIB7FH3awC
Mszixs2qVGsis8ZVovEu+8uupi0+1J0s33ouuUtJ490CaVyDbXqXIWA6OcnSxebJzkDumhZSS6e5
ABolv7AHxmcpFjxVgYoUnrjoMzULtPuaypGEFBifSQ6//6HF5QUMFdNoqmIIXnVMNMA2VZW246hT
iL6jozFhfrKpQS9nbgKkapezoGKA5YzM9iJj0cX05ySkVL1Wzgto0CrV+S5CaP9rDECLDzrvDqjj
k7x7u17iLVNPLfV2MTe8TFeDdJYgwuYiHx/4RxT/1Jgw5hl6UJIlMxHUKt8ZJA1/QVz48pRHprQ1
jeApSGq16YX/5+vN0JCl6KR+ChxIRtAecEMqbTLI0LdK1a1nxh0g72XBpU0EyIrHPErwpkgYCwUf
J3lFL8kNV7K6f+6V2dwv5YfhfxhGCVvtSeeGcD8YC9urYWKdZBP5wyIwCqAfWarBuDEh2f+7JqkO
fJLCehqEQOABLEaLNvR/NTfrJ4jgRWXZpso37UjnURd3E0B8T84UozMOBsPVoxGi1effzn0iDxii
A2/NnkaQZXYdz7nxpJJeSsHUn/wyGnfRWhYCrJRTVPHzy63qR2osuZFpKjhb0Mrc31ZfAJGoHwdw
EanPb2XWIIlWhOi1/GieeJRZlnwYBxTkRYLjl2dNcAuv3/lQzhRaMtz6bHYtAG1mPWmZ0JfmRbAg
8oCR5lmt6GJXsEAne6LyZHVsg+YU9By7kWJUy0jjaqCy9VN7fLEmjKed/DsUq5MFdcryllPKNfoC
4Y5wPIRsteJxRw0i5m8nis382+y8cGgCypmRDop4zdqm+Ib9JStGiWcFjFg3w/6ZQxtO0xKTlQhk
lGVqTmyAbCeBddaqZxBEbDPf+oS1TO357C3HlHMncRHBQC8tfS98IGaBoJo4hZr2O2tdw/NdUv0n
YfAPCnONxZB2qfoBnKWbLRZ9wfXdUQ69x2yZdfdkMBhXGhjhG0V+M8JJ5sKxfva28/wjgCOi5q/t
4V4bK44tWodVBc6Pz/s9ciADZJWlqBlilh3wjJZns7rcalypiZ6w9Wy4iziuc8UT+6U9GLHZvwKf
axsitqkgLbb6aiG7ti8hfkOQ0PyCib5VmUy21g7+nPyT1+F79p4pqmTMMK3uAKN9pC8UdU6ox8on
Dul5LxG8iNDduG1N+P8ms6fkWHAulT7cDOEw0jCpj0oWoL0+gBrhwcoHcaRodw+H9Shh0phe4QAp
1DGDF1OXJUrHO2ZtAaKn4HWgz4Z7DrI7kI32S3OTcub8mA8TygOebkrGt0mgOB5cSYrKolmM1m9m
dncbGCZZihlqcr3E72nltIOXZ0KWeBYlCsXP7Yvu2RsvJtt6OoU1CzxQx7cW/7SJP13lWujRdbsO
+Z4EacFKngDMhJhSSLmTyW2MrL99N/5Zec7088i2E2Xdgn+8LyOw/F0C70GO0lJE69UgJ+emgxN0
R8SNcS9rDql3zt9PaoTZ/t+NA0LIhKIitIbck6Oe+F2uSE1tb5LUsD6AZEdjitHw2rnw+cuKTqhX
1g3fafxAXSH/uPKAPRQnKhk7K1o+SYooV4G5XaWIVMwc0mLdqK8+q4XeGBmU1J4csDGtu9PKKzE2
ewq6nDY03XCBC21kyA5A6v9pJKgw3XAIAK+0XdZ7BlVq//Nr3HjqsenkfWpYXCl583tpoUYeZxUx
D2B7MtDknD+RmqFm0QxOpc9vQhXf/BeanS8A38HD4MYsmvE9xPRXfvMnZlF/CUKS2JM1WrmddPTM
v4DGPG8+jKtfemCauL/tw+S3wNNVO2Vtm63kk0RtdRyep4ZzLvDIA43urK/oGts7SLs+RNwTCDK0
P+L7NqMtdc/0qOvO2F/JOFaATfkzj9LNj5YC/LJUQLA75zYKpV5eADQxawFGrRsdS1prQ/MQUEBj
d5aLbhL7aYQ0yxwYy5y2Qb1SXUwqoSNYXil6aH4dUKWYPHQwRLS8LCPUdNBTLfsHau6ofiBHMqQY
ZaFN7cwBFu1Hg5lucT/ncVPcs76TLOpH6LAnk/HSFmOiVsuzg+YXFNtrY+d5PoNrPVGEccIMEpGY
I6Ree/JEGBfiIU75LanUHvkzICFLpsUVBWMHmXm+pInHvxAZ37lObEs4cP2xgexabq9XbJt+A6gf
h9BpRdzYUli2TJguzHYeB9mclh04gZQ6F7yvvEZ1gWZjdJYiGGlF8wput3uefkNaWKr9eOn1plaB
woTdJFCq+fpuPYoOd4foLaDovHOoNL4Swl8PsU5UhGE2M7FJ0NDbeckm9rCLEJw1xe4ZwrO+n0WN
qegtIIECG9KAm4nO8GTfO+q7rgdOU9Fd11zJyPtzsMAj75k2//PEbD1Gp1HD/VA3vOQMHF7SvIwG
akW+uu+XgXxBBMktl8IwDPAYAQK7ZOzN17YWkGrGObzTcotWW39O6wp8MtXHxS2hGDlBqfQpfZKU
99JmXu3hIw8ECw4CE0x6sLW7zT/qGBS5XiAUJJKJV5nKA1+kaSz/aiyZSs3z6qYmV1n4SLecfPQG
gAEht3ZOd6ZUEwyBejFwvr/Pq32HSrOL+/fVYaetVQ9JP9DIQELppKhSy6jNSVwM40AZ4a627FRV
8tb1xBehDYDOy3DM3jrigyp6ydw9Wx1ilasZn9N7hG5il3TMRg0ks9iNpx9Mf7ecPfMKhtX/Jero
SF11PKpYEJq7cOVsCWW7cTB2wLbwUxmmTTHCxUVaRTVOcOZwPyAZJslHB9ydtCvgld6vHJmOKDI+
NZwXULK+mfqnPC4ABMiAvEVLOGIXjwpGsuPrXkwON5vDfBeTCBM0STm58etIVyM8JaE8YyuK/CX7
gbwMS8V53Wg8QaPUYJrxbICx/iRHBri5WZ2lgpg2/8Wze1Tpr1MtjpG9QvJgGjNrvwHj0tsB8XTx
1ACZ1N8yal02zenxSiE/ZXzVFZoY2ROY9AUROHxnaL9pYbSnM0r5OkQVhNGUHK/KFPFt+kJibijD
iqPQjnelzVYxk20yPro307ZSqwyEKR8YLmdbhBh6O8nnsF8mtqudLbCACpPpSwpqNIoVKXIYcHxu
XrFOB87GoNPilSQIerzYyuTdfWOjPhgIliD3YFgvYWBHChpZsjec1JunL3uzg3wFLP580xYZlHaS
wxXqUgF1a6DkpeGIvkmvGeZRjaVQ4zrMtddYXD9u++T+OZpHqfDrjLsrWZA6syl9ABRXPe63loqm
ztixZfNPe+Lr8UQxAG0Sf2MdEvrgtUrdZr1QqD9PnwEVvMkOf9S02o80ooAdjmVDoXPQ3/KO3bNE
DW/tSNW1VcSLczT+XsvpG+3jNsjX2Nswenm4HKdawZlFY320iyUVAEFNw7He9N28DdgB1wnrJvAG
i96RTu5VPTP05IzG0JG1WpTaCfETfDVsFkNF8lznHIgH0ISX1KG6EWVmH6VHjs0/QrvXYUH++9xc
GtboTubZFOIlVaBod3gs/kEFUoN25m83hMd5tfrk5gGUr8XOEP67pUdYaIApw9Kp/rKcNat/o02D
oDO2zLtQN6wS8qlykuZ2mIcOnJsP8gt6nMfLOMzvbI6Pds8LcC1V3pOsmylYjYe2h7AZNWYakuYa
tUNRy8Xvhi3M7Gk/cRdfSQxWrixwOb8S62eGMEPfvf7jMk2LkLXLyGDBU7lcvzFBjf0lcu7zOBHu
JsmhY7hNTa9IjIg9CQ0lnYCA0a/RgQLtH8Y08ZEePbXSHk7Xe+Rk97PznAUFkNSCY/v5JrewI5lm
C/Ya/0+mnJlX0QnkAH82Vj/gRigv0DzAECOhvWy4gkKCIg2uXsvY2ztflOjFqDp8zhzcxMNy4KCT
T5f3BYvkmGpIMwABrTgwTSA6r4L+cnnlljIQ97Kqfkg0W37Sn7gil63UehveShbVYnCQdfiztQFV
STK2PoPJVRtbZlxkSLJL+iWChZEPZlAdqZ0CGsA8TECkqgZLTYDpHkaXp/CdZUzbbqIcMhRe+qhP
FUBeHJqfVA1+WgPSexYM7td8PJej9WLqwm7d9sMUNRy9WHn50hcy5fTDz74ff5du49vilX9yaXT6
QOCvlVqfUKiwbdGTJhCORGDwH0Bdn4N/seHxZahYTQaEET9OiPLdmptFDMCflm9be6pPJMmHwiW+
oLh9NIWR3LzuJhlIMuZWrKBYs62M+Y8Nmd3vvci/iHDX/hR1inYUWWopavPqatF4KcxWJZbygWZF
PpURP7RoqVz4j6UdBEr8shiuM3O6acx8tqooXxLB6OZlxZwXbksc0WDPUB0xPMo5PQutdFr4AVhr
EVawmA+baNevTBtvHH6Oxj2h5INV633Y2E1gpb3UbhqKi07EzSxvb8XfWHTTOaiDgDyf714zVgMa
ESHCEIkNAjs8Z8AmVqNKKoQ+xWEfTF50aeI16BUok4mzsp9VTCYquYjAGO9YGIjIfIxEzO/PtM4g
rDUHVywkqrAscSJNlxAJUmrlszrKUfDZgLY3X1NwkarT6mE7rX3SzesK5u7kAMNFFFtGTqm6rzco
iBpCzXQ11sd8rpw65o/Fpf/nAfWBZe875NkkULEiSS3HyhxuQZFuXsItDZIbrpEyrfiecnd0nQ5M
komSzpChspeqn+WRiuBxi9LXYfHAb1KBUwZy3T8zzqPUHiJy/0xu2nr0yatm9eu3bQsRWhptL/55
O6VFNype1v0YurV4i34VtnbyVQ1lI4ZwYb7I96y1zH2h1lymJDX3st11ZlOMKAZkvvEs/r1VHt7u
98TNaao46GgKLGoNunvL2y7//cxeOosV3q3ciODiUTOnZTrrMmrj8SfO1pozguxZvXPyzEpWf+WI
E0Y0c5/paCI1zBgAR+hnvq31K7T/Q7cWdPtQQ5gJCxClux4pI5i7gopHf2gHdCVt/sZAJ3rM9l3N
5xaibP3NgrW7YzoC/ymo3A8+Jn5Qp6xFU+of5VK7zPDg5n4ORZYXZ8Kj2wZzjwkgIgKh3H3KrbRC
7y6OtEnKvK35ArUw9LxJI5jnlWEetIXJnGklttp7tWENuoOVbxpXI/eekOpg/rCdjMqT92EGf1Sb
Suw2W2oqi1wcQtHUUzPvtF9Bb9r4aPiR+cCOcsZA1IdRgcLuxnjlIKf4JLjrFsat51HQvgA321O1
D8nR+EZ+ddBIqOOQzbKsr8GvWpLONny2LxNBwq1VoTNyIUVmg7O56/CDfGuHJTQaRMtdrriHfuhX
TpzIBPtGu3amzuyNPYBnlRhMild+YEkgOP6H/0HVkl/ndVZjGFucCASVCaScH6SR8kjbPWqY9JMJ
yC1Tqm6SU591nTnBTpYMtNwj/YyLWzAUnb4d1ybXjfbq97qkDj15lYM7qf8u3kozcfz/0dK65zpU
vAkL1FUfm5PUH44BKfyAzFvEemR9k1pp2MYKPzezGAsSXVMf+DYQs6TDprNY4jCekUES0zc2Ff9B
LpNL5KQ/mO+ig07NKWRdoyzym/Toa1Toz8N8QnGmN3tpnPr8K25fVoZ3ZCu8EVj3tswLcvIQakDk
sfuDi4mV8O1cETxovWiocdtlzbNq/NwjQ0HWjjL7SckoJuknR7IbeV38O5rAT5SYtA1px71AMPI1
pytv2siEMxq8QxBVoQ1W+ra6f01R9B5VXrC3KM2UmQngtYf5yNXobOh3DUWD3tp0Sg2oCBKjPe6A
VbRGNoUn49KtQ/Pqs1GXGu/pWR9RJ6QGQm0Ic+76O2yqya6Hl9OGTApeWty0pZaCfcfPeY8HeLe6
qG9WKi3ZsLfxtiL34nhUCW9dtAme119PYrLQmkoDv7/JQ9JOsbOAFLxH+9bZZ0VbtkHW5QnJGTxG
iStfRFjrpAhIsDawnPnqeVmyDki+5fRWjFX/uzOuaoGcDlJMtFwdGzi7aYNtC4R+hoKyXQx+jWa1
7Yxd4mSNpfZJaF2TxgmdEX+seWRvE03s101Xt9gJsAOy9IbmyE5GaTBwsizBz37xQcoWgim0bUj3
FBgOtIUU8guQVcQqu8jF24dK6WYMS4tJB3S1uQ9U73yP+NmU8HRoLV2ij658cG63yTAMrzNlcAhu
8KBpIXXx/hJz+n4hYE84eX4E+QlnFdU0YdQciZNLARdMMmsWkvVIFl/iMUkZOinJnKc8aBCaVfF/
b+f9McmlaMWqQOPPfQT3d0ICO63UfzlPCDUeoWzMGN+dL6KWRAlu5UXsDxQRltz3iE1Zw6ozFSOZ
71CplMaw69P219lfwVJwGXCfgSd7V0KuqQ/ppF/6dKpPSN6fsushccvjYszaFNc6eoHpMLmz5IsQ
LoZ4k6NSk2MH9lcnzgxAkspBw1nj5BgHZwvzci05J+Yqd/Z8fOjQFn9CjXy17EDaRfZJR2tA5THp
YguYKsDjDn7I/5KWP37wpNLp06NUoZ+D1LCfFlISGdvW8lNPDtMMZZ1ktRKdPNfJf5FXfdw+yZla
wS/vo850CUie5NIcZu0UuYM+oXB5a2SdZ3lfVCbKkXJOf9i43Sid3rHfuCPXoT/l/MBpv9JYP6FQ
CfmHdjcaovHppARsuWrW5us/dtNVtZVdYwyY5NS17YLspsrqP0OsVUMUIJlp7uwV61MyTwoezcC4
daLsIEsMFq4TXR4fqoWLyfasClS8WEQgdLE79wsoBaUlwJz1RKkExZcu/yOnD/I0la5FJpI+hcBm
Q//wBO1gi6gsz5jaahgzsi+zTRcyL+H2txId5dmz+p7hdRUcs7R8fS8De9AdcHgWZbqVtpQ8W5Rk
sLzPyTVm+sAf/Ri+yOZpBZkRuIH0iUXXnBEVdiwzwviHbxJgBdUZaNgH52UeQmNNsb9MTSb3rY5g
yH1lfe9x9J/gTC0E/vifOLLxmvnKTL7o7341S4UGGrEQNv26DjVHXxN3qI4Sj1wQ6qepJArNOJZJ
9hi7xWx96NaYJ/3CdOk2WvEDViG+snO2qfi0B9XBKGj575/kHMAFT3+rtFR27uGYEAlf/leajbXi
Z6Bj6sagKUHIwFrfFj1fkswmBORuE7hlr4LMuPDiNb2/wH6GZPhJp43YxI2/EoFgE9yd55GwdSn4
tz90STO5nHosVksy80MZ1xEHiAn8qdLLQvB96z5abRJ/cyzVy3jqN6Xe5oC0Gt3Nx94f0g/+Hn13
+agd+IPwKQIhF8nL7VJ1EOueiZ+j63ikaydCOnBtqW0CSq9YsWyAscypGQsWyXu6hQhlA68BuQA5
vMUcKhO4CKfXOndxUhRGdP2PuOEssIhG99WmI5pFPA8ItW+OU2YUFvvnHx2ls77y9TnHs0F7+kOa
tGYWEUClfNdReC2lSSUa2w6QgVr+2iPG2TpKh345wxB9l1X8WwY3M1lk+VIkgzE98vUiCugtAYPy
gRTVYpUmzDRvKROzHp0iYNpnjV6G3BBOvArMT6CguNogDLB3Y9pwAAX0BD2aaBbBiGScKm6WzMYT
heIqTFitgppfgROeF9WwB/Q1KrgvKQvS/AJ8tqUgshkZGDINucay4VeDdCneqaJk0e0mH/trnk62
vpv5vSkIAUdlqBIGdhP5N1ZVYg5awRcxZobOrFSwjILI9Iq/FMVBBOO2znlj2OC1wn08GyiyXQuF
EGlMmFgehDzwayMlXPN+8jD+oHZakHiX12mh2OnswktbHzU/xFSxy6/KjHX1WGC3U06ajHxR6EPa
T282y0Zp+QSMdXhXYA6wKf0PqhMQcxRXve60mCHBAbYvjK2lJT2xRj1fHjQHrZRDYJ1yF7IzHZod
hTARIDml+IGYJjdTbRMIT5nnu4r/X5TEso3bACmE+NhqjhOMmx/VOPbVvqzYJHRpKW8fwNFakYRN
nZnCbyQz09G67mPa8H5zfptehuXbTvrxwbwImX/FWFo4F7lkAY30wsEBlef5Dy/znf/7rRaj4074
85ZnNwhBpvuR8cZ0GBPnrYK79Cu0r9l0022J/rlu0mtcfSV7dtzNoWUxPYM3fJ1kTxRlBZiZZT+s
XsY+JL3QCYDWJSaY0+cfIztrugiV1QbTpIz2YRPlUnFALgjp2rnyq8psmDLZxJrnDmlLCnq9WWKG
t5LAZa9XeWY9coz3dIL203EUvVnqCHSHT7E8jBN/v3h5aCCXWV9cULOEwqp5srz2Rz6KWE4kDljf
nCNo9WOLUrx5XAjWpK8nR06EnnieSlCuvoJ4ZxFeKPSL7/+QzWvSv7pidB+vU1wcdYM47w7NY54W
93XDfkgFH8/JliJ/+s2DL7c38eyNrWjq33FosPpzJ6ryaOw0RmxdYon6IQZzuBQj0mJ9uc7OyuFK
RJUZySIDG049gAX6ZzYP1+UKUw1mNl68Y75AaOmdn3/bBjFI36LWG96xWkzLKGrOFT5visTWD9L2
S09phQcx5U3vtLoBGzgnUh0m0IbBcdFSSdlzm0NgvP5Ef5Na/KhjexpRiUKhoN9XF9YOz5WSGB56
aTV6EwgR8kNjkyVQuucL4jSQ8hJQeQRpQ34+aLlZQlUG3pu8g0arsdKVCSksFGoGIwTFNutXbgkD
O7XrKcoTEgM38jqEJmyu9QeIlrYmQkv/T1vWu9QPa9ZGB1+/OBjiPRidyAEDZySNgVk+c/E9nuMs
GKDD4l1AC4gumZ6co2A2RznuZDtVVu13/UVNFD1ZWDFlejJ/ZgQ+8PRDjSNNmqV0fg67XRj8PQWk
bfuErCbb+1da1qv5+65QJevd1faWWVyrFhTHSv6wuYI6MWOVVfnNcT5V6P7RtBCRKUDlB5KCqm7a
XJ3e5AncOOTrg3fJkHo9suAYYxCeeUikLjYhbNNmVsi5DnWYtww1dwlbR2LHQb0lXp9HQ3Wta4ZF
zIbcd+CNLIj5A7IBUNtYf8fN50rSVDvU5CBKBkL31zJoCYQw54EEi9YV7+saWIFSwopD16XnBrwO
U3LaJYizMQgRNJ8afP+SeN2lCKRIOL4+Qx5Q5d0Kyc00eSzKXq/X+jWaUsV3odvrFdTfYPft4WY2
R3YR6ZlHmZStzWiYxxauhBi1yGJCXiDg0gdPVf1l+vIS4b7IelXbDJ6kLOAgtLucM/Fk2V2tEYt1
YPnuuFXpYv+3cMavvrn0HmAVZuTJWXOsmLtvOpwACqr5eMfqfvh02L2GYNk49eK9DhcN2ZKR8vbI
oglmI3mJPXzA8facKmQjYnxyAsmwgBOaaYWdJm9x9sSyOTsqgP/JIWAKXDs6Yq2KfxDkv9MY++ky
r72AnA6CbzndxhQS7TXh3/cKshDnhZVLqFk4/JJnzTxkzDDC47QZ8LucqtCBQfv70wKUhyF78V5y
Qh+cJmmQC6yrnkM5KD/i0RPzGnVzzbmlymrUoAlwAGTIT1PWDrOHPrnDZmbpFvdeUU5fPA3AVXfm
MXgkGOqGtXA7wKLnvM7WRsBdvQCuYh3WsTud/8ssFZVjE0GzGPSoYgaEScLBwgdL1Ylxgx/Ufo8y
wXx8BtbvWKwFNXk4bIdGcHKd+Dqvnv2vcOuQ3nwjYdIo4VbKMms41XfWExRNyJg0DQfnVYOjlr5z
RTbuAz0+sJts7rA4TfsBB8q6IF7zEFHCjJEfJniqk+kUi07jw9z3kOpZICX7cZYPjPhTAoMI/4z6
CbAnESr3OmbVnMOI1HADWoyjJqFkvSlZQzawUbkvzudbVCvBBbKy0T5VZs2iffZkIycQKriS/oJD
sinLVOBRov0XBWqdxbdQYyD3kBHbrafODxuucSQrYrEmmF0xD64hYu+KonExeTQzLI5LRSkW67In
lvxr4zDStIl+F9RSwMJF/AYTNAvyjsUardRnYGZ+q9isgdG3hxeL5OalH4dXN8UWFttu6OyEhOBL
KKlKdJFKgzBzY7GXG/VQa3EKSuI5S7+yxiHa5jwk9sV9JJJ3xfH7UTrPOXH0ccAtKTPJNr4fx02h
rfmwF5okKe5I07tC064ZAbxXmhYyjB6brSxEQN+Ht1rd36JnuN5KV3nf9Zm5FSSZbBrwU0lI4xiF
5RWo1K1bdZ7PnMVWNEdceLi14z0HZHhyysqcI8zMUTHBL2IUloBc9rFhXuddGP2o7hsjCImbw1F8
Fjm4T1TsXcV1K8zYCdUP/Fs309dFRbJwJEU6vJvUD6xNl3ixRMkCt1WidIVzC4fEn+plnK7REA6d
ztSr/0+Va5t+z6KyJfl0Bnu7fWsOPkO//HY389akIyZmOg368N5i2DJgs08668d0MILPdJ53qJl+
szpRcYIOQS1/+DSvvOyyPsxt1du/qq3txhieqgZWBkr5iiTalAZSnAwpByaA5Kc8FSsAD0CCJbWY
xLAtyKe3xBsrzsSrPvBLDHzxD+yAhH78lGA99gbVH3Xrsd0qEakXJHYeSmuaC9xWNU7nsWtk+0pT
NQA9Km71AT2w9rVqNXpX0ODRuwfI7V7sgN5WLjlPsWr758U1v2JYpsrUg0XE3nG6snwjXa+nwOBt
bSyGhuL8bxxQoFaH3ubIFjrd1EJ+iqfcr/IRsiZ+wtB8J0KVxJwfBBPEVdyr2CfmSd9e0HZjRONM
4G1M333i6WCHXulZeMgfrDSHtXzf2G6mnArk90bmwKhvP8rtkLr7cAQddCOVaOTIDr1ujTXgcMU4
T/ShWx1OpCz5rsRZpm9ergjDsQVk3uTPiy7oLgDbE/lijU1lGgI6fSGEzYTrAgeTRUOckypa3gxk
eeuqA0yWpKquIIvuvl0P4dtGfLqVEkXxwoThr8Hf1SAJjunuD0jm5unT/TgtTzeQJkiKgWWXnycj
2zDT9yT3EN0pmcLRv181rUWSjMZ2OlpVXFLGd7fvl6BHPjqwTfcf5jM9T513jXt8/kvpllyIEKvA
Gya8BJJdcuT23uryzOWq9D91spBopv/stCFQcZr4Xrwcb1JjgSe4YiYk7IcgUEYtMhRK3K0fFBLL
OwJ6shMVbCoGR9TvTQrm0Xwh61F4fJOyWIu4eJLn0tE5MKJbQIh3sw9YZB5pABsG8Fn+pOLwCooo
sA0/b5uprtMhBPMu1QyG9dYjZWsYmIkmglxTBtIzrz5AXvw0dZk/NIgQhTxdMOqhQGfqS3Ya4Gnk
kTmapq/zdsOePTl037CEi5ZQkDSUXCAWOELeNtTStBk0ffABTp6iOj21ZhTUBZGFExfupLVKbQKF
+9fxDVtrdfqagh7utn25Cy43v2RouMBH6+adTbd2xq1k9UdmXEgAW6T+SB5pOA6Op86V5V69nZIf
pPqWwlZHyTNIsBwJj8Ik8Jh7PJg0bivdXlZ0BCFiY8VpMRG/dFtzOD3iH6qZLU20xiLXZJiyM/6g
848dNS3YgFttpbADBRYN1JTOPKjp8AvJGbzebHt/hvfL6fF7i9sjFR3rzBLtZ2/Wz6xdOgfaAp78
2VsMnwb6VHkWAYj492tWfqJrr29SEsXWjnCMrkokALfeU27lXOwq1HsqTBrT+6jnsU7GbohoTFn7
wxRYHZZFZyCsuza53hxj497DQ1bNXW+XFQqcZDkoihst7VnntdnToK5X8QgIX68LfWs7O0NR4lX5
ZynhINLqBnPQucSKOAl2tUjbDRWTPmFUUIMQlvU7EmtkxyyrrNarCM4Q2yPobK84EkL5ZGmbBoMM
or6DaYdi31s/wxhfRj9rwbEhEURs2qoiyWrjP670nBgT2Zy4t75CHKuD6u2ThZP067sj8QQocZPp
6hEXfwjWFONBbWg2+uPjMrED22VAyNzuprj6F6JXHPgmJBxFWztsAQktjOuy42CM7DLw7FfjcAqZ
KbTinbuFBlYZwFJ4e42gYTvuqgGMWozIhjOsLMtzxcyQMAMbuAg70H8+AnKkUHCKz3mqmykMnpLC
uhFMww39TjNCZh+L2U93dSa3LK3DqRCa2rOkjA76Ey+9SfRAZk0oiKCpJZLh0DDITjAdB1N9ee+t
4nUIz1AzjmdaXKCai5cuYi0moRizfd9jAqs4cz6H7JwuQPLVvEi3JNsoN4EiWK05elrIOHmmYkNr
X0kf+0tQMbdHB0fq1Y3DVS09nJTNpUPxue0441NET1x0p5wUOvHIPQgihZ8H4iiWUGu5iUm0Iq7I
5ltqJkLIeyCxyPnBwaOz3HhOoQ0uFh8kenOK4E+KJykexk37bQBuSbOP92+JwC3LVhfq8g+zhKDf
7I6XygCUBXefWqP8RWqx32pebsvuiQgDIHfTLM0lOkNaSF8YjBtyeCv7QDNfD7INsEowP9K6hhsD
pB3MNtLdfMYiYtMEzdQkFZejsyfcO6o6BEz4L7QhU8qTAp4goZ3sGF36fS8GtzLgKEfuzZnDixz+
2DwEaNjnz6W5VnTy2YxXeG+RnQaXgRK00yHQId5ZmTxKPssMDiaRcyt5+SJqnAQ4RxDpwNpmUYk+
u6U2z7VHd5hF3bvFVGisAjnsbd+Ti2T+vzY+2lsoim+hKtyyaRgX8B+YxtMhcLqiubmkuzzJy6VA
866Jyf9Q5kkJ7Z6FIgFhy1cXPRcNOsYG1a1iVWMf2912kTpE4DzbRwUcPOLx6nd9YB2RkcpVoAxd
hy5LFP1NKHQp5ZvZgBC3lpzrztMTXe2VvQQ+Q+n5Vy8z7pRWwQGgJTc78zP0W87w2dYITPnp2Asy
WzCLfnUOrHh1iIE3rohBJ1sV+efv2toZ1REqSGBCs/d4bE3BSESOykxe62s2s6tVvQcscVmc0rPO
aG3HJZ6aM8BTLPi7lTprbEiMwgU+UdC/WK+E3VnDYTv81woYS6L7GbIVDWv7YDFeI4QfUOYhbrxR
rvLTLvuM2acBLr51zFUFwixGcPjBBo0Xirb0gxrwnHnNN4wELOu8cA1FmVOxAxqQ3xm64fT9i3s8
/CAjQsPd6ul1c55Y7xjBWddULrUQ4TOALH2rN1B+n4sHJzZS2tuBEQerz7uhxuzd/iWfrtab8V3U
gSKJzcoG/xxJlNHGUMmqPUC9mnHefvVMthgAomIvzpPUV+bvV+re5YwkZNelSxlWXu3RK5q1bpxg
GVgEShmgVvMpnjvaX0uEBiZDMPuF6Lyl3Bi7ZP0hVfO4MpP8dX/LnU9LgHIKDlW+K23LbZwMZNry
pCsCssia5yI3Wv2aBQN8cK2Nqs1UuQB9WrupILWpSgQRTf0CfgsgV5TNMd0pfFOuzA65+C2kizr7
ymbGRSUFG/VO+9psBAovyW0e4ty/As4B03tm25jxuX8tksQXmHFj6M32ZvBbLm5iNpsGhiBts/W6
kWXAbNarpTy4uIE5z6v3fmDO13z1Ysy3OnjsrsErxHXUJLB0SGAzVySBY6mC1dA0h88zcBnVnKa9
XAV1L8rs34SF0saTtbA7KDDqI6SW/moUhRJb0tzbHuKEg7/gYR5Cd4/VcsGdf3ODlYuMbajVbCAp
rJNQAMaJLN4BceqEzad/3yg32JNRtwsSJA9Oe+LuzMohauUeKbk7P83dvyw95wtbRU9m4PPKtlYu
J6rtduu3++GQLwJmAgYnlzgF/aLLI1QmOxRAmqLXS7hG62OMnbYb1qMz2GM6VB2IAPGUO7Edi+OI
4A2tMEtI8CBIhdfbOlIsLRMtCIgGqFrfso+FVKQryas2S8B7Ca2ByPTipY/+uQ8KlKAN4HkPD4m/
YloXiECScMSFar4qxK1mvWQMyzOqWlEMsfoxd7Cr/lozlna2PgkHckrgEnuKxwgsAJII44wZD2y7
juEO6DUtzv47o5ZRx5GI7Z9Q32/QYcjiTl9Hf0tCGfxNJfIcda9TNW0dr9irM5G4KAPbQWWLKjud
tXEGu8ns/w4CzSyP/7eriE4nAySa5gtxxwzf2BqNQ8WOmdbqo88yVQvElxuWxvbNjZUyH7hfVihX
3lxCUMpl/nY1neqjUw7q2g4dkOfigxIU1l/edx86/xCLmS71kO3hDHnxVZJC67GIbZlLbAgxAhTt
nSM+Z+cjHD4cwwxNprMbx8VCtqLwaE3ecI+nVb+5xOTrNivcxa1QSbO1G15Woj9BgP7Qdf+LhepW
q3f5LulI52Ei31cRwzfuY9xsRqpkwJc+tw6V8ZlynpeiGV395A61cW+hFAX9f80Fx5ImUSwnXy9v
cp5sv22LJPy+I33OGMVbhB16wl6ExseQkFfPPCwMsirlwFgIUaNQJU2OE9kfW61GW+m5/6dPnRuN
ZLTlCMDZycDo1EffQtMOdY2pJWXr0zD8yEW3ezXRLQoO1xG1eATOau+I0HT/SOJqPMrkCCtxUfEh
gVNr17sQeMILXDkTR0TcJUJwn6nigh5bHC+J5O1Zcc+lzxMQ8pP1CDRGOors6Db/TeHl59bRPMMm
ZxpnlPliSt8XXsyleAA6OxqH3b54k3VFOCRsLpC/Fn+87xf4+qQDyESXF7mwzfAoDaJyMp3r0Rla
jG40P56VvaY6ily/N9JcjxuNSLZY3mRxXzd765SD1cYfGHkKzmYVKZR9YXd/nr62AOVyjITGB3Tv
iyZo9jIKo+PA6LQxtprOJJXXyYrRR+MyKxDH0gcMxJb/KuzqNr48/U92eTyrYseZrTQPC4nrdKgf
QeH7Oytkf8WpSPEqiGQwInql8oQzkMVPIi4X6oTr3AQ2toWkpqMrXv1vOARmYjNJ0Ic5RhfdoUpB
vtQvPFGQRinmFSWD620jeLoSYAbf+SxgOwTJaNzrbjxHcXRH9PpqmsBA9i7IapHoQIJTO5yfHt2u
xH7PvQvizazVTzAVOnc050ucU00/P13k1+n16pDIwU/wFCrhSPGP2stTe7eWl/HDNHQXsqRDnJ63
q3IsVWr57zt2ZN0AKWM3Awrt5eeUtg7FYPFqy/hm/4kNQCUth3zMX4infe6vNUpjP3tUVxMPHF33
b+sYc0JoSv+CuhOwj94E2c7r85xYyQzSWVsTKQ/BXbVV+CQXsEx26sACA/ZoyfTyXdxuE0Mlayoz
M8uefNaJeANnmCZbqh77hklIPrCUpZ0xj7/wF0k0QmtOfOiEkjqnJRLVzWSJ1/Ds6DapHoXBbaz5
sttyPm6ddkd+QD9cnYr/YOMAyabDeaygBV4z1KZ9YS11hwbGGahz8WQL8JwXHfwp9UsauukhDRnA
07HInhrXLTRYlsaIVqJ/YoFZzrcW1jT0LxL0JxCtTzmwhVGL4nERGnhugLuQYRw9MXkyCrJ74kFl
u2wxjH0dSReYRiFLeC6pzV8Cj08ohyTy4cOCN2cujfbD0MZBLB+lpk4asLkhGUvZsWKtTzF18ONp
6yMar1QQs8Hjai/KjSD2s36li+gTb7MS4sGEKOn2nHNKCu+08xoI0eKPw3B84ONm8Oex6jd+bQOZ
AEs3g6P3ca+tSCEfu5AUCSueO33YtNSV37zjWI0QRtn3fIgEX4hiBeW63+JVslzftwJwVYyR2e/D
j8x60s+Jvs4P32yd00TDfN1NKiIojCYcwUE6pBdIr8Gy1vT6YMlV1V0HRH0mYK3igc+IzBTf0a4Y
wiYEvOKG73I2ZJkFknn3RREGD7WQzcyosruldpUdMXXqAFosFMEzHubSo0yeqRYm2LxVhowhloZx
jqf7YY2drPL8BEZVJDrh9TWDtx0nleyvzHc1f2aFcxSH8mGET/uvxCdAnESDTRw1Up8YeulBWLrV
VrJ9ZGvhmFGEUiR1OnjlAmaXQcWf+FpjjDfd6EPWqppViDxhd+BI1enTQtV38/nQs2Uq45mcdgHv
Eoa2iBkCrMuEDBiDY4Ty7a5wAOI9YA6+N+31kXjtkua3HLkNYBXP7BpyK8Y2jBcafq9n7zKgsiBv
IvDA7Ymk7C3HuvpfUk5Hv7o4YhegsZBzslFDhpIVeHWGQSkYpuwudVRykWeAbnhx9Gig/Y3HFjQM
N4soR6xV4cVWyR5abIR5YVP6Ghv8gqtJYvqDUTxgWxN/BMOcZU7PBZkSk/dQ1r6kvBI2Rl4Gonq1
qPXHRzddl8/mhirT9d9hhyy6gut/htohCV+MUVKQ59RKdujlHHyfR4i1Pwidt/3l27KIAeQBqITq
tHTcVvSkPwfUXVl06mN8+Aeel+vAy3FhJgCoZrAiF06qBUAgKVth2uOD0WYwRsjx07pBpLt/oFkv
y5ukwcfD/FnyBPPeUY4PHTP+gY11789fy4N9rgYn2OMuVbcRLrGa6skGDxOFJRmcC4Uz8oSQ9vPP
FBF9xf3uyBItGc8rNo7KiRQ1Q0Gd5wapuPq5DTyZCRlDzFQH9KRxIgNVQnZz8x5j2ds0Jc13dKDC
Rh3w/BbWRSZf++U8Ex+JJazbQ9BzWktDtucCrm+yECfhzPYeOGmgs3iJZJuG7lX3ABwXX+WQ1HIR
FZOaS/sIsWOetgowbKHf7ZJqaGRyD60bOp3UwnyOJl5jn7fsB50CIf8kgltIHo40YPRjkmxdRMWI
Tp5WnmkA85rno5HeieppKafefQUQpn8dwTtK7ucLw9ffW9KYXw5N9ijj22w9iWt5NRm87gP653Cx
sChgqt8ugbKO7gK7J7QDmL8RCdwwO6cDzkjJkLKhuKQkBSHZLVK+lNJBZfHIlzzF+R2nUMJcH0oD
01Xm92uZpC5mKVY2Gad1d6vvnN/I0IOtMf8LeBf37D8QH4YPUtMYWlHL2Vz1LjvG6H/XNCvH+hgq
5Q4uW4ZaB/kl8Cc9NievVKt1qZO46H3MAnwvTiYzLMpL55p0e7Zin9qMKFzyD1FkwshBKhBNbzBw
8WBpkHcr4D8vXCh8S0/OUNPz3MLF2qL78dKuZfVL/aBrBe+jjo+KpdPwm3WaXLRkhGoqjgtYBJgA
T6aTSkaYwHoPfe4wHL5teZMok5bHaPvM4f0882oa9TbgpeU3v/DjUE34YdHX8WsG1N0KtbCFs2u0
qDzW5ugZHINrQM6PfpV2KFJITE1YXytSbtrLBDxTv5E8RvP67cYsNLZVh0ysLUss8Onb/S2QMQ/X
JgZbtirhkGXna6+7FoXwwXTqrvh+qo4+mbAzApkCWh6OTeog3uuSEdTKbk2vKNaa68A/rmmW+tRS
5EKAN/5JureXc19AcyaGXma168yk/9g/6qSbuvSmatcMpHZ5P6Stmrj+3ufGhVajqWhxUyFNUzom
KBRAG1wjdqbu8MPjCGLtlukM94vg9AIgw6V/qtYY+l13ekUZDa+11A4CLivE1IMUZVIwYBc76JRb
E5NLv/NK14PRF3kUbOC0PNxxun4PDLCWbYtyYABeOaTy8hGNm5O+Zl6qr0EIywri7IFyvt/Rjg+T
aaWzrg2S+ELGXQvqoHwRc5w3QsrUaU+w3u/6Q9/jPCbn1VMvCpuk7NNJyEIaTLg06Mm0aF8Oh2a2
3VsW8zy0nkH4aiQhwOSchYPpOf7o4WF+doNfGAlDh2ZZB4OGZOTG7RGpYhDJc77cuYWmbWg27RcH
XJNT/NeiJlZxaAQSIilHha3vW+gtGd+qn8eTbIez8h42qfRPyN3CKGpSRgMSbXo8R2m+nEMRGP/9
0x+mRqfHrrWVGU38w/WzEFgRgrApZ3s9oFXSwMrvsau4RYno3WMWV20PPnCqMezga4clMQi68uSN
C3GyGSxGzsjjK6T3BokcGYiMshWoheZHw9yYCqgjyqEAuxmzfHuRYs4LsojPwgtdwrfKLwdJ+0p3
t7LaAmKKwCBsHCT70Rh0zNipvqYtX10PntQDVznC5m+kGwMtieNRYbSxCo/9hSjiGZY5kkAd4dx4
tXDEVY6bLIoEomDg8Q/J7GeUuiG+7hO7VV2SG11Yq7BHjEfQucpdSFIfegQkP4+MtenD0BaZ62Ol
UzYcP1IqWSEn3HS0aXX8V6+AYcdkloBs9/GHZwIKyTchnad2eco7C8B03k9sNM3jTQg4lYmQkGVG
+wtelQn8QN54vyYuqa70K91fHSbocV6TdGFAUpVyLZV41XtiqP3JgsbwxpHPuiomEBaYAIzex+yx
JQj/oMD0C44qrXrQpex70eyFGNHP2NP2mnlu9nf4C97teCnwYFYEM/HG+DfZ+MxCg4ifdeOPIyEw
JCTwKXlFOxvKSQqcuoDIudE+Y5X0a7kv0w9FUD6pcNfPEtUjuh52iYiKh3b99619p5rsfF12jhmu
QbzqoP42Z+3PT+EjhCq5HZtmodlboUndhvDQ5uFjm/giFfM+m1O8E68XjAelag1T9Q/aZ9TIvDhi
b7xrNP5uN24SYUbcWMy2UkTJggsDhzupXV/OLmt6FNb1s4kTud/VkeD+/j+cvfRI3uCXQY/bONdy
XT/uvkT7Imv150NHJDgYa/n64mpVwdZIuhktJzizSd+zyEQYCwzLzDtuumDt6jtaJvfaLkEl4AdE
XKCZA9jAoh95B0FC4UZgBTtH0hZxO7h+MTOUdRQtyD3SJpmTW8bw3GlPaMSDjPAnKHMtyY5vusYH
D5/HDa9lcDkrffgbqIwrmzgIYR96aBau07B2nM8iPP7da56FHgjX8p356Y4i62hDDLagXBbm0cWl
VpMp1k8yhov2gWNPUblTGrcxHr74niKQEDYEcl221AkSjS+DKGHUbu3zIQa9Tl5X8IAEZsSyDf5b
CCpbpcGSCtEtngWAXzKgrdl1OU94m1+ZpsexOEjulyvo6vRd52NpttM+vQZX8BCvvM/B9tDJBNVu
0u5ou+h6cqG6bhNZMF0h2HtE7ZExMLkX1074FligtjC1rbXe5uSvjGUJ/C0BSydXblY4+Zs7zJLV
8H6RUpDoerZRoIEbrs2na7MLIAtcbmyO/0v/IXvwQ05OAdHs27BCQQmauFKbMD2gF7/CwGdj7xz4
e1Co5IArF0dAHrAa8Mr//WtLMZOgCux+Z4CC/sX24BX8EOm/xzX/CQuaWeLqbc+zWPwcy810b8qq
aK/RtAhK+OUckrk5NHEQoNgcE3y9MOIXdZjSlTQ9oMt1X2CLtQvsJXBppuvN2HctoL5Wwp/kuVBL
t7m3CvYsrn+xmj85bC3rIH7m99+WDBIDqAHzap2U6LjX/OVGGWf1kR41LllEqemIqGiG6tZqR4t2
CugABiKtz4bqfMzHYPW5imrmXI6swuTJCbVdeb4AWdVVpLfwPvamSe+mqubjAFuV+klMEBpbY5gA
/7LEcxditxDK+G2RO4UzjoJkoM8wRY3D3fwzw3ny9vmL2IdMVfdN12iPDwwvRezc3TgY9Ytsvq+Q
tCSa5cIq+duK0NBfYTJQ3+YsHDSFRmiVTA7v62JFyd1iNfWJwb8FLQfYukwffW6fDJlZFshvarCG
V8MZEWIDLfOYJVskhPuXoXSJNl/0g0pPLoYcPoTMBG1gLJLRgPBYYCOttAcZIXxQhRitR4NMYb5Y
5qAtcdAhsSGoT4DIRrdeddLoE0lSpcdhAADOqYcxS1pc2c7kWL/2QFy0QBXR5/hhPqI5TaCD6Buc
vlyhj2WGAhf6+52w2Q38ntxJOop8E7iEJ/HPgabE0jeYSey//6ytJfVC0N1b4cryQR/l7t5AVrvd
jMkSVIW5osW1eezxv7TaKjmDPgaQBiIOyGt/US/jA9MgHz9I3m+LjkaxTaeduULgbdRSNP0yVB24
IL/TG6+/4QSKnkMbs9BjAo6xVOhp/YnmM3kU4vbfKb60mDKblx4sMlZhfHWHFX2KpLCjnC/+EDPj
unXuxiiM6Ue3ff4SxTCNATdRUKO3iBTeSUqpuujbUQfEh1w0kU0mY5IkPVDw/Tjels8iFglOjpp3
RK3OV2/gZFvY29ab5o3D6w1zW6ChbUFp73RloXKGeAr79hFoncmqEAf9SCQR3bqEycouL/rjig/h
cOnk18Rz1BJkm+uTtWxRw3gsrhz8xqWGgRNm5+kSZ7V77ByY74aZ8BBkFkLDPHvSwpM6DgF3DvIe
xYvcen/q7Yx3TRgmbGONE83dtXwU0k8otFnCPT2OYp0HuA/2x//kN7z85H4fAOM6QNwiXOBNp3uK
ZZPaKWtMlCHoNdQDA9Nd15BMZ2NvXV19fiafNc8WvmQe9vkCJxUCvhONc+f+SZeTe7XDqltA91QM
1k1YbI9LD7RKPcbVcphohxruqaSmkfbXQC5ruCS7n7VjKeA3Hxb+LGrxoxveTPxmsd/3qjmtZ8N0
Z8uRoQB8xD2nKgyZd/jw2mpPHA/Alugrgi93VdxyntNDpiY75rGatCFI7ponM0Md0hHeuciboV7g
LMKK1/mJIpVrtaP2Y7ihq0ZI54U3akR8x4HvKpYWERTfK3nYTCViMlBp5mrUpz3DSKgjy1HDYsG6
YtNH9kCXw6/Rqgr6E7h7l/Fh4TwLBMFImV+NAIHDpjxkSF3+1TkWUSyQB7VAcqEl5bucj5gD6ZgC
3o91V3JwhC/KCss5w7x1zfWruKLOYl1Q5Kq6vBbOrWWkv8Xvlcu5gKjeWxhPwUir24d9yYfyQwqC
yJ6VRRDouO/HgVaGjDFaqOoGQEYqDNG4noN87ywYtyks0NMPh/7zd8ohhPzBNprGNnK0au3ikaaY
zp6uTGrAWvve1VL3vkaVMru/449gxL6QiGgtxCSHGzRtt2SpeF/gXbXKxQmC439xhSCtbg0k/6PV
H32podl0AmI8PvB5QqTl5gX08L/fsOF8T6DeANo2WoYc0SgJeQW/jSm/KTFig+uGoJnWLcAaQfkC
MrsKghPKQ3awVlU4QoZh7TJm6b+fgABtvaj/8I+ZRqmnwxadZmDrkpXrzsBLAvnkLJNH6pmq/rTv
0xJzqM8+K85qsTjkd8QILRFiAnuS9wSYzIz52TYl1ozx+6ryfNpjFASUrE9SNil4DFTMrn+7i57e
IbxtXPDqrUEWHemwEKPNqOMLUNg1Z5WLSodIkKSXwKD2M9IQDSieSPNl/v/6M3kPtX/gqovtbLMm
WDFAv6m18IOcC9wfklNhcDhsXKe1NSJRrF4hWVmDIjfQoYE2Na09IP0iOf8rsdRn7grjGT4aDQFT
EDMU6mYcYzAoBrWzvreQGIcbtusANNixdR3lwKubIVAmqXTTIM5x+M07aU1umY6smSkunTe2sdR3
2Sd++jVieCRPbEjsf1QUrJlsVzL5NTexZs55Sp+JgCarIYkY0ySawiMqejJMxsCBG9kCJwHGHhKV
pLvqmfx0cCQuZ9Q831/avZ4Sm1iW1DzfWn1u+0DUMn0HsUjS4OLX3Kx+lTeojQpqiTCSBL/zaQem
Ma5ZpZt9nHU5JDvsJfvqEgvclf6Fm1uKGLTf7b/4o6d/ofMZrX+RohO39NXDsJ07otN2bsWDyXGo
yR6Y5d+URw2ivySaZOHrZx+fgV9PtTiquZ9VZoMpSZaSWgI36fd/q4f7c8xcDO/e22IOVCGw2xBC
7kIx+UJCX/MhC8a9/k//vk7j6b3PCFOa1D2XeUyCOng9fR0kCjOo5tI8MAyez6tobhtVVSBuxM/j
ZhMgKGuqGGgJsQNKSUJFwSFXGC6cx1w48Ft4slUYo/4AJcsB28EyMTyNkEjxaXl3PFPAFa4ieDzc
X6JZk9yQ1iicSNAWlD9L/pEd7LvHikJhCyVvovT4GTNJcpc2BKpA7t4VRUuHQ8iBJRuAZOCMGi4R
2zJ8pe5AsPEGZQw5v7v0rA1XGf46/XtWjiHAOaJvhn2QgxdobmCjV0zRA+SMDqfVpan4MwU8J2av
8vJJwHj/Km3EGWmG1cxos9+JxZvk8TRcjFx0K+DDzrdpnXIIugfisWF5BOhqd8uIKgfCNc45DjKy
q6YVn8FSYme2bYY1O7Kz5pTT/mVX47m+NZoJwjj8W2pGUuNwhEiCI62WgNUp22hHA9CKB67WNZ0+
eZ+yBM4Jleu0s6mRIUFoC1ypreRkQxviKvTAIeF1qho//a6QVVlNCEs2e+F8N0vtq1zQsV2Tr/aO
wtPaZugsIRrN/4/0YqsyVRKMW7YCT4e2tGPdmCWDndpnWpL8tLZ9ltGtUYyL12w/yzq4H7ypeG7v
TLyQjxA1QUlQ2MCxhHSVLv5mYELIXH2Q7FA+nXhg2pnUNuZTs6SVmIhSrH2oW/ibzTKw+Fk4RX5h
gYOn5LAcvEYfQzWVhEWypF1YmhxzRcFUoiiUiXwHxBtbQgX0GZ6ROhBgbmcOMI81CEpHGQj/OS4J
LYtbFeyCvyn60KDOgzoa/CDfH5rOOL/aIlCd6Jn4SNWi7C7/afXyNaWax248m33YuOeeRPKvkuEc
QHt4DcIqt34UpjKYR0XKuy/2unCbx/bt59Aqy1BEiohXd8NnRCfkhJ5c2XsJ+Mhb8nrLqVsgwSQi
8B1plC7GHpjC4ZkN8C4D5d/3VNBRDHFU7KjDX6s3UXL8CPf/3eibnl6QDNZjsCgjbXYUQZzoXqiU
UJafpCryK98RlogSS6JF5jnmtVnpEdpvbJTj5HtH7A8WeHIpYfLIuheX1ZdYKHRQPsaV+n7Fxj+V
vsuhAukE6K2YahM96BH3tQTA8frHcN6z3b3XqekXVa4BWTBAsPyWZGQkaoseQHjWsOh/pWC/cxQm
5x9bIwyEh+IANHq94A2MECh6oynmRGFAChKNrQJyoieVyByb7R4WLdJNSnuiERtb5JHVad4mfQPR
auZKSVeG1A7OTGIYNKANmDn5Mzt8yV4fg1WgfiHs/hlPWoo7I48RiLOP8pIM7tHcUuMtDjEn/poa
JxMYQg7k8DwZXeD7REV5uPxymWlvs4WC1zeIKzCGsfUk0jXgJhudik8h8LbFFpYDgATDsmvfS/O2
55BQDwxxLq9NhS/CcvAEr23Pnp3LPuVoXcH7lzTihX5oLhK8e1OK79UOuMSPSnOtFJ9TkvDU+YFW
QadeDBXqthV/glFWZL8Jpb+jPYM71Odf+gJYvuw2sYL8NLCOS1RI6QNrORAgTIvhxXsbp57Y5scM
BeTALenWnGxX2jnKTOr+Q8LxgNKb9yhpjU4/aw25PIgNIHcT9tPrJGSiW061juDLKlkNcNvlON7q
UJoc5etEJ4tafrGVNEjnttuhT7rDUzAM1ncheUsqT3089JqXXGgkAGPRWWouS2amKnlXAq/g1gwy
H9SCutWCwIY+MgpTLIoNXvC73Hu7OpnmWTMsyC4ajmPf6fBzyNqUuh/iQnEilCL8yopXNBKTmIb4
OZG9kwL2pfvm36CrNAfI3+QsLdigxUFR2ieNFYms608Ul8Drug5KUYbkF2guLMY3XgtdxpBZHTqz
9lbF0pyyYWVsPjN3EDwPi2Do9053DIQL09+OZdtX8bqI3vvDvDdtXHHEwrSALoQOvsdfff8IUZEz
3oODdDXy7WjXYdTaUOMVHUoFQ2hqqoiyIm/npIdZUm3H1yOHSire7ZUvqbqpxluROSB3H89+kCvi
exSkJxS3K38fuyyQqVdrIbSkO2cCPHK9xpBmjPef8v+TLCNcY9h9dZoMu2zgjyWvwmjf/2dlz73D
HyKc3UtWLw7/2CNrQN9fjO9L4Q4Vjs1/1j3oqtBFqkIV/lfYh+1xBcIEI/09BEAhARk6SxtJM5ww
XULnLHnn7KdkeqXfsl1mZXRE+c1202d7RhBMNsWoX2LubcAOTye7lMsKS298ENkFM7ci94+dU65q
2qgYaN/XWGPRtw+k9qYmm4GLBpUdjo0zw85cqy7SBOiLjr6mL6M67/F+GKTwzUbOM4pTUfwfWpuE
WyfY3eioTSlY73p2jOLb0t2Tq/10jDeWCs34W5v08MjeoMUXY6RoEDPOFYgZH6DwT3yJNK027rwK
uAGxNrhb6vPIiyCWItU/J50oIlRzJkgWd91UNFeaZoEI/Q1/EA4VDQHQEvOcMin0k7AvgJRlqsn6
ZjAWIKUgsy8zuo+V6Lw/TLBV4fF4wQHmuzlXFT0M0OQJWsu2yh2mS5GsNObVmhbblVZlHdhGCP+r
NMTZxAIA2+fg02DDJnk+EPx36CQ2G9WuTmLZefrnH+NuhZcnD5bCdEoZ1hFUnZY96/kDETnTcmWb
cz1S9wiY8AflNdPkH57jw6X+LxH/gee03JohmcKV1Y3ro2sUbqrdpaKR3SYciRdcAKhUKtTJ/xVQ
f7qu/t1URF307zJdKppKiRBIYVuniMsqs0bnjRyhLwclMTH5IXhEZwdBXUPAuzkfpB34+hkxZmv0
TWODAYiJO8Nx6qg6GpNDYYTgSgsXwK8hUiTcHPw69Ca5LpZd55g1SwezvzhdM1HAYvrrd36x+1OU
RPiZ9u2/CvLVTqwFpuxA7gLGqThBgdMk3buw4S+BrrC4TRbGrQY5UpYbb0MpFNEzW/5FHX/2o0eP
oiCYlUCztT16a08kgCg72+HLcM26iMOWMze0x2S0CArCcrX9v1MtQYA7H9Gw8PlR0pkC8wnnLlp0
1rQwgd31jG7VZbfbuSIgN7IhIvdQq8lyImuxF1rC29YSgZe+57YVxo9hRKvJ3Thz6wS77wCqyp8l
pNfnH9UoqUYYubfQt+CHYspJ7qcjtw1TogsyAVzTUf5bhnY3ymafPPnU6FZh1Xea1MZ0A9tw7a5m
HOuB/BIjyk1JSDoUAExyZDIBuOxf41m1Twlnf2JYP4qw7gXPM/N9sSeUbvClzFEYm5DQJULaD9td
IIEbw9X9Z6gN0RiJJIH5/oj67khXUY6Pq8uZXFRkQoOckZi5u/9q7PjSQpYIGFP0yVGbiXmsTKaz
tAiNVqS0mfn3h9BR5TsBl6Kmx5EXEgRy7+7n3hZNkcUEQpUbkwLOrC+q6l4BwoXEML3MLUZFd2Rg
MdPE9NsHGORnrfyBxR3nTNRHWEGhZvJQtwlxYNzXa/fjiwJBJYkd0iDHuI09/j27Eme2+57U4Fty
I2bo85xsm6tL1yYKSNL/IMsWVYToWdGBaIyjkK5frOLiYtyAadGbUrXLQaEuebp1Q/BOEiwcZ5UX
v9pVMlz9Q7CtAm+w6pB9RNPzWa8RY865MHLi6/lz6EEIsQGODPgX6Vx3trNSVSCLqUJ2J2OOdlah
Hh7TCj3RYnFD688jLCxwcxLnrfqEela+EtaEkIL37MK/QkmdHTUmhE0xALGLBdVjNBSRwSk7v3wJ
IdfeE22R6mVIDSgP1sirJ2VLi9sfastJcbY5Emd9UTTNajecNst8oMQuvUnn1wdGxHP8WshqU8k+
DQ6UN59zG0o0zKfbNAntU6GzBmpXKjUajxiif0BJ38qBaekXKSQnDpNJ+3lA4BNNaHUtAy1q/dn7
lWZNswZavkA5OQXCVvuBoUdkq0wvUZZNfDhOVaboLSJt34VUTDnKuZz35Q8/+OkKsfiRh76TFe17
BGijoU+K4pxXWFnPH0NWIZVQNobeh2twIHH3+4o5vLwRzRVEqEm0ykZRPh32zIwSMqplnvlxVDsL
QnegFtx30fLDO/noEefEZJHYR5bUM6cu4crf8hNKa+Cnmlj9TSOkO4eMhpqnLAcnNGI9r5powv9l
+VifD6d0LOkmvaXHJTy93ey/Dh+N+hBmLM8FulZAC38SxunBEG2LXk9XnSMMnZRvccoFY9/VXTnO
dOmlw/wqzRr6Ot84WhqlgcQJ/3GdxvVKbrl95Ob5mDSCP3CkDy97PaV5wImaajL4KIZJ/ePl1Bv3
s97ZyIOCkbm6TGy04WvUUo/E4g7mViOCp2wqY/OBDNMmSO3XeNVeSiKWtOeHtxQvYy3wYaJ/waLK
kjDMT3Nf54xVjMWgeK2iR/mK082tZX0Zxhd6Ey85fhyvX1qxNd9+pM9S3WSGC0+2q2MEZfxt8DU4
JjmRoRioaBk0Up09nqfoYqETJCyw5+gQPZvnWeG8feUeQsuG53puy6F5ZgLfKlXxnj01+WLMZmbh
Xe9Rfob5wzDL5CTYHfjH15uVDN+VjnmA5Z+gKrHFyh3KD3E3Qu1K0+/uoNmW9B5FaLcsGphfpOMF
1A5VbaRTXLLzdH67c2FZdSsOrRl8/uV3bmCEUfBDt3uXaQfkfjoHJdqVeq/FnrEKOE/ztBgIrIVM
l26ajZkCLktr74IH/0CbjXB4TOBhpb7UeW48TU1wkNBktQAdiEtvwUYrdVTL8EZOhv1IK8Zv4zd7
lRu/FHNjgoqPtIWFilqBYmIhZBX17YCbTJdyIzagusetA+HTwh8FexG7G6eIFY0+1ObIN0Kt4U0U
J1vpom4+0IJzxBx55zZ/ZYOv4BQkvRCzy5I5hqZbYM/4fny8iJ+UT0YykBVRJbtln6gIOIiXAaqX
9HeUwC9aNvfBOpVlp74fj9+U0kD5btjpv4iIFv19l9b+owAmeFXiYfvl/sXFaB6j5ghECx+Z/Eq0
OStLbFZHuvWA6MZPGtSorQg+s/3wI5avbdRwyHaU9CNsyESkseQsrwKwFfn17Q2latJq0vmX1Zvn
BR+83WTQbQpu6otR11Vn1vebGa4V2oGsU9Uqvw0kSCFtf13WLcneBRk+X1OTb9ylZbdxkOQvGHIj
S1aQQxv4JOGVvZCWz5/Hjh3vGoCdmBxn9976oyCi3I8Mjfn6xWY1BwLn3AIEMPqzQEx/qZZhpt3A
XsX7GgXAdwB7nGGhlty/ohxFBX7arpezDEiyZ0dMzwnzvAlsN2ccnbyEDWuR6N1Lz1ocfkeeouY+
8NuFZLBjNvYDmhLbdhJPtescQhTW4F52hVAPD02GKCbrAGMpl9Oz6tVXK7Ica3aY3voGQpO8Pkhf
Vl2Qn5VSlMpAcGkSCxultiJLEq5joH6pfYKXrRBb7hErQ5o0zmdMNsgu7PSXA2lIgBhRRP5ovilH
AJqjIjYyCDypaI1Fns3BfF2unraMEVyQKRYjtUtFMIMttfCKwGWLvG6ZpOSfXMZVPAjYlJz3dfmy
F8+9Xgwet7TGtX5JKvJXdhOnMeEGeH9CqmUATnkQJFWfLDGEARpWSW1WVyNm/poY4oOuEXwEpox0
n/4LXBcfr3rBKlfYMn9RoHhxSraQvH6EFtTq4fQxFQAfguUilqgXxsuJawSqvQe6eZtrcCTgLy55
nKGyFfBgK9DLu72Q6t5SxrrmfO4634ARoAgD6IJDVStR51yk0cnoP1b+JCrgOvjKnzuispHvzGXE
gTQpMvAPuG2e4xFdCbLSe5vjPOQFIp/coH+zr2YjVv1X0MbfmYj3r5LH02Lfg6UUi3YxTUPgVzzq
pQvKwiza1BoVa1QKAJcu1GnTwqM3ld3Mbe/p5rs51ZwDHGpHPgRrfDCdzd4FkHoif8R5pjziP74J
4Bh3bzqnb45mjukA8S89p8L3INLBakLRuzdyv/TGGQI8G90hAr0gWT0kBDSfHnLryc0lvk2jDtuP
xql1pQT9miCvJk24coIuI/5H915ViZUAm8fbc2FXvAIelyFphN/9WtjzptyHpyAgBQfkQsFKsh5Y
jbMMQ4Z0ItTt1wrkjB1x75qp13m2Zz8nFqHoLwkcAXYUTUqBBLd3YUw+itXwYr1Om/UIl4YbuTBB
OgRGQmj9fsrT6yo21Qz6/uDIkJ8TSJOKo9T++vEoKojJz1eDmwsXTxK8Gf4GGmU8KKbI49CaUFP4
jIjKwcOEjNFF7ImA6UpGPh3LzcjCoIE8MV7Hp2QIxKH7l36ClNm7U8VB28YiVzA69rbvt+o/CmLg
gxTmjz1RyJ9EZdJKcD9jfXy/fbGgMC5U/g12ZutrEwPwAGsb1f28jQvwAUNXLjv/bX0xyhR6rPdq
/Dbsk2c73r0l3TzRy53Lw2dwNdK70L4bD4+HY+/xlbZsWoLaE5UU53Fb3R+mUd+Et/PbqowEXcSu
HxAcMUpqgiZVswmWJ4P0b5wdWb/ur5Ya1IQHBPVNKpooFDciFtWSUv++nhRaduUBOVsQtV/NXtYK
xrHsQOWF7tHF/HF5dccUHeORgWzpO+eLXyJurdlwf4g8IKqwyyN/OLBO0kidz84R/s9Xk1QYxFLC
+2Ymsszmyoh3jQcYWSE26EzQ4GauQXuJtHVimrzGfvomRxdCx8yRps5sle/9iO2N8TKMSL7YeOSU
L/7+pz3Ur0Nom2tb4X/g9FLRxUUzan1OWDAILOo4mZ4LaxWHGGbFshM66KXkd/Gj5TYI7IBipHCd
QwiNIWqPfPG01QRhnd09etX8xxOYxk1OdBWk+0WCIi+KXZolExFc+IgnGi539VAs0tDcWIawQJyg
VL5KHRgOmD/B46wcozHuekzwFmNbTEr5c5M4hLkKq1VBPAov62tSIhti6pworKZNtK8r+36tpZyf
COJB3nMOBkcy/no9fnIaBU7+8fUpSQFXOwtLNue6rqZJUhbTkJZgscLF+Xkx8ZXc12qgrxgyJ2Dt
eLCs566P24DftMGIphQE+9310wEu3MtBPR4junG26Ttj3KtlWTez0uS8KQBm11DeWygIwIL62KMh
G4rydgB+bMo3Fs4rBBwQNMb0Fn3GZQj/AGPMEHfslAUXlReexZz9AmsaFsn4KqNTP41kS+uejqsA
+KjNsPF4mgtCZNlIrIf+IaC2Rl8d7gbs+sJDtYWW8RDMsiEbhyvr8Q7DM3K3DjZetJxV9kLNSQyD
8YwPstZqyZhGml0o8orM08hfuJLx3MGAhLQpdp2Yxo5Wqo4ts9xT2Bm3HLA3wMI2S2r/XjqdpS4j
gm3LbwcDYzBmN96LRs2S8MbnMK5ut9cr0rDAue2CTyRcEIzyMulQP/3xVXdLcszbSvR4+NnxaLYj
eoxdKHM3koR5N//btEgPrO151yLkZwLjS735d6MZD66fTPP7mY71Awag4TYrj7vGg4PcrAwTQiLf
myv0Sqbb44gQwbs+cTfBCgKEXxLPTNcm1R6qzRiOJpspVhELg9HwBCxrQUlrb8dk74Nt0SsA1K1u
kjdfk60A9H6Co4K4K066pYryNjY9UAELmWEF6Wu/K+NXm3pnkbVYf8Lvycy7J+rPye32kcw+KLeq
O5GG34dL762hYD1Fmv8R4itftefwghZC/slauDdNV/CDWSE1CgJDvisgtQyCf+aX3yBeokMNbEax
TQk1i7BRXaWqYGI3HZx673gJW1SJ6LWR549h9TjHi85f7VxB3FnX817Na6X7r0ysf7mAr1hZFA+j
CXKI2WxZd1uO22VthDxATG1Nuy266VmTKLuuaiYByPipAsWcIaSS8IJkNTLVBGqZ+qbPiQv6oSsM
OdXCjWVSpni7G2/Ok1gH4ST8eAgVSBpEWr2h450z3R/0p06U57ITYGTayJ2nUGaiWEcFqZ7oJRCT
YG8uPEf2JPPTVWPanlZn9aIUSDYe5JXaFBb867OWUFnHfmATeHVRMxrnKU1gWBHVo3O1AF2XRO3b
PUoSfxcDfwmyVViKrqNYe92Jgq86StN8JLUrAtpEmZLcolBEugIepr6n78NnQ91ACG8vs9Ua/Sgg
Feh8HZWxzO54cvazSNfrCLDObbL5Agpv+DFrkynHHUMr1N02wDhKXmnrAcY+udyisHUJDr9XuGHd
UBcicX566iRnOzR2DX5MQ9N3z0tR8fYrSnvndGsM6jEdwI4konGrwdiYwWMQlLvVoz5LFwP3/vEK
2KwRg4aVqH8vgl+8XUDFzyAZ7guutnh79usPF9D2LUI6YXIPTc6c8Oij18MWgObxmuaV/K+sxNDf
r4yrcJYmO1Do5LjwXqLagRMYp1B2BRP7W4Iv5+drPZMKxMJYCW2guzKSpq+okyPOJqWxDscdek4l
QIDhPcgV0X/sR9fPS4lHNGvgXqwIxnrwD7pB+cPi7b9Ga5LI0u1sxgHsq4PJZQI9517Y0xzrzeHi
Gcfqz+cxSoRF7tXQAElZQ1cneqW8OEBUmjEGjPUhJHgnfXkeNWIN1uq8CqcB4oWD7eAakyoi0ch1
CyTIc3w11qng6Y71tYwK9adfn/Uv6fowGiOQRMPFJw/mTA5BchTpBmos6legI2RAflJNl54fwQyF
9TMvP4DBd6pKpvJ7KyKRIJhABqZQebjk0PW7Uk5d3i+W5LknHZicn+D0IaIqNEHJtXS1A+mSwDCV
bEYv48msLYxiY4Es63vhb5K9EVWHvrIC6wOFocYhGUT8S5DK4TmMVfbaC7Tb14BP4k9SvEfk0a5l
UTb9VsKkQhnn0+QUcN7pLHOeScowlj+mZjMSw8T7A5/ThkqGe/v9EaqY65GM9FFFcjsHlF36C443
S7UQ0BaLEgSmFsaDqPiwzUFGwqUx1fLjK+/aeqqg/DXi498oL3rdtwUoWzYRZeNwWJqFibF2eRJf
UzGgRniPSN7k+Tdi/DC6raXatThecdp16qyxYCUV/rV487dlhKHj8zXr8onjCpSR8fPHnI9cokjr
7qMWlGpJ0zPQoKZNE6ANGVh7q0Go6HcGX2voCRNWuvHzrnUa5ZwkN7lLhItZpDvHltn0Ep5yTaM0
7+U8vFV+tDQAXwN62VNH8XP4Xcb+pr75kWX1QryV6ElaTwpUNRETb8gSPvtNqeREHhI9AA+r56+G
ORpHGMIm1k2pfpfh+B5TXVF/1/1xQ1fXkBDwGP2YBkWqCLlYGaZi2A74cDm3QeLKX4a5KOhiKT5l
dgjMDy2aGL3nXCd4dNTOuqsNql35KdvimCiJLFIv2AU71IQryNoZWCgG8u+q2tA5IBkAtb610pQx
EuHym80QJQ7y/0lEEXGFK8QjATvSRpi0r6VV+U2xM+wM2QMfpYC0FMdmXIu3JbBUVu6Zxy1eDlOk
vPCYh5hCyHIdCkiQDF99RvCyCpIjz4BS7Efe9kdT4WDGssWkklw4LSTJTJqqT2xbK7w9Ku+ypesF
dEeZHlqoVTMojMKVf+PL/TV94/XW01dYeTKlU8U9ccaRMLuy9+3/ymEzcqtfDzmYXrVPOd3k0Lkb
8sDi9T004yqBc9e5gBypwlg4Xdxdb8WZ2u2yx0FZkYd27lqiCMNnpFd+e3RXbhRh+xecNQFl+TEX
l2q4UJ4gYXDZi4HFs5Jw+YolDBbh7WYlfnNGO+ne3uaxMOxy0qgbL/5/Y+nnjx2heGjp7bPwQ4xk
TKgJmIWfmsf8WJvyz7AKWezZ8HeZ1OU/p3k6TaGiOXeAJX5n/HmIBtzZRD8vhczqX6Q189r8enq3
IlvDtrYCXvJcP9N08VyRt/dyg80G05X93leMuu7+f4pobLVxXGlCDodmsFlrQ8FxP8P3DTjV9TEe
xy7IRSDY6DcwfhcFBTVU2fm6vj3r86G1+IKunmAfLdXZ7qIMgQU5c5YSbnuu1QCbqhcZnVczQIt3
ZtamcUd0QKc5OH4yOYJh4gcN9NOyjrIvgbLwWLoskCzEZBrlaWmgk3vzyhWc586DgdKjn+ZZe5Z/
EJsZDGNoa0JPehYUAKenLXMFWZKPfS/5qp6H1CBMBAB8Mb1XkFtFMHD6QeZpQM0yzNu4D6sRBl/y
O0Snq64fFTcaR2N2g5rYYcxkko0xZyMgikjYd2aDhsVv7V7AH2G4fKJHUhVD2HloyVelCMdWNutR
Lui8DtpWitcHRuw5H63QyfBfbCzr+FBXQSzIYFjY855G9AyWStewjy0XBeb2DM2jIMIegawEKv+K
c2GeuLI/cL00euV4bF72FxmHgOcPzK551H6cBaUKnYEULwehXJF2iXnVXZqcqY9CXhzxD/fH+yMY
yjdPMyrWUO/2goZ6TfuLbwcpCG2PbW8gscO9LvFkFVd9Igui4EF0678xlxldjmdUVjnfxE+A+pal
MrCgL+YQv52AGBk4/inv8NqflIqgT231J4+ykfGECzEglJJYDSn5UxAG1/E6JHZNij7fIHgewC5q
zGO1I29mXArExW/RpIe9ZobqdKp8O1A0rU0KJFAyptNim0umEFwwiGHCsawdwkVGDH4J+UEwI1ab
+YkAmDWO99R1G3a8nJMut6hwqyuxsxoVUv17/zUXUxFll7CxSBfi18bOJyGotdWp9BW4hrpkaI+X
H/NmoqOB5YA0GfW5+HbUn0DEMgESJafNOX116cbJap2QQJ5bBRVWCdFOyms0h8ml6014OptH2jgZ
PKaCHEno89UCjoNTMVtOX3bUKpYwRsXaDw5Ryl78HPceFzzOjv6BfsdSTAPj3xU6aiTABQuo14V5
evG73sVcG2Vb/Ke6ECr5D6fQgzrYgfJ5/EUjYxLC8jOX41Stvqx/eqT7TJvxY0eP3tAGFu9RrpEZ
tv63B6dlVv31lqoUqVDzxzO3QtR5Tjbnle0RoGL+vKg0nMU0YcFKJ//H/Z74u086gB7IHufa7jDO
AlTSY6CLTmKYgT5shytX9alMhlujhIZmOzNK7tKkWqr+FlTWwvUeH0ibAUATrBhVk5yidzrBcVzX
UY8rY7WL+06tq563nh01kAJOPU0LvOXRBqXOLG2ta28C0qDAafkv2DCqgQl5BVRdvtwOwp8PGUtz
nwi7mkXA9anFE9YSrVFGmONHFZnC9YZ5hdS+/z+mROBuOTn6Ct9+zw7Z+MDeXm0gl/zYVVnOBK8I
4JdYt6YVAN3GK53/WTXoYUob11AxvA6tfSBtPaaq741QAPQSFQTAYzGvHRl4oz98Gi59CopZWOTi
uFfeLmgqMPPZcB5IZ+aveMytfgbeV8gLRT4Q715dag2dtm5/A4/8/SmUHeg27d87tpinP6ol60Bz
Yq/zpUbM0hCHpSP9BTuMBcCItM8ufh0zVkwkseP0gSEPP9jmkBmFV7ZpVyktjTGpL8zFt1PnhWhf
MdRnpH4MYT8ljO5uTGcqdMsDOJx8mjTgrlsRKvA6DZFL+QAdW6cYIYqMvpkgY7pQk/X4Eapq6IZh
i1x1gLAWKIZgP5oYtqzQ7fzTnmzIWoShr4c6eL/flRiB0lEthBigvYiQl9gP4faYAVS6bKsmf9NJ
JJ2k9pIW3hlGWGF6P0i6KffFTjahZaYfae8+zc4m54I/zGGHGkrwZhrvpys9K9+gT4NbhinLMIMU
GbGTSFOFC5ex8/XhPsjWPzO62NjpjNKpPTAH1mFP+pj9S4KqtjAnRqmZYN8VxON4yrFOLDfS1a22
jWMeRHmZTk47rN6+Uowa+dMKCahSdbOoEz30lIQvIxwNzhXyeeGYsr05b461g+GVphz4iH2YvoLy
XNJ8dFWUCcJ1ZRoGYJbvDB9dABacW4pwxZIlPsMa/vtrl9N6TVtp3x7RAf8mV502S9+7890+4Hpo
lq3Cdq71nBokst6zMibZF7SFfcZcRvirQH3obG4wrUSbv9iCd5bHvgHuR2euyCIyeWbkfUxDg7U2
aE6/tc11sDgnaMHtPYfDo54h18QVP0zMgdxhdM98CUyI5GHmzR0F996ukcPyD4LIgA3vI5maYW51
7K15sallyvrAbTNJgZ2Dh/U5ZWe0OAyOf3Y6jjvyNPz/9jQf84+rE8zRMSFvqoEM9FIbFE09oncJ
PzisE2J1SjKirMHnkAcCU103NQeRVmo/LQ7dH15aV+R/IaLUNd4v0PPS3B8G2RvvJekXB6SyOXHo
1ACR5heOjSEOJNT2vq/qqf0SrgS4KM1LCo6h5u3z1bbD/1RsRNpOAF9PnASVdfqwd8vrnNRZv9Gt
zLxcL3lHR4sSvh0497KrCv862hAFwQdmwlRk4vetCGuv4v7V+ShJq8U3f9aIxpvGTzfkrMzVAyfA
1RNS1lUYXIhEfYZpv6VJabPsbvajLGkVQWTyKzI+dNKBm4mX15Pv94d3eEM4h10q+b98uUjTJBgR
Uz4Al1LVZc90Tq6NJHsDQljeMdcw6FeAdJkJicQ2s676YU6jTwPrZOVoV0N5iO9GwnfuF/Vtbz9t
xUZMVlZ+3qpdcEEK84X5/k2yEfi5DJFC0EXN6RDTS3DuR2e/Dx/eb4aVXI/ml6XlN2PTRhbwOLQc
Vxh495KsjB3k6jIaJALLm7xY29wdjOKVU8oBErmdjoKcJygPEPv64B9aZmwCIyK5P+X99xbOQTFG
aNIXWI9Dyk1Ue2KD1zyO3bsoPOHzoep2lfLr7WnCtWuocBaidGr+4cdYSjX6vs2MI1X9Kah4FdVB
EoL4B1/hSKa/88mwNyNRtc2wNcGSG91aFMinunztoX4mla4qPoxXB5jL8DqS9zNNB+9GNMR/P8lK
BJqpdo/R12KMbi2D3f1fJtup7JnF0Rg4Ui8HrM4D1fQVSJ4Kq5X8dYuhVWqYV89dMizEvK6Gh86F
KKcGA0Hf3vS+YWliQPGqBVqvEzRva72/p27WlLd+wBVjEnSmjRJ44raZuzpSPKGYkrbA3ATspf4j
AD73A0lIZS28G5L30RPDHi85KnF9cgjgJ7dXdydYroYud8/BLbkJ10jxB+YrHos8g112Tp7V21Xu
sGE0gp0zNYjt5zedrYFJUBqXDi5rl5lOIEuYNmTR0wPFMLZPRAjzFqgTMDuxHXNgFFnHrjKhs9T4
xslIJubTON3Mpmnbrjbqz0itoCnQaoOXj1rtp1lPKBBJxG95mhma/uZPHp/cMJV2eAgxjHjKAGjZ
7xSHbr1tXtbri6NlRHeVPYeOKvPbeOsCqe4YlgiFC2MH7k8+dM9uw6n1x//OnKhHZo0caAAs8+Xh
Rovo2FpAupILL++MV6+8P0KLJJqSgJzzPcHupJhHLDk2qBCqxW9ebHsdoXQj2iO4l8ieSw7tocdn
IRhwKx7zvwc866yWQEYH/HDnWEkLCUSTz2GMRNL7t2PDUWD58lXgfUqgIZ5+a6bCngltj/wChGSl
99Q+4FVd/uR0FVppg98uszxNKhDAT5xq6dM9GMe+EVTxtutW72h1wVT74zxEt9y0siqWdzyRCjeX
I+QjbudeIFmHbzgEKFlQTRbFDaEOW2wnpJeXP1G9VZmXg9eZ4Pj9Z9cfVQaZXliDMUDuh7VXPUuA
hgjz1KZ6SRD9/sFIad6IZ33ALhSHs3kSmS/XcKm21c5QYq11ASzkyndbqgUj6aiaFFGdNRMwMO/D
c3YECPxJ/ODpP0qhO1HoF5pJxLmwvAfbUlbVdpf4alfOwqLWscnErRoIKmgiAIhZBfXipE6kdkZo
+t8E1p9NiuZoD0uHni8Ue75ahY1LWSovzfic7f45AKU4hh0LJzG/AunWdwdsPQdfEHLUR5X/bkvY
oy5DHe6ujoDVsc6BrNDu4mBYFuwrbwwQ1PLMhP/iT3wj6+COEfqL94M13u9fSk8aCmeA1FSmnMkQ
wb2F3CovTxaP229VjoQa6obreuuERCwtOtAd1YhV2cxpHANYaOsdRIuH+KZ11aCzT1pLRts8p/qQ
czvFaeW6VAtb7XBpdr9h9rDVqtz66rHUEipzvGScFmHd1XCyQ4T5socFw3L8Mk1pJeVNRV7SOUAy
NMeQbeGbcV7FMF6O/FHiz+hCWe45HYcu+CdcobiC6EfIDs1XU+67MU0A8Q6VCKW4y/VXId9HnSIi
VzVoUgIxgktKQnQMh9jYQPGb0dlJhjbLaJsQSxMJpkdGJ2XX/SW4ZygM08uL9F0KeLFdlkd/XUSk
m8EtyFQeBuZZHAtfhb65G1AKvxFWVm19CqanveTUCL9QoVDubVvSBURe3H2Bu33VOBLYwxQU/u0q
ROjoAaS8GCvQq6JWOzSTh01w7coTNcS/TqYeay01Mt3Haq1nTHKRiJITz0Jl9PRlHfF54aFaSjln
UtJ76LIvMLRuDtBjmjqpJAtxtmI1hEC07ZFJBG2e3Ku5E/cHejdEYb6bXX3ZWu6B2BPq6TcoH8QU
FAHkTOWy/3lBdcgjxPqeBCaedTEcyGXJE3zzBN2uaLFwosJtsr9/Mi82TXl9JIDL5tQHbLoo1bL/
DP/n+pMy3W+oo1cjBKLFgm/DnGmmjzj8CS0eSkKA0nh9MSQiJo0wzqQyGiF5D9UchZUjaTCyyv0Q
MGAjxXPGJmWx8Pp/NkBUa+1cpiSFwaVrHZhMN6MgLqOUVCfqyBf/Izv9bylBnKePEBV1RNRIiKy9
8YFA95Q7vaGHEa8PlPZrgybjCFFoZB+WnFs6BmEZHKG+KDrZawreKL6BBeKOoF1/LwKdmDxJkiLp
yh8dRmOU2gP9FAcD6ZSV7XWpc7VGyju8FgvBUhQ0kS+XmIGECqDwoK+Q1hbYdQjfIaCpkt7s3Hu/
w6VBypvliz3JoI+jvrkjrBk/f8ZlR8OsY1GXOqOpyJCILOXBU4wtF+zC4org7PMeTOFIpLoxBmwl
gz3hOBA6dzb4gKYfED4GUwPFiSwKe5PBsKKd/iJMbZwhY2W4DqcQ0f1BFhOcyBz3wjGZpz14c6k8
6BHQQDvFsIbvKIXwdPDTg8WZlmmjsTasmWib+yqfIqqekxb+RaMYKIx2DJdS+9iNBRC8of1Cu0uB
7RaeEnwFbwDtZV68xMfxN410FDlTSJU4XKiPL7IVpBSYn58ESWxuqRqdYx4+XLOPeAW7CBCd4H7F
8ZIEs1Y0te0V1XRiS8fJcZ6Y55JvEdddb6fpN5ghcPPVtn/1tSZcx26iKsnwId1RD1LQk23Zwk7r
RJfKn/UIS0SZFfroeWVLycAeEY9/6BNBKDXq4dNkvTuGZ3XeiSub2foxVzCq5eEMbBsGAUipX9e0
8kNNw3FPxYa5pYpkt7+9ggyRwb/P3OXl1QgCsgSxAbSTSRqMnk0MghPZksMPOLRN8pWMPIgps4rh
PvN/6u+1Yhbm5hqjFJX6LG1eB2bjAfZhPtpjRKbIOQQnfoOQf3/K8rZb5Wt5b3Mjydgnv50nlfQI
lc3DB7aB5FsWl2LpBW8d+PG7LWBNLi7BiFjnr48cAp9TmbrbGdYtKCzXRTtmYz05Os5DJ7UGOED/
cARWYKAk8fXYPclgYlGuo7rhnFppfOJlM7bHADyPN5HxNZQTh+zaSe79mFN46O+x56/HHP6SuWrH
kGftTU5Ug9bi63fU5Gy7AKLMWqC6/HxI05wy3F6tPxTHPiu554iEc/jSQ41sR4RC9ddJQ+PGFx2h
D5rymZV/eQQbJuvJgDKA3sc9CAN3PJ/7H3pQQrVBUtAUn4wTkHSujAuq2K7KY8++aqNfSwFvMg4V
2qdHvHm7a5HxEF+Koc2KgQtY20XO0eb1wFGngJ1IkBRfdd5eC/yo2a2EIVMKQj/bUWueUK/OHSw4
0Gd/GLh4TQWIcBs6G72f/uOMGOV0U6lOEucZwsTe7xJ6jI5Q35QYK0qmLo6l4a0HhFvH71mgVtE6
38npjOIkFbl3HYDbUvxqKnzyuEh54ix+g7eNGIyWjcm91V+QXZtKKSik1MyKkl1QjMRz2FsgyZ0C
sNKnktejG9OdVN79A/QzSWqgr2XRcQ4OTAMxYTQi3Y80PTZA2tNGtSqYmUUhwf/bXiaUQKkH5gSS
ynFpFbRqCkgBQExW3oDTJe5SkwpzQBt9MEHiEGWhKNRf3hPUPmc67qOPvGoF+y+dEW8seUhBQsaO
Ud14geRHi295fFnSpGCPpv6lQWwLvwvFNCyJoWlVZ0KZumtXjJi8dqvX88BJNhAfyV3y+ylJRJcS
v8XyWSAZuM2BL8i8o4XiU22aFH3DGfTPyRyoLKPbi/4AUq5oZUA/5mnwuDX/YdkE36GgagltLxWy
Ju7FDa4+mHFQZCaK2qcPrVN9CHQyUYyifzHiUzTQSNI+O1LDhqCMleIkZRVbCfKc8Y9K0sy2b/uH
duOo2ywXwqOCWqtJH8CV8zg+b6cTg+lovYmYFYYdLXQtJNlFoo21VxxtZlVZ289zrLEt5/xKVqov
3i+5+hbmi/xRvDVlDf6ZxNIUPNvod7sxX0IFwujNmVvjZz55acnk8iX3JyJFXuaThTtYi9OWNqg9
FwSzp1Mhj73jtPL1aPb6PkAXBxP3KSpQkLNJbujtKXpfv9Cz1lRa+v2bVLrT22VXKaqo0Xjuhbat
tlG2HLkqywNef6HNLZ1BfWRdjawE/OrM6AVgTMtUTWIQgfWgT4mnTFZqeaf92pphT5meP2c0RbQV
nuG3srxw3W1Lqe9fBH6cnzch9Zk2fyxEuegqxw5uZOTh1Iuru+GUyjVO6UeoajawibVvqL0fSk1D
sHLAIRM38L7QxzzeMbs4TOF/Mi/6iT6dfI+f8hZj1ly+5HbpDVFbj4Hjgg0jfP3fBClicriI1Fcr
WVpydDrdVTIku22+BTRi+GT8DZM1/xdaG0gUt2EAAshLk1fv1A0pd2JL3aVQN4pkArT7k/vCfka5
94fXd9M0/qzsPQWCT+gQuOPEY57q0uJnMTPkogjbK/wA2cV5pCEQ66+vLPzfIKlXNo7QlqX+lygc
IKk29vD+kmuwG3S3sr3fIpjgNHqgB1TB8KTIjavaAl0DRmpG7D5VWY9ejNdk4GDCJP3nW9+m7o5T
yEE/MI9XCjA9El3ftmWayIEFlwd3IfUDNlCS1Tm1fGCfiNSYITHk+0wxV/JQoIOhu9eoZ5bkHZ6e
JkesZc9oBfMqTd/6irITXRs4EO9uGJUPZcjcTe2d/ARnV9/GL/r7kTUEN7euSn/XKiWJKv6cJJGo
qexyLkgjW6dLvbX0WV7arhASEo8LKW8pMoLIbfWgvdQZXXHtZiPRJg7g5288RJpBUELiLcdasZx8
wax/d0Gdub1wrqesLwQxKhrv03HeVvgG4Jxtnh23pKGp3KaHCKNzIpyv8UbM6ofYKq2YUmOc7EFA
4ptyaLPfkpG9oGxTXemZzGA1HSPhhkrdWgyAxJggEGGpRmMauOwy7iggWJ/40ZUBH9o7GhVlfAwW
kU4aLq2xlTOwnsyelltnkXsQQJTzcV8aht2kuqdJdFaPZxt/I6xM5Cg+Q66TF7GU4q4ZgxPPLSBZ
6EDT2wSLwa+qoLRplgSIsH0DXzfHum2d0cj7lMwVgu1H8wByH2OIF85tYijfP+YLvvgmpkAYyvco
JIFqnZUXbC6CA/Qs9goJJwVGDhZRgYTYbQBZQB/rW6XDawlT+FxBjxqWlMHWzn0tMwENnCWJwe2X
IrH5xTcUPLehnZIO067PFHLWdtmZSGF/WNUjuPzsilizCe+t7kRLbAOUF3tlI81LBkQ3ttQ/vn/A
hX1jT3fMsk9ZbRQrlfanydtsSoXrxtYXEQLnc20Y+dMEHbtKNXBWlBvCfXQJjC0qqCyQcslCf33I
KCa4/Ig3Bew0sNe3ERn6mzx0idbsFQ+ufijqHrOoWUikhorvsHGGZxX8PsbPHP1Hhz3RZgRxXaGS
TYj9Yxke03jOtjpMaRTRvSHyLLqzaVgFnbYY0zS+yeX3COV/oSy1QHdEtYxwwETafi4cSz0lENQQ
lFO5mAJIEYPILNWw+vQ64k4fLd/u6RoM8c2LroAE+YimWUuqtgGOQWNf+Rxngr673WP2SnQrvy1V
AZpf0nJJTxqPE+YpWvGVLQt5iGgp7Qwa/T0iOrJ5YmOZN5WHXB6Xkamt7wwVYgv4ehDn2BYg/9EZ
rdH3H2Du66Q83IHQoz2Jyxchak4tJ5n5ivLCX+Vk6/v1fofwKIOsZoXtLiz3IEzzoap78u+UGTmQ
GbUt8Bkp7zLDPaRuxchbbkZtF5z9kZ+8khLBogOA7FXraAPEmrNwLsDsc0Ia45HBpXj9lCJaagpS
BNnWuaTZX880V4QdDmpWr4HD5sQAAz1Oe5VJqDBvgNPXjgihMWiSiP1emqX2FDrZBZoBk3zCX2Gb
+h907gVgeHAisC6cCHQQA+6LK0ulH4EDKCd2bJKePUGu10D0Xcw0LtA3l0d0S9RSX9h2y7dQedZ1
3FXGniX5LZpZ39zLaCuFg+n2Rm6Hl4SfkoS1hM6As+oC5ZuGAJ7u6i4tYitDCr81IXMZOTHZ6QhS
VMbbaRpz4vy1emCk46CDVoysSVccdFucYNBbWkdsbrXz9Hr88u6WyDjMEJTjuYfBkTdr2srUzJe8
VdcVirXcvrkJxbcTh4KORtIH2lJoGy9prjJhPfPc2M2SS8UAq7hUtWQkh7K2LDCwYqrjnEXqBfst
Z9V3xxfKpp6ihyrR1jkYFe/pJTGEtU+N1tHW0Ksu2r03Z27rdLSH7JVOmSt8fL3mRQSy7T+uI87i
QKFixTJ02RnfyUA7vVszI04eySz50QuKpzGVworQVH5ZxrAi8Xt/UeI2/Hz4lJvuAwUuti8r9Vwt
Zffc1usaZA9jtaINDQXYhBAtlT9PLIWA3FRtNj7LzjpsXj2cbB3jzrbPj5pD+m1NDT9AAlOxMKxS
oEKX5UUk26uP5IeaS7QXCqMlJ93JV9QJywqwJZd0Z7dIlnJ9vRsPchpQyYkON1ItiFsbgLYGui+p
oKDSgmC2Qoz7Zf8sH7jPSXZ2dg7yaxAkduPV+Fk8pHNfOi89MD0FDMQUChelVMLksEuEgEaOZ/U6
TmLBta6MpEOYK1VsVBajvlEuzNWnBFPmzUXrrX/thZ+DpkktNa7+u0AiwY4EjwGtnAokFan+UM+7
eLwWzKDlCeLt4fVkfn0qRmAREmgXFa33lAakQYLAKarm1SwNKmlmte0J2785KW7V3G5+cMPJC2+T
tg8x/G2UMhuEXgNGMqEx2KVILUPISDMyUu8zRUzifnybFOCVbOqT/b5fYwmofrBEkORxYi/MTcZo
O/ri6O4ct2SaSaPKXQozb+eck48pysknjfKRJmr30npk2O4HfyR4QM68rLE0zwUaB5XIFQNn3FNq
Ca12TdYwml1UvCpNT8atgK+VzrF97BvcU8riPeLnw6NlB0UNfeSBAZStVXcMyMsEz7QfKYsLSYdP
zhqOu4eWNjPQl75uQeMdcvHK194LIif2R5LzfbBc9PLCYTsrUbE7atoAT2EavfRZNt3C7b3XBvIG
eyGc5NJEzp1Kd9h1AxUUw5cfkV+tkZhElFAoJCvbPIWj7XxfLGKm8yZh43OdiLRGuuyAd+J0E8PO
4wmSXIK0PbSV+BUYDcyPHnhz697by8+m/mK7ePEQXf913KBKHGrTxVgZVjNQSKJ1Yv54IM98T91Q
9LxoyqN9B0Axv8RolbVpy+tvTsXCRK9NupjgkGVt3VcaZB1kdweJKlVFLlcYy2dv2Dz7OvPpfW05
5eipvTrga3h7PEWjaw6AwCXYAa8lvrubV23p1AJqMkAFZtUz5nyVIH94nIse2a97V/cM9tgPYWhv
+s16jf4zl1lz8H2KnJEcXa3JSKKhRmECT1aXuJzFUDBPVI34dCkx0DhlRnMZ73PY1k5IFCtiGMbq
0Rp6s8FZ9UbneWvKQE02oZoDbuO9HINHFe8h+30IJiBH7WE9kWOB3R9U9TFZ5HJETlXfougOfwTq
uHEoHueetfwpCK1hic1VuGCaNVwe/vctzMUVZZm6T4uAhGmG2c/VC0HtsbuKBBkyNxpPGWfiLvh4
xaFDdgsQJhAYCuv6hpc51oadBzPgfgmnVVhHsSlD0bpTrG4vylkmh7mCixoJmKdNOjMO5mh2Lfei
kxteuolBfbWBNh7Te8KP0qR0+oR6swk0aL4qnqpRIDqQJ0QRjJw4iwN3mzzQO5ARr8NS63dzYknu
zftcIiZKJ68UcfhMFqz68Bb0FgD/fmPfLQMxfk3YSZ+dw6MFmECHEmre4fW4ZwiTwps4F9idDW0Q
4FXBxoY43f26ObG+883z6y68h3i0K+ka4Txo8q0O92Mcw3spAPBM/AMytk3Y9r7iOVNTN9hU+QGv
Urpmda+7BmhZ0RhBHfkD3Zu8DVyAd/LfcN2+hxJHDLLMgFvCECjAWyuAr3jLVkEwEdVZfvzeiNV6
vCicaBuZ6nRymB0qNrdwJUu6aI9fcZTUZL3flxfKRTIbjqbdSex+/miFC27sGrWBZc77HzWQnQ9A
QBLtgbKYsFENXwotsml4p672NRs8PdZGZ9aAgY4jQE+ZhDsQvx5tAA/b5Nml2xiuXjKgBHjbacnY
Ys/cDQcgxQmx1hlIqBAV/YkL9AxPUtlMyZGuTJhiwKRnhKpO0L4Cu4LFO2eGUuHT0z4Shy/eM3Pn
UIgjuvUxbZM5o1tmfqsSNwZkFt1wgqxXfgqJ2171Kahlb/p+4uYuAhixJ8LDHSxbTusAlVKzybSj
HVIbFhnjdtpclWLYCzODZAw1dw75LcEnSAmlp5b9X9Z0YBR2vdN8gGdd70Z2kf+1tFsS+IL9QBDC
cY8PLUhMgCHiR04lXJr4BpBQdaZ9z18Zw94WKd0q4+cgKiQNjqfgi0qsCObOYXWIJk9vF/T2AU2I
j04e8bVEnl4HKH1BoBb3BhMTzOIDpR3LE//McmHdVv0u/Lzh9vVcqTibQiJGAkdD6tIsl1FHHQTz
OMCVLFJgYZIDRdQ26/T9v+JdnA+KqUuNNaLH7OGUZ4FaZ383s0+ZkhL3DtcJW2Ag+8wot8wimaCa
FTMuxnDk7daKGGZVN2/YDp36+k+4TLK00F54mNCimQX0gNdmhA+bIfCE5Vz/qnsIsGWsgKH7RvJV
glhPG6kcC34pSnYWNLRWZK91CYAcxW+JvTHRiwLZ9i5qhZj+bUQ1LEwPYDwJTwfNUI2lUvJwbxRZ
viLgiYd7gCBy8oQFHCwtIxG6DQtYNV+n7xYnTn2US2+5/iB1Urny0ljAzo13VYsftOTGNjCIUoMK
IFE2cdRPcuTohNVC93UW8RwkQdZ4bNDLobYKCr/EujTPhDawttQCzPCrk3JlJFT2nJRujW8JA+UK
cheHh+iNxBUtGiL4nqnv8O1aEMu/et+ekL6aueY4oea+xJhXXxy8UNt9rJGEEpXhtJE/YLjfkRFV
h6hnDAB6alPs8Nhff192lxE/F8aWq8xXDDo/DmdZdfvxMr9UL6kE5KYxkL6F7lB+8Mlw45zHsXe2
V7DN60yPV+eVCr2ndyXNqBz8MHmMi40QqkQbv8A/v8XVqr7j4rl/RCFP6W4RJ77Edcq2Fp9iIHqw
bELAODGNMfady42Lcoza4AhisjmAGFB771gOMsWdkXB1DOxRbDnYywARnfPkryEqMsE6Fqc2aGee
04J48uoccaJ/aomuRj1b0EGd6rb2EQSb7QaZi8iS1QKLByaKmNKMW/2Vj5nTeyP+nCTJkcEWPNRI
t1Hp0c8pWp6czdv7UcWRpydS1FW7He860rMlWMOAKe2bvxTqqMaVnX2OjFmKdJnTuzwysC85LOW2
nW0sCGx4f/uhOilqLkGId78DTKTb/G2Xo8gw7pLYEfy5DDyjo/Oam4aqjKQqhKW7fa3F0+rWATz7
Hq3g5SnLATcxW0+TcA6RjONl+TGKd4t5JFWat5GRpsJUFf9t9Vrbc+hlXLTsgCfVQqz+9Gn2mube
eNie9+mkJnCMJJIrbfrA5kFAbz8T8iHdXsS74UtRhNyNs0/w/HGzOp3BIT8BTJdbjusN3k78qp2G
eCjxKjXqd5aemzqoicG/gCcanK8YDgk3AL43nfgqxQ/LM0urV7ZNtCi5Ld7jZEZlpLGz6vDRocJO
IBx6rrbUR1dmLr5BQ8w8YJkY7qELDGprcJZhqQ5hPibeKDsEGoqaYwsJlqs/Rp/4523tjKkwhoW3
oE/dJaOR73kRgAnoBPmvpWCM/w3nAaqIDTeFExgqJYTRCxYL62kArsugeugpwyRu8vBiIhsw/mlv
v71zfZBhLQzFWQ/tSGaDFMZ3NrvqVEqH/fnKSqLgSpmd10rh6deXqGeXVGWbrPRodlatLPzNatBz
ZH4qAA0L3mNqcDW2C75PYq+ifZu3Tp2VhWnSpUCXEVzsbYJezKxNHUbbyW79kxVNl4q733xqLMgz
LbBmR4JPckpyK3peiEmgDPw6hjP9aOfZgx+9bXND7+5EKJ+cREzZNmBH5Gk1XsNGHP4KUIazQi1f
O3/IRJgykFI458/hwUXT0yJKFeJYSie5KqPGOhYyfgn3oAFB+PaJFgJjVVLhgad/1pJos2xnfbwx
wIQznf1pgryxnVeCiUgyv+pwFov7ujjveZSKUeWq4XMjUim31qg70EXNzjJY4Aa2pt0onZR2rVRL
wIzXLDTzAroZwgwh9eZZ1j01eKqJStSnUSheNESC0XZmrSueuoyHv0I0KYoKY/MksvopwnOT7uru
DkK4AJbt6Bvy1MXTiPp817CtAcjJayhRUwxaP3UbyyJaWcFICcf0fUoL/6Rl64hVTrLdpMknFpaZ
EnGgal5Hp4pYOtSplgGmMSoTcOXibWkqPlgXhzvHE7XE4iyyXhJEqLNNTstW+wEdxpsF8xcdbtIb
v0favq4ejP2AEQD//ilQ+dn/Z0yo3JWQE0d4FAKcpalGHXJhE70OzZr9Ho/+QYJ94ZxE9el+jh1A
59R8rMNJBCHroRypoP6r6MpFYPhhqvT1vO2C15OJ3ryFQAO1WRpb/mvf95qR+v3pQs6ZxaNdcK1y
CIgW/QqYL2Qon8l65Q82yDyBWtZ779fe2dAtr++vx4F1Jj+HVVRYvu4erT0SRZ16QoEg/Sdq8mJe
0kXZb8kMqejzZHAyL2b08MEFG42UYqUFm0XUlwUIl7FrAIvHsj5ohOwRPYyiM1OoCcQQ5RcayWxB
MCLjGh2W9+GquWMOKkEuvwz3df4TahwDO+CFl/O9rxLNk3TLlcLB3etHZVjiSicufISL9MSWsMnq
cyEbyszG/i5BJkNeNLQZ7NvTmJJ9NKOKm609Y55060u+wr/3Fe8gMMtJEj/wa78coEo0WyR+HQX+
E5mEu8Aw/bpdy27eiqEd4A9UyXz5YH7ezToOBg5oT7ivZl6500mtMrQzOKP1YaSSfLImI1BQHEVt
Rp/YEy1rZoU8vFwX7f3wHuzlwwyd81AO3TbR9wOWq/J5FI8wQXA6dUJyuctrFTiCf8ckG3O+njP0
Nt5TUVxkAQN9GK8yQ4GiGDrloLvfrO5ukXkCHqHFh56gb3MW4AnazUVGdzSKUqHyo2bAChf6EeGU
kmg7VVWzNm6juaGeC7KMkOorXdmxGcZo5ik/Iq3RMJRsYovXcTPX7EE939yz8MqqjvWbh5Z0E2xr
f2L1xYACdoevS27qQUqJ7TUDCgixb9tnbnixHNBBnwAU4k059ZCakP+M//42PTkhRE8LoR+cS4xt
KgVcK5EAyykiAKWOg2OTGrdc2gtjY+0O6gOKPe2DixXNiW4iv3y+Q/Xtl8FSnl47mf8ocbpTTqpl
pNKHOyv8vmM8ojBsj/Xby2Keh26WPhy5bD2l2n4qvj4FnbF6u5CYx/rkM0JQm/Wa27rXSsZnbb+F
/8gSB4UHL/VuYn//DffV8tERhVEucQO/XsW5i7BNsw73aJaUZql8LPbZyR4AmLaPnP17rVTAfUpl
TddrRWL7/7M+KI5G8CNPTGO91shSDp8IGpEdyOoZzxWWv2p4IkU7tFUr/6xev6bchELO89RBHV0j
V449C0qT8wNf0YJ2nQ4zOIp6QGrjKD6hLaCKzmq8ifJuGIh6qo7BoMKJ733PC9/FCkrqw7tOPQln
fgKyCbBuZAaGYIX1Lndx59UAfzmHXX9v/5JCzOQgUIOFwJ60Fky8gxHnPTljpDLmhLE0jrA2590V
LK8wa/Smd24WmBTfB7eFrSi7VPOm471U9DMy5KD5ou/FzrVExoIDafTVeurRa27ZkfN4x+vC1w+7
hDmQU1at3Lb1FsYhGFeIA+4JEKWmNfUiVt4i118b9Ahl5hOah1fhWQATX2T1QV4BcAgJjYztDJIh
Ftowf5pTofPb8lbljUv0Ow3c8/pUMRD4gC+qr40Lbs02fmXpq9JG9cEUZjPusq9cfdvC2hXd28f7
FI35w7JJGG3SBCF0+3BGxMm/Kn/XvAW2KkLlED6ocPil+zLTRxkID7Zt01+C5LDPs41PqesqY88Y
FovVhjeEYmgfgI7Ly/gtvdlJww6N9MUGKUmsibdAVUSgQMwtzJbyjtaBJR5lzyLeqrN5mTByUnCX
ccHf5skPiKBzuIprX2JRgPm+rHIIriL+EgRDFyojCmfEaaYfTTjLIlicBvPDkOxiVyHdlulGIlKd
+ZFQoLAGjtZsXrkLTaZtt0HZaV5Mq73NsjtghPmh61K45isgtBtjJ0IWK2HUkTZ4yU7mabwtfTxw
i8jcirppaGVlCOgeryVj0a2TeAzTiw5wJ/fLAz4ncM/4il45q16Lg5xFja23nlIMksdr05bf0dF3
4R9ODpAqEmN6Lb76JSJSXmRv47PTHz9oNr+iVAzPG4M5zeaWBbuZYG3Hfa35dHHUUKpkJ/U4+KQY
919anFDwWJejLFWkosQJN4RL1kAkGOJ6YEtJEXknEi44MJhQGpYxfz4msBmB0u+M9GBVIrlqami/
JsCSixa7KVpEAAMbCjgzH1gsQ9j54SdBGo/FXCn0wK+k4OMYXubmBGz640+IEbnjNUeBO36Iry33
9eFdhpt9doIkHJ+/wBlzXpedRbqbpgV8yoFYA8K3gwUYqsBHdB3s4yl1E7YYrD13celAhUo3GDeg
lJUmNyS9YkSK6z3cy9ecVoG2uT9ZEQjQWLEjIv9szYByI8Vok9KgPjjhksrxNRLzkSHm/KCrtf0i
rY5UDm0EAffc6PpWkc9IXjwW52u1+zvJ87KyTPD0wqFZRrVGkpT1CsyycTz1czcsKlVBGZPw9EHb
Kz2yax0vEMgcFonowUSKb21Y83KN/XFtgDP3XE8T3vp0/kvQWbt/dHX9M/yCjx5FGGch4wh3WQtj
jRBR5BHYESfuTMo7jntC0r6o6sc02Z/NyT4lm490uEaSZvUUXDdZhecMARSWJeQE77lcTgB7bG7A
DYDsidaxL5pzwnnv6JQFQb04kvOexxw0PvhGEOVSHUYU/6flqvk+NRBtlo4Mti3dQmobAZvChMqB
XS24AN7m0zFv9ywJoDC8vuDyFRue/15TxS8lAyKdc213kWQCYooX6oEYwdY46PdTnG4Bwf7xBjQL
0S6NXHLREB9XV4btd+uPqEVEzFz25vV0iSiSRxiOr3hqw4qij/nklVP0zsJdU2qGsAxp13sD2GqE
WFOTBgwlgOY8PD+0SWScsBt/JuCjbnWwSEQg3WRfV9EzJBOKePo/K4w8rWI2u6ksKnppFiP5mIRT
vp4Kw6v9E6VG0i247YfkJ0Asg1+yhqZVmFIAgvXhqPMBertb0KIAkg9xNzK2mpt3hGTC5nlI43vE
CtARW6YQiK/91O5xvdqSq4/bW/uRoEz6shPAb/RKkjp3s9iOJV/hzkuouW40Xy3SJkDcWs323jFd
tWY7qkJNVdBvOKxVVazF1CLYlrgeyw+Cf/jKSekHDNtJVzTxJhYQKB8njSVZDVUFSbvlaes+MwrO
S3X10gnknjaGdh+uvuJ02qL2YfFuAPC7HCdWTWuCFCD+W7fWruoAfIrmL0EWlWC93Ns8pUOpDcMV
tj7xitieKAYyXSwQ1AUg08pjwubSd1eMi/U3r5es0nkwbdDVR/6vH8RfeBBVBJOgLSSU2fU0RRKL
ECC6W6lNi3yDWzJoCKmKQ0UOMXPG+RnbSVEKqDfz8qPNkZkbDRlLWbTq3Zs7erwnE22oi/ERyP1j
UpgLrbzFqnWFHDFvaasqVpqhC7+LqkLzEEZPrqcfjana0b23L7OUmcPi+tapTQHQIcycwjfLRpP2
xhtl+CznGspPvXbdscCfUdZeGw1T304uhoPuXun/jX9hQQ4S6zINtW6eShPTYIHYdtFcAWcLV86l
L9GKQ6teTeAY4P1DpxRwBq//Bt9Xh4xoGEPK3DJu2zE8CSKZAEEToOTRdqM4FyhKKx+vXzpOQ0WV
5i6fWYpIpi79j2bMNFWH/vX55xBxEKqaK3AeNyXfDAaPCSlCpWptBmvpwvGh+T8p1x3whEb/3zes
V0WKxmnma2ejIWWMU+UKThIZaU1xWbDJaIo1TLjiSq8BjGeharJEkv1bFZ9DQ9LGC4+icWUlxDSD
mjgUcJ8auq3Xnq5pAp3LPGrW+/ZPZcc1IblXRCDejr7IYdvaCEtDg637cZaOguC7vdJbZqr5pph/
aiXpGM9z913Hf5Tw3f2DLt7xvYREWMzajQEgStfNY04LMXJYEKRz+9xKBg6a47GJTLBnk4tPsTrg
ed/fmqltK4xOCwQTts4EBnEdnDa00+lvARLhaY2yO+ukBlnABS/oDh0kPHagUi3egjVwvKXsy+wW
a5U6qdoSAh9+yLQ6mdf3aYk4RsnzZEt9q49LSne+Z6kfZQnnVfaa36829pMTuY/QvRJBkavsV3s6
xfzw/775selNi0E25FoRxzTGIZldCMvCTyI1eJExL46H0JXyGLAGXVFRa8n/hL2V3KKQJZKQQgJH
FayojUEWoDOXlZ0J8H+QOZFVUBKZoq9oe1QJ0JPWwco7pnp6NDFyqWwMP0Ff+zANVhprj8IzW/pr
NkFz4utHpB0eawYbW6Gg3IGF8jcy0qNkMIDcvPDv9aTUcFZnQgOtLnK/B6xIEShc14AKvcdmnhkM
PisJ9TVh+W82wiH+MPgo3AHdh1pECqhwO550rhVl18X/6BJy2DPxeZN304ksqczf48MhKRqSsbs6
bFpPMLkcJhS013OIrhZRtdsHRkGxWmeRcRwU4k6NgBfDtAUnuNoS/7iedkB8mUqno0hKHjGb1GXB
TemhjnDzriOd2qedZY9lF0vOXCg4s4umc/beXaySeSjj0sDG6xJ9dHUwqrgA4ZTA0EK+m6Xz1LnF
g0kj5kyYFYAC74KuX0RT8TNy32tipSfBI0D4z9tzUJbbtRwOWo3Mao4qAESzy5xWwPZnWajU44ZJ
HhRB5xlRwLKAZ+SgjwYlLDruycrBDRvF6zpGGp9UjOvWV5WL4Q1d594Ps/LRc1e6UUXgqmyqL7+h
goflTISN5/fYY68DmohpGmC6teok0BrqB5/fEBBr3UzOFCtawLh9FEhqRdZwpA0YM15rPX6BzwE6
R7kDave8c5QAagL05y3K3IMaUb5fVoia0zx3NYTm6fUyuan4Hkxh7eYpMkXD+5JvYKs3ccPbczeZ
PHMZprjObaB4evTZdvedoZp3ekx7FiJ7pUl65Fhnaz2l1dO6z7y78nqdDLjDlBKHLikb94MCni07
ki/v2Cu7CQBL/FlVmOAZYRL8shqX3/Ff8ARe+nVjoVZ+McPi4cUCSdauYnHwpW50a8OkG7Upmico
QhaWbYDtmMFKEYqAjicd4iW3/wx+XJfsjjqAX53OkUSqVJ/4ubzsPYy7C6d5Z1XGw84Y2Lh/LZ+n
dZm5MOw33xDOPgv66o4sL9hibPNMz0feqsR1lRhYFrgeiHV+pN4D5lHr7Q2xIDsh6g+gdrzvOycl
wYFaekPTk9YNd5xYvvYi0lWPYWk5PBm1Cf2Xnu3NeHja/GSlXE7BfO4KEaxT5Ep5oo8ekGI02xJd
wkZYqGNacxVomIcj2ubtfAg247vEAYOXIJnqcyW38atCK0yLUPzh+8Tt/Tu102Trft7rJccKL28p
zs/qxLzbDJFsLiAUTxegYiOxIkOr3rxW5qnrqkDbxt/ZI3v4AjZRBj5BLuHGoAfBlzEngm2+gCqI
Hmpo1vFkrh+e+i/Oz7OFW1TBQiK/Dgncv4CeDz62BdVZbiopax7ri7n6c3Oc2wuaC0Bneli1Lmte
xbw2p4dklUf5oYVpuKXJojjJ4yvua9ihy+26SW6bwZI3rSqca8n+uS8z5nJN48ANCwPrAlOz7ZoD
A1fA8h/p2VMABXC+4WtoPiOfoPwZW7OVcTO3N5SDd+jLq2i9tWbHNUJA09/Aj/sN2QeFROHClZoB
FnqK8a/MblXDEwMm6CxVgJvkjqCO7R7SqJRsfrktKHmxLGIcIwv2yosLwuHF6TKAd/DjN/k4oiRq
cW33WzgwdHlEI/KKOtUXllMCg+k8JG/VrpIbqHKQCNghNK6DolFtDOWiM10MqX3J1To8Pts5W34Z
CriQ4kp7phdj4FvAiUKNUKNywtMJBdAk1QEwJMVi8KRNHDiBfKVMB6nVjjByB8ZoBFinEJ+16C3u
eG7hfme7MEx11bnlqchZlKqsY81weinqjsJYt2eXa9UH5da7YNDUISv61BWx1HtFM4ei0ywHNigV
7RQu6GTO4zoQMye9JIaFDPH1VRWAuu+masjntj9ZTeIbSCkaUW0qrVmxgQKOSDZ/+Wh8yjTtk80e
+XauocPPo7KnOhPffpd0FADzO5fXJXaBvHYpqJZbE5qbtjRazsjIq3bK+7Jinrx7IkvyPW8CgPT3
3QFR4EDjhN/Oe6kwEF7RotezblXCaWZErX9jZm9qw1tafNDh1O3kLHXgArgk1IWjXcit2uwEQBKT
TH/vuypWuq/lfOJof2GN8NQBJiSi31S1z4kLlaUPg9tUfLrDNZuR86LqNw75dktA0EpXk+XKHW0j
Y0LNJHQCqunoKEPB56U4ixHz5BxU9FbvukD4CVBQiyZWiF4tn/sULzG88x1reADx6qg8uP+eVwCv
dToBsS3OQZW0E+Ss73ysZgD9TvTFcq3lsOcEQxSl+lpI7mfy+I79oRNjhpSL209TA+W/3okORQKK
ip+fTURXaX+Rsz/DgaXodqVladrBcPmbFYnp+m61SG5Ptmv3j5BVjntkLVaczQmQJHxWuf68z0Gm
O5w6ZA3px2mAwvq1ap0CIHxedurJbZEpiks86bPWAmJ0bkY9EiRb3MrsD+ftXAajOTfh9AA9Kaoa
VSKUjqXMAzVSxD9AuUdN8owFekhD+Hc4ariRaLSroeQ2E2fLHBnN8YKvHoeBiVt0WRw+X0L8w7ay
Tat6TsuwVYLO9g6qZVPq+qaa3wNu0xu3vY8KtJtsL/oqX1zUUO6ojFcn4DciNX8m6wV2Q3hFjhpJ
oWcdP4GN+zM1rCPODJZtgEDYuRiXJUT5h07vjUk0Zzc+lSbBgzYLAkHt9t+IIaA600KFbBapdl+B
9NUu2QzwmUrsww81uswJbOMXwKaBPsx2K0FrH5ZEdE46ow8R+G/SBpqvVp187CYgg3xGwrH+vOG7
cz1qra68Kadd+oBf3iXW9GJIUhguhFYmCKppu3qjsdJHT1ttCucRNMPmpgvABTe+5HXYOI2KqvcZ
3bD4KpfyFK9OX3wfmMhCxI0iCDR8UtHRb3ZI3Zhf7XDtwgTcs3VQUiyx3NapIl+ewJOP+p3wD0sl
fecfPW4Sj7PTnidMzjYlVZJz2aBZrhgYSUCKZeYi0zmKifBN2/KRifPkXG16JjcAHQU/aPx4AJnw
S3HqrNwi3AmHCitPb+PX3wfzmETjtYONXI0PD7VcAZq8ooU5rqxGtBTE3HpJWiWLovYWoa+cC6Cy
28B85ORudDT2U23k8WG89TGiOO/zE0M24BQHOXJR/7BgcfexT9f74+UXlAgm9LSBdy4y6D2BbYbi
7gc2uAqwIecbksXWP8dyLZuwrRv+CwdwVGEZpNebRyi9/Hqff2X/EK9WRw3w5rngOrBXMfvlCjtn
SwhBAOl3RkFRW+/yVkYcIWhF/ZpNeXAWgyw533IsmFTys68MxRaMeFyD7n4ZLXBx1W7B8p3GuAzo
SUiX8sp/tjZuPEDHLQ2reXlT+yIabBUAXGK4/uEEbJnzg9mtsOfyjbbke6IbRgoopIbUZ8H3OQkT
vAka96LdLGlHhAl25Ezy2LSW64tNuvbCxJTcU6vYXd+583aroL/iV2uqfLYJT94oEiEgPhp9NgXe
XQJw1oR6AEmcfi3ujgDkw1FJPQOI4z5IO3oJBWfhmUrXd1cocIdI0mEkJm1bJgVT6ljklDpVl0Rq
mO8lfPUAhEYvU0uRB2zkmh1N5wVM/HrAsTBiEzb41z05yJed5PnmU+E7ouFGcNR9H3hKhPG79ZEb
JQ5xd+lN0M+XDpT1OWAeZArPld8sH91+sLrcDg+K+Nji0azjTkhmW3wZJynupqNlTdhdJb97X08w
t/SAu3R2wrGT227aP01d8yERy2dLSeH9LADrqV+RN2k3MYj0MF9/1B93TjsKZlVVrJmsHUn9e4EJ
iz0O6X27i7MzpH1mszEct9o/yUDulgT0dkEttT/jUxjJQFhurE5q4fcrOxz4+45nUHqs5ZLk4EzT
1Jysp/WPdaHdZeZOJm3HeHcNXsSfb1gD9xuB8l9a8Eq9vTb3DpdgeL4lBGBbOz7yqBzRPVkhmYnb
9ZKqvp/J3ICQujZLX2rSTktHNN3fKInqWfvhh3fM3sIa0zjZki/0x8gOaE54aTldi5VmQL7saBYD
Wb8qqd+QXlGXOZHs8BH1arGnh9Hg9BHkxXEZqLBWFnGYq2X62AOHt8rNQCBAtmCztCY97SiMFJm/
87iRkco1/cBSAHTB4Z1nHXgd7EmYdK2TYzKvPV+bwqbr4UnGZ8DqD/04yi9t1TwubS5ygi1464R8
jDCVm1Rkq2nLWiawpjBLJLMAktCRXNZ27KwybVT0v8RnummoY8Qnc1FyQnzcOpwh/DFD2yZRExWm
9nMP4gCfB14F1NtCQKD8/SUqzzzJzIhzPNDRpb1jfbAeRwZMFfi0MyZ7/WZXZcr8CJtJi7Hsunyd
xh/O11RSa7r90pWy1NbTLOAaRo6L9Lh/c9U87NW+YFdT5CquJNAwhjN5HYEbAHKkW1mwAibkQZg0
aNxePVMIMpF7vtf+HAziCmcoaEAyz7bKkJvnhA4wyDXD/fambxy5UAtivfeCxAkkQ3PGfZDyhH0C
JTBCtAVjQ33c9TD0RO+I1uS/vDgbXcI3MCQSwvy8hsS2546vvmluXyeikxa77vdJ6PuzwyRbBSgF
XnaSrjJgObD+3TteFbDj6UU5T1TbQRU7u/vFl0+X9eJ2w3NypCVN0ema4eE2hn9AFhM8Jwd9wFNj
wXBt1zYMcr/z0H+bx9gASybtm3fxAKmO3r5pvi7UdUgU03fvSxgzQ/EE8GknhEUSWzhHPUUUZ2Eu
CA/VMxd0EWJOjXthg87ThSurchEApgSjczoxbCtl+msEAwKvDT+8Upq+VjRomRGwQGWmOVbxrx1h
4B2LzWUTN9m7ADFCws5+vi4vqFndfZn5nsgetTF/Za26xZnRLex5vk6YmHOFqa3/Ob0AR9yIzYeb
GFGYu7gPQKPxTIJG7n3TfxosKJ2uGrhJWfRGeFmi5R1tcYh2FPfmMPGsLstoc6npVsFiYgr41Yds
mlga0n12AEl/U7/Z3aZLwebyEaxOhfwVhu3bxDew/yDkb5UBd+NCt7odSQzdabuI0SN6FLC4MkL/
UyOlWGc7HaeFIY4uyYTXnfqfrLTZ6RsJO7+hTOK7wx26xBMxqA+6JQ1rCzxSkkZOPoSCwRcTm/BK
H6Fxbjt8L7WgMpgYOXoADXWh2ay7Wlys+UQQ5QI40zNWXP0tDt4y288goWcdW9955S4cqXtHPTdA
jlRjQFvdKd6GkezZzlzPSVkIRyh/w65LUufvGPJet9wuR8r784tL9wWro2iJeB4+Th1oCz23VFrz
BBQtTFttRyXH3RpJGEpJ0bEgu2bRCbsHtUcQ4JB/ocHoElWYlerTRKAfbr91YVhardf3FgoTlg11
O/DvaVammORLPZBQ7GJV5achAZzy1Kt8k9QZYFVqPAgIaCf7cJMk2gSiAM88upJUMOov9StlWVP4
PKbmNSUUzrLEr8EZz9mmp1cnBwVjmjV1hau8rbjIwyR02exq30LG1f0qT74m+KvEBCv0J1Y0YIWG
XaNsDthWk6GStilAhX9qxoR2th1/AJcm6bR4zxGz8XZRxYw8/EXSAf0R0ywjmK06FRU4qNxiWlBk
Zm9+nTvgldsEBxKwLkquYb2z2QNqQcwxF46cLQXtYxppuYhgM0xJsExq6JjOdm4YHv6GLR3XEWbS
Mboi5MkGGin4iHvGNQAvVO7ujD64n2wyyI+GLdBoVJ15Hdfoa3lmypDBCV0OQGHVn4VK70dsVI2X
G1AOX2ZGOfOTbaAQ0hxD7XM6UEJ/PDLiVynUUtpVPmYJ9TlSeM4NZsR0rkY2UEQJ47gRGQGTGLWJ
0GLKj44GNA4foer6Q/QKD89o1dAWYbkPWUSzNtRisTmqfN+1P/S8Krs469DINWpjwNboHHdRtw9u
GeZbeTYMzckc8+M95wxJld63cWwKt33xGWZ7QOqjwwEYWxTyqIi2mKaiBruTUvvLOnPmncUJMCRv
Nquj2Y8g0uiRqvZi/8rB0V+6QMhRNjNiM6bkarctF2fgsIibidVPRzBVhEK3m1fYZa62GyI+oAjB
kuUG/jbFgjwW+tT+3elz6yptc5XuCnPi0ETj5vkVoe3lfCENlMT7uSaZKLB4SB7kjvRKG0FPsXdS
OgDgR7gu5aa1hLY7iHFP2qXf8HaI9Cc+0bjLTvFvjnW9zhvHOjLNOmZm79y9uQRzMmuHReyK4f9I
Gn1RYVIg2UnRVrBl00SJKniTiwHOpe7nqapYFKDT2qgaI0QwtJCNboRj30pp6dptkbkSypRB60FS
+8g6a+LWLV5CzduGkeAunYg0I8fczaGomM7mpGRi6uN70wMkFM9KdEfn74DJxKMHcRVFeI1SgUcd
bVqGsNXAff68xSDfd7+bzsoKT9/mac7q7PJg4O2mfUo5bLVbijKxe3tqPQh+HpCT9Cs4tCxHZJoZ
pxu94wiPPTm/hgi3Yi1/hysYgKH1c/O8bJuXOAYNYSW1A2LtFmZrJO3ourMgtQuoOTn66FujxFdo
DYOFPzMMjLe14Dqpq2DPmL/7iB/GKkF4vYY52GBphhTi+7pAeSNN3ClFxe9rHhfo9qTi4rj4pmNk
qx/agCSd3dNZBVXS70wOF0GayZX889yztB6+139Xktu77CInZiLXAhB877aI229vZ2Ru1ln8TSCy
KhEbqeU7juVm+Lg+xLZ6iNlvsiP7eMIg/KoYUF98O/3gevpgOvFyqk7Tnj6I6OW+UWizwpS5iYJ5
NbxK4yO63Ynveu/93tmEcxgkQP8a3nWKQ9lmtLZZLJ98pPlOcD4bvxCaTyUKROCEVDW1jM4Q/9yy
q0C8rUrcsyzJ1IU9XTgwM7byLj27aSKJwBdDf/bR48opSStEsQqzgywM5xFp6+dQaebmk1Cp3kR+
z0vN4KTaHjxEjDfsGkMsKJot4JWen25Zs3DGHodrOotDnDq6GPwEkBTpu0FqGovlRao8HHD9rt6z
hwx0alPhLH8hTlP3d9rhZuQm1s50PRLqBLm1VPqFh9kcz8JZtNsMFAXdjyXVbxEqtpsUIjRJWm7O
9IybyTPtk612SIxVMexhkMSw2TaThf15PWnGl9dmXOJnVrT8YYlu7hbgwb1RhtAbu6XwxBWwF22Y
dGfP2CPtXl33a533XjxCnQQnw8T/qaG/52OFKQm3r8AbJqNmJpvE1rBkK5zwlm++SICUp49KMr+s
JiU5lcrJzaZ/l+w9FyiyfqLyem3v08LWUKQoczB0DK3B36fokL+OoEESgRASToERlEvxI+lOYJyE
D2f53oG0NzklYtASyS3Vd3/4a3Gj7Sri9GWlppNdB2F6LaniYVyNx058ItWxE26L0U2gP8UO33gH
c2n5kJJ5nhcUrHbJuVdZQiddKKDGDhRhr3t184Gb2zbBC4CHeiqJadG4Myj5vtKulYGPscM58roK
xid9iBEEoDGlUn4qdgq+VMLIFqQnhCMF3R8P6uFrQIijChjJoCR+isFDtq7NQhPoFOSIoWk5mUHu
4Gl4ez85Z3Kp5dqFfOMfCgku2RW7YrWICXkQ8S3TFBy82g8HQUVl5O3epS0KuEwgrzBtKV2lQPOx
jMj2UNOCXu+I4EHhfvrYeeRGpay3JENnGarW+FMf446ntuAKnxFysShD1/EwNJzUKg2uqUdKse4V
jonD4FZpUUsWJBpt7UX4zPVwBohNi+Dc2QwSiVuzodnOAT+q61YMmatjEjwJ4CJud2unH57pATFz
NWN4VqqXIzmm4xhKHqtqg17kll99nYVVzNnjNWhLaW0fiujUsgYrxDIKtbmKnfyuTf7my1LrS6QK
JP1Cs0NTc31Wz08hpoHpWU/z9cW7McRnqdE2J/sQ0PIbnJjihNOplWC05yADVfPm++oJ6zR1iC72
Vpz53VwODBQIYmmmoZbkQSWlDLR6LHoSjth9kw9FEbmvR60Dtz0FUb/dw/DhdIw8U0iveL60kWMg
Mk8/uhFnnLWVqIdxSpWefOmZ9sK/kmOla9+lYbMS810tLWSb1Xpl+3xIdxIf/k0KmeiQiSbf1b3M
b6+Z1i9tfclyxXd4yyqYRu25O3cBprsAsqhTwWJzeaXLO3NfWidvw8NoghbvnPtDpWoSzpIFAGWW
/c1OKTy4hEawOtlZxLDVfEBR7AHs2THhkONxl+7LwFfbbds7DdIeXPmDH8jQm1QQPWcTwwrJtlZG
ZEp+CpeiH+EDQgf+0Sat3Okz+slTTetU+QwYNmqiZCxEJqisMQ6APw/YlLLNjcdH0vAUjG/dr/xN
d7P3lQ1oURMve1helhzC7JRze69nx9rkW1UUmlccMwbLNZMPsuQMPlebtZ4EGBsmR3sE/tjHRBUI
oKKpmurQORrsk6yeX0VbqwM6oKk+P34cNkK15k9tnmOoYdy9pHbB5VpeYo+v2CZRnfi2uhYKn6AV
Q1vy3tQJMw0kwNWqIE3hUOkEOjZDdn6vc6BOHK8K4dwZVqtB2SKsaIBqdX+Qy4y7Gpu1ZuKfz9ua
TiUvEgBjMz8Q/PtKG1WjHDIyOTl4jf/vPcMJ6CubuWYk1iRwh4YzWr4VNcPH1/WVJnJbRXHvJUK5
gS8w4bSpxRt3k4I2iCy890MCFeqq1chfhKWupfGTV91Bv5zdKcxIPQ6/N3pXKnDWQ499mDPpsjA/
0XIm9ikhwy7rnbdV9m29fLrmSI++NoJ/Ia73QRuVlJZm+pm36xifk8JMQFWlQ3sfddOhwMyEM3KX
WBtPZqZRRFRi4C8g5it0BHyhPmW+GJUZgYOJ9SqwVLtEGTvtYW+U5gLQ0FZN2fdOXrRGfiedMfTf
zUPNkAcYdN8yhA4ObIsFzrZYENYMfSXWr6+SOpyPFbOhDKyh5K51D/smU5rsM7vaoNzhqw1645z6
bI18j3jFRTdt61cRaq8dbPzKTNib710u15pK84WtZw2G8XButmSOLYYTOV0H4oOFqVX0WLLo4Whe
H8+jgv7nUBl+X4wie52Ebxr0UGArK9SKA3Ttgy5lSXlL08LA1YZN2iO+WRQEWu8fS8JX2Qzo7L+s
1Ntx9UIfikp+cAIP7mdqZgEElxVeIg4jI9gwciHIfXfCOfhEskKbKUP3we+KXSNZkuLUQnW9Yrf/
dGjC5wG69Ugq99VtTX3vYnIVigaWwLGJcsFnW7GJtlRsN2UaBDVBQQbbpbeMaNDqFM3aoc5n0KpB
sIA8IG5kXy03ismCTTGmWGuo/fEIiohLQo1SX4HPtONuuv83GK+Ay8BXUQPXJK9do87x7uaV7xVM
D49wjvrmG1CoQnjr9A9SQr4X3/iCvIzgFSsl2aAeqozRJwvSM5ZOMKZq+gjHMZ1mk0XKNXje2I2n
aFOsKDj7O2l+8m24d5nrkXoc2ck7VwTDxWTpkVk/AnSjVDmf8GL1mPACwgEL2YCc0jEvS5QyS8tx
YPsQVFQTOMt6+5PfvQ5fK4+YIDXMnqZuSgX1kmLo+yZmCNQnFqHoFfqUxT5EmZ7ZCuAir6035XY1
CpB/0YIsc1KDqS9pdhlUnvv/7mBwJ3J5stbUoecRvW7xgcdMP6A1iDeodSFCywGRzgYgOqdhEyS0
+EJmYTsKVCbjw4KlU9Js4V3CXpniIbY93j2+GUo8RnUOUks0vVqH5HQiPbBMDflZzzpiXhDg/C0n
HtF/d6aom5vOnSRb3wddPj0nIDiYil9WHWjgF2nBymW8id4Ll5AiNCCkBwAAXMHSoFNLO9yKPtzT
TaRydlxtZ4EhqIUiPB72LU2JvEwyEr1XHnZuyPw8uzendsMOPYFR3rHtvDlLRUU2nYDeAcC6OjTA
VXlgIW5wpaj5qUItC3H+Dp3ybl21oOfB0DJx69f8ZWjV8ZVea0wci9uVvyf/uiY7eOZT+7zHWHYs
SGl0rjjXvM0mvOTWHjFwcmbfl1fzanB+sc1j94ASx5YJaYrhDOVzw5krOBp37KoB8VSgw0F8Z671
LI15FQkARgNS438IMbNxo0nynescgYiV//jpBOCDah4+nwq7IXZLOGaqvYJa2vegfyghmAjw6VPX
xMuxoSswLRJQO8EZPgWgQ8/Sn/NwGS3vb4sRhnzZJtc8brj+KZlvH3guBATQKlTzlZiezWgbXIff
Iv2ZnBkckw4Wkd5H3pKZKpkmkZSD/F4g/Es7uCCYSEqhaxETsXKjp19AZwV4BAxXcygXtEcbLImC
v8rUwZ/3wVvvx37JX/0YmomqT8PNGTUup+lnDWdE6oHGshQFd+syzNqXqF5KrDpRaKfAVt7hp+Ug
YH2+jRfUu8Y+TMbLQuuQQXi9aJrSgB2dNSQltbAQ2Xmj/sAnZedwHL9a0D1YGyMf1ivfK8m8BZsa
exlv9kp2gJew1F3DlrEElt/mwUknXRnHZnuBhi6kkdwyVR0HW+0dRbHlfsnUB79/HxjXieFHRoTx
r0lF8a2sK9r9DsA8BwAbWkQDF7OOLgh7v0Gws2eJfxzbfC8kW59r37AF6GVWVEXu3RwVFzEJVYWG
O7JXt42gGA/1/fE78fyshMCk2sH3bLO1+DQmha5YsYg/LtcZAn7uIExENfn2bknHVHB0VxjoWHU+
6OMG9eMyT8rQluC8SA6KCzFrBOYYXQRU8Z7n5MwLG25kHaofUFG7K7r+OPSn01i/h832VXOVdMbp
vLnS3E9NOIhWveo+Y2RQaFyvvadbuRpgQeujCkBjuNxDewOBIbkE5yf6pjxmtKluhL5t9vtXuKs3
tH8p+Pwlr83dQviTrHmM8BpP7aGAeu2ycRP1W2203APitgyuyFjj/zaBkK2qeOcgzRoDm6wiHfvk
2A+b4Hoa3JLTENOBvsriMG2rN55VHc9XKrbGba3zksqFBtLDSdachk8L+bBJ7BhZRi+6fIWz4Ly6
uL85mp+LT/5ytEogltvilCC43sDIUcV9AXfZaZjJ/ImVx2V+2u2ItEv0erWR5WL2C+m30T9HWrAs
GPqwD3OOY3M8dMstSYdak5dpNweICdXwv5hbEAyfCNMBkY/doMlbKyg5k5O57sTt5DPz0gqMqzSG
LVzdp1uEC2/QhTutvELdMT2fHiki61YFdrVl7oip8kTniC916Pv5VCsQbrSvtJH2RFU1VDL8G8ng
33bwOyHFIzSW8X2OzgLFTPaylEputhA/JDFr4aPuXr8W1TO0tT/RbJTxPvryz8wJ2P5fIszZb60E
Z2RpLe0yyJWdiVZzu6gaPs6N2Z3vEPlBm2W6kVusT8K5cdHnYYg6YwCIIJ0ldJDgrflb8wlpQ2c6
z8+TTsgeAztdjztUrSJAcBTqUd5DOGVb6v67ssZQ1CAaI96oP1BCcoBjePRzjy/C/NqaSPiOKERV
6IQOH9fvzJtUGrcSPOzvjL/mCPK89zIEozxDkNnNwKuRDJ9lEvE3mpMUKMlu+RXhE4aDPqmFDNa0
wPILuyajxL1WL2E1f7E0zRrMDTujSA9QJSeZKoqeZ/H5iHh31D698BTdomZ+aMgqaWmChIpAvdN9
BsLCcZgXAstqQPDm3SwKibNe6p/r53eYRauaL7ltXdDhrJ5XWBrvKpuRIniBYaiavXYLkrCbzD/k
e/8MiciOtzlujq1VwwNMlrxbTyldT9EBuCAhNpgCsjC6ThwDLqrf1PeZMhapqVw568pX8wSlMMLm
Q3tEPvE5RZCjlNPX0MpMSfNYVKdjbLyNCUIFKlAGZFioq5HQmAToZcSXDTCD5HlVPZpTaPZdDJW4
rN7K7QZ3O5ehUlJgaJQ2eb5k4zK2jBw8f1ZVAtPS8ydIH4sGX1l9XDMC7vZNUqJJuIXtUBY1vHGl
a9uLF2QqFf+xZuEgKt8GvSamtiqrBBttr7lDUO14+K/kAz2s32uQ4bmuj7fS04wdeuZSv9fwswhr
OTfMDyxboPW1OtcJ1ffdwF2qV14tn4+iKgB1yDK/3XovzDKyWoc4NyJ9heuK4ENWiVQrnG7u9foH
NlM62rOTcLOfxf7svprZqgRNL43yP9lUfySjcO3K5xECpaMXEXBj4AkMnYbmWp09avG0oxI6oC2O
y7OaXcbMUIV/PuCgnnf5/HWZKPDn0okpt/x3A4Az4l7wxe85di7lPpSx4gvJ8txFUGs0DcBtG9B+
37IzSkMFaOXTMMqUQYmUYT0VXZU1B2++D0tY75e2DhdyS6+xGnBmajySnOA3E15zrmNh2B5EOL6a
DjcVakN/njrqEoaviJtb9p5CCERmY1VX+bj1/rTIaGIKnkXaAfojap65gAGdn1cI181WdoJqksJs
7ISIjV4ywaQ6j8SkB5niyqNpg0hVnY4ds2Anr+eg+lnvqMrHDMToIXHyu0e150Vpk0s+wCPC06Il
qPE8aQe5kS5J7HurqnZQdRLAr79+6vuwR9X+Pk6/8tMa6SxJQC/3adnC27HjcbTub85n/qthRg8Q
at+gPpwbyKf1RClN1+1xl5d5XbseUZh+vHFOrJKeLX/32K5cLPlFWnu1BCIJGrJ51JK/qNDZvKrN
y1a9RxwbrRaJmI60+DsGAqiFGnWgCYEZHfIXI/fJ/lnGfoAPkxJTU8CDrOR5jLWmIxarGaF8ZKfo
WcGlZqvJs/7Rc/ypSRVT/sn1Nsq4YkzN8bRuGaOh3+sD9Y/Jf+tpE+vhXsAMMmL+Mq4F7eD4ejEy
sZn2yXWN9h2CtRZmDD+R1o8SOmXc9R+mnzkSQYIs4OiAdCmpsrfQ8sgurFKSQ7isovR64gfrnvrO
Rb3KbRvm0Sa1jfgkC6HyAJAIB1MeewQXq/EHzvHk2WSr9faKUKLcKK4rmnyCP8gL+uebS4X99GkP
EeGIiII+AgA4MIlLMBSKccnLeVIHNkCQ4ku92VRRjCUK2PzuoFS7xmbcuZoRdfyGsH69bQNm7nmL
B5OOEZffx2fPU8w1GE23BE34K0HjH4pvdThGTyZSbqDTwX1fHa4y4M1/IPcEl0dp3Kb/RErzAZ5j
ltyhG3v9mM+zZ9WwoMHpVQnZxFnWjUHR6Y3c1rmcqHgw/c1iLU4bHYyT4P4tQcwDd43rVty/x2xk
SFsXKjWVzuvQRqQfv1AJ0JtLo/5fe3CKAHwWQRO0cfIxG1TZAC+yGzmBhBmSiotlr7GXu482rA21
M+/1qep8ywD30dvotABk/TYiTVBD01ZP74vv8XcuCBU5E0WA/qyJeWdVBz2fD2kF1Pd4xDPBANqb
gLA96vjOEPDQwFgbLyB5qDjDjc2K4t8zTozurLgOJBZpktqGfXoprgzT+fa1UFmf4IxfHl9diVzB
jpJ22Wr+UAEOouK8hfKsWgIAa9Wf7Cj9eZqinWcbTZ5102tQdIGlnPGhqHtY2K8N6fu5mIkRSd7X
U6melU8IFJbILb71gPJMJwYt2lOchPz5Vin2S1ZjgCRJkXAPe3nY107HT++VAdqFBJMPw7J7yyBP
F2ojRxDbzV7IGpVNLnS7joRrrN9Cs6a/uaDP5hZPodzzIPVA0Yjxk2/gPcKQRn0WdGKP7x/2QjFN
R0eN4kWtNH9Jzjw929ka7vn5r5xcF5ZVI+uWkhuT7RiziC7w/fDKjyOKebVBm7OTUJB+awTnTzNb
uP3sxWmzV3IRawbgdWWKU5CDde2ZeGne+0jRqnSNEdX3Xttk0H7QsqSVpJIqRXvDkGkvElJNkNUu
M7s5K1yla+AdzeWMfCzxXMUl7+AyC1LGxbuvedOCS4z49Wwf6NfU2OOUnVux3gMb8A1Lz11WqJn+
vkEy4QjP+7UcexIs5ADmzvqJjaret1nyV8YHk4bnlY7x3qHmAV8K04rW474hJo9uml2EaCRRCGLv
bfiZ1L9rQX+NU9u800ViEekbGjwL++SvyfWJuI4SjztRTSmq5VweWGPVWXH2kBl4MGT0RfPFNN6y
iB8EuLR9hbDeRqFnc6mH/WvFARsmPvzwsgA9aL52w/9oj3tKMpEuEW+uLTUPLhcMFD7+9+f5h5AS
udcvhFtduryxOriiFwp7A9aCbigaX6giBtPhFI6HD2dlBfGTUhnOTZbqZOvjq9fBnDKBOw2evOM4
KMx9qRAZqinPvFjFC0yLzfff815CfnoVqQROmihTaLeDUeozdw+bWueJ0G9qHeJ0Dq72VTmpYVUF
mLCUaPEIxPiaALTfKiRG2y3PZ9nTNnwg/9fjeQ11TD1emFEenY13vPpjgDKqA2Bc8TDEqCY97pjp
bOPD14IhmQfV1QpJBqcMpR6w9+45LZ9swWh8GQCrCnHNNz4VOb+7C5orSwR4CoJZoccBfGWVe9un
GDznB+i0KhSkOuWyvCfxVtfp1EOWZcUsG0g5OR6eW+vu1hSfVN0TjXt5dD8wNdCC152qvo29Xmqj
Ttu8Qa4riyWGYoMJ/AyyG+y+9WUVWX/147ucMB/U6fKZxcQc22feYW/Omvqw51JdRLXHp+1nrOBA
5gXyilr9bBMJCMoKdV8PSC+KtMlAhE9L5sNPI6WnMpXh6Et2QK+382eDY3bkhFi9zruyutCq2mHX
cuHWAfxc9o8UwO3PG9cO+0i1WegRVnt3brxRlP42uDOzAy+vAyXckzfs/SY4nE6QiukhLrF6TBtA
0rh6dsdLXa5WEzhJsQhjoYL0vv5C7icorbrB6kUeUHnRYh7Ze/A8DdBIWO9X+cSJ4hyKps4YumwS
6oo7yHUr7rL7c72UDE+u8jU+bTnFn2b3vybivIP53whodoS5m/cFpj9Tkca31Xluzz686yWnk/8v
oUBIU1Rd2nJhI9iqKR+EQ2/T/ut5MZSE9CpgC2lsKXyjE+aPld3oEFRJ0n3/TIyAzDgzhrYasG1w
Wmsl/JdJFkLvDPQ5UQltuUDGYV+IG4KdHJ7mFbDJ15mWG8OTMIz+T7TJkZFO2oUd0rVmLJssZMOy
cKLegxnc6D3jYXmi72HsR6TqXxPsY0Ajou5aa+2ELuzGnMXZsjKEMYculeOfkcdvZQFnltk6+clt
e7efSiG9csYrhDNu5brG2kwU3KOHGX+8Il1VwyqSwo1pa/VluScdk3N288bz0xIWfEaUAnu6t3Nx
nnLl1MKmv9xgPPnM8vsK4euWpSlJefGSy8xuJkp1u8QYpy54Ry3QZV65gOnGJsguQXgzUBTsTwcm
AXXRXVVOhQQZpHtGum7mFBAx6v/mayaMk4AzNYxHXi2cDucRWF4GYZ8POgDm3oIS+KB4vgwqdcSm
MNeHvmAiBg9z3HIpwSByhm9WP9ElwlDVbzReJGfEA8VZSOAcnZfFMunJUl2EEQ+mDJzzWIoEjHHY
1dELGl5WwFh+jrKxK5pJEHclqqrTWOX2OVUbCY5jFJlzUb7JQvApUGBvr2D4TQe2/2GFRHgUiE86
phATTfh7pFjpUrnt9KuV/JpcfZLxVMTTjxtzOOE7JskTveHavzGyb2Ia8DZmKjSvRjcU5mzNQ1pS
eAlPsGtiGH3y1A5CKC/Ie+OnEtwz5riyG1kLZ2vCk18W6Ko/g5TsSueqjDHiSnLglydhZeeetg7u
5+6J/3XXcrFUKeb3vxgDHsp1F7qcAXcz3ZZHAHoDCqi7AzhH2q2/6QtReYZAt/mH656LdOfHV77g
Rqs/Ik/4t71ga7Zjdf1HS5TdOPSHksy9xF0zZExAfCk2326cCqMmGFu+a4TV1uusY5i5PyA0LsV0
xd3kH8OEDFsZp2ZEmXl8VIVVxlR1409jpzybX6ToJLaszsN4vthS6MtkM6C4roMWl/EUE6XeD/Yz
bXg6zUatw8lEbQFF3Cj9F0czeOXW3oB/QwnvU/9AuQvuAKte1wEoxN11PXHGI0CqZk/UtUoJMKV5
JzOGmDIUkN+8b3pUM6X3kfLyg+HICvGZrq6Maio45ZL+3SD2+0GO59ZQwGGupI7ofkArFFrdozOO
MQDqaPfYIDdj4cVCuTUQfB1DxuTsGVP8PXBJ7l25qESZuABsU7wuhuU+p6jYcauxc0WZOqfUYITm
UNhRWzkaxFuYHmIxJwrbuSsjX+l1TL3PoBuD90iWRBvRZubQzzo+KJygMjtAW3JEPCbIrfyQcYrV
8tn4cObbFOTgwQgGgtW7I7v+DTk/gDdXMz0QncZK1i06GbIBmmaKxryR2xqEOg6r0AncgdSw41Jz
xEt4xFrDsIazs9IgibiY5Huqh3RptlzJsFpgh5Bsnxz/V+u9C44UmvNwDAF8KzvZrrL7xwaXIt4H
rIFJvgQIXhc0Au1/Lqtnw+wPHeOtqvhz3ZUnFoskTvVTMi7Thh76dI70Zqaw2KGHo8aGTw8nylz0
MQ0KTsMilijUhca2M+G5zXZyrpnDzCN3K++nyYG5eP1U+bBJhBvvjDzqhNf62lyGCYcaMZv6VqHf
MSwzBndX+5av4gtcyTBIWEtH5zXKvvxWGiIEGkgOSKnvBCMgnO9lnw+qTm+k6WblobpZk52YO6m/
1YcMte/ALJEoYhNc1U2jSn50VeyQCUr2g8Py66NoefCoeRaSIggfLqQhlWTYoW1c6vyB8cvF7JyU
AwgvuflOlO/6LKoEAGGJ936s6iz/q9aoo6hvWgMTX7sT0130MpIrhq60fjBcwM0mL9JXPuN/w7o0
nls1Yq9598KYUAQlj1yKMOCFMBLaXFjSIt/PcwXv0M/3VcbyVFqnZ3AEUYMV40JaRgAGAdtKnM++
96qgYs9SrglxpCSg5abldznjMXihg7hJODnxxCbLrsSmVovsV3scYA2SRrlC+hHBDSU63w7jLlof
5z5hvN8fTSRwKFs+CWXphr1qIOOwzsOp4afmhb5FxjtYAkdB3vD9YfktRvZeEludRKw+mgDYkoL/
nj8M9GbvgeNXT6MqnEgEmjfxc3wUvM2c143RhbHw5zmh3XafA/RrsZUSzN6S5BLvoWl98A7VndSK
x5rILy9O5fH1Sou4GDechHr2FaNdl0zocYJ628HS4KZvsOVyZP0NdEfMwU38VdjBc1/SXl9WBnva
21TpR3zp3dSBkNr8bPJuHhGG2kRWCvAS7BgMjRCMha5MMAx+YI7RNm6uyfOnShxDt3Os6N/hfC+X
05sjs5DjEGkqodHZJ8XHfUNC5XhgZfCuKnrm13rorremcdROmPq3exSgWv9qtCEXltCSv/T4RNFm
TCHarVZQBDSEIHRTbHGff8vnubiEmaN5nsmEfLmaSRb1XHZdMZjW/N6cLzl7UARf+qedsjxFIwHz
juSx2VcGDlL4PcUThDt9mD2OZFyZAZ7YTBB7F2IFziIXMrs3JL8iMPHhjvw067MQN6LaM9EVXN0N
DWiUm4/uPayFqRMEbzfHbw7FpRRKaOpzHYV3xvQ+xUUBjAbItBTmGh6faFtPr/3zaYkPWqwr7AMe
SQDmpZMcmOTkp5tyFWWy+xKLW2XqwijtMIQEqsGgMMpZ1srr2zzzwBk56Rf54qiGuoER6D/AZYBH
5FaiHI/6rmngYIK/zEXlfIuQlGHDbZ8aAhRBIEndESS/gtXUzCECuPrXVMpJn+gUtdohkBBn678O
CPtYfvd3im8NEOAyXdmA1XKuOTZWcfczxPgtFpcAt77VM0xRTJPTcws4JOmkcoM8ppBhTA8PzuoW
/E2xVslB2MkWWcb06EVGE6pKpy1dV6l6tYqeZ8cV05ZG7ZLf4GwY2tQJUZzXcrorn7wzuRsB/Rk8
1eh2JMM4slBBnc65QjRExa0ccnPQ4CSSuRWjKNTDhe4r/QitvPDnhD0W1lzyK5SHOvRWIFnruHMI
C1yYtWbxgZJUcJizpFHS50Jfnqs9hPo/taYGgwFxHwmtNr9EZX+SKrx+5tNy1ChnNeW0NCf4norQ
vENI7GurViGrzB+Gc++brRKW+f0Fp5qh7mkMnEo0Lb1k10xLdb4x3AxC732COP4Sj9bvoWfevlRV
NfN69spD873NnTjJQlQNPYypp6p69SJSp345k5sTtS3SUBclvM49c0LXSyrzVP+t8mwnS+AkEFax
E/Uhi8wduM/wxk3/CAyJRUTDFabcm9PKmuFDsJC5Et3sKlGA5GtanojnRGduck3xxbJmF5JWZnmA
hyuh5HUEPFH7mnTjENH2dISiJZ9lYJIFyPiJEWM8GRkTDBPRNdQA4C/AEelYa8+kIpzTT4BHJuyf
tGV09nRra2b/Nen2STn7ULiyuQOmF3UfNzM+xyimknutKAjTNdBKiz91ayHzO2ifiU0u66R/nt62
mnl+4uZ3xMluXx/FoMqhgto5VDFV6tJS36j5ug5y8VwKgpaFQ5f2jPVhxV27a0UJA4Z2/rdmM/AD
CyfD3odglmrUWtNU19r802A4j65/s0G68k7txmoNeTQFZBholrlgQQAxKcyED1ZgrhE0h/2FTq/7
KAYbRPk3HdS4S43cK54Ksaiau9l6gfT34UVkulaPRoFM+BvVgyrA6ePhxxNT2X/KZ3KOY71NyBAI
rpPT/tEigYJ9Hc87tD80psAA8NuHGbl3/qC0OWDzCAvJBmYXF4PnLuh7/v/KFOSNYNPdGcF7jUgr
pECACUlU01ep3ghW7CBr4aH9pyMyR48vpsduWwlAkgCYBItEic1huF72tcZjFoHXUYQyIBS8fyoR
AkrzqDijQ4Us2mQ7HaL/RlKBQiTaWdgn60hShU5upN9Tlm7DFMj/hlvkUVOJ0P/u0l7/tkQ8PCzR
iVpC4s6B01TygvZulk3xe7sP+xw6YDFcgmVFi9JEMhmajJ+RJJ6LcxLWiir1IOFGhap3aqcy/Swl
EsR7YjwR/PBEQg6Gi/85pexNYf6jPp8OCj7Q9HFV93MoehBbj9WA+NlKLyl2VNTGW2R2WD68KQfu
bGVERBY4mnWc0+ad8rRJtBi4QTwQ12PZOYXs8cMH3Gtxr5E6dxtuAGADX223UitOYYixTT98Z133
EC9GWJjL+ZT8Fey496/yt4xiHVJHfAnJoSryZqHMAvZbBCN2BAUTeAd8d4H+4dDboBzYfXv4kjTO
qmm8CgplfgaFJG9zPQT8gs9vIMAw3Cpue3fwj6/aRUQzv970CUV3XK+r2+X8IP3HCxD4IySDB8EV
9nolYBy2B6D0+nexkHF495+3wAtjqWIfOIfsVW1Ngfv/VuR6aaB+papc+rQQ7fb6HEHUkvRrfJef
nD0jpcyflA07ZrzGPR9r8SwjxEz9SO+csXope0Wqbnt9/ZakNGi596sdyb93T5cGRiHP5CFuy+vM
1NvwhL5Vyx79qGZbJUsBLVqCXK3IJ+zwcQdXN5g9J/hqi3KlH9W1UdvalnAgupPY722PmXPbxqkP
E5FrRfcTz3qW8Lrgp+ROepYZBTF6Sqy60Adcrt3t+e34AJ3z6bz5ziMIfd6srRTg83hFoXNA8QX8
mhRYMLGWMDn5dN1+g2TAvqA9nu+W0Vd2pJI8gA8YCh6mMdvVFLSUxmX8n8fjcT1FoZrRsDUzBqIO
FsCEllXplrDi1I8+9qrx9DLlxekByvH0tmG98o16CtsWLWrh89z/RMVmAKqH/IS511KrJsdwjh87
rIgtg8fL31S7dBpV009uee1k6tasbz8qUCWAKR729scZRZeTHWGVZYkQymXsG0GQ3KPY+P9J2xt+
3NtM6vtGZPpbEQA93C46+t7V9ijs93DBXiHg8Wg+/1RMccUXEtK1cGvXochxYmKZk5RKFwdE1aIS
TfhP6Dr5MAr0klW297gcRTeC6Yrq149y/hK0yjHEuWVo1bNUSNM/wWSEKixQeV4NEkuESrmwTaxa
VfYAuaGiZH2qjFicbbzY1608XGpX/tRmIoA1Z8sYVzk37TjMp2epEbIucUOEe4SPG2nL4n08s4+0
N3+cbvOw5cC1X1xR9ZhisN4eu5NLOEDllCfviX2/WaJHw1JYgcvWX3ypiGOlRn4HyXoHYnGFP0HK
Mv/XxTN6y+AnVyjnM7Zwk2LnstN6vP+pTehM05l/sDDPTpwvrKZNXljyZSPqq6aMW2hxpsZIQa2u
DLdZ19dXMC+4+RXcrwNysD5KcJRUXdrvhr2Sd0f8m96cuvYUSJmtntVBuxQi1gSi6o8s48GvE7UL
rhnlUqzmuuHq9w+JpB0EUThjE5VeGh2+JOsi7SHm/B6XjjX43k28RLePFw2iNbfXK+ajXeRJ243/
zSp/gJeh4pnS0kchDXQOrBkp8qKybA2N/j+xmwy5AgyHy/i/DOa4sCtfcIzMrkVo5leHZTWpdIOY
KpjhAv/FG7yMwaR9X9eS7Xagvy7EPwmSdVOIuxa7+tyf3QndbduvF/wCK8S4K6vDTqPaBDwV0Iqc
tXg08JlsWgtpNO0stnAW6NwIIRmgLNkIjfBW0eF1PZx8kKntouGUpxwDbSynTJF972/b3CwQUenI
BFicvEyEkZ6cgze53Td9ImaVwBjkmiJ7o+XFc9fGefbkvwKaAloMzt0WefoRBT3mKHJgMbI2rA4q
Gu8yNgQHLLnNcfe4yBerMnhQ1VQRw0DjS5atlHzSxxooFu0iEBqlaYmAChk0rEwViiHq1BYYJPJz
GFfRlQXq9U3NqGxFIqv3fsH0DbMiD9wxEMaEal7rU7qG32A2VM06RdIdR8dA61pJr8t0A72IgbMj
la51qxf5fWaGCjIGzn03jgvr7eblI2lkRchNGzN1y+Tt1jWghSC/8Dlg93caPJnLfg3tbW45QEMF
ovuqSxufftjbWFssy1TwWCO83zQPKpPpI3c9nmw2hbCfSwLmP55y48E/VzsRk7x8gJAK9W7k3Mk2
Jdzvfzn4sppxXo7x/2BqJ9jvzRzeNPfLlIOwU9cHQY8ruB2z53cgK3LdEc3coqv3F3kXhhHFtSYz
xsDgLG+iTbUaLuiQNh8AwoHJkcgoG7eDxGHEdPty6wPU8O3Zm9VmSgVY8ifzSz7XaTyKDy4Coc3m
u4nVF36DVz9JXAwnquJ6qz7Urk6LnT+6MYoShYNGzB9QlIdubLLSRNO38GDZlHsUvKOjlpzg6MmL
KF6ZyGMl6EHlONfnBZWU2fiCRF6Au6eG8TScawfBNqVfUPNHy7AOduxiRiWVaE1T/YSFDI5XnvCh
pBHDL1BnPkMCt8Bjk9a/D2F8dZJn1orr9sJZ/t9IH+xQbiP2UHVks1x2z/S19KhX5Jpn2DsIjxw8
8Z/gzsvj8iFKXLKaFu02rxA1adSHJrTkTVgeK0uPHOF8Kne2mXsBwDEph6kEafUvHZGFcQRLb3RM
O/pA0av4MB7EIjEmuL9Z2AyfZEGSO+xljy9bY8YsFDD+jDb8n83bY1vmuvDKlVzHpSNpesAAT9wz
90XcZIdgKVnYa8uNAhd1FGPie1NsWLj0Fwik/Dgq6oVMUKc+0ogT4YCsaVpYrWN3TsgDC6d3Hx6M
MFEW+r0Cra266TpaVy1VsGJVD6lIng7cxWJAKYnGXtfY9Je9beZVwRvFNjSbej3jizIKVUhAzBmD
iDNWL97CLa3dRYk5Bj1BjIeQN/pS/d4O4JlwMgpkRW942atRLSKiWehmmmYL3WsE+zjI5Htx2QBJ
y5iQsyqb8EuPFcoJAsCrWznXgi73PFg8UWskAu4I6QuEV+rKSDlW/Y4Rg5HFTb+Ei5B+Q6yCHD3U
MLPHq9x3lR+7CwOp3ILaF1NDjExfgBYXCT11ZOL+iw3nKcAAK4sXlPBZNqtsPTDmXFyToOmF+9xN
bc9KTvlQcTmH87JtD/ao956XC6tAgqURmOUxTasAhtUwjd707H40gnTYOH5veM//e39F00AX/MU9
iKujjZSrOwCRgi+yuYyK6/+Y/+Tkg/WcCGcdswvAsUXJ2ALhwAJ3zaS5v4Oq2nOCG9OXwIVY3JZj
lrWiCWRNpEBBr2YbHJB9SAVlJ7+GjLtvptnB91J9aYzlYj/PSGJ8GfxLZrFme7x1929ZG9alKlEZ
nePKrWHfYAHw//DKsV9t5h/7P2OXPVqvn1yPY6bAjI4uG5g0KLTcsnWubxEsFUjW5yRX2eDvYlgS
TnMuIYis0D0mKFen5p8H7vlOro+mRe/Rl2uW+G30jHhIQfN481JG77o5qrrzcbuU+lHal/10AJor
YXZ56wasTLqQmLqgJteC7STl/aVMyPRAuo0V16A3XsTDT9GkpG8TgPeILiM6Fp6KLjIUNVdmh3ts
yt/9Ve7w8pXzi9awGkwI2p+Qt5pVobzt63s6rfUNPEpT/UeI0KdEJcYW//GRZXQ8rwtKEpg0OTa0
bblBetNiI3RQU6bV6YfnBgma/E+N/D1MZG4MFVUmeWfLD3/Olc2bOIhIsVXirVGE97P0fP9EtPAW
1i1CZ2XWD3M5WjXgzoqUW7nm1Sk+u8k2cbJjiGHWet8td0ctFsVlkvb9KaQSXRWf8GgfsBy9L0GP
jrh0fYS9rQLs8BUfN8ylH8cQqZ+E4xW2H3EL53rm+xSeIDajY4zURKrD7p/ptAjt0o+ToL14iXWR
BiQ/kPbW8v3dIm7kSIgSoaB7pNE6F3cdHQW1EhgTpvA5Udd+nmFxxn8snrQVKSOh0faEqu0yEMa3
VrDV18pB6eEuB7l2CSZsdeU+35ls/SNeV7oGqM6xKQk55BSCCwAWhNbQDLSE/bcLquEcyBP3bQ2O
ekLiCJZKI0XfTJIayTSpHQqYjV2obnqJPZCQ5Vgfz+EGK8jOgMxBGCPpVMU5Q33jPPkG+knFMSB5
qxnn38bL2yDo6/8Vd1qdwS+95XzMcI8a2DN0QNwcbxOHYYJNt6J0rTDloFtBX+O7yOigCQ7GCC+x
n8y2DMcyICyQr4JITeNOuQ+5bV2ir6ebC190efhJZi47xLLd4bBI1XLoi9NiRmy8G0t5ab6mGPts
nvYw5tzAsua8lP1j8Db0+3kCGXO/lpvsk3U7mso3Ns9GPjE0isaTOpN3DhIX5PWSSH+h2ZWnYc8z
Bkad63vjb7F1vPWQ5cdNUPtlB4XJlTqQS2kVt1e8A/iT+z7G3Kab4HYp9v3aLRumiDRl60eNa0NX
flw7n75WBfs8/kkxkJMHUmW9aWekrEbVcNIJRdxr1rKBQd7dhHXX1ayaG+mLCobteIoe0nP6KnKp
50joQoWNfFJfvW4Uk9Mg/DboEqS1vIzpmDd6gypkELCVVtN2v2dzu7VTNGVQPSMrjWX98gT1lzCQ
v1A5ptwZ2JlYsIcJRilS0bdCCHsiRts9YS30+0jwCcmXqDI7ZncV0mq67FBPbRQWuexYNtZ/2KhP
WPuRn9oNv5g+R2ATFx3lGxeaK3tzw6NlXAGV9k/xYeiB8FchktW6PHeXfQ7gJPkSec9GvKlDZcKa
qOFSRYgLYxDnBAvUhcZUY9/2spKSnlXkw9j7Cksa61r63GvCAc7y7H2zfxcv28I6ZIRa1aiQcXHY
NQJOdmWaSii8w7zHsio1BNDaystHJODUTEW1PmTuwGsOgb9JNEvh02FU3/XdGUJY6xzQCut+5MP4
vfJH4hTB3E8GTt6hgEmN/LliiLXe7yDXaI0ILTzPC9Aox18xAfEj5glSaGlYX1hFTQ5xNYCfpJSm
SPx7uhtSHEJNYu0MX6wbe40/Rzehd4mZRYR/aoKKyOzzbG+Xo1mzDeGQRVt1/nKuks9W9SqttMhs
TqtopffW1e9V0keXldnmjcGtbhAbx+bykjNtjM22zGPl5sRvC31gnnHvjACXpdeDeDi6JAMAOZ9Y
CZvBRmBp90DV99IO1/ti0srbOU5AI07JZKXtpiYl8jK9o7cq7V08UfK5A0h9O1js0WugCr5h/HAL
NZW46evG9js9yVEjlhV4xleTKqHlVK5Sxdam0C6HELuvKxz/yRf5WEri/29iCWlATl66qRSV3xAr
b3kXI3RXJsgFOn4jeLXM+Z5JN1b7CsiIKUTj65LXPvEiNawJb1DhNzonnDJt7RRBd7qIDnZq9cg+
jY9STKYsazP4WzoIc1L3aOxGraD/m2T1aMB56v7OEN2pkeQMvh3nnIvTJPpx6AhokObjmxNnRcUB
VPwGpvAqUvtVgeRaPmwm47oH7QMEwjEQOmXdgZ6f92LuDOSZ7xAmZtkVF7mPPnSDtQY/1Qs6Mh3X
b1XfLvj5EOwtACF9MvmUdsBMPL/PIRSxQjA6+8yJsSAgkDXsnrHobY7Z69Zrrle71ouN+FmVZ5b0
1CEf3aV10zNuCHPROoQ/nCV8/Ce1kr+YDlp8CzsdQrN6JAvzdrvAIJmw8DoumJlLd3qCWkAzmf85
pHdFK6Cb/qEhxXSwxs2rAQ6bB5vmhDV51mi8bE3dl8/HLoSuXZc+auQmLukHVLI4rWv8UCp7VeR+
V88knpwRAMPWO4OYVy1KPJBN5xyEpSDvoujnb8+UvDRTnc5bVAriqfYSqzqRQwUCDMNDgQYgGK8S
yhnC/80vFfEEXGpMzOxQa5HO9FBkCFB6HcgPBE9jdz2suL2jqJ/01YaK1RKyoANAeC42Zfmb074h
56KHJqkVVDNHUWx9fN7N1gRmq1Oz3X4Gd1TONu9bSJ8b8oDp4donZuteq/3GCKL6uXxgVeTrWZzt
jRkXMUGvYzLVKJnK0Nim3urNEvQSJpy2jLLYkqUcxXw4GUPIRiX5glmOSB9wovJ1Y+PtD8vGYwZ7
iRpQZJs6H81bez9CZcGsV1Vgz/BsNHkA0UOtKQ0TQbowTYrUO01ylsf8Gc0bjUWqr3rV2WnIXY35
pjpg0y4rjRVyo61fOA5q8XHvRxWlbTEEiUhMcqfj29nfGKezN1qJK7d3jwOs+pHerejhJ/uoCo7Q
XmueH1jcAaogYfon/tGDTT8Y5x5fyUVBWpxwk6o5HpXJTFn6mh+Spk7qudHJ7IdEE3tE5S+Z4AKd
qehIzrAFbg4vF/hC4JUYdbT99/HXJAU6iUCHnN0Z6VDQsPTF1OKKLagN5+Cbe9yhbW3iAnSDZCaJ
UCtjaKD7CSIpULXQ7AtkGy5GGOoU1wBhsHSddy02RSAt8NKopgl3niUeM9yXFL4anf2qj9a2tH/f
mNd5giMStOGKbA6iF7Ss7R3yD3S4kwq0Tk+3O9RTDSeHmPIlt1a4s1foGkarek6GIPtKL/g0mXHi
IPvp1qcd7Kk7j2C/5fOUqjWLCinT4gCQPoPUv6UlVENqI+joE36bnIiw/s4WvUAfDUsYIII02J5f
y/kj4SmZmR2PkwD+kMoDxBkYM46luyplG0im8Igf4qorDeBDVHHL0PcgjLL+60oqRJ0QmK0awH5F
CQVw7GA243alpb/1D2KkObY12O9hRBJ50/5RcSvG3ApAFYGynNPzk7zSQdyfOD0qIH4/LsoSEfSQ
GPei2+7jvxa4rm5iSAHkEcLdUoJByyNqNFnhyrhcQqLjnByH0bTiDeYClzz0DXeZvl+cTsEomuOP
jhl7Vx0R3BoqlQVh0pZGvQYHWPXbYsbvzaHaBJXchkINchirTN4H+SC028Ksj9zrCMkmdrst5FK4
ro+ZFmDvoRmYtb7Gkzmz1D1Z/PJ+qy0flO7V5KnrLNCdae4NmdhCchy9XHLEzA+S3xAC635Xo5Qs
ZYAm9UCEIrwVs+fh5IhNhql+o/3ckNgbGVAlmmNPswrJS0n9zQOrRf6GUKNBkcE1NQQHCStGX2AC
iM29i436VJ2tbu6sQ7z/qj5mUjUK2m0H/jWEk9YzdwLLec9dKDF/tixKyK8EH07o9fo+qx0/3o9I
iTMCT0rbKPP/h0mwjXdX3Gh8rPVVY9bhHKbBTzHGpeas5CFD4YMmDR3YPsMm5NqHAwPIEeDpOYxD
SEGXVjIErfDNOnQW5Xxi8WYtKrNozVZ/+ab9KlEyzW05IHe9KNH0JgYaH5nZv6JbEH7Po9CdMMT/
phrl1+SuN4QpCZhHArBg1eklOPF+u9SwIGUQC2WFikUS+tobEbJQ9BG6aJFBPz2EB5jK3YxhfFkb
/0G8fDY1BMz80GsKCiDO2JrNVTU0MbTBsg81HtfnKLd2G5m/gVLBmKlcTb9TySg1b4CDLIyM7Lb9
cPmHLRDYrVCG/n1VNn2m11P0Rujq//NJKwvxC7O6hrueTlkT9UZK0WDn3Ng2DFypFXg03WjsCTFi
l1I0M1LohOJzabzudlTogtIjTsCVqn2HRVFbKmTn0V2cScCWW92gcKQaBoRn3cPGK8N8+UPJPrbU
BhGni5+5mTYvuk0Gx0yzcWYOjEwmzGinbmQq09SmUO0alwg9bI5sLekOJHi31yDV+8vb9zxVbjb/
A02r5409iHX5Zjj/pDw9mJubOxtM81HEJGqIvgnEBO+XsKbZ2tPvYIqSVCLHR0Trt2PSkEWEPVFE
g/3iGkiRRtduqLdOAGn+rugWOHxOCRtvP17zckNHEA65VMo41NwRIdXHTx819d0Jxm4gNGC170XK
GoVCcORB3mnFa8ZOBONMjzmfVqy/+Y127PEKZrSwqrd8Q4vgqZh6TFNd1ZwJCkROvSCCOsbGDIxc
YcSjw5BWCoI+1RbdF85qnkANZHK2Po/ZufgmzI6d1MGJr7j9K7UkVx+xIeI6lsE1VErAo5kUxrk7
lNRW0BSNFjaTH+a20VkkdQnbFrEjdd4eR7pXcEN24rHrVV00aV1vgt+m2cLrOzJVh5o3OPUICUMT
awS0STBhuLBA9/dCq6AZgYagAWNM+M6ue+tmyW+U4u6ZkyI5m5Q5P22413NfCAUmybsypq5eB8Zs
REgV1tj7IDVhoJDquXUz0vht9oUpTJA/cyU4xoYfqMxQrhIrQ6YBkCOaVxRfu4ESIZxJyZGuy+s2
wTdDdZDYvB9P/cNEie5VNtadnZ9DRxYlPcchx5ZLDDK0vXTQwfv5LEPNIVPlqkxm24Pe8+nWYJoQ
IUB79rIu4ObMD8F4eAQmkWLFXyL6sfmQiFDdnC9EnOTmVPzNtxm6eeSX/BY+nYZy9aBchDjF/8h5
lscuBgfIpECEhv9BHqTv/oEnP4TynEd/77SJeljLXGM9NU9CUobs7CzfU8sGgo/4lgpUafENYqNZ
lgKigSd4CWH89X5zWw30OBtl0zckJlOsrwfSrBnslKxFvgnYO+iVPnEGG9Hi6Sh20P+brdOnG9yT
olXjm2qdYAwwMhCtPKfZjkhh3o6rAPQgoJMzVvkdlLuuuVRPGnVtjOEVA98i0Ck+V0140P3ivikF
OJt7g82UP8Cc9Ppz8Lw/ruz2w8z4gzUBqOa8SB+e308IL9zhyGme0JmzvM4YG4sTgzAn63JGv8Cj
ZE0veJyy7He14VlPFEMkKlpRFttHlh43+xFTJ14rGScz4mOvGfGr+B+XBPi7sjZ6obYTbSBt1xy4
2HylHI58OjPUdnmQxOfM444ujNAtuw7dj0O0b8SKlxe1VB3yev4MAZnhx7gBMTQNPYX52ZTF0Z63
p8sFUGctPcufpl0ZoTs3TjltC4cUfKeP30zaBsaFWogy3S6Oy0EjnM7UkCHA+eQOUwHVzc3B+A8X
Fe9RofSRxZ3zTzZElLw4JGpxEDDdbg3Ec67jicilySpnd++tnLPJZTgPt+S9eyf16dkOSjpC9dtG
mhg+a8I8fnTZolmr4Uv/y5CWo9ypdzJd5PN7bmKjDFga2z34i33IWezMur70ljMj6QfnRTj3NdPB
od1tAtVf/y0PPm2SI2Wi2MKLMA20Qg+3sXQhsd/oi7ZJ3J0PXhGK0aU+B24piRmxJZn0l7oKR4Nv
jXGKhN8eojqt249HI+JW8jpCw6c0LEYBu4sffv7nfQrls8fIIdkggM/k7FhTvBPzYgIY7C068Dpj
uYxg7WPKDeCRrI4brOVctMsYxs0p5P9DIE3zwOpiFoxdWtwWirk1IoNA9rOT3Yi8XY6Ka6ekzDdC
pfzGUjPZ4ofVkTWyPkptqnqei2nJbJVV9cDfQ+rj+20czSM6FQjMsCeiyHUOlgjDTQCCAh8HjHof
7VRCG5OSLP76xMdW7Ha0uo+LrBk2OonJZjOoAE8TnHgTUtAFFd+L24FZfv6ltIS3LfBY8Q06QQSK
w8DoXpSI3Tg+y+2AGo/UwOqf4/U1E/wurEZ/AnzNlSkHoAyUMPEA2huwqGBqwWXabV4EvR36lPmw
JHfXiwthtlFRS2Ah6LOmaODxS7878yUc0fd6ZdUSQjDiBJyZDZR/JWBG0OLRcUcJ+utr49t5WU2h
dIjihRC8FsMoXG1t+oYD6Lq3lgssEe6qgqR6eaZukC+O7agqYZuj4faOKd8+g6BJBsplw4h2VFK3
6Ka+eSQ9t8RmNrr6B9XAITk/weZP7uYb41houCTFzbWapbZnO/Wo+tuFDKJUlcBoHto/pM5gyjsX
l1oMrk8w6OzFrf/w3/p+mAoAMziSBGPZS13r96jby5k/4p1SKF9Yaz4ZvrdXOO55JEsBdHOHfdTo
gl4WGW9x6OUm+koLvzjKj7NwW0FxBST3vIArIadnjHioyXWm6y/XIGmsijss1cFqB9Rg1AzEK2uw
9HaOsm4/6zDnawMnWZAiXXCLJxzUgiba1QywxAf03RoK6PzkbV8V+0PrDKl1J+ganU1kUEycgC4z
S7Z3pfzEKu9zgFkUpxs8Szt3chE4A2VG3v7bN+/FpMJkjcLpdPSfXsyNuvnosWy3gkL3/1CQryqt
v60Pyjxm5wLVIe2I0feRmYViz5FSR0zO1WARuk5/sjKU5sRUhyffPfLu5E32/bEkrPonZgZwFR94
SfP7mkKWt8oWjhbvYpcdlNZCjilOzAs+GYQ6BRUgy8DT/9kVPcF9CkYo7IJIVzIm23rA/aD0sR0A
fVmDZ+Y3pCUnqQqmsq5RUZqtTCTU41tr3VwY07EHm1NlFIto1zCNr3joj4WnQcAsR1QLWbsqatne
VOU4qzOYlagvBFzHyfKkl2/W3y1WeBKTA0vUw2JolreEYyE5AJKMtaTlY0IB5hh+sgdQT7T8Ww0v
MPRrhNSIiG5a8deTYLVUGMbMxvlwTyGVtGMWOsTmzWtVjxxqEeyxh/35uh7xBPDbihVZRFrtgoNR
nPPXkdLDgWv5e44plbx+xAQPavKX8x2ZP0Nh8kFSqoChPNLavOEQSSZ/Ku56VyFwKT/8h5AKqtIQ
wtel3iJGTXnk1wUI3GMCYlhFaaCL0eLMMhqLtJU6yWZi39tj3t9rvxhmv/fvF2hsCF4rOszKO4ph
5Gv9lu/IZaTCrDRzHwi3owuF7z8OCv0wWpfIhC67BN5YPmBiyhgjJyF761F62ZwtWiV5vEjQszbL
G51FFgmQPwXam9ZfVjan//lrkyrEv0Z1wkEgOfHIKU6gyfWFQrCafCffuMHykGeunc1ovrDQIa4p
1ir/wgmtJLJyRuXl3wVnDO+dGfk/NxsyIRg5EyTJN8QLHe85iKTIWIQAzBlQj+Fgr6LQs/pVN1FH
Aj1C3JkOu5zchRswDKe/4JEY7TUHhI5eMugvxXs6bJ60D6QqwyNYK9hNDzfqRkGt9sQTnKGZHRFf
X0aRkUNlY4AyE+Tq0LfZQyXsPL40Ao9I1IPj9ikmacpFaKIroW9y8HgqGgRbd3RxAa03EXOySWW4
NhHjQoOe4pjRoajT17fDpqNaMvizpfIjAGU7LrS5jn1op4g8MwvwoiS2GxgUJk/ZJho2HRExd+cE
nHxrmqtJE32tV+oSc84mGx8dMAcMMvzokGoyNZ1WD8V1TCDN6KMzMJX5YWqFeYqA8W2DlVXcFygn
ea8OY0wJw30SGMlf/jz8snx7IrKPitiNt/gg0ptnmsXfJWIXPl3ZSzS7Sx2UFh2+7DSWToRImfF1
8lTwXhmRhnF+kvfhWAvGjZIxfEpxZEy1RdDVs/ia2WR6nig65rfZaAqFaiMZFPFxh1wY2tmHe1Ww
uqEytWBc+ap2GW2DuWE4k8jKeG846AVq82L7t+nuVw1pWADhwKJCgVP5vkRdz5C412zLsOLW78UA
78lBTgV7zWslWbMSCt64UhYkRQyt5Nny+RS1bYCIsZS4uyN2IXVadDjRbYaLZZSnh8cNLctbVBd1
qAoyJf5JrUE6ym7EQYkkCqt8faAVDSEb6Lllcjvl+HeoZ7o4X88oKNarR8h3Jack1fMluNKQH2YA
UzmL5Az2NRCEKtD/7XNT2GEiitmRzxQhOC60hGF/6O0a6MprTKIY1SknyqJo0xN4eCRr5BIqnKA4
4zvsCTpMTlmvDDOIccfQNsmn0/Lfpqf/Gl1MrvvuPxwpo9n+MuqHyRU9AsYHRbKobZ4qwQMecr88
iXKfmx/XlxzR1L0cBPmyaoE1oZLML5fKfBfEugPN64GHKv1x1dHJalbzjEcgfioy3H5gmnpIDRHI
zslHZqxuenmRFa6/24jpcE8WNodgH6zjL0lYfXob546Uic1anAaH7ClXdVBs9kJJvHMso8Ilo+vP
VRKbbliz+JXVeIMsKrcX4rdOpJyA66rFbdRhsOOpMWJtUqtJaRO+XNrC4VYjZDZv1PafIeNe4qyX
udVyvFTQY4XzmXfChdrwGnlWNjhaQ4kALFe8jMSrDKs37rf9s+pN1Cy/QaBMGP5nynS55QR6zEuH
eDuseWOe5eee+qUYGSA31Hx8fNaPzHvtrc6B5ozm2LvuLGXiIVKXeMeJxCxzvtjI44YlYqz0lwxR
u47M40Rp3TxjuECSIXNrOYcsalhZPBNl2bZb1WbTfHuRYB5XlVo2mXL1KA232oLximVHyjpFdn5x
6PFxbtAmGcUPDvYRTqHfxygzL89tep8DT8p0gnYmuoOuNkKOEZod6Yfrcj8rZSCfgmHL/kf7yc26
cXz2i3dwSoOtFbtRhSoZNaWap0p+A+g6ZAVv77USWJgaD5oiHPSr4N8IKf3iSuboG2LtULA5kHYg
NEDe/KSAMQ9IYlc0qwLW/hc8/3wJWUZmEJ5cY6LUCHKnsQ6SdJmWdvpRRTEq3AYUPIokmxGJ1Wwj
+R2lDxKCRvQu5xmVQGbTYuv8KRe8aYSi5a1lSPDk3ilHecLyDmzw2u7cudicQ1tSL4x/xlwjxG8W
mET9lUwkpJ4oqjM444j/fqgg8iYK87EHq0lu+sRRIeIEFIWRoIMpeshVTflCdhzbx19uf0+wRubs
11gRrdDlWdN+d1+S5Oqz52qlE0o0Ssl9mGaj+5kUxqIX+I1A663vKBWVOh+ABYTdFsGY1aOeoYFs
8eCAPnLxScSeBKadW7x0A5E90j1okBG4o8bmaR/OvsoQwr5Iw7oLqRlL5p5JCZIkmiuq4c+E5hPb
sBdqS9RIwGXN0VbD8iMDX1FqrVT/698BNXpEdQNOlGPIqWy8+O9UeMISTS9MBytN0PrBFdSlgEtn
1/s/eon0SHj6MDXXqj4fiLeGSjHbCxVQN8cBrZBBGudtx+Cf8WPaLkvYGtxvmgNC7V+vv2oai3+q
x71/pp3RKSvIAuwQJZlhyPjBHjbouOP9InxcDTgjTrUZEwPGUQ214ea3XNMvGRa4z9Bmase2so6r
ICetq0QUc3g6bqG/DawCwxRrLGWkLzt3ArThOIUpknfCfcM5ed+THvv7uM5gLrjSezHKGQasysty
KiI2xUX7GjxDT1aiFNjHj76Gw9YugWBSSRoER2gJrHpgE7poLwPtGqt7Mr7t6TIv5OUBBYpCkh48
pPM40XD3grERamZs51pU/EBRi4gStWwt4ISqLmArOkmqfpflPY7VXXtthABJ5HK6Ge+dYpsHdJZe
ZBBB1YApitMlzcOxcrG+3/FrMB84E+n1H6lGi2H4hyr7GYltej9aWyl5NI5fNkcR+imOh4QK683i
stKXnh7jcUhqHpAsV8ZzlFqKYZW5zAE4I7V9srMHTV9Td51Y/LxBmUZv+JrRE5LbdgwkVahUwYU/
Ge6UN99emHa63CdkwtgQVB5J9WTr+k64YIAeqO6jHVqiOoViEvjLsFaNw4HsTwIBIQoLoevJciNp
drGy+58qH1QREHMmU9nGeWaW2m8FFH8w9cPRQen+b9rfMBYBJTg5a7tcaDwMtiGp9xyG2NcjgHcH
2bEXejlhHItRBnKCk5n+yYaaI7MdXqLNvBOgGIQaB/MzszAhMuLHRwc2rhYbLmTLIiR6EbomYli/
o7wUS1prhUg+b8BBQa06ylTzO4Po/p/6TASSDPSmUgyXwOugRf960k6gjLHMvpHQI73GADRntTkG
73IiY7bYMsDWfCZdQDAnQZcXPvrC0TEvxdntqSblEDvOkBp2LQQ9Ubgq5TFYqtJUnSSRLSKCz1aJ
MD5GfUZFxifjqJyF6P0+q9Cwg6mzIBsC3BBj29d+K+JIEWMS+KvR0nko+MLS1U/BbNDzsV7g/Ytd
F+4ZDtvvoSpL1JmfJ7mjELRDexgEVk+HbZv1T+TkdYDL1A6J+GXj3lJ6wREi3ja9hZb0T2qGxfRl
BZimodsfndEYb1XWpIod5gZF0L4hAwviZLjLlQ6YBdxxrWlt0pbiaYJe9HnRAHMcLdKJwquEdtQl
e0AkFHQ4cTxoAg+53aw2GSWnhdLXgPfyapSdePaX9JMmIpTFUJT1l+2ZUqW8LxGfPT6pKKYTxQlQ
2SwwAu5N8WKb7SlviUBlZLxBYb3MTUELEfJsmoqjHTVc/kf2HXjc5UlRHe9orcUvPk2M/+paa8L7
xwZeaxolRJmWBUucst5uUIAKThBOo9T0/+o8P1rMo91uIun8iFnLKDoluBROnNZNZhDdq1ZDhEkn
LclDR+uB0OJi6cymkPisFUaBzY/yOYYVFgcRG/NjSH61u5Kjff7gk3paErfSgDOWDbesuFzHVsDq
EJ3dQNWQU239Spz4Wb1cY5f9FRXoXcagAZ7XN4VOfj4ctbHLTTZSah/4MH9xVWgK+3nsz9j3voPV
qseHjJs7oK/xYIxIHcrdCh8AV4EIH/5fWcoQ/yQTY4Zvu5NQzZ1mIV0+Rwic4f0V3hDw5RaOPpX4
N8bahJ0WzJWpqPIilKv8KCNPPifKrzQnQsi2l0HfGyX0nrX4CZuZ+D7FCBr2kM/p3JcFlS5P10w3
4FqCsvGgtKuwCt6GwtfbbBMmlIwZkF7+ThFDyP9iOZwK6lWIOoSQXZRi0Xmbpr6qEErQ8XFMPM5E
P7v7zT3BD2TS2W/5zgadEx3H0jUoMwYoqfhhWMbn2aPQWuqEfVEI76IpIRZOcx99R3loPY9dgX7E
8FUELBYnQg/7mxru1tDiLEozrhkV4yIYNOeWtFYGu5yXarYzdJJFoFNyFds5jQPuPnN182dBnI3e
jBlfiXD99XMwSYrsVKKC/Qle9LUDsL3GQWOFwcZwyYkazkB3hsxu5UWY/yetSudb4RlBaOfeGhsf
5FpVRyKcO1zGBM4aiH5ihiT3sN2HSA5Luqh+AuG3w3/4TGblAjJht79C4CF5KzyRYxjsYnHk7FDp
GDGPtYZ7VMg+JkD36bNWgsznNvE8805uBqP6ZjujIJAys7yEPKYmF5R6kgSO428vlGTHbFhwHREZ
4eEmKBbUl2LKfBdVkhKxLyFBJDgge65yp/6BNy7tOu3MgdeEO4dgdI4Fc7B3IuMGeclUdaqsOvnC
0IOQDcftTzLyCfJR5iDiGitih4pHdsWyP80gybVVPDVH4DuSU6FfA+4TzmQCWUXoGSGWckjVKYAP
GUkuKV6q20Gqx5qHiNP122VfQRJQ560plsD7x4AaSv+Qfk6DuRV0hiQe5bNdv/YxVE477hXiDdzD
30x4He5kv7jPtzX/ncHzV2CnncCqKguAdw3b9UmMAPRIPfxy3lenXps+R1BWeFVVpw/MCVecYyTh
5tXNVuOu4JRFYWT0ZqUHAlaQUqR8diutzqwM0QHAfQEMLz9gSao0fJA/dkIEmPLIoeGnWtcGDCfT
pa+uPWHGiYTmkog12a/v5Tihd5fuZJTEXPmWg9ceWb4fUi4FZcz1hkRHlmlawUeCTbucvsM5nwYv
Soi4V+jsXd/9/wCZSrWeiom/w2E4vVuurEtFqzfXA5ZVZKS8qgdBRZcfqrdBn2p6gYcSBs24GYz9
Ahnp/qHpNPSfnrtp6QTTW8yklj6S33lD8+LHQxG+mDYLbFzrzP2Nq6ZNMu6T6lAF9MZk6bNeU4RH
AO2hNdtY4r5T+WQeFzBUnbYJgXZqUR5ohjbmBR5KH6HqnxjYBmF2lnrMn9xzFR0mRN2EdtYjHg/D
ditKx9CiIigA31y+KZ4ZSzsS4d0JghwnM6NSKindFoejrEKM3GU1ENKQTnxpvn6auQ5KlG9qTVUu
982shVNAlsLndjwVTRVO9cY4mHZa0pTskvuzmfcVwRT0P9uIK3NTOIzBRxjdzn9o6y61+dop1HIq
zjs2q32ekwnxKc9Kos6qPIIURkDf4kstz+syP5qzbdvG5n1yugCTgIOmFKvHIGZRJ4PQXyg3kAdC
VStWh1SdzLJdecS0rWhL3pK9b4+4aPtT3puA7ljAYo5CVinL0tGO1R1Y9WZVd9MkGT+ALp1bio6D
ScyvYsv8nT/NT4yR/kpET6BorL2WL5D5q5UmJLRnWxEhX4nU+4pTFmkouY7w/hxvkGYogSrpCowO
6cb6gNSfttDY5AsPlHltdYdjlIG1PypOG1JRv2piV55mx5YbBIhzXyj/nbJgEdDgmToxeIt7ZdEX
R7jRJ3OdyHRY6BmtPPKq4ke6E6Cf5PmM7GY2WvKgl5hjhSnGmD30Fw/OPxPIdaN1m5RCJAVkhB2L
SxFG6J4odd0coDn29mRCQr1Pa8tHcDscn2SjMDW0jvL16rmqX3wOzlZSCa/zGdcJThlJaGjEMtLy
UINm+LMRWYdznQgrTy1UhOn7/mm5pZFlWvR7Y90EWHxPYQkVZmq2LayJsDPBBRSRBjeX1H9sq1qn
G4QIY2FCp9Sqfzuvcng5zF67T3GoRzsjcNBqUtii7wcxdihkQMMjRvaWhke8Z7z8HP0tNy3LQeE0
33hSPSFPFDgNvp+v2zfIg7RocZlKM1jzVSCagfXObtRlb1EglJfoApWDx7CCbRLzYm0LtUqRGBb9
wpM+G3Q2Kgbs2/KnhgzxQ3+8bCVMjeh6YqyIIlYO+gmarXPaIseNZxPxyFM9G1Gm4Fgk2IPMYlyx
BlQsezP3R6RcfEoWS5ga7IECqnd8FqvAKk/Ngmdgl/hLwkQp52fD4o6wt+yRhIl2711xiuCgMVvr
GBQkVvX4lqO7hoHfsT8B6QfTHLPStMMO+EKH82WQHQ+Vp6WfiodSYP9mnHvlefb6ADKRCvyvfRS7
3D30qLvqfLKg6J3PCAzF2CgNZ8yOOO08a+z6eRpn0q2uwXkV+zVD1jGmjT3hFZgB+Ff+Gs6cbJNl
kd0SpxSA9WMvp/jUUenTfj9+WAj4qTr29LE7UJ6EEvcVOCNSQ/f9LzCXGxsCdMVOMYG9YDCCSt6K
QMsMnzx1dkaDGPVA1k8BCPeq/umcHkPRbWLEshu5ma1PEy9o4bXCcywHgNP6C6B5OryWsAoFxrGl
t+lTEkyghcEu23FoyYFlbHV0XItyZll9xfvGq7J8GpEti8D2DhLqOUn7ymkyZSneTsegaW0Rg4aG
GYBslwHyNBBcflHnZIxh23TOplOnYf77A+M4d5PnzCRNuwdEUnn7qs89pVNnSdSldGr3XM3zmjpL
Ve9HqevAvtKJ4NZBNqwX+g95SNeDG28bKCXafRZAiDDr+NQKwi/Q2AxIeUZR9vNdKkBWZefKOdx2
7O3CzQyeQdrPB3J5M/CSsfRdoKelMPOUQ1LgBg4GWyIoHS8iudvDVryLNnEY1D+yg/YEVOSw7YBy
+wJuN2Z3KbMNQiIUy1aTsDnez8Dv+C17IlLboAfdj19gzOAay1+8yzqVaDNroOzK32xwFxv6cxIF
udP6dtbpRiza+15kvyHXe2R6kjEYXwhY+JZCzrWqeoTsgQgwiMQQoCnSvz1zbtRvXE2XGg+ZHWO3
wFmqg2E5sGADfMCBfc5D4M7QapSndo95Zzif3SP0LqI3ACEHpLPgQG3pO7MiG6XWA+Bybm874BCW
3hCRfP9ntKoHu0eqva+HkN1WeS91ICX6JHDovydvWzPADGkjfulC1cqb3TouONmHdm6DYWS9KWft
cfiZVSeCWQNVZPLHlPA3rV12kZbIPMAQk06EdTFSWm0jCt7Yscxt8JmCtUbHNJCYU/NcNOtBHtC0
bg1nc/pO2BxjYxiDRiBPrdc1uvVs0HsF5G9rJaFnuYkBSqMKpjTKWhIU8b9s88J0aoFwHB7kBB1x
qEnuRXGdnRC+CXtka3DLbJ4P9k/44feBNxL6DR4EoqgNVWgawzle02ZYxsr3ES+a4eNJm0SxE3TZ
Zy9FmBUEAWLmRmHZ/ckrSDml3EnQ8MkCqu+PZzns2Qk8SjVOFNQpxDNuddQphqamAdHIGr4lC4eq
rl7VgPYpOlNkCneA44WR8oOHcbl25FPzSPnTJ36AjVTdM5mCL9iKilCD1eJRXsHVr/jl+ndAZjNL
qnDTTeR4iOCCemF9HZjZqzMglXRAVNFJgLeECgPYio6y6V3FesIa6iMLEt/Gwo+xf5KKE0uIlYtW
ysM8voukmzDXIRCml7Nx5B5QGxb9r9r2yRUis6jp78T/nOYTJVKnhNQxBEnyYh3ReB/D4E/4UboD
eliQSBB3zO/9z4X84WJVhF2KSZO6Zz0ocxRGYuVLXT84JbAlWn3LmblUwBxN7Xv5gXfYyizS09Rf
ijryXJjISHoAVD5ndeAYdmEBp+8Iz8YJjkiCPFZTSaYLsUt6qQlEMFKK2y7wKeLgD1C95YfLmXmW
ENuSqF5eQGg/eDxm+D/zOTdQzyuP+q2DvaOXs9dwB2s2PgQVJokPWBNvkmtzOmR2tAP51aOF0Zf5
HCTrwa4PZWtmFpg5FOx9TA7y8fKxqzcrbKBb85+RBx6VDCQhOExEeadIunjaKTW5hsH3o1BGH8rV
qiPXT32IBScP4n41H2DavrDO9O972yecvGR/nja6nYEtMJdXH6Q2uVRyWtGqGH6HX/uRcgQGLMRN
nabqVIPOE3ft6kqCH9tN0hjN1rQdquHCaVvCj4LQ5klJq8fVIdeKGJWykaBdEzA/hgwbHsifaQOS
Jt0ZSBOxyJ+q7rQlKMsPdDDHyEjeJlGVJfwGCEU4oDjtbJVM9Kne8qc9VTtYIPlX/Aa06d9oj7L5
uiSjgKzRhgpxg/Gszy6UVHTP0IhKz2XSzPKFMsJc0lKbVC26f7sfUps9D6LseBrQbinqelu13Bc9
JakPHup0rLElHF0RHsPn1L8fGqqy+fJotUSqboqIWtkWnhf0/8L4pMQ2er+HHy0abwZRr+zvkrCR
IYgVj3G/gtW4l4HFcr1Q6mymIz0UfcGcwLvztE06VBQk2Pk9IIIyQON3xwg5nb7BTDE6WvOJ4xG3
cfgj/+sgo8Aovder5gaMGmf2PKbWOW7A50LeF5fcDkHaKw5M9qwkTDoVaDWvU6YO+0e7BVI1FogY
L3w7rCx8o+2gqtGrkS9cNHv5rZ8NHt+tktCXKBG99teCy3hi9UGhxoBPVgwNJpzFug4NPPPUmMJ8
THc8Npoi+3xF33KivTS5CocjrrQBm00u2bNg11FA9HGMLAUzIldB+mjoM0rCV2f97Qq5pXl1tro8
ekLu8Wy/6PpVMEgn7CnjGN9+p9E3FFOffpJ6/fRmo4k0Ol6qbhXzvGXTgo63BomkzCum9PI3OyYk
N+4RdMfGHh9ioD0BvRNjWOjGf5psWHFf4qCHmDpxrQwFjxeNyN436qsnN6hX5HjhN6Q2Fog+KniN
XTv43yyaMPqF4Q9ZuGsepOtDL/4JYZK0QVkCJPJ2cZOjSSAe35hElWaoZ00SavDD8UcwA/jQ679A
LrCvpxAVIQjjXv/jomGLn5VpwvVIgegtmVT73sSVnjyjAthCieooGG6PyGva+AP1rMueu+P1QVmF
bTw8mDBWRSz8rV/BHmc04WLpd73lCPPbtQ7P1YStJP0AJgRwZOLN2POH8EFLEBo3jVmIksqXShd5
HN8cKkY+HaaqX2UkhC10KAwwmNY2AvHCcmNnHrTZQViLcuZXNyvf2xPZCDXk4aamqumFto0p9cSf
rDu4MaXivBJf8PIuuNPcy1i9ODrDsJXAZjL8uqR+ouWoE/PKOVVmgugQ9LSYjQc7TxqlhEdqU21F
i5cqSdMjiET30Pf1LGWeur3LnTOhhCR520JnBUqU3ds8Ce+qT0UbVcXEI9iM/vlq2y/xgc9CMoNz
tspPYlJ34YwBA8vXdokUTh97zCDrz+oRSZrG+PNqCIByPHKijhEcxYlHrsU3fZdPXH/uk8Gq3XQp
nz/mTq7FfFsSpjxESsg/L8C4fViQtpR2csJweuOrtvqQWJewz/gNOYhpyGHE0Qm+Ga0JNZMvCR6t
L0yHHArsmwJUoUBD40qv3FGH49FgZ6FRXBbMS1y0VmrB3of1NQywAoE1L0+RPp2V0BcmxBZVzoOw
rTMnUTq9KyyJ2LcMoENmrRMgX9FK5WumPnnqasQ3n7cNJdhsoB6aKRUATPgGWVuiOvztlnZlqvWW
Rsq0fJFVogPD/sQDVtTaBQjIhaukLKu+/5vrpwSSrS3MruILwCleRifLzCk/g9NRSLQO98ZlKJZq
kgcAYn7msE/A95IX5wFw2D9BtiiR/Rkk4zwthe4mLkU0xzq404r0JT4DQHEdW4LAigBkw2D/ITVv
A5crgg+cz/WQ9C8CWMzauugyY0uVnFVZxQRg40j8zAVGZcCsEhWtnilZOehXHkuhQZkEQf0D8V1Y
i+/8wHajHxUjJVzC3E0elwLaJflVerwTj2Hyz2eUYkBVmq9zSNthKHhgR2n+izXZ6cS3VgZ6fMoR
qAlpjlC0h7Bv2bvt/YO6nuEoUnUuoVtSna1iowjCnWuoTPOAXp6oWxLswcw8TH777LB5V0VdaNFW
WCLo/54ocGccOBixmS3//D1vxOesM23YJpxpA38th7BLFlwuDxNBWHP9QtfFFg+l6nrmurNxF/y3
qDCbWoBUGBHRC1V9cP2PscZo6PjDrfnrpG8E9W5eLXpekUX6XMiyWuOAhozKpb01xNWAs2lsqDbK
1Rf/t+rdUz6V7bYl+8Mi1Dbi8JljqquRwK/Y7r3TYf/9FO5H1LR1AactJecmpvRo7s/+eEqBYg1V
qQ+jVIkMd6sG1PgXiDzp/qIGyu3uun4vY78Zd0kY3jkw5q9Hd6BnhYs6uZsTCjU1oy819wpxmrdW
P8BS1I6qV/CWfGY5XA39AZDCJltsuyq2mXdRmwZUiYghyktpjhy9E0IXWjiaPLQhwZ+a0+RPgiM5
SjyR0+c1FJb5ac2TUlvBMEJ4aZFFd10/SGD5tm75HLLt+7qUgD3Zlusyz9Ab96iVbiWDvXK0XJRN
W/7lZzkW+MGb3TuggfufJCPfnBJk4NYTzbl8x6ErRFDroSIAGdbWR7D1U9GEAi/pwdc6TyU1mj/F
UU/TLC2SzyuT8FX9Mz8xENCr5VuFJNGQw+Gt2PRT/XjNT/sgEQH0ZRzo4bA4tgIPSo1aOtPpRdfr
F4HRDDD9z/R9zqYELTGlRwptB3iCKL+FgFw51mpEZJKxaxRzy0ZeH2kp5Ya8tGg/uSAxdid0lckz
9PEPKN9Ii/cQ+T+rXQAVAVlVJ4RRvvr1IBLJS1NP3yoxNvKbnW9dsIlg52Q0tqK2mBA8Ww1KBch5
h3Hmp48ztFVCwUQlZbYS+dhTmHM0sxKDeMzcMRTzo87VNvJ5DpzL3tQHET1duI2OfWnbL3rBJwmI
0QifIGw5HOQyZn7j+cjPqqpM1YqPEVOOSoamPRo9KOBMgeAQjVq8FogOgibTFJ8peev0dk7piRVL
PNVlK4ZjtP9B4cgSLVamUluKb3sY3RXA11oZNuDDIN42Mq7Cd6VOjMXkNV+240U1vouE0Y4ttUNx
/16y7R/+wwV2X/Lm8ux7gHx1sRpId0zEescgA22Oxs4ppeg52w8OKv/UHUOMKTOjzqdgKZ5TU9Ea
68u/EOM2mQUl/NWebIwWz1PGCLpq4dwzs23tQIEFE4NpeIoWgIdF/xaAB2gFlzTZzPIUlWEKGtGw
hZ+tr3R8GUSJAFozutjzKFbC3AsIyFSCznJdQDa4QJ3KCUouuguunCNvHSfBaPYGITw9cOHfrjn0
PqU6N2kWfwpuiYz5aBU801q0EYtXr3zc4ffeXaSNp49RKlM6aaVXNrC1I5hNyBgOiZi2a4pSu9UE
QkPku/3yIT4AKFU7FnZ0vnKKNXr6Jrx01Lg6wSIUYZM8qVDbhNibqL8inKSEnGOR67uqzOjwDI9G
FwKcKsQOGQbX9Y+iwEwE8NfCO0eoevMSFU5+TZzxbHOHJYWbJc31LVdu+tUyjjDR7lqoTS9CnwkK
93+qxxSwigQnpR+qtm2xwgnxFoOGvJaZ3DkI4eRlWEjqSooWCmayssw2PBcUvMSFhxH4rZBKYN53
qT3YcsCvfnqFSzHBj2nO5DktGhwANMsa13v8J3X4GigM8QzVskvW5ZcFPOAeHVQDRqO9opFDMTZK
svw8OHf0j6aXBEsduUWdsigKTO+8p2+pns0wfuGuL2bDVQfZ2AB8JQutJJOeuempBVDa56Vyo5xR
QQN2xLrkLFF3tmOYaZfndNT8Z85rSbW3lsfs3+CFnjzVgtUZC7Anuh125XnQ3JQxUn8iOdsD6y6m
L874s7P5/EeX0An6X+ZyPG0AW1UPq0fSOP+71I86KTLnJmGqeXgaVZglsTgju2gHsV8XfX09Mzim
7HsAobyAyH7031kyWpnln9xdbFOtrjtCDt/M1tLyHn82/kiafuBw86k9ZrdlQbaQ/BX2dtT4b5NH
3/7T1NdJHjUUaU5R4nGlgz2iMtXyOJ+4HplGqPSGWnfT+8fdYxT7du3GhuBaHLB8z+JzNmFmHqcw
YqYA0gw6G/oVJX/4Hm02Bbtg79hSKpdkqrtdlnGrab0cCO2WQVDDWHoKPX4jevrbiCYEezdBdXnc
TOY3nCqSTKKHZCSdBsgOvmTIWBkK+Rf9OAn82bTQTPYNTjeDt62ZlVWO6em0MKVC5/gbAmqTFiKX
jDNPf3XEpoiWBWRePt49YlrEqI23cKgJwJWVBRmKkAHWLDCJAwkzuSD4S7fKtlCN6VYXoR2ZFAo+
cDGPoqDbGF8W1uXdFivxnQi3A9fpnBEbeJYj6DAqFs/2U5HfqVZLlSEt9JSm6JECSeKMkc4zfMXY
hSOvXh9c8f1i5njaVlNcqUulsRL/VWlMao2dX+WyNh1s0pAkO+IT2JVRgQ4MfvM4um8aGyAPqpBj
/MKTjBDH4Ljf2YlVusmsDqZ1x2pdrVho20yA87UXCYDX9N9g8OcaM3mIb210e70yb/IwbgXENEY+
QtWc6cw5J8bdyRNuZE5PZCEozzlUkvx4Mvisbh8zzuVCNsFZr7vKxJCMUVwpe3ioR9eANmvGbzCu
cuzsXOXOU+UV8z8UUv17q7LZvnlnFMyZc3n7+HJa3qrXQUd0G2leyNwYuqI9HrkP8Zw0xHWpBcjA
wXlRcxm3BoTZ8Qv+WAmIwTy+lXCWp5j77gT/Sh9slDnttbXVqbu9Fmi2cuPWGMKeQTTTR5ZqOjqY
GBT/oyZmq3old4kunyrTvZYZP2FfCNiTtyfg9uKlVjVPkkSr8XituWJaMLoABJ4ssuENyzQDlPL+
9QqQtBEVPgpi5CHHMQV25wnbmvLm46JYumwX9JW0N15N2UFD5ta1+8uXT6aarwDFsDXkIa7wGGfF
hzycwCR/ulq8IHPGIVoTrSse8FKU6rKPScOo4JSULiAnSz6vZXFP/TuGENCHpLfYAGpBb0BT7tlb
ek1VRADtee2s1fCjMlhorK8ju91S8UiTMtNrgZ+22u/XjCNCeI6xX342uvVohcKhe3SKwq3vHFQ8
RHhwQTXcOtPn/w/ZLfLE50cmWFhGFWIymuxJSlX06fl5yArljmejLSca+c9i7e8yA+LE0YuxYodM
tK7tZW+DUFsg3s+Ffyphok7I/VitMSrHQZBD71pw09V0pU7D2rkOdYeRuskALhOian5KHpkl8MwT
MSKzYa6nzxdq38UdrocvCJYQUgQb0rv7ioC21dKFF0KICSHxvvn/47N3sgW3BpIWxwRimbAegq1s
CKzWpyvgT84G15UQZ5icnVOOEYQVa1Uq8NYqVn/pu1O3/afUGhw+cqafhLoqNTgAStO6LSV1brrg
/IAEgpqWKcDdBvMKG+AyBaNdM/Mzy4MTDYqAZ6XscwiIKwNmpJlOU9aIdHemulGDVKam4Jp40cxW
a92sa1OdHccZ0wut0N0CQmHXx4ndZ0e8uhecjVgpEW8R65jMdpsyppEcPypbHL4YmRHxsFhBjwC0
9Gsq+VQFtg/Vq3gflfqJLQZou/87A8H5Xp6I92x+VayqaWjZgJWxuv+i6Poz6We8wOO36ZBBmxXy
+HrRCiumFuy6Fhwum43Qw5vTaR/2YSVGYdq+T3jGnW3Uh1fRAsKUlWrtHtOoD057nq+OldVngQlv
aRzawEuuGEx5br82/L6BcvaIkN3JCSPcDEty1hUZH4L7bykRml2j5KY5sNOUFzQgQA1KTI+kq8L8
mUg8/rcCBhFfMT2nDwi1FMXP8kMMQTl0a5i1s21kwtW1vG0AfUED87KaQZ+OMA9ty0xfdgG3jSbY
cLQb/puqRRYzxfEUa5mDIvQTl7qNRPS+hyTqrFpB0/Smxqoga5pF6vym0s4QUCr3G2l97JORZmVW
jVFuIpNh2vP/yFki0Evk48HzRAOfQhW79rrPvZHFYKMgZpHX41sBEs3YHRkHG4hObXvpNJ/K6ytJ
qvCMuBzm22nJuNLcDiO5RtWsj0lxoBc/2O9nhCu8fNUVHXPARwgvjJAu6ibBmAS5qd/bTSVG6j8Y
lX7hU8La/Htm1+5GFT+5g0tYAh1fcjb9rpQ9Pq9LJYfb92056gUMtx43RC3P9sqMI8rET8knkIbr
FazZURVhmVQC9JAt96Y1cR9+rSitt7tPgTsvAin5TWHY1oF8TD+sZCe0FU42IhDoqh7i7DrZmLB5
Ww0vtIXxpi+jy372HX7voKGXaaLguFWDtpzed6HTOew1KYQ8GkeN4CNRMMIe1YPEWHl0uYmEVq2t
CxOf2e5FjfAJ+mZyEVGQQdk9096TMpkETB/JD3NlJTMup4UQ47fKPvWPdgNshkhGIkpKPWAuzt/H
fOytn/H1BcFNnDORduXgO4R+JJH9SRuh0UbeFM/OyjdJF1f/d7tkixl86FJAHdKc7scBoPmOvPNr
T5EKFpa2A7RXLkXi5pwGPIwP71nkRNmlWbr08uvgO8a8xmHfLrcaSGHXv5YWSvTIXQT2S8wDDJGu
ydpy8Ul7GZ15JsZXj5xR7WNWXvPqfEFFAB3pzpHk/dFi5SlNatsdg4KWZdHLDobe45WaNz9uQuam
PzTEk/ZitP1M/s+Z8UStgM4FriPHSSwk51uNRTF4gGT23ygYXktmqviLAcfn/6IpLU0iB1JHuNyk
iiRF9kZZ/5vhsnjrQCB2vxOBruLBuniux+TgS+eJR1hhni/peuzpUV2yNPeEtbcuJBCZzmFFJfTr
q82tZBRfOFwhgbZQiOky9NFJi3BUjJ3pH0mChelzCif17yBw5XQirfcyDYZ4m9l9tfi5Gudk7bws
SU/d/tQuzQf/ADsgTUZZZg5UKbpG7zqjqhwXQwWghT5j1pu6Rf7JKEdXN0t+AsGrQNSYeKEUQqEX
2IH7jHuWgEBYB3TkTvfJDBO9pvNNm486dlrqFgp04elkktKLTO1/QQvKj5mOBzC7c1XBzmdSVWE+
WUZlHboJDogzi0WxKyVjOROnGNh3ccN1plLJgJbkjYioCf0L3qXnywG7D0KkDHAsGw4C53rEBeoo
IxmwEwIm4kQvBYNZ9FR7TvCt8JkM9VrjcDfJIeQJ8AdBw9jdsA9by1FU9TtwOnjqiyPkb7drkkyp
KhuhlSThVitLuQ04iqU8xLRzp/oSY1SNNs4Oi7HgrV2YaMC16ZFDlsX0BSpRGeCgklBBt3yzfwJO
PUgaaPBdyUAWgRkRuzY8DY531DfY+a2OEmL037W9S3Rj3LpI6DG4Deo9lcqvTpN6oQ3hihi0fcnb
YjmfhGHkWdo95ZxlleiBZHeaFtU3KKFGvkXkiobUgfSDIUA+2/Hevtbw+WTccqkqI3tPe+31Vkdf
+Fmu5b6//vk+RSViFWoKJ22+3Ii1a68yOVYc9RLV0j/JQORKCrvMJ6IpLP03HTTuvq0B1FXAQ1HE
ymTStv02uoFP170nsaqID+foKZZ3THYdjHs1pXBqQFvaMaG7tcuz/9H2z1TorXcrtPpXoOn415h6
ppQ5/Lhye+aP3PW5pk1bUMdSC8eS8yKooX6nGcjsimofi0SUWVoZkVIe/d8iQ8o7kR5WY5Yx2zKg
jqkSGKTV1KuStCuCJerRrBS5q54bcRO1ee5zk/U7i9+CeeH2os+FO4eVK1wYNKCcx38sed6Gin12
bns7DufFrdW5wMdLiwOdpcOo8eBNBMbChf6X0CcyS1DnwJSeaSU7Gr2cwETTpMvlZ12cD7FgZ1ay
IKWZ8G3ysjeDE0ctKNQYw8ipKSI6fTzVNsbk0VE5ntZWmUiu4xOdwB76I3Q/kR0YeDRotLepWtxz
ld2JnRh5hmaa9qhVmaBQzuqB4MZCOjTZlP6kPdwYgI96xccwDtaHezYHDD8Jl0VsJTbAqJuTnH/p
Ir3UcQW7XQ0XTB/oWnTT+3j+xs5cqwp9xbDATfobuLd9Wq8uaUwEbLXK8WkYwFWyEbq8D9US+nf8
Lb+uzijoitT+0pSCPXLDCiZHQfTe/UiyrKVRZJBuL14UHp/DWDViheeeEDPbOLj52K2nA38WE2L6
GrjXznhTqK8yJuGFDL/NBA7xSg1VT5/ePTmI5brfi7ynHgThe8KbKLT+cHNS49XJqbyxgnHpl8UB
PWp0wSs2t3RmK0dYYWAKUlV0DjLKR8eYCDD5BM1720xfjkPbEjrI8aQrBwrTDTAiKUV4tkaWf7GC
sJRKhkMtWCEsJKpf701oO3CYw6BQPTfb2VdtQuGTkp7/Wffn+hMRGQuIR/TfdMveUi2JXgW2g79l
gWXkU72BOmCv4T9U7nBRJB47Ys8Tf/JEgLPreJZC6pkS/Ufvw4pxbNGcgC3u02dylDKcb7M+9YeO
lK13jyRHnRYCTQJEJGEoru6OF4DqIjo37TVsA4/KD7ugsHc73VYeHk8vfAby8KYHYq9OlR8p92BK
RGcPwk40FuB2pHKdUvGDu7cQNwGs327WDEdWu7i/eTjDHBrkny6x/VuKwemSaNUHp2G6U0t6qpaq
qloxDrC6+99tdRqXRkVb15jCGSNiI0U88CMRbEUOWATlmVvwtCLfAhKTpShvSrXkKlg+wfNRo8xW
zwK5Svak92u4DqkaKrPTjCXgyXY2J8nvwyvGFqSyXJGLP65te0CYGPFqiqgSEzIkpDHmhT79Pxa7
IVCJo//q3Ww62ra6SOWnbhb+PYjNUmChIYL0t5fZtDxAoSkaBxpbzuj0owSa5R1Vy4QHecK+92Ma
tbezDoSCr5tuEQGElUEkATbg8kqLtM1LBwc3ySf4NWGU490zT1NrlwwpkNcS2AV096d5Tyups1Oo
dwv3m4QLiFuauRJP/JxfR0FpBS6lcOLUdsABLKDydgqemncfJjYeoS/a546wz5791hepkAu8whGW
js7Rv0d8RCwJomA4KC7lEBzQYxGRLS9sXgovHL9NdSvtAfnuzI4PeidwGLfqAdz+m8zusrI2Hw7w
qHZWQNLIqsEdtJ7Tp0L3JldPElU56l7Yb3VYNUSg0+ClYd8AmIsLwdhQRJgUHCt4KPoywSBXjWvK
l0BXES8P18/4R2J5OwLkDfd65uul7SfuDUtdfv4p65EZHvU5kSjeJrnaMtRMwYwQd9b7SjqemN4D
Eoa7mR2UOR9TINRs1IQloFw/+jzmfKiSOH1wi93s3BL7+DW1lDJ73nqzhZ9G1+MMzBPgGnLsUzA2
0BcooNFPhjiFgUCR2h+m0xPS+JTUr4LUGmrP9dBkd4vrOvmHeulcqY1hHlNvcGXPaqEEra+JnQKW
Yl47liFajibkCYbJ58PA1PyatlCcVZDH6XMyprisr6XVPppMNcMRBJwfQaa3kqcvCrBF2Lje158i
SDgIl2YNdbfjtlWY51K9h3pVVqRUdPpQVoCDVpzXq7wseOOkaKfYoOgAqJeYIooHlmYqIS0tyB3u
0lssz7ID6iV7UztAWS7D6HMlo2+VBYE/TGleh67lEGJcXfx7hJrgKa8MyHZPCsqcYnChxNBY5S/L
3lw9wK5odUEXXEy8i792rbZznMa3hlJ1RY/moLiLnXd42F9tIrqV7kTExLulz6wdKbfBzxr5GUip
ttgnJ6nycSdF8i0NjXoem3piweCa2vPHTPvW4qhl2Lqj1a1qtqGupjW62yjOzZdBcdC9UmmOOHIx
jngiKzp/ESIuK/bYWxU66CxPklpRwMGDBvP8U04CSzSd/7Ump2N3o4YWqzXXFlJoATwSkEFTW7MM
f2lHxvuMi4e5pzKW1QtdZmU1Cst2u3CEYQ/nhm44R23CNNVTCdytpyHbZNCVk132sKaSouEQxWTw
Bq8vuuCyEKDy+9Q4woLXbBbzMcVMhJ+qltAZqquHo71mIl0W0t+Fu3dEFofoP9kDvpa+V1BpBnMb
Arn5FOfASKUuYhJQeFo+iSqpwYNnO1OpzAg57BVPOPubWqVWdHbmUbiR7EHyBvfxyoDssT/fonr8
GnyPKQbmCNGG+QFQZCm4pW7eDahviAyxHxW2cbLUOIWX0oR/tmnlyGuheOmSv3VIrpmaD9JDNRQl
BUmyBRkziH3obnvZ0MBAsmfn77JErykZd6TGX0ylDXT6G1QpIl/ytIXEoDK6K4fFA94XFIhPJGAy
BUtu0Fw6aCh4NCOSzqwCsFMIOacZtWjMMTTcQxjWzgq9pg8h6ENggMQ13zlMSjVVaiCNeD8WOQrn
NXcaG0LnLU61QreXWuRSq37XL9EjkSeubKipX9adOn9JLLQudxvA6MF5l7EjrrcFxnw/Vu3B8WEB
Tiny5qq19SMWEHMy/7z9DBb8zXkVKMt/l5O6wcSYAxT1bOp2menLJSB4AuDa7D50gr2/b/dOi+mY
23sCZmiR/UgRLwnN1E3d6R3WRFI7/Z6hWHEuWO+e0e90hl9+E14xqikSfu7TyJNWKP6t+5Q1H/oz
O2MSLhqQgfDA2hutukHsTpuy7jXdMQ8QR/mfzBvXNKgpvZLYq6ooMBJlzOOlxGlD5pjzZdLYjKQq
lPbFv1Yb+EQmuHsXclk+OfY/tufPQ1hK+2MQTQC6aqoaLWSoa7FzNBSuDEvPUYBeMb5Q7e8hw5e/
XrN4Ukz7GMNrAGO91+KrKe2rg++6k4P2zLYf8YlBS1rswYpN0D20YlaP9sPfEl0CHERdGf+ir3qu
CEXvATSZ+uAo1JtbT3C4nQDgwuwOCIGcc5LAZPLOHfLhDH2jbwJ7A3dv9awsdRTtGQOnZL8K6lcs
/0CxdfiotI4eF4Dar9/rStUevSqdGfme2gT+mw1G9MpDAUWDfxSF0awGbJgS1wUHXwSghrV/AC9J
KJB/rTNFObGY156XuyUfbtAFkR69ttlemrBKh0KZIMjyyNo+belbCccLvDL3V6xRzf+MAL04r85i
utMk8wYN4NX35pp1lO3mhJOWTveMMBrLu5Lsjod5PVtz9pqbXdxQ0s3/7FeAnD9RLgZVV9rKDX4L
Bmluh4FOG04S1ELn01QdGbvOPXuPGEq0SnFkga9ihz/O4pwcP+LaIxWx6umeRaZrVDNkCpgYeTpI
3fQnwKHvvaOpc6nQxUoO3n0y5MBUf9xVZ3koeB+bUOj3HbjzM/iEY/3TCQrnl6iro5b0eW/u0/OY
UQMvu3WGYTghIwFKqPU3a17+tSf5fr8c986Xodww/7cwzasVRljcvvtxvMSDv2yMI96gvZ5uOv+6
Fdv6a4E4xbmoXxaApqt4vKAyhNrP7j5i0PWmTNOGhaIxWMuG8RMhtYad+0LkJah1V5wcLrIkV9nM
jv2++FDlApGDfR7H4ibYRG8xFGEy/0XfEoXQG9bCaPawro4+bUTob/NlJfXFsSsmUkGu6Wgd5lbg
j6Jfxeu5K9Rbq3nrVm7PC+QB7ZdLPQtL/53zvfHzi9skkcsckIIcV52JM2sZ7t08fPKdGxm889Sx
Ct1PubH2dD5bisvCZtYhsUpUVSit9O3g9mmQrq5u5QBlW1MXYKr5aGBfXQt/mjciv0gfnAvzv354
tIsR57QHyrAIKpPWPaSm+tELlOkIzctVjE4A0Ds2auArRpyvhu5rCtY4Tq1w+L5hDFPx1ti+/CEA
jjOV99oVHOgJB8HjGmnSYETsjiyb4sG+qA0zbzKwVXwWSKJ8/xFB9ckML2dHClfyD/Ko/E/wkHE2
KrWRGfYZ9FINRaJyNevm7Ys+ZzFrpVTLj4SbG+HB2kBaVLkwwkqaLUX+EG62AZKnG4fmwbwtf0iZ
3PvfaVffMzlc47QSGXklqWykSLtN7XcrZojA7tIeQF7NUCNZP1jPnWNMnde8FaVdlieWni/oCMMc
EjQ55MOygyVsupcVGuxoV6DNT88Kz1hrWEQFoTaf3LDesdvDDHuJ4yxV2gFTo1oiRbVcTM4R2EKr
Eo0k1QR87WudNmrz+Sb7PWi6xSnd1H93r7UswtxBQXTXrpdNKROyseSSix/ggbL+0fKzsdV5fRKS
SQDxLKbp9Krvgex8ESg9H4NczHEMXsC5dxXPNENZ7uLyiHbu6Amh9SxQ9N9AJjp+8YlhHWe43uib
DidJZPbyZp2jr5Ih+Tshut3aV5GBcYl4q5UI0qiWXdqsXtdP3hAoYhz87Ahzyl3qPzoo/3s8hmrr
x18JAEMtlEfmAs5hssdzrK9OiwqyYeBHFzVq0d3rkZFz4WENLCpOSMNrtrmffPvS4k/RB3nuKf1N
9607DDGu5YQWUaaMuf/i40oFT6FiOCDooOQiJ2hzB31nwush06KVKElbQNnIjE7rq/crKI0dveON
7wO1346NP+lb1/bgxO3Ez2UpGP5kGe9Q6p3KYvyMVgSKw5uCsOo997YfUomwwhNolJ5X1MlwBrTo
pFZdorkItPVt9HFHKGseoKAQSK+XROhdvgtN4CMYUspvCZGq3ctP52Oh+5WxAH/k325kOcpcbnzm
PcN8QgN+scKU1cPFRi6yxIj2YiZkdRQ6IVXP4KM3BaL5wQ3kA5PWQTKRNjC6HwLbXBEmT6xwLDNU
GwbFCyrwOdy/Lqx8ldkiWtDpkVDI2+cWXBqEKQswYd/OApRSo7WzgnJdAl/Deb9Xob+X4c0trl5J
8vGCuBclj4kkHZKwyEggvVBvklpJNM6PMkHdbO2cIxeLREmFRDZp5Xpm9cEbERjZ/W4PaRnD9+da
O/JcuR+U9kYhOK9aogG3V9d/DPi355neA6M2lHzILhfutxFaxdU+S8ml5DTdn2D3UD+YAuMraXeo
eArhWf4/zYdFLPf0pjrGM6jpfqI9/84NuHKRVBVH9gIC6GLnhRCkJSZ5i8xcaydjwLqdO/uXBCap
4hKjKTkGXUhVZA3UbrIK1YIC97Tp1XbwOT5dtj4J+fA8ul6qOyS0R2H1+JKtXeLRLRNeF7MPjTqn
21F5jeq5L0G0x873DOQTGl20+946xfrONU2OdXWC03kBq+kbWuQ5tHHMTnROIkkjUVw6J/Gjdgxa
QRpvydri5d8rP2ySacrvfh2DHtOhUfAlgx7W0WxZdlLDyodnKfGIWyOGLuiZydLII+028HQQ3gye
7f4rpsleeEbUJsAjMXNWX3zHPG2xaQ32fOZJbuSAvUVOLTwcZKYtO4FUY7tIfw+k7JUGUhhJIr3M
PTNtFMBKxGRGx64ZV8obiQSNbgRVN7S3T1Wm1e0tuk87A3QXc8x4/5ZOnxXn7ueDmzPSOIVAObnc
/xz/VukcHfoF9PNn6/XkPjwAh+doJ+DvAQITLV1IlLRFgSV0HF7qmyKleFjh/Zcv5yzuBrtw4jye
eum4zOHW0hpottfj62yZmmyg1ueNqrWKN37rfFicblrwkeidq3IWL9aGBZ8rHYNew32zusk0eFQ+
3ZbJEulYN7+68m0hoFLAgtluDmmlCLW90kby3F5/QQSJMZmse65RBzKSveK9NyXTAXDg0Ta+eIsU
7Bv0/WYjSzyCP7gS+QLTVitPpdebrEJIOoaRtWfV4wojzSJbFx7reSnbS0OKnLxdzE4ft6kaYhu8
9t5qDEXrh9WTRQ/8QOqW31xJV15TyftlqId4lHqwxCIEu2aKwl0vEMcn0qT+Jh5mJ8dkq5R0jFCx
ya4T6tRdqv963KCkhX6n2PvHLNnGsFDPErvkE3i6Z30Cor0YNwZvEpSie5kKm5lbfr/XsmPZLKnK
Vn+b2p8DUlLDixx1JWrQ1e1G/sR5gexpjj4uPucHMMIAhZvyd3BXaD+fIKz05U2IIbjaSbcyZvTG
IC+3lf3L0gxyMQn6IEgHmbGSC/+5P7pxepvXtjDcwDeliQQk7csUS+T9W3nxMo/b7BBj6DyRxfb+
wmVmdM2z9eEPUGZrmKh6Ubmvrt8DcobGE3iLND2tUQG16gokvYhQUrCq/+8LAGBoKhHgycofqCjQ
H4GKg2U4R3lVkw/s+cEmrChJJyyhm62WsaEwJxU9k62ZfWROi4BhIxFXtzOTbgGnYqa5zr+ih/l0
FflLtCIXo9/iyiFa8EPZruXqa+1S4iLEdTLZkO8AfnbcTRVMHekqodTFHneTIOjPRTJWG5KwRbsK
oNIleAycme/UenE1sIvcIMdxZbuhQPFmI4WYsBAbm1S1vDAP6nOf/jIRGzTBJBhpDDmRW+K/F9yY
hyCrJyULbWeNieiqVSDYSUfWVLbz97RHWl5BVaIo8c1aumcHgy7pY86TNB64i83Om+ITx/sts5PV
wI2Q+mohs9eKq/NPoE4r0fdtLWW5Rgnj9top77FideYgY0cF8hdydGZgbJuT8ybaOOC3umlFOLa3
18m7S+jDf4bbbuxuucztbL3u+rDllMQO9qZF3dmleMjmO2NeezKGTL7lgn8Zd4xov44z9hTzmBMb
4oYf3sRvJCEAE570r4nsbo2+RGIvwBH+qMhwsetygt6OhHNDCTag7WEjy1rWeOp+Qkq5RSPKREbz
SulcDZJufqWmP6Sk7z4UnhSEDhyWDQDZXjFuCGsNvO4g6vGMI9RogFAvJiAeIKGlof9/5SQICf/A
Lh1csn3T/H8hD26kHV9nCt/WVKKfGLK2ll/Ixa06lcMk0d9lgGWxuj1JIZEqt/m1T7w3YOHtlsSc
tsl/anYfGO4i9/4O3s1fyNNrKcZm57HnJ1rST+0bZEwiQpQz4cs24849MNt5mpMk2GQbz8StMQte
hE0qkmExbUWXN9oSyZ1RJ+O+LRA2PdUyifQ7AOuVODekjybUdwIvFdCxdrb/QrBacTxubWh32gzk
2gblGsrpCOvB6qz+xlmuAjCXTTtdWezGo+37DD61IEooJPZpck8cQV4bfY+pBPdXODTzOD6cJttV
CwPXzyro4KZ9l4pX4UvIbk7tka27qoLSxsIqv5SXhx/zeUSNk7paoUYD2kWBBCYBqcTRctc39Wao
xUvADJRVso7ioCl2/6j7gW58itfOQ9SX5Ap0jTLoASj8SdOvLW4a2eI+T89vMZwYdPL/ktfdxv3+
ajwQLgXPZYD6LQNoZuhWjt0n9hF5mFuO+ECbbEo6PJCi6i6TKGup4EYcEJVMydylQoFZF1BKfDvo
qYgjMkdBVVZp4AXgTqCgo4fINpqVGJnSwdH8lVOjR2GmZW4G3+TjDazTEafPUZ7+LbM8r33OpoxX
I4mODu1LSBK/VX9h7VU0/exrmnfgOjUArYP7N0WM+QvaI3+hKcBTCTElkbOY5YXf/dZEfR/QDHPE
tvt5jdSr55yeq6sd1eAHrONKoUkYkNjJc1aaA6bksHny6v3n7jvSXHbFZJwZXZEksUkCbWpUnj8N
sc/EWdQTWZdTr8HnVBYYcIUdFcUCr8btckRM/7c+Z191OIeH8CazHLjTtZZlYnt7YgEN7H44wT4O
veKuN+PKZch9o1Q47Lw74t46MVxyuKjNhmly4UNDZoHyyU8yfgGdjkyK+Y+Pmhg6400w3KdUwk92
9QPu8jNaAV/5lknHPQIPKhEkoknnTAiU8qBvboo3IyDGyVWM2fYaKzHfL8T4c0G8dk1rNgDmDKyf
KSiL32KJTlAni7xAEqhOu1IalXSRkF/hXpUzKYOZE6y2I40GnOIvKhwx+pA8wV9z350nQexnfhRy
7NvyWo6QyPYRuRjV/6DEMW7PoZZ9xM3lcMefWiiVVyf1iDsM61eBDDwrCPLTrf4iaitWDSXNlHjq
euUDUPdRvA8a3iBGJQbO1yLU1VqdhIzpf6JvpFZdkl51S9qddtEoAnhZbgQKyVNCXw8k/qV2AOoO
48t1T5qEwcwkjxK0KwoJaSxXWE4kilZ6Lq7+AW/mJ60qE0aG0ocWTYBuNHvS9ht8UskbP99hFToA
yDc3IM50eHs9Oz3laZi0U9p4NiKu9ClBTQRzsldbJNTEJp9cEQCoeqNT8HdNQIjYgpt9hMGEcjwf
wd4sgygRJrWBq4RWBBm0dCJvqKpgi2NNorsoFxoEFDtlCqKFGPExpUZTeNtH7zEYQ84fQH4cjtWu
0B7/OnpEkhwV8n4A1Agh5mRyztoeo2vq6eFJ6vY5DYzblgPRQ8L8JgIZbDlPsyZiYDdjoUTI6jok
dXtvNGM3YHcqpsRrrSVqfWtwMEEENG6xBcyU4YGUOdeXu+3LB35KtjFt7nXtkP+IEoC0yAbS5wn/
Hnb14JrXHu+4jGp8NOrfK47c5E+7St+0V/e35RG8lJv5vXB2lPXJoHlyqtPiDtwPbFUH+7xVqzh5
vxaQ9zaAaWciG7xuIRyxBZ/tYTyAU+jF+bkcpqrMPVzdJYhxs0L639yq4Oj1yIyJa1m3hHqkjzj6
g/lzqFkp0vjd9RqXJ73498Q4tMKC5pQ1HNSNwphdB4lVqr+pShRL+kDqDvXkRMxJ2lkvCX1NnBj2
PtcCwudfcNAoSrClbhaGsBoNkzXaH/9NbPp9ZqXhNyhq8ykVmrmbMxJJWWqBdehoTyaQTQwesw39
YpHkodpM+nCM67rtzDVJ6MiX4j+HUxgdRCq7TiiTdY4fi49Q77P900hRDNznYQSZVG4Y+tT/IM56
NjFHRNPZyH+YWVTEU+e8/7nw5npwHnyVyNBo+12C5E+RzD49xhxFVS2uAVwtrEokKaQsM+kL8KJ4
PYbEH6rEKK0sRPWgfEr3BKs0eiGntYwgZ37eI1dMDJzk45S1wiQVeh9RwYY/oVCgFUKq9rQ24Mpq
7GDvLvayRLYE470aIMD5wfjyY4nrtwzbNHwv27JbvkjUYqvLeVTMpvbzZ3AUhwXFSerTlmlNNlc+
y9ETUef2XHCGyO3xW62uo/qV+cMh4Qa/cZ0GXMb4atNK9enKsIECWUbYKHhHv0fx6bX6iIipZD+7
OLgzkYaPYhLstwAH7Jwz5cszYxPCh/4EM6uZe3wxlIeLVpLOEP2DGhMROMAjREEdN9nnk1pmsvy1
NrnODooS5aS2fN9gl1XQWA2FcWls45PHAddMmHjswtvYBQv5/uUE+IhQfRDk4mjAY2i35CNghfVz
SxJyV+isTbj/5KEz3Y8TsbxW5MSNBzM2elDS9sdY6sRRfQfvDslpHKvryrb9TV6qT+R3UNUp8L8c
Y3ier8en6ZJmV3fjMDpTOh3dEOxYbHjAfAkyjnYaWN2kW8OVAXHlob5HwmDOIR2zOfG60TYtMvq9
kRXYSIQc5Sf5krf8hvwlrbZnbyYFkPneAxnA/Qr8eZc42wLCuh6llU3AUdLobEkakrOZwLJJmM0e
9mFuqfwpZJ0j04CrOEVYb79c76y539GEHZAzpx1vg25tB6wv3mAVCyX2nfz1gC60zsZV+2NXYOLp
1p9jCaeVDChRtqJ1bv50B/P8OeZISrqIoexu5zM6DvBBg0r9nVafOGNSOfavQSWy1YW1/GFU//qW
jMCKU0YLE3execYKszVkFOIU2JSfsrZNw+RU+nnj9ZdhKEx/lOZ/1p5hmvJfWpNT7xW75d6DVGTV
41PngeEtr+0Vfm3e3HuPLLRY7P74HfzjvDgxMYfNj+KDi8k72NC7A/tMU7qRzOyhjeUNCa6l7Jc0
PqOsKhSqN61GcITX9aIUpuYa/1/vbaJfNchU1HPj6UWihETfW4DvnFZozS1tjA7U3Wk9fPGBkHdb
vGxls8RLdCIRCxR0c2hN0OnQGPzUAcAk0YXD1pioiim5vMA+p1GrdFVGnjMqJdqn8/qnmNjKEK+g
lLxJAPNYdsnTM2aMHrvxzKd509p86Sy5VN5MoQYKYlhZIlVZ2C3v28HidTY+TNIoam6guQpFlHQp
pYUJ/uP2fJSIg5lh2LOpmkUHw/y3eI5prfEkepea+Xfp0IwOWS4ZWffY/b8G0wFoFpWGrgoQlA0e
GqzTgOVGab1v8m4evtXgrfP4dL/Yi1tfG5iLZoKzYmuOVq0G+KCs79JHezuavYpPMhFZ4iQT7BPh
m76vx/ZoiaCtUSm3lloKtQiDkBBQEbb6Rxhxn1pC5qBpF7gORNT1kjPMRQhyKNIAta/Ckx7U8IWt
RUoNTWId2EFm6Xe17WOpbLFwCJ5qRmF9+vfVmdqXwQIcuSCdp4p2ppIFj0drVDAL+noC5dLTKRz9
dCKnajBlj4dU77/8XkRk+vkJ8Dp5kpkfC7quv3iXukLtT1zcXs2r+yYpx4WwxMXszJ11rnnmBdeK
nA0sheuE3JvrSHz9Ec42pQUWx9GnY8m2u+PRQQfMvO0gF3CoF+YqDzHOMjHXF7biAz5xxrR19WwZ
l36jpGZxiIlBzbn4xTCYj2QKMbYT5GgR9gukeB0nig3FTSJCyHdzD+7g027oHjyLtAVrelR+dULd
NBzYoCBnQICWSfSNbfaWNjBF6zJAyCNxNToGW4TAxj0mItHiQWpgx3o6S8H1DuecfP3E4mGPIqrM
4J/EDdbVa6U9R53TGf8sp5AIl9ksdzve8pRUPa3WGm2//hraPav/J6yDvgI0tjIiPJeXtlRpLn7D
uQvMGKSoFo1DInrGfjS1KRuS/OZUPgnAZbxVqzeR5KvBNGrFKVOM30GmmbKDtR+Y5lQA75uZqR/Z
fJSWFpOPbWO2GNqyaGmpvAXqo3Af+feCxz2Sk/qnPHNbj2pmrOf6L0Kc8uU2x4u7JkxL7eNoEfos
fIQoPovICTrrYgaXk2A2BHd0dHN8B4vEGZpR2Z6Ffj6qB81XQmSIpE4ta41CdwDobbx/Zh/BiZP+
6VxD8xnGhOYNFBUDOvBKNprM3PwKyKEy1OlvC5W0X/azY7KmZm3dpV6t2fPTS3SxF7v9E2FMpPNu
0ONYd5iRMkkMRGy8TUEE3xBnPHzfBUyF7OqoJJtPUOZh/JB6TpXMwcj/nqZxbEYynSdUAcqDllXk
9prIMP8DUreZ+VopVJY6ZtOqWd/qCJR6rEL78h77WawYc857BegyYgM0qVc0SM7y+yUzsbQ3GUh8
PoJ2QYvMaspboQ9fN4ctzD0WiX4rAkU+mqB+dGZyxKydQwq10mLKtX3qNSgaQgWZzucq2ZU1TSTt
eyfIiSIhUXhiNh2XovfZFx4YrZor373pW63SBsK/NaWf7LQqEtckJORWczd4wUuVQ6FygE6c1Q7w
WDZQUkq9bSqGvhKxPRDvWkG5IALsO9RSbAkVErB0bkh9QAPHabDgyiR4EegvPtwa9eyTPrZvaWo7
Aam143Z9KNCX07/lHxUCg2//+mZRmZoSBNJEF7SSvPP+Zp9CsPlQVp/Tgp3uRe6kzoUYGSS39OJD
m168nTMC0GEOXwYwP0UCFBIdrC0JJnrY7Zhqn73IAyDfJroIcM78I5RfBPs89MjXXNdckRCFRf92
M1N7CZ62edVFAUDdpflqCHF1tLu9UqaFzXvRXqXkSIOrqWSwOOxpR0IODqGF+UwLfjsOnrSQ9hJN
9JV8dez3Wx26abnleJDIsLiw8SwoGiScYxefWa4Mmxb1p2hdXwusCIFw491xVY8LFCAgtHqQLpf+
8KSQL55LV9Rwa5xB5P1iDjoNBMrSVsNTGnDDSq1089Kzr9PHAjTEmxLJo4DaqswICX0s94Tuv9GK
lqgMeCvmi8H3BPuCqGYhh/WIwWC+Shz356HGxoZNBqwoD3/pM8qOxxwp8OQDQ1XQ3FBQ2nSZIIQj
290JN35NWqFV5WUpDnHMfLUwW8sXh7Z1HAVByRCt76KZunzZ8Xiwv+kZGpLlN2rWpxFWIjgismut
GLgbwTQSsdrxKBVh+nMJjq0oWkCucP24Ukvgd0iK12F/ZQGj3V/dJkCWjLQtYeYJkh0wnA4bxpGz
e86zZ3P1eEdjsqkZYvls6pBcxKj/K9dpkGFai/GZFpKWrdV8sJ+spTxFBGjqhvO3PaXfba3CydCn
W3pcoCFc3Cw/pVnMEhdIDZSJ+OGFBNDaS1S2hzb056ESgwxHoNRiWekCZPOa1qliGuNLG7RfbwvU
Q21mdxYF7gWWrtZT10y3LP5RPJcRYadeZBUUxtBm/uewU0nad38CSOTfP4NSGMAD3mFeedaSo9qU
ZhsIezAhvNJkB+2XjfVIddKcuxTxUcGW/wpAVI2qusMK7DKwoTXahCpsaBf9cQJZCc3/i2ZPPPcY
ASLn817+0IHRhuDCSDYbg01owTaMC2mrae1fzLETh47Rp+SV4DDfGierwFWAL0MCsmIQwHclbxKy
IA8wHA0KhWDUr5wjMKGwBq3jfdN9MLoOrHMi4Wqut01w5ROamIAOweonNY6pi6GUpQR6wP4Zikru
gKoIfhg5wCHa++MsIBTdeTbGntRr8GCuFsYNf9g4ce7chApxgfP0F42kI3NJIVCqTHCRboj7O05g
tz8/LkWU94payY+yzJ5NkJiTF71MC8cXk8WJOiv7PKTgB4/cVsUlSVOvDA5nDSNJSLS/rundNtiL
A1HPXw0UP29+7LnusdZGyv/vVwGSvBqukpOR9pWZXwhYbBc6vSGnkk7w2aeZOkUAsiiod6CKyoq5
X+eAgRfIWoSjusnq4R63tCAf14X/ecn5+nKqix8WvNs1lDmn5rEt3Npww5+uf5SoqTSUev1sTbTg
AXwIVoMqotyxHgsBVrUWj016ZzU6xArBYR7ZutvkJh+OjLxiok2n1HevDxSr7TEe/Gza2v9O86Kv
ugY8mv0v8OWhuSNyfhUuUFDckCKohftEpG2Q8XpZIm2xgRn1msLnFwXX28bvW2rys/lYJkFUb4Md
uVwpScHDeDqt9q2GF5xPiauFegsJ/gNuJbTej8FNE6bL40aQBKJg48JiXnu2/P9ApiRM6PXjBPCO
sk9g1ltsNP+isLBIPxSGdKLSHnPovJ4GFaQQ+W9b3RtNO1fn5SoYVpCV3lRg3yKS56HshgDXw5Uc
md47ryrDTIuiftdFZWybvmxHQ/MzDMKg9xaLrrCKaYhMl/g6ahe10HrPtYzzaWAL+gH2ecCnSwf4
XCDbV39HLdDMu4Cwcy/oiFV7oRlDgeSIMOAWssvurlPvbE/pBlKv4Y7HiGDRUO8l49/b19ygL6OE
uGNSlFeFsRAN70j0WlLxNzu9iRRKHJDfJZtch2gfNv6jnP5zD56cHTER1cQPUI08/Tx/GSIjukpc
N5pRQ/RZJ7wceVZVn2f2Vkv69ddz02EZFxujZqgmZaazU4wu0w+Pw4yKgb3EMlmTPDrjHnVIB9R4
8UuZf5jhz4Ikt/b2FhnJU0cy7hDYbOpdTLpMHIwDunHDh1kB7fI+OXIvoeDclHOe65AIbkp2lBqi
rcOpg7qYSo4na0af9FSnq0uohdOZ1jv1jH25S4ATZBWUc5sRpNpJTGi9QiGgyjwKSctbH42GtIUH
Pd8q+ZX2NGZlLUIgHOob2I/bksIVkOzmrhAxrbyUsD2zg6NIYTvDVjMvTGjtXfPukrI4E6O4dNQd
N3e1xlIF9qBDu7WOlPoLySmfjN6ryOifpIQ0GwTSg/xFYYp5cJ/OAy9UfPjICmE2ewfd1C4llJNK
co5DJkp/xJUE4/9vDjhvTnB4nUkwDw7WYbrfvE+pe7A5nmQwOjpaU8L5pa5/EpwOl3xRJhfxoiiT
S1oQheCf7+YChMspO9Bdhp8wmyeRZiHbq2dI8zVdeARAABZKLLk2cBoHNXMuM0ZwHjFcVWgKd+rJ
daNHK1biT3gRcyn9K4u7quRSuTpTae+5Ap8FtKzXl1ym4aaoa8LZXGU6sUG5AXNzi/OSRBPeLGQx
blNGdHZSTic8Wal1tOQ3PjfofzXSO0EB2HGmxmMgbkZxoVQzPfJxaqo3aZR7FCOqI8/z0ZjsxiMR
vORt9ch4mqwUY3BeYnI/u4OjMeK6Amqbct8ucvzek3It4iIKmxUP0/9OsxeqNGNp7UY0KLNCikgL
JKKtG3yUVT8n5L8OekwsSg592PrhjuUbNn5cFH0b5DOdK5L8jPnxIb0WzG31VVbjjn0uqPcvzvNx
rBTbqESV8VMMG1dNbm+gvVbr9sK3kS1nSn8rXj1krsToQJbja7pJjoA1iH2+bsx8R9rR14DJvFuo
PwqUSfmum5o1rLXTpt4hU0PLrnl58mtQAvF05oCNibc0Dfb6Fp7ZipiqizONRnuqsGHhU5kh89f4
Hy5Mfk9kp8pY/BoJyTFC4fj1pWe0ooI9SsvMJTXJhDjV3jAKmy1Q27Eu0Ri6cXYsSqAIeZ9cblrF
xkCfP1Uu9KT5BY3tPRWKbfPmaFzEva7VtomrNl256OlCT4UUeXrQZoiMjRXkVOyqUXfZLnpLEIkS
AbILoRwLV/FZxa6qaZi7h4/0bxQle3tXq6a5ZCg01iUOt/Zi5HX5pZIl78uB16qYa0iB/I06O9ep
u80PanYBO1/4nhio0+7xyQ7UIrErmJNH2xjiGNch4VqCaWvU+f9DNDaqpx0OTuZajOOtGF/S/NzT
5ah5vNb/EEjSID1Ejpo+ls8kJKvWdeg9sD/NWj7JE7UAMLWyB6CkI2bC1WXqa/dmFaii5gJUVFh+
7hdXvJ0XBiGmiaBzwIb3BQacausp0BhWbN4xGduq9xQ7x1gYtn+0SFXqONVlUTpPP5o+Ow0hZqBn
jLgD7+pq1b3WNWhBNhgVA/qF9eT4czbeGPXtNoo7b6aHb9lBXAhYxJ6UM1dcKBaBfbOaC3ttmtLd
3PKv1Gvx+aqomHF9oFAs6sckjRslDDOm/8ry94o5hVE2NFwPMkoITOerKv6pZns7Hx1Zn+Oo2hWC
3YhChEZ3uzsM2/jEOcbpPt/cw+CLyJt3FzexZZacWXypXdgwCa861yo0SB8ax2pTmQd1/S5uZSxP
rJRbTQ4PzM7YGza9igPvdm3g9PgKEAy3VElvVAgd829h920YIdWAruWLFHr/O/iXY7jGm9qOtbF6
LeiGcgjcGl2wYWwp76XF4jjrWbYzybZpBBW2iM+NuWnhJk1F6xfgfMVUnNqFB2CtU4uBhFt8MZeq
dc6LGac0BwClGo0dobW/dAOgifD5msiXKWfbWa1sc5iTQCCm/YtJTcDYLtdPs1qxKS8QfvJbNW/0
rKnQHHFoIxXeisKssG3fkFsG2VS4tKs5jBEeoRfdfddBOx7qbsCBKA/wr86POVa+ksxDgbL5VRdO
EyrYTEc2LdflR/wGyvQZpCq+lKouBkj9zMiozlAbk1w1QRiqIgLt6WqtrcA+xfQ6TQFO/yth48iM
YzTr17oOCx13S7atpcYdWYb2ioDTROnqL0Owvkt+FBkWxJfNraxbnxMQNm+0/XEOcF7Orffwsu9k
azCF7XVKVGc7Lhzkeiyu93Q7anyTIt4VTdIpGEiPLlHXyhp5klemm3kggtkLpyEvSamomH287yK/
RNWQhFNvVi2ZICs6ViVeM7STKuFj2OM/BHIBrjsDb9CF1+u4C6kEvR/wmvW0Xvg662Ok6lqDFVAo
yuRX2UgHyQESJcy3BqmHNR5SJ7JPPvJxYF5ue89XpUMfVgRhuvvz086Zs2vAuO1d+CcDNjNtTzSy
fyG6M0819zSrKvJuAG1AQhWBpIpur/Tn4E1Im7TjirrPPpSA9l3RtJN/XtOroaZkrvLtjdcij3uI
vuk1L784hGgd+ZhQg6VilliWnf3Uv+e/vGrTQnQqWRucPM+Mbj5An2xVg78rACitf8yUtN46kSb5
g6iuO3s6qroGM1XTy45UHisrTzgf0ciccMKWbowGi5KPBcb19WIiauFR65TvhlJXeLv8DxkrcWcq
1jo1qej/CKCZyMd3w0D1FjIGbU2BWYt5B7twdtpMImNFRcJuQhlLDVJjaP65weEEnePjcymq2+Ws
KNxmXd/3GfaCrVaDp/BstzgbVBlbxDm6h3KVNRnKg1H3x87Mqg3O2YpkMj8671VUlLnNMJkd4hBh
Uumwb42wR+pljUz2K04wTOOHxEXgwZ9ipadUdUinZm8IEix0sasELlyF9dVTI8ZuhAw2+CIbt/As
JyQcI6WzQtDAS4WCZ1rRmQ8flUwP7UxKmngW7PlQuSZ6ZhaSSgb9Wb4vNYeeF567sTmJvBCKJXdW
MJw378t/G4/YUaNlyo8pM7mT+ya1+2Y8syPjNtg9jbYNoax4qP637nTtPw4VCqbtWN3Aixw29DkO
W2JoAz5w6DYagRDQLcz9tPAa9sxYflhRAfIrIKBGpaVOTbPSgcskj6qOB6GQiciNCCzPf2r9jDfP
phrwFMDb9lppnatwvSkQPbCDNHPnoziYG8o1CjIh5oDf1R4DxzNbeJGz3eSJIe4lwTOFuK3Q8HXI
uBgXOdBKvIt86CQLpp5yg+9HXnnN8u9VSODXiLTq11omSgQbmLJ+qEwjsLzTc3LPU6FMwsneZ1oU
71NnH4/rNOp9DsQmuZw6CLaTceGt082Jxov8yk/hnq7vpOztbXUDo+OK4BxjDyT/5mzMEdBgCVOB
WQpXVpfn8fflOt7hHmlBRy8t/XvPwSSf9+xbdUDhRgl0U/0XjSzPr33tR6PpNtxpb4LgqdI/W8l3
JlJ2KUBEarNAG+zij5wbe5VbrB+3+CWEpw/FoHLApFE7MA6dtC2qmmt0NOiRWyTX2+JxwDaydC84
YtG4xzglOWk6J2wjgLPPttYKUsQZb2q+CHR3J5TlwD0vMFLuDCdFKa4AIEdkMRRkF3WH3j9hlbEi
7Ov2dfEIgBW3MjT5ZQZMQDy69LuFFDXi9mwiNhoWuQ+02wICzcpCOQWmGFYbxVN3PgS/HIqYC59f
BPcjIrz4HylrO6YdUOPmWQjsalaEyCiudFplghNGdRqjc7L9V5U9i7yRhX19HfjPjfAdFDM+6w2W
Q7klJxPRPM8vXijjSyAAYNDPjxfcqskeHz57h/CQKwbFcypLziJy4gNCsMbH8FXULt+gsT0giz39
iU1FPpaE0c/+AU/MLwzFPari4FC4ovyZWJUHEQMcj+jjYkCQE36Aydj3FQii0JnShC8IZd+pOCOm
4d3hOIVM399SlMHzlmho9f3MDWUaGceA5MGddQloaOKyZThGpc88aZPc04zhfRRp8g1AJWoGquNi
+SYT3uHlmU8oEv817QoHFgPmGluFsHjbatvWY9fHpjtDEoSXhUrdcmeuJJoH1TBWWQ+HkXfEwEDa
CLIgWXUQrWjqqfzCK7gjEwkyPhDK0IqMl5ArFY7p8cLN41jURfITDuyujCE70wVDB1ReTj8HRIFT
arjCatl1CEvjkiRevEPAuPg16N9GY9vDOktPCWcioV7PVWyN0UKLBi6/X5IzZUBYq7DrEZEMsEP2
C80mSoNrr0/X56CKOA5OL4C3OdLy1T3PPGP4HojzD5KA39wHdvpn2MqvTCkvf5Kc9iNuTHtx1UC2
vOGXLetSFPh3Xfl65UuN9+DY+iPzyvx0Sp8woF+9qcc/5LIjE4Ni8br2PJdIq79ymvzEjLVyvsD3
xv5mIzUKid+n7q8d7aXLIjwSE+aEg5Umjgp5RHMXYat7tS3ZpiAFeOOK7rLnPyU3ZqmarDTPw8KK
nWp2I9nyK4D/pvcAuJeHbzjBZ9cunUx+i/drcBGxlGiQC5yFCsuz6/Neg0WUFvI7lBSQUNdXZBHJ
gAPJ3mZodrx7eArel7MXdCAnqNSHztRO5LM5IDy/q0UpIf8pKkbXj9qQqXwiqafjpJGS6j3Ze4sy
JHmPwdtnqtubPcIfsA40EreZRKZXgYCBAyka+Rhj3L7sAJF4NRjgpPoDfkc6quomeAbIH05qoL10
lQMGEiivKPoCrONMqrFwdlf5cspHj/2AK6mTJTH56MXbVgmCfVD+vlZqzSY5ou1zd/schZGM07Al
hxdsrVa4W/lcvVP/Z5y1+nKJ1tif2a3MX8irnYIAW99upnAPZJlrLatuDiuMDBHMZInlV+3MD8y/
L1cFQHPK7cnh7H6Fp230o31imZtxE9Fbpp2/KB9MuuIhWEZSXaC4r19tLtte1gWh+0YiOdTfQzdW
E4V/VHKKUO+ZTXdobJcfyUYeryRtus1dkIidrQ7Db88UtJAbIE85sg92mXzD2Xw6Vv41rkqAB77o
vQ4GrbJHpbDRHU6NvrH/qciVVGVxhvNcqV1a3ItmRBc1XfrzJC7kbhJXQph11kWGyDwvNfER3lkO
BMHc/VhHkEXSvXjjB5hetI6Pl14+VztoCvdlUOhQ7PgmKxnQrdG6mLdWgt/yYMXFbBK+/CPxPXJw
uBKKoiKZ+s5V9Eli0JrRYRn4r5G7ESfRLSedURZi6sb/KwDWwcXzhcS8tjgF2auc8MoDV74Xz+3w
KEtyAgyA0Nog7SihUOtqr0IZmdFh1oNrbkF6CwTCFNIIeylS6pCsQdwJLJ5I5UdmDDU24kWJxIyU
Ctr2gz4QHr+cugUQXfW0PjrbUXyGyP2ArEFjc6LrmIZPfUV6TZHyB70wGMrJeiRYGelAEa35w5F6
EGMn5EdgimRkWi2wSmrdBZkbYAiQKt9A4ST/CM8+Pq49d0nOAydeJkQcGGnE+cvldgw+sEMtN/8B
/9UzoZVtAlBhs8DQFfnpbcQrgNsoXtRAsZbRLICli1fYgzlLZ//BUET4xkZqaxIHxfWWXoyl9Kre
+bSIMf4gWuwVTSwTcAecA7qwDPlJx0XIIRGxYqDeBTiQz6nRC9hyTknRPVjgXCsU9MjwR1QrDnsn
SwqikoKHBdxbjbV5F9rcN/jYWBBwIxnEZ3L0vy4YxJP1UVby4Tjj7CxaD/VP7sq+cqkAQJHAgynZ
vAen8wjZwduFGUTItRXZbU5urUq8LiIxpK8797G/Bssc+N/bccU/y73tsQLXCNmkterCZ1VmSMQ7
7ukEam0qvwHcBziPa9TArBOl/5ZX5ssuzghcz4AvOKKegHBmw8s9T8pVfeCgVUb2nHRsBBrVgiJj
Jb17UjwyeBT3R1oMOxVJsU4DZWAg0mNEae9j1eEtlvfHSuKit4srSLGeqFwNOj/8edBURygRE7tr
zApQfS8a13OVt/av1tIcFPzUicyrPnH6duOe0i7h8W3a90BJt6TBrWq7YoyNU3pDkrb4U5iNhecj
gPL5ujQZaG0eclHRW7JV2jju0iEq7YlH60vnN56tRITITTlwV4r8U3whHlwlrdg7Jk9onuhWGP9L
AOBFNwMbWlqztJQZ2ac3Y+QA+q1UFNNMR61A8BHIVCvHHiRhpwnQEVd/RAe8OFmnHDjkyA+8+ZHl
XDiGLVl7ZXU8wg5DJkEU13Zqiyw8eld6D1g3c6yOvicsNK3DIr+E74J8C/uzGDW0ZIPZyYOUTE78
ASQsflGzhxluTKUzlrGw0++7v8dlXAqXMrimfB77uuIq+jfxhl+1eM8MG4r7wmdNksqF9K2XCcM0
ACcB+ezGc+xDpHNfnFXl0QdO0jqV2wFjVL15588xXPecWvnweaspT0IEYlFQBWiDxMu/ntqn25rC
WHUfBAar/yzBY+FkijW+Rpa+HMWEaYnmu4g3HoRDZuHe4peRaiY8pkCp652Q6j3ofI2NsbYwodjj
sY/TPLvym86jEA6Ng6VauVsN/OgIm35JTHVH+3OgNPA9NXoesh5Hle8GIhWArs5dayHKPsePMZtD
Im8zOwC78tUqbvzgA24PKshvfmlfUdX64ho0RvbHvCUh5TwTd7Bnt3boX7fovVPLW7+vmUhVWrnX
OfKQ0lcXUf0u+WZdtqwY4VgAvpsPTNvbr3HEpybrR80KYlE9/Z4xp/99iNF67PEid/aRvQ83BXoD
3yfDOkVaB4o3EXy7pneGcDzCH3wjeFgkP8NEDIldcGYaL1/6+q9lIKCQHw0LkDb2L9gl2efbRpUk
5FbjdeywKGY/gFOvtZjKudUSrrDxUFFLkqr+ZqJpchltZcqxTvFVZk+v1zreSbmI3Uvwt9ekB/vD
jrD1eCiAnYX4MUhDmSzx00BjBavMYXLs3NsWSfpRHt9G/7ogpuf2bwtGB+/Rq2ak4lKdFWSNMCeA
QuiuDwIe8OOyegCrHBW8g8TNMf6tpHLc3aj7XqVu5cCoEOra3oQoNsKCLLA0cIdEdK9VQpzgMpp8
YCyQPLx5REYoie9di/il5D6wPBoWV35Cd3g5HYMISbqWE2z+KuTYfwS8R2GIREmHOOtTDXySmC24
F+J2QreHMt1Pvnw7ibrKSimr+7Wb2/mH5KJ4y6VMyCq7wyrvqFNLEjbEP45LWC5VJKMGwxJSgZWT
FGN6pvYhBRKeARZsyWneAYSYeuqV8qISzLTzNx16+VVe6KfYIdvx0u0S0oOJo/Z0UPRbaQPlCeQa
fYny2a5ymV4VZ18m1Ep/aah3/jnSpUUW7gtgS7o+1nJzUi99R4yjx6P+ReRlwLi54LtEbLtCx+sm
AfCZM0XRr3b8GMQFtXYw3z7dwMS+bOA3DNRBKwlDWKG1MgV9yyhxDV3qZz5heeFJKF4UXFrOHmS4
3RdqDPK/33Kax5Njh4U/1Vgfy36P0dxKaErnI085LwRogxYOA7eK8EhvgKhO0J9yVquzZp+7ZtWs
Ix+HIECz0AsF3ZZeN8H7AwKekZEyjcoGKgsgffmQ2k0NHml59XlddiCXf8WVeclPodWh98prcHXj
BVReazPAO8bfsz0pW7U/9f2RcFwX+XacWOcjXEO/4rdlB1q6HOF0m+ZMcvPzFNIGMk3PMalyNqsD
WHbiDO0bUrmeHazNyrwKJMf3/yQ4ju1jqYCJpO44AxuiHSKZjEMW7eD9s1OzB46hQ22PcLAb5KD9
eC4DT8C8R0zL2vFu7e7MrBGN6X+QN45UuztaRTADBsCm5MddC2VTmfoeiJ5vrzdNxvNh1n6dqvVB
8qF4RCP+GJVaDHVXnqWuA67vmVSPuGRWwcukqXNgllaLuTknopN6rlaJlsfb8zur7zGAVz0H2Dtl
vHvf1Do5EYzeZkT7Vov0SXAFhqGJtQTf1QjmLcgHUypFw0gNisvJfepT8NcazV2a9E1b3YczN5xL
BUkLfBN2J7zQ7ZT3sOTO8zsNp4lIcpkSES3HCDD5CAfLENGOVw08mxQuCEYzhQ+Fe59xjKu8xKCO
0PFec2isdDlVUl+8Ht16Wm3gr+r34Y3kvGriXqSr86k7pM+tGg2z4jggkROnhZWVGmf326yoF/x0
9qZwfufl87Z9CjhXYDqY7UjTlEzVYlF4SjjcsFtnhYUpj0Qz1oZXBrLgtD57zvQyAKTXHejGBrfK
llNW54v+/RVRhxWa8DA74IoxgqxDFjC8fsfiKzlYrj6k4avuXhREyrbLAVReJSB6sOdCLIOW9X7W
p01Okf2TGV2fVVhcK0XEvmbfm18fspeham9wXmekeUj5gCGZQ10oeWQb3kW6u4gkHVnOgO3lhWo3
OBbfNoTfAooXP8/XM4C+GYxvjpSlUSQPNFqp4kk6KxAudLMdsIaDzORg60UQ8YR3yqB2dMHFQCnW
dwXkNGO2BC4oKhdYZLGpq9cWs7Km1HnTttoCQOsC/RWlebuiWw9nHfcFudcfLdPAvNCCLEl5Ly7s
HoxsR6anxcv7j0n10UexRwShDCvBC8YV1WSwCuVuLuhnYKN4cRDfWu4giNU7v2GyJ1BcyErcEjHA
Ru7lKqrR1uOLZ1njQ6br1/ihhd9vPvy+FDd0wMtfzT5GEJwBkKIlzI+FNXQ2Qx8/ZpdMdN12RQl4
WEO/oaw4QUc6QH7UEj/tu6dzVfJyjMjKYvwIXLoecCarK1hN0Q3JT5d0mL4k5nJNzBO4PLMKD6uC
0RV++l24l95vAvnwm7HTwQZCY1JYo2L5yr2IZllSSsG31smSp+buj26X6eX85Bi/81Ciaw9kgION
DbcIoU+Wi2iR/sCE4EdlduqVj9ZSsvc1kyQert7DoEmnwZ2Wl6JMqMPcVBDVtOcUKso68v5vE6Pd
WWLSxfl0V5YXp1sukXOX0IOsEOIhZVXLfB8oPx+SzWLAoLHknfSLnf4c+wHIVwH0Prp+eRCjbzTD
MZ3FmWZY/UZCrx02lZyGsLMNIfHC1MrcJJSkB5ALyenlVSaDMQ9yfPNIC/WvspltpgjPZPzhoISN
3BoxqHoC0rNazf5P44bSj/iyQRWSBdnm+wOcebtTaodoiSBcu6H57r+ZlcYeRflpF+315ywmxUy5
XGf9TiYlzqwoTtcFiAbShYvGQJa354ONXf1c80d3XaO1gFmqZ1GTzEU474tFhEgo1hSdCDhNui+v
qX4zSpmVR4a92NvGR0ZjbEyuWdg4tPPMw4ASWwdS1mWShfjEvKBN58JT1jnnA+bK9yS//5bTIZ+4
uIrelc7Auchq9g0W7OY0yXvf3Y4KupMAAU48VrrizZeF8WW29QWsphXEDK6pDMXjeeV6Vzdu2x0m
nAL5RRysMU4Zw2a4U1d4pruS6g3KOiP+cy/6xUwkW8FOSwpid+VHAGwafPsg4vQzifCdXavo0bMB
vPJDz8Lx1tN+WoC1na1UxeJJ6NNvlr+TRb6Gdj1SqX44PdpqSlTdW8483sqenyJVu8SuMNa0fuET
O+08dPmP3IGHJ1/ai8ldF4noYJtPMMjtxeT2LQO6pHC7UQukw/Ymv+5L1PwWGsqzYrUHYJOWJlv9
arwf4rmE6dF5BHxvhE6Uw0qKuQsPR84OA4G9MKCz2Xq9lUCBDyIRk0flqlfG19sDOLn5BCnKD7Gn
XidpxQSmSOrYaSGgrihk9SIhfvseuFRVl6aPNSOWuk1+yH3UzB4kHO8TdMdUj6i27oNRwyp94Tdu
jBlIp/cKt30Np9a8awB3qs+c8DRuyHXocDYL5pCGarnuTlAu7vv6FWbl/hpDgm1CfI5JSGz4/raz
E2bNpNQV4kd5plgkgUzsGho96EAFDfezUqHhnf5FLrNxGOQaCe0SZj5vi0o5JyJ65tgxjvomu0Ao
DJl0MuEGSCYxrDjC7y6OrZ3vhMNUvTCypsbt8zVrfC81a7jb3yQpDfpkVATROPoBxroFABlf4a76
miJO++bvP54VZ08EeVBKi5jbVQILxxF9AmCsL/CipsdsDj+gsXKJOKw/VOOTlkHmgyhypNyTBH2o
sWCxEIjzGu2Ux8ppNce78qQzL5WaE9Q1OebhaA4XOA2cSz7EIWymCIbrwrQcEsxMSpcF7lqvLkUJ
Cg6tU1DgHWxO74P/oSe0VqrDcfzITzlBUXQMxyBpN+/jk8vw6cOtOzBp1For6Yuuj3YNhwac3hXa
dfImT2Vktr0Zz/55vkdpQmtSMzIusP7Uh344xkm1evDPmtCVwtmdZXhpzUGGA3MGucmBrKCtJF/H
h1H8D7+eTZJo8ZKrrtdvu55YPgRCKU23H/bcwo2w3xPpb2FRk1+H4sKYKKT0AdNohN+DC9mBfcng
6bXjsR1J34rC5RtS54Kx0Q3vMOn47aaGJzK9iHK5FluuRlVB5sz+9e/S5beqPzfQKt9Xb/xxnbyK
MtdKGQUm6ryPY6OCz0egvTeJP+K3J/LGZheABoIuPT+TLfh4CnyY4v+e1qjzlcjWeTGAEtAX76Yz
k/c2spjiunygWMzqHnWAYBg3bVKbA5ZC9SrbXpEPtgRQy1MVUSM8PiAn3xkuM1vu9dRoXDG7fOEe
JTs/EV6NZ0OgyXQhbvvTdqtwi+IlnWj7NunCUHwBmjIlMczAHH+3UwgTSk8LYBjbqQwpujSS79V0
zQ+XsdBq2Sq/YwbQeOsBJPIDFpWhr5flGq3ThpUqcjNhUYgdp0HRNjR3NNQe7MdUh1JplUPReErR
EPfuxwv7mNiyDWS6oMEKCRRejmIGeyvacnnuxaoAOkYnWXayEjNJPsvAwtwROnj+mH6e6A4vvOM9
bgndG+Zh/k3mxmIgpC/96nnwCAL2Rqk7LmVIUovQB2KK3Ou6FKbRr5V26X4gVUduCX1qPzduTsOs
dChskKl+8RIO0weXCiQelW/ycS8sYrpducy5ok4lCQdnzznaXystUn6y3ygiOyq7JkBb4g8sR9zv
RriFv5JNvHDtrlKi/NI/Tk4nZDHDcJESepXUxzkTavPw2oDCnuTWAReys53ZLyzxD1fw6pYXWnv2
1nui4NAH3zihQ8VKfROAJb4EfobqgIbYSFbALFyU40ubM2ZhquLsHSoi0lC+/gSZVDSGga34bAMX
+Y2YDw7Dt2FYY7KAJP1ps/TF3OkxnEzBGL/R0szJETq8UzFNN7QMJSon+s4mCtILYV1pK4yW3YTH
8eeljW8OZRiziwe+zUqX5XzUCPvCYRQ/ALh59mYD/JT7q6tYSLZ51IQUJTWEppw0xzKsIU3OZB7B
nboOqeYV3nwi5ZahQyQqtNuz3MnQdzbZaRT1qGwdNhUKgB/1X2ZgfwlY1+ojZtRr59w0Y9wOj/5J
gbhQvlAQcKjlBuzoqUzAsta7rENoygr6ajTowZkIU+QhZOXtpQQBNoqk8OwPKwMo6i7RvZImRkfD
XbEiqAy4Iu+ZcQKkUOBDvupvx2Mbbyy7B/FylZM6wMz9CNNL4qQUIRyPKpNUWxTNQE1sJJdv07jG
FEbSafn0ecVN1C3P7lcsAQAYtZEDzt/qAg1xeHIPS8Mwz+NDiWZa3omVObIw/WnFJcomkhKS060n
r739sYo4r0bCxsX5He1i2jwFp3tIx8XuUvfgJlJq/5RjoEeLzFPZq9RWhq2tbfTrWalVqgeUcy94
9znjtePiZjNn2kr4FqzajS99z5JXsyaUsMS4rLbEQRwJXbx9hcuBkOj2dEiF1Cv9bI09JU0dFlvl
POcDrsvXJoneJSF3c4CxDVAO0sm2+Y/fW2Hp+9KFFEzFJhVotXQ30P9UREaUHDM+i5azjOD7Z9OV
6QWbt7vrQXVRgXXwG8L9P9marCGjtUhb08TIz1Vj7OlOPqd4739Ntx3a1cnDVAb+gWHzF2rEHUDE
dksiXOkk4gmtB2+2TUMGAAIRrWZqJaixcdHL9dyGzGZPSHLxULUk+ejJ8IyMZfOYEDS1zAqOiwKi
7P+iZfV0Eyo32CC8dmywWHDNpYUfFd+V0rgZR3FgkAWk+ctx/jS0BSXj59cYdAajKM9Ae+PjGuGl
R7JdE8BMNBftuQmivCB10vO8QyfY9E793xiZ1LLX53X0RFrTbtr/XF+1Mg+eUP13wcOq0uPhtVh/
53e34C2Gf90i/SQs2qZ/d9mi/8AG4bswXTx0af6JZ+DvT64LGWCViEzA5ejtYD8SFqgPofIhcNyT
L/Lke2uRpnhQ2w1IQYCo/0eXwe/+/j+cU3Jp/O1l4+DN0BA9OYuIF1eBd1hmUS1v7DYtgnhRP6oo
g6alJ51T4ypbbNp1F93PUvzfRD6dLg7ohKkvG4cxaSMdmk68aDN25HAeElxhVZh2a00CcXpCOSSl
gxXlu/CyZCXv9bTsVKA/K/IiRbZgVWyh0hrEB2fF+EjMZV9aShJuLeid8/5CKiZzTU1f34yZMjzd
xp4d/5MGQcUXXw+Xdwm2/E22/o6GCEOiSbIWw2OLUHJFYAvvKmuL4ZYczeFSSlvQK+p7uu0XKq8z
qLEfT3gwMPD5y6zS5xrRmfSoigZhRakM81cZ5aVxz2rACozjkP+dFNd844EWE5bRz/FKtpAtryxl
XcIzyJr+3qN8yC2SEMyEHeqAgfqPywyZKPmTD5QS6I+SlhYDdB5no6K0lVmBLudFpyXyfhjKk7ws
U9tPUS3+i0gZphxcI81ffug9nia3tky0/KECy4ewE/ItMTNFNACFGu2NhrxXgWHCJeP+vhU9t2xz
Y0Yd9ZcZRBngK/q9dft/o4cJgvkjj5e3UzNXhuqJp2lmlQy6yDF45jHNcKjPslt8PRoiTnnWLPh/
li02ObPyO7ur2wGyI+0pRfMOOh7jeD07BbIXaTuKPeEbjpUYW/Dwoff6vWvRgeuCvjSiihDdQtEV
41qNg5UTmSKcsmptvC8+W2Kb+QLWhD2H+7JL2smdUis8o71ZfD/HDtKK8KlXY6wbBdHmPBFZ8lJV
u+3NddHa28feNIVJQrd17anpFGJbHC6KWGRXUC18wlT4z7XEUr+istQGehyhmLY6tvDThqXnPJo8
ZFxpHt2XSjcESsQMzmj/hTCQFYcfrK+Al8x8zK5mP3czynGc7cHCtenUa+eoUYQtjFGU5PyGzrRO
c0pmbvMm7lp7o2SgLyQ3KNrku53W1rcR8tYupmv0PQlSTbEwnXr8bG90iz9FLLldSyp+GuTP4z/Y
OdfzWpTV6asuFqwHcaCprTdTc5kLZPMMVMxVIUm2bb5Id8jrVbCPL8S5A/OmMzI33rCmRtP3nzI1
VgmugelmPe/te4+SQYWWJyeuWnZ+QeDVnFJQLhgk7zLzFmmaDCe7kQhfGAqD0BxPOZdvYV/4XJ59
ynBYJ407UNkdglkN7WizmmBn/VXkkISRdrbQ4LHBHLfAEaM4BRaBOmeO75GYel8zjw49P+ox8F2k
oCuzodYIkXe5hacoT1KUXq9NC1B7sIo1ByRl4Xd2a7vU2wRWwbDxT7KcZdX87ARg25hnhEUBJHlx
4rSj/+BzMPeDEdTSLGh6CXb4gBg2A0iSiOPbsokyIcZxRpzqWBv8DyCSiMGFk9xqeC3vdQEAK1we
S9q3oVL/x24tnoi159gDa9yKETyIGNDqWT39CFuOSFRl12/se76M6t46rAn/qfGLrHyydBTUjG7C
ALaYEQtq+1zTIpcEITDjFH0duH/Aw6HA67V0BzogGK5D6xvuekjc6oB1sdw+lY06oeWqNgpdIN3M
fSrU8MzC9hp71c4oeTE2TBgLaFmDuhI/PhVCSJWhHaswMJ921KowwkhMrVjaEXN5r29lxWRAkDbG
2QdYSPZz3gVDKSqHcKlPy9I0KldKRDqahEWRBFtS5CWqPg/h3H9DuC9Qbi0FJ8otq3bMQ9uCTUod
g7qV0Iiu29mX6tgNTdczpxlsaG7lGIcaJylfvnqtmwqr/J5Wr2/2B+rNDPGd39klYomvgRnh6syP
kwYLgozqzRnsT1lpETTGhqVRMGgHrG0/i0i8g0xWkBnkBJkQy7r51cWlFKmlmwO6a0lBIpMk/rlX
6Dx5p/StfU5mF61Ael9wrQ4YEDIiDv5avp/oQF9j8Y7ETEK02zdKf9fxDx/W3YHx8djzUzaVKhMc
0TJSORLXzHzm4/67Vt0zHVuWHQDEt+WoerDhmIsiov4qJGzISh0mK3s4vm4QERTqZaQTDGoQfVpn
DKuVe2iqnCjBPmMDDjLCNuJTKSNujLwCgdIrUETX/jZHA1K5xdfezcCs7hHSi9g+PeZXrM96dfIU
Odq2dBurWOH99JxvKn7FHffetQ88PRlC/CE6sRMptRZDrtCTDK7QsDfIpe6V7XeJ6cJLySvj4LOJ
+xLgsmnjDSxv+idZEZCR7/z0LhqGX7WycbYdoFhwqW7ouYShtQ8LKfhySW5l7qAv5AxJAysCFopJ
FSLmpPcrLGoVk0+sw3ZkN/JJ7nTHVCwZUz2TntvrTCCgPpACR8kuWY68mMd2HsTLtxsJ04sIlLWX
K/kaER7ZlhoOZoCyfN9oxCWM0zyrlKJykkVN5hRITqJyolNQUNFb4WxxEqtqUY74xZaf0GVs1NpA
SA492g0q972/l8YmkHqFbpk31SbqLUHkeA/ARkhl8TceCT6oqO6MsdwTg3b0I2/FGwy4Ur9gIaku
XJe1Y5HOkMaBwV1nAUnttwzY8mn8P6IjDFGv8eNQbeo7Vx6adhqL93hTZ5KFWGJ0BqkpTS0Y0pM8
ZIrViCfrMfoWGGEor+Ij7FTqw9IdKOiyOkIXxmtxabGPp5whyT9Mc37zP0k63VoAQonUHVWQiTst
4JxSaXBPfDx2zB9i8PHHR24iZPRer1KRspBuz7G4XqoF8oT6hJuP9Twg9klsDuHzr0lnFF0L7YxI
I3jItHf44OxYhntkkF5PDCoLE+clLaKicg5XYACQscRGCMSVQXQVZiLVFlKLhgf4KtlgZ/LsfXPo
b9hmSxcYQcujy2U5LsxRfz5tIzeEcp58XBBkvFFjcJFFllmAJmMjtZEK7Go5zjP5FUir4cO7Oo2h
4j1FIkgImvOMq3s6Bce209ARHGvIX4iXPe4QkPim7eaQ+VuYVgfZ1ZRjDTlTtY3TwhhPQDcKMdNW
Rib8U4R78aXGmkiEz7QKNXpr/RwqABNInftL1I55CjvhBeMrgfLkyLo2UzQOyQDjlzSklu3ST/7y
aGqmEdd7MIP25DD5DMBNF5gBpz9Azp8wr+VV2gi/P2wkpsGvqVzzc/2ieXcasG74j7qHKMB3p0On
lI0YNRELnwTOAC+ycbj1egWByZ6LxLa6nM+NF/6wfRZMfMWvE++oGmjwSbdeHDwGXJyYg02GlM06
8+vL7sqQXVcTy7+uNeO9E6qhT8WCSG4jv7wneYvFmbcPBva9MM0LfZ0BclIfFHDtqLO/0He0UVA7
igUnDRxSJ9c4gEdqwdEIbe18STnEn3Rb9glbeRMuxLdgHiahvlY4iFxopqfUeIOdHWQ4b/8GSXX8
xKCNdKd3tkYTMzVFVtHckIH6Fp86DOMRaznSHvcPJLMGxdmT2sTGOHUdXKn36dM1SlUTlLo8Uo3D
j8SGkJCysIB+SMRiVvrsdptVYBrAzz5usdjLffaCqyhAqDhIVzOAbsxD8WnQYS1ftAy3gBp2p7s3
+YwBBaD+IpT7Ho6qQJ2Tv6Z7f6+Sd2JDpYyQdg60HvOj2lJMbPvn11/yzSa/4rf0HzdLDzlurYSx
Z4kYihhRR0gxIneKgCf/9LGt39LDeNDbOJAU6osph/qEPduYJzDDWp5Bki5PqXwbeD89E6MoceXn
jevYEf+YQQGcAPMuKFcpgp2t++0pTD2K80xFw5n0vn291rH4T5N0GdD/mOJZ6eJblVbFurLDadSn
NgC3Zyhv2WEFUr2EfWOjyNpt6WgQV07jcjyAC1MT377bPBXyEUFsKF0I0hgVY90NxSkIMdjQxels
r3bsQNguRzX2YyGa9seteRLG2bwwnLJRh6cF9z+bnfUyezo62uqX9FGVFHvJXMgyZkoGQYxYc7Sh
BUFiCIoFhQsr2rmt6QU9P1/IbMZoYoMvru/EXbM9URVhf52zFAo6ynwg/tRZLqS6eBWek+NrmjW+
Kt+aWagFv7VrEWJw6Wu8jRV8CU3xFYYdDALCFrFtiSrx0z3J5kMSX3Ro2GjDnPgRmlo4GoK5g56r
4KgQYe/QLrIvNFkZD+hZxRWum3rbFyFQf1vPJim5hEfzyGM1GrhKygsRkIeGeO+z/e6aDXZ5++uS
qzeeVP+8WGv6UFPJKQjX8ffs+sO2r6sfBTQNor9eC3pY5moM9o/4GZ3mJ+vYFuCqbeNTuxzkLhr4
Z7E/ATQFL0fvB679dnYWTZbfhmYSGTE6QHyHcbvmmTO60QhrKR9K1iuFm6wz0mvcgAfmtuz1hSC5
sYJ8VYkQogf8d5I9iiKEsVXG+yGxcB8C9q8Kj2GU/o5NR1Mkzubg1izdI/3JtrIsNzL8ePoTu/ZF
q58auv7XUyaDyylpjN1VV1jlZ3kDhwIgssaVUw29g+A0j7VWmljQQtS5FOIc1nYIPtbfgHDdReqQ
bN9Y/YWF6eZIBDwEYTPUlRAodcequPokRLMBMtKNcvxRzpZS628q1dde0uUwapPJBc0OgzlRNmZz
sTnmPxFog8+sjCJ8R11/8Kt5ZsB8YleASFtD0ixSLmt+HS0OvlgMY26GBxlPCmHL9l/EjAuI8oRX
QOu1406q57qyOxevPWePNPBTvRRySUMrjlKP3T29VGkYXk7NSdyi9zBNANMscSzhheFEQGHojawZ
g6pggrTKFY/D6lvjfj4b3QC804WoZ7OevP9qwWK5v5FSL8VWBhY/VoVPbwaAdfAn/yNU72xcEGMB
eKEltyZJw0+hiLAOK6zK9pqPaFIPXtQKiRQ6KF1tJ3doCDU8u0Zu45TePwdTP99F7OsIlFjBXj8N
+8kZWVUadD92qLxDmN9qKYs/TvlPCtTGa+Or6IRkBnhIuc7G4DgDgk9U1TEzdGSKAIk/W64nxCsA
27h+K4pxCB3ekALH8s1MRL4riRPk6mRrN5sopakDnsqdKC0nHDnfYYqzjOpb9p5QMvR63hJ5pnRg
jbUtnkARdbpAuqcelQaIlik7oLGOd5UiiFrvrQIaf+JDdQOWfxERR8j7JAdXX34VDIg1PpOsMRCt
IIql2zU8GUHP3LhV/8GiXw/gUyML7KlyxyhiHRvm4ltCSRiu4NM7cyQiDpaUXS5dmeAGA6eSv56k
aT5i25ySrGQpdsyeCBmE0APdsrOUtR1EYpgVpRLczD5+DnUk4zjd2CrTE7nliHPaMJ2OHxpWKUgp
UL9ZCx/lVH99VNsFYjEY8VXGjILBvi54VrhZ/PK0nFd3LjzEwy3Bbm5BMkKiJELEAsybfab/Ytr3
W9o9OGq91e2u3TXfD79W6oBACy4ouFWN+aZENrQyBehEF9Bj6gi/R5buQ4UcpJqw2eucqsReMql6
QUfNmDgcRIIGUiRBGArYUI8SFAHLzKcWcpbb0C5XIkHwFHE6glusWhxWbRoXVXXsVW/KxDK4Rx0n
aZu7siuxEAZ12axFgnCzv0T7LZUItjq3rKiLl11VycA1HlZ3f6GCDnFVtKHR+HI4TIcTSS28H3e0
SdjVj1sW/KfDGWH81XFwKjoHpObe1i+0Ax6GaOBKy4tpG/alUZcuZTdPRVya3V+MNszidEClfWmj
IQN/R3rE7XPKRHRFiXS5mOIouPVzasrAyokFKMEm5pYWDiS4OM8GI4v4ZCRc5cEbXcEQRgjBsJqG
JSMLmEG3RlQ8yt29rMNzUKsdl0sFCgdYlZ/0h8fPL61HUw65u1SS027SYXaYzAyFdDUYDDMQ9kfh
JkGEASBC0PdRPxttj9RPF0vvWe+PBRjgMqbjThFjYGHuS++DyQGSg2N0LfLpRTQL3gOnVRZNzj+C
m4OD7AC32pchZdc3bDt/ZBCyUcKHHVy5w5oDOKJN8l0KDNtGMKippOxvxtgCeT8P5uhAVVrKji2O
/0d0tBmKyUmDilWW8rLs0ldAi3ytwZ8BcEq9k27YROK7Wb7XK11txTBFt5OEstFuiSyreMRHBjgI
UG5d+K25/oMmX0wo6SQb55IIQZDBjMCDH6QW/bbriJdR64m0PWKc9h5kLY0UqP0zvuC2i074o207
X2x51RWWnNSuXGBXskGWl7772blk5cEqiv3uGcuuKxU+pIMPlRDsbgjSlOXVYV71arFQ+0+2B8g6
bIkvAWJsk+1fwtBwt3/tkaGHTYh3wOhVlrDOEzyOlhItjhNMYhu6GqiM6MwmFKtv73MLsn1CRJYe
zz2w2vd1VhY9RAKu0Tx10uR1mBzRYGavG32b7abRFKBtwTNNR2sQufl09lM3LdQrFYLYKZuXwjHf
8bvD8gFkhFnuvxLvJvv9PuUU77b6w3ZHNzpn5malJvtxAFQR5Tn9UdV57NVXzlChTwZr4xEoCbz1
SRLu1bkZGiofAKZlj6M9hf7qvpRDoNhms84VCWu+IX1dph314q2mZGbjl8trnpRFWeXikX1UUpx0
7yguw5Ly39Hek3ahdioSHyhYFcL5fAH5ye4iS6P7dVzUTHxv7zKPreLApuPUAzFu6sTPzKQMaEC3
jb7tABxZ2dBPzbUUT5JP4Yl8F0MvR3Rgng36Z3fqJ8bh7+1/yabEHaxesIjUiCJRWLkqwRdGE/Ul
qwP5rQBQEysD6NTZrBE1goohqzdUI8KClM7UI0k+ZJUZrOv1SR94q5JgS09pH0yeCXWnIId0w/WP
K4I4aUy67SsVKVl748vFIMmJug8rhc7aY/3CtOBGU/YfYlFqX0wc3RggH7E2PmHkAipylt08GjPQ
SNsNVi2Gqk4p/vktK2m/oY6FZPBMu2NJA4kB2IjV4v1gSa2rrHfcmSenxjMmkxDeTXEhw1aR4cr2
cmoZLcvV61V5l5EMATC7isBHusZmMbmQobF8u25aDoqWQu5X6FwXFSQlwjd2qugzPiODCujUyeeN
o8ljQnitGh7tWunV7Cxi4o0UdsO2EUMiiESfYR+5ky/Cv5YIcuu7QO4WvJGJ5Rzv5OsX/+fBMSy8
eb1EzmRP+Nz1RZCkTn/4Nx8vQCzPjiPUn8LI423AE6FjEH9Hk9QWev2Ef/1bKYsqELnomDsybZZe
PrQ9gE6kCySUZ2sQrp8nFysnBm3vlgQmaWmT30Yi8p5ZCObU0k2Syhze4rO2LrLkMR3h3yD0RysE
cxX+HrRZU5t0pdF+vziviVQijy/Q2tJ88/r34KcF9K0XGyNpdPumN6Gi2DeMyRvCT5Rqq4ELtO4z
43vzAMdlf1bl5giwjKQKu3on7FGesryqWXm1IxIIZopax9zC3N8XG8w7pem9GAaaXiN2Sg+GpxOg
Fjl9veh0/da/Fejy7TNVNYNedNMXpQcm+uGMg26bdbLGc9v6WpMoiYodEfikLShVO7EolgsRyFtx
gNe74CZ/F7GoolTkWjbC74F6ay2HUbp6+1RjPzW/9bPyJnCIOdCcXTVsulzxiveBl65shbgqpUdp
SigPYv0KScUm12iQ89jsvUTRnALz978esoThIGlKSZatJsg2cEYNer9ywvTLnDVRw/ANFnM4xW7m
PD7eEg0jFUBjyyXXRQJsqDwHKoTu/X+fYdQJbEITRF4qQnTpdTPNIDjt0/3WKVKEhVJmWTk7Lq0G
heuhDFPV+NpGeD57DiBGH4n2PtLwSnkbGCAMYFIDxne3CD7A0biekruS7wE7qn4xP4N+l0pyCqbU
xcYwafEES2HaEisUSZjVnDZFyhFlI8g/xJfiZDHklbMqmqmfQ1rYtsPc9GaCekbJ0swv5hVQHhND
CWn32Nobw93oFg+4d6tYJULH9+iBcYj+wWhpYdVTsIk4Fj9Ifs9vrFRotHQHIJpkXPccmV2YgOSv
yYcbqtl1qEqhJoWwIjzgsGDSkXlrSM2EU+hVVNmOMaeWL7FrmD9nuCXhIGRZIYxj4t/6FHyJYlnG
YiMswcQl1UB8vqYH7yLbYrxx1y5ML1VbdoWHyqMtFQ7FZNg+8mTs6/XNUIM4o93BlXUXbNWU5eEe
/0OdjzymV0oDv+ixV5XCjDS/IDGs+6yzocQeh6gksAa6HbLl0zAJczxb6dWKQAiP/2mJw3V8agBP
jEPm3EJhlmFupS7zs1O9Bn3mfx6p5HayDwI+qXyWYoRTEsUmZgkbKEc7MTQg8+V/8KprVJHu4/cH
/SRYQwwZv0PQEAs7RpqNH5FofLOmSbZRI1f+shNJK58DOQNssGvy6NAkLd/EI3O/32gg0kishqyo
I4/V4PWSz6/AW1aOga0p4ckNfLSmxTWJlGB1xoAoKxaV3sl84nmdo2UJWplbfgR5z/8aX0yuoqzy
tU0BX0YyFXXq2hBjC9iSd8yC2o2u0I0mU4+kwcmNeExRA+j+4+vGsJo+xksBrFr1ryCziWWV9cZq
6gOpEB67bfuRExeJAiEQ4CAkEEZG9/GiQC+gqJrLm+SI/B6pPQUSU6Wxch5FJuksp7F2LyL9DtgN
eZuJlP+v190td965K16MNVxQtgRPGS1Pj3PtYDTOjCMWYupn5DYt1sNo6iJY1Vq9G3Q2HQE+xKOn
+wrXydkJq0YQnh9tdF+3k/YoH4IwKtQu3oSnoAz+dTPJN58kfrzpZ0L/mOkhv0YEresaS45FxRg3
g0tXl9u2nbkP8nRJjG3pQ5DeOCIWLOEz2BEbd3R9ZCmbNR/UjFqk0FNeR7d/kR2+a5nRcblBoUEp
Kzip162qcSvR/vSrRdnXNn2gjXkaubojg17LIFVCnzGRUapd00iqyg5uZzMashEEN37ThOQ7dqSr
OH1DeHWWUJlNx/gbPtWiJS+b0ZBYVplarFGbT3JyNxN6Hj+710nrMIBfniC8qCZvFbd6SIgTX13Z
9QNfZ433Wbm9AwOTTKpMbO10QdbIc1QSJPJNXUKw0XjC2wV3g3Z2RUpAdp4f5iuIe3p2JUh0KLvN
ADGPPMEtZqQhIaA3CDy3WNjJOB8usYXM6asotqBdTugtyCFnVkBxkYr+pXQ7i6zUVUUyF9Tf38YW
LSviw1QpUECpg8w0kSewbPApQA0U191l8XNRaMI6lWz7xzGdc72R5ECiXBvmE123pMAKshWoXC4B
OSPdCZKLb1fgiwrYRx2P8TvWZmCG/0X0JkrEGf+R3HA/TZvMhAx8X1qStUIFMhDJLU+DPuHsdlWn
7SqYZFoC2im26z+y4myc/vpCm07OCpwivFI3L7bNcdoS8byxXq1ocQ+31/9x5gnxfFsvYP/nY4xJ
UQlLm/5FIivtI3mTxowaI6CObYa6rN8/DIv5eF9tnhjCt+vrNXQBigfpJsvW7NlSM7sjkB6zZpMh
6eg2YxN9QnBwjIdtrIErBRmRLKwyZ29wJL/olGuTPUa0uz1Uwts5DFe3H3BU1ni3vL1ZEbp5Y80P
KbHrCAT7rwu+MuttYUFURuVqsdd98++oQbvP7axOFltZyd1gk1e2eDfUZdRLKbogBgWso48GSgHP
q51tq325Bve1GO3SLpTFUEf7M3PtAdvV0a7ZVcW5LAfOJ61T+Fcf1tm5ugqGF5vAuIapkwJfLiJH
QP7PH0b88uuLmbml900KYUZpKw1x6Ju5Zbdu72yWGmmyjKap8glYzAAGRYxrHuSu9DAX9Pd8s0OG
YjT1bsNykLHdpBfvN7oxR6P/6S4ALg5bMJVKIiyLGXq/W+HTyy1K+bkEKk2OIQGyls7yIfH4XkPH
diRb6TBaGkwwpAzgJg70M8eJcvjIIKBnwqmrZk+TdrB/C+3QKOWZIqoeYamB96yg4S4vrbgK4lBi
SM93saRVUBbf7shzMVKEd6QYF4vZxM+RUj9ZhjUOOXY5kGNAogHV27lf3ufBRYTiC0TFIBWVXu/E
Te0wHidwPc4U3tSNH5sH31UDBcYbw82MRYjI6dVzn2nDcwtd2uISu/MD4NtpctfEj9mt8Hec/l1N
fdH5ZEWVVUnzSJ/jp20yXFrjkJchtztNHMrpLMmsO4u11jgPJZ7EP37SQc69V2zOMQx3dsefmWLk
aFTBoUXevxYGwBV+pUz53LWYa6Qj+JG1Slf7xpi6WGt7zwKQgX3XL2FUs9SYdlmrlJFMwFNEEYvA
vEOgsRCvGq9BrwuTBgxL+MAVbqXIfDgJ06yOKL5OTi3QR6RlL0SUNrfFF/74L2mfzaFOQlsJxyWI
fuEHy9/95LpFODlpOSAIosoWB2x44Y2Z9up6hKSGZTxceuD3BZdeGoOxpoXmaRoL8Asdat6wYVVB
MRxYCu6j8PxdHa6zNItixmeVbni+fP1J8MWl4PDFSPBVqstpH5VYL+H4kGGPvvv4exHVPJIot3Ds
btryxxBvQOOqolcLdkO0TQv6+pWp//ZMmw5I+VFXB/qN5eo2CzHhBXJhY/Gb24a8+RJfzVUvHv4O
Rksyz7S2M2r9kfvcz/F769PVR+OsnS1b8Hw9n50Wi/yF3GU5/8Whzb98S0KM7mvFjSdTwQF5tHRB
ZO6ZSuu1Hb2A1slJY3YBOjnK4zKk8poTOs0ykbW5XBx5D66PXukwbJmXTMLS96fU2BGPesu+9T8B
TthW5b6Fh0Cak+NlaidDe0ln0LjS2ZRrA9DBSyuuoWrUPS95JcNP63nNbgGvmTsitdWC5RcXmm/G
2qGTHjAI4LmwJKQGb7nA2/zAwiOH2XcCSFrFw8du6CMsaCxVPWEoYxJCvG1jx0VB1CQHYQQD/Raq
48RXCs300JlQPM7bcixtSO7xHRUfFYlQIlcGrFrnImfX6W+2uLP4fwnbj9hbKYVuZbQ6ObvMsJQs
8nxP/zBFr+LGKu/CWGpf7D3xdgrextp3cE/Z+VPqRgUp5dSmV24c5IFl9v5PYpZ+SPZj+OA8d76S
C2QU54dkzZj5N5wr2I+iIdnqVoAbuX/Xpvi2wB1Gtnz/gBKbERjpX4VhIlriPhF/FxlC+jHl6hLU
LVKXIw7w7fRe6ZREgWwZ6//B2F8HUQM8MdUk0TVKNvp6CiI4CW+unbFMTaZ7pK/sihqv+mW39sAn
zpk94pnicrotlu5DeS0LQGMev8+R5B+meh2TFYaDaW8wKVnlcfUPw2KiJg09oY5+QyGVqisbd1c5
faLIYWlUYgttoh0tuaL3L4FoUeJ210o27w5C+YEye59I7DPcWWavGNrdrJUk8Rvn40EvKr/xDU1E
RxTVaVyAh6rl59lc8I1WYsDghhkvvXTIEF9N+B6kwOeQJ+vsfzYUdSr/hMjJyfeBnR1QrooyqsXC
CRnEgUHQBtjdbuMXLDNwhzbe6i4QlKioNJCCQkd9Aih+eE7nHsXM2bGdgg9Ab+65zlHE9wXgBTIi
vl26JeroHy70uPo7ieT1KHDyvMsm+/Aj1W7ixygzU6yS3H+DZlL80LBxExWwanXUdmgZDlckqMS0
mF8srOVAxI5QHYVq3WTQGcrANMCIVMVIT+Y5QkMQw7RaKVwrEd6+8kQL/zU6MUkLEMkoYOFgD9RY
uFVs05E9fesMCnnDDG59mdWlOzxYKkgueAdaC8umP+fnLg3/+J3GSeRROkuV0WlDCM3D2A87pMhR
HIll/vQVzC2mBq2cXmhfxDrKqDiYfzcqcEeZMqo+epYVX7g6l0h7AJmC68b4V7DEmxW7hiHILwoh
CJEMfaOZDkIgG/kgejbp38qzjhDBVcTN89EcAuFkiRUnj+7/w+ry+JcDcmxV2+h5mWurVV/8MmMx
ot3ys0s7FSHNGZlxU4cdiuV1iYvd6zk5wyrIoUst6x+TDopmsx1j7g1Glvon40vuqNAXB89v0Zye
QUEpLNQxY/mcuhiWkPabLZl1iyC9R+LFcUvHBjrpMQkJo0O6UxDFSpzmqiqAiuKPrhcG9U+7Dp97
nXNUY7KU3gpVNn94SY0y7Fs6z9oFzYq77bJMngEWYLPhmv9zinbwZweZltrxTlmp3HDEEd9h12qJ
j5Ra7vLBDMrrPfWrnljsZ4gcyEliWdJm9uK9d1y9uyOfsxznE71jcSaC61kg5OVbpEUJv6Anhx3q
csmxeWswvh/yAx0/x3ln+IiA5jfi0w59PDhRz/H7NCDvhKNWBcCVTyFE1SW+OajjPiwW4FL2DZjy
Ph1swN78lINv1qGSl6CAYhXSseXGlnxhRxAhaAgRr4L8WZBEUkkWo/LH4jm/NYlIfUMDtHgdqqK0
Dl33dwMzLtncQsRspD/B4o2TW0LeBcS5UVewvXwVqtMFUIlfbh5orV6oUgWlsFEt/2d2HuMxi6s7
zuCiuZyTvhud4dt9MsLhEyigJkcUaeAAhNRf02zWQIWuy9nuVqLrusa83VIPRdPIetlq7GhH4EbX
MBnTaFuUUsk42R6KxfgITS/uLh0CD6DNQpT262/VpHhGk7Om+N1TYIJJp37SqVElAOi65vj1G1hS
VFMGbmHZfG/LgIx83AN97ry5JhJeuJkeKj/CIqvWvGt91OlOeq+4qHlPvI+HJdePM6KdKgFywXe+
iX1G+iLycX7r+PdKfww9cp43lxSRomjvVQBfeyg8of2NAsNh5Atq8myNx2YeUFgqtJixHXyn4VLA
ZcmJ7et3f+Db/lGOZwO6vSJVRvETifqaVNwb9aQgf6nW/5Fo6ThGnqjhzWRGCHO03Omw0gnaCzuL
FttPzGqPQ17KBW92WjM893jN6WbLtvoK+GYtxI0sAffzG+aslsVFg2vm4ISu7NhnuPb7aHWI292d
8hAxUJ/0czNHXhqRjHwgTGxAWw7czD+zVUEMP1BMusQWlMHXWCy9C3dUYduMDUMx38OxF7e1qPzK
CPBRiJiXcKbGgMukNQITx0JDykha6Tickfs/rItSi9SwFTPSYjXQ9B55TAE2GyU2spaMkrVMF6+s
ZiI0A2P/UKsVjqcG4tgEQDbhMMeFLcFuhv975rPaylG5jgNoJdKn5wQtD+0Xsx7yHJr4V1aKv+tF
7jcZe7iAm6vGms2JeyGZ+JP2RaZ5Mokd2jr5KB/flHIhZGv2cW5uVSPVodF7p5uL9oJ4ynhFgOxr
Nu2AmzZoV+bDAvGMMQNqqHubULoNATpkX4RzdUHTzlCf/2v9DLhynaITz1ANjQVATytSUttB46XU
nyPPsnsvn0OJwiufPXfq+2WGGRsZeematan4vJgujE6COJLjngGFo45BqUL6YP7UfyN+Qq1RdJSV
yytO8HObI91DhCFxdudUawRL0MG85B6LWFtKH1tOWl5sr2dECHE73Bbq7aO3wWqKpyBY2SNTFrlP
dAtvigEaxzfsWiuMRjabZGdIEs6M0/0HBk4HVZzOTZ/9l5/WTgybCu6ZB3BIrpK0y9qQhc6Ikw06
V+mVe3CssnGMGkNZf16Fsk3/si3QAsdgxysBqPm5rQOiMTWwXaH5xYuK42q0GD/4VBPCxgpOrah6
gYZGiM5PumyD8ACKi9eXmTYMIR/4S0gosLk1FWYGcwzxV6nClFpTKFq6ng77GmpxndgpLvDEMOF3
ZLhBsdKgFGl6Jcbkh4l0AQHLYMsaTa1OZFQ2vnC7lOTA68+ySPpJOXycEZik6WEnRZ7N20nsu4he
XBhaU/0HqegBeQdKotSr6hVlSioi5KYhPO67fEz+zSC0MfTak9sak0t/aJciSQf/DunGRc0xOHQt
nzLBBA8UAzbvSBqZoAscs5GNWJ07ELV9Mi9j5I27vdDygp+TLjvzhZEDf/3BZoxZKDeg1P8CP3dZ
k9cn8hRHQpih6H3PQufCrYuEQ1PAGxWBncl2khmKuQi/9NdZd+rTdi9gv6ML6u1bxW6nnzwf0WA9
XAe6py2kLBXUnREFU/w9/uboLCbzp87NEnodTqN05o4f4QUXgtzckrzJ+oy7MmvH6ndq1c/h2tDe
y8K5H/D4H74MbvTCspB71jdwxEw4D9CrUPAy1FRHbdVUeR8JQSmB0ZBT2X5TLOr8nk9JAfkUWeUD
VWl+DiLuO7P0Ahq0jahD5PiIXFsY8Q1T853PNAWsZAou8z7ETrmKOv3Y50ZpGlfVtEq3HotWa2kW
hDpdbG2aIBMWvRIFgTsIX09jayWoYcOOWeRoB6YgH2XQt4k70ZGI/LDOjGHV9FH04vuSQz1JY9O/
3AieWJ8R92uBu003p/66cwjaFM3+lfY5tlwU+k4b6i1xbbfInVZoASrLjzDaPxUpybTwv45S/WQD
cZF1DRBwc52VBxvoZb/c80EigfvEXjwwmgPd9OvTAQomCxRuP4jov11wi9Gn3edLVvv8qCtQMQZE
mdiVx6YNdUBHpTD2wvrBK6BsW2pjPeQ9ocDvPImwJ0YJwYgNeUrUEsnqoJb8JDvm8HNErgoYNQmd
XIKL9tWt17uh59CXXEnbHTly1rjLmDrp5YlVAqojaasXJz9vEqCupaVcvkq8Ub4K/2l0u9TFhLfE
DcLAatcEVKnV9MpfVdDEosPxQ5JSxint2ZzAxCBWc9eMVFKzdDPIYLwHHwdOwp5/CtrFwreZk4q+
1Qlb/DmsI9MedNKfDHAJc+5r//ltTqy8kFrvmVGLaHY7M/SxdeYXBdLLXUjjHaZusBT4KGnyXiZV
IMzrwAKiZ+go+pfILw3Le3lvPtfhu5MQ188GDr1h854M4ZCL2Qvo4mibpbQ2HhF5JrAsO62y/oXV
gCQc9nQwIDkimFIzlduRGgW9lT03kfvJXHO48KfoI1BcPiJabAghQKadhNlrVwHU6SWYt4U9b/7n
DLTxSuMgEw9Jv42ufcZY/oxEzNWZXtieGppR5HbFReP/k+AKsRIdCjo0a/rXQ4s9ugwrCCChERzv
Xw+sJHCn5FG5pjDMAc4ZR9A2qva7pTtGl0FjzOHZsviuRq6BEa+3RwuLCQ+itgAm/tDOlhNxdGVq
9yN/6EplwRH86+XGkB5bQ1aevsWaQRj6x1KPcZH3IbAFqzypKFOLAIDWN8jZgGI0Iz7pgCrnVp1V
ON1VXwdHigvPpj5Y2KxCC80v0Jj4QQNIsZuR9KhI4tr4fMDbytCHea6306JwuX7+My2aS4ppq/yF
2OGnAxKytoAQk23F7Ve6WbP7Tutf+MtNIm7BWAbOWKZ6X7tKXVhCd3nP2BYgrQr6s0xtQInG+gUQ
Qa0R8lZ4BvNXsZsceg0NFwcFhDv411ZKR65t5GCh3FNMCSc5uf1TcxfGAfAB8Xdg5ULVxkVrS0iV
4zbiSGDsEFPH+EzdgzjPp5vNHUyewMUpUk2wLuocmsEBg7/ZbnZKSAcY1wNaDxc9IcUaKh9McQT5
dqk8w0Qcn/MW+TFUX6G0UxshfGmUzvIX5SXjV4LDbj/+sXrGFBMS9HxTHnW8C1wc/Q6BzjYjLErP
Uu1qVct3S2A761bf/+EebyebXX+ROoUYNKsac6obYUBKPPJKAjtuq5h1OD2vthQ8wIs4l0tndyXQ
6pXQsKKPFd4lXl2V47XOmIub04tZMl6LqX4U0PQJJYJT+S7bqCaZmJsxM0AN7rfnaYOwLvN0f6uH
oWGc8lsXASw/8H0TTnb3tZyMOLoU5ug3yscl3+KAXcfVzbV6YqKZ/96E345AVYySljvaOF7NP4pQ
JSub8tXgrhUOuXyHOgqnOoD7mKOupLuWso0LcqOzkxws1OoW+YKavPi1OR6vEf6BHcmBufz2WKPA
8tDY2t3wTXn62bJkTJo70sebF3q+vHU3MMCoIoclGQPaNwSu7wnrejYB+iiNcGcJ+Wl6xoAQXdRE
mc2HmvjYrXQ0LmqB94gcLGMyDlahqfje7g881yRtw/YHliTTU2czuHh4CaKU/f6W8nlc6zcoEVii
nKOlG4uxfmd9vFgtSDeyV1Gy6tETjUz2q6jnhWs7knMIrDe1tzPUX3rQyc0q0WIdTi8rnNF1zTY7
JHaZA3h9aTxgxZtGf7KbY6uw3tgvSEK9Vs3weXYW7tuT9v4BqtUgPGlbLcM7QqRgA/dkJ6wJhcnb
bX5vjn/LmRmPfZsy9Z8+zliEw1Cx1GwR4x67C8AFVtVK9V+URk6oTW2QupQLmUoB2BxoDvWOYTCJ
EMtGh5iOHUmHFVN1YVlcc5ejgytAQZ+xkpV9I4cv9hoJAZpx7h1saeZgWVI8gqkhSF8ccO7SInz7
43c/Ze4A12fCoZKgyqS5aFP3UMw0DlIJZLJU/KGVssFpkUU1bRHga3Wn9pkUpRrkmWnjfYAehh5p
wSzCzayf9k56zSeF1IE67YKGqMm8hsEVgGWuE9zPwlTPMT72LP6Yj8+08CH7MVaJDuhq25ZG1WOD
iVpQRm56GW80N7Ds0xNtYBbTSF6AYGLHYoy/uVEeBrym2+IryJsUhSEvPXV3sR23dn0UMf5fe/AB
qrxDB57CNBWaaSvGWRMF46jfSJT29J0CF5lYSrdp0LGiRA9pHnTkhnUt6RG5grj70iy++NnjWDC5
A2UPBNIwmXWnWYM6memp9qF6epGUxS/BcgPZLn5iNdWG4CnnAt3Rtpyzm/9DOarm1o5cZ3/2P0RT
sYJMuW/hFTs83D0IrVa9fRDN8lGs699EsTsezPeAdtkQSM89gCVp5BDfANdNEK3YK5HRGYp3G17d
BA4fkFMdVNFLWPETlJ4/JcmrnyueOTIOGoWF33gwWBskt0Nbsg+G46PCksx4xJjWo4HWywYcUkoR
rCS53x2eMgOsr5WM2fy1QPdUFMuokbiFom6Whv1FQFeF3RCjHPsdNYcVca6ZTihh2LdA37SaGjhZ
t0DxJPKDk6VaX0hom+VmXvv8nCBxpvGf5ugiQ7qNZ6X2Lo1Hhsdl1vd8H+42qpooXytp9n5T0y0+
09/hkV0T55ceVSQBonSKgsSStJ/k5oRA2WwdUEI4m8tW3AIsahY2HItcrSsWc8fQi2KRQrpstrnX
zrZtHw5cHydVNwo4zOAE8Dym2KuugrHq4RO5WLzBFdFzrM78Wc4VYDQqIVwBDnrWl4quFq5SWcwL
zGY0jB+2xQtorFXNTeqpLsIZaEExj7mjwClv/lR/liivx8ZxqKp9+ylDX2aSgENqfhqoh4Fm7csU
AvVbAiXDRmnR8bIp98o/bWKejsMKF9A6dzv48TttHSZrhlVOlWpwITEJtFD4keJKJWti64RbVCrr
GVOAE26f+BbrI8+vtUJyaL8r8XcmOvNdZuQAVJbZjV9VGN76v/cvyMQmdqmHy45YKK0Lr1ZnPWNE
vwEMsMVMfZ3vNzaKWOqqF41UQ7hNqjSWC0tLxqeUgwnhcDsB/sgy+BLwPeRvp/zHp+RRkXywaEMM
GrH8h1BN9u3PXzQTHMNOOQ5b761VcLMk+6lu6AAc/80mgwuakepsGnAkczYJ/UWRvezIx9U0bSqU
bmyP5NYATr9vR18sshelFfyf+vjFgCdVxT2cea8rMYqxhVmoWvlucQFmiThFk1/84/5ifJz3gpkR
zp7OMEZ8KgjOs8zsBaNDFOjjDNQyoAquv8KLXFC8ggBYud9oWpAh6GAIvJGtJmgLo3gitGkvJNVC
koF9ODT6wSyrM80LCQ/I+ayQn57m5v1wABpU2wkeVlniFUPGMIkmoGPygan4Rb4sT8uxqNOfcuIY
zcMXNfbuatnTeEjeziUfABd+18g+TDxxBEmeaq9XlCi0/5t63CpJ5fjuXqmEvKP44utjDntC6HFX
Zn932z8sSE/0vLX3bcYrIDvxnurrTxmsAb5HIFoZ2HdXExnsFXmw45oDpQG5GgN+EXlx0sM1FjBF
hmyFbofUz3ky7C8k11HZCsH5uPJK+AtJDTssybLw9Uw26LKhVnwr5808oT80Iz+u9tKXt20dznSC
kFSce+AhjjBcCxhZUlu36w8NJrS0gZLPXBlkjDnmM0rn+WtKBGRyJff3ACNCH0XIZNoXsqsh9Y7T
tBgVxUQbaugn543Tl+uduaOXLoblmqGUEP6IWy/U7Hanzlxa5D8kH/CyICBJW2ZU4AuxkPFYuZJp
IusjAB0hZPAM67Dt92Z+k0rxRqnjziiSV2iQ69K+4qBv4Pbl4GJizGhmmABD//1oYE0uxywiULx2
Mi8uI3Ij5W1Z5gLIC9RstP6YdSuzy8lLYhSFzDcd/W4HSVzhGUA/egtyXj1g+vPDAZL6XSTA57et
wtw5EMSpFJOIfmDY2zrxUvzlAxt0D4fVKYXqMPp+9vle+9Oi9oa3DE16oMqXvtQTrCKaTqHQ9FXu
pIYXyUwLCOnNLR+vpP4QDYZuJrA1OGncsDHODmmRXpRSV+qzk9Qb1zt2BZ5dtGCemZ3oOs8y5NYc
o3cFHpxhoOHJFR4gtxkhn6DPYlr6bWgWhIzfFu+2kbFkwlfLmcRCquQUkj3yVg/MFBRpU4g+bg14
CsIbYfVz86iGqCvRgkk2Gypjc5+Azl65NjfQZB3g1msalKoaxfe4EEVRTsRcHdQOOKUpuNm64KF1
FPa4vvhcdzLbh+/4CR4tDN8rS/pNE3Clyt8OyudPXgMv3JQrfy47v3m0utUGDjS5As4eLs1PCGhq
U9az+X47uxlIj1lux7Rhz39eWdRQ18WF0T0JQAkjxiett+5Zv/T0ZgFhQkzbC0JK2k3vqK9Cllt9
coMlM1W3E7//LrwMiZ6EyvPhm6vr8lxNArQ1YEkml7OnYMk9ZK9/XfhzzSkznxXyViU+O+5hb/2s
zr/v0vusqeuD+nCdk0VVYrrd1t1Oy9kLkfjwaLk3CaFUYdftdW5+9kQqoV96J4dNF+j2Hn4EBokl
BcwM/z7N8QUG7E1eUGE1/geaMuEfXN7hNtw7JvRY5FJUpnDED7GPqCmthceDDWiG1zHjkMXnNnE8
uDTitWN6rz0kfc+yFNITXDwk2D/HHzdSfHu7V6mrXr+sCjkv8dSYuaGQ5dZ4bapfGMuIn//Nl5Wi
peOCgnLvyD5mCTWoI0TpkgGGHpNndoq3d96WAeDMMhJht/YnU+8FDbvlfWqC2FssCpTjX4dZUiQw
vLzaeLeNCnLM4HVu/QyzKIQpc6nnT57l9FNShVyMHTy/vo4ncWOrMSfEhqf8dlt/N3VUKwnuS0IR
Bx+G+dzFZ5UtU2uyvZjNcReByqdQjjfJ0JNmDX2Hi4tZznr8BownmW2ENTJsyJLv6IMJrH2QnYFB
DDGDSioA/I2vzNN9vSOE3QzUW0NXFVkblp4vv4lpXsF6jLIh7gyfg4lIO7ps3SKpyxgqP/GnhuzS
7HejPham9/bBqki9i4xtpnB04UdpIsh9lpsGPa39Tx8K9dHjKF+5ICNnUjLmJy+d8isHM1IG8N+u
qWi+lNJi1I1L71yfzqvNF3EF2Q1w32QGuToDGjQLcSyVOSOGSQqYkk4hW9vRi9YFnwFzYYV/FYLr
6TRrvFloA0TFGjkjMfUIrx/8+++Pm4oXjaq4jslgRNt7M6hVwzbqWVfBIzQynBraO4XAppvNoUo7
4nEI0BeAR0b07IyRUJuYQWPwyQ6dU9gtgPWvJ0gCzEgzdnT96fWNhCsMEH3ZgrPKEEwTRs5jl46Q
zWsJHvCnu1koQHYH2Ft1uff81TAOj7fLrxI7B6Mvx/ZxpWmv7KOdeyMDUfVP+iwQJ9VfjFz22nzm
lPy1Bkgt2l2Urp1h6VPfu8N5QGD5C6+2eLUCfc/HwIC5PK0lTuKNyBD7KUkW4qBaPWaGEaIESbch
BCFmqWYrX7XIqCXqvXRv4JPP52+U1kh0IIoEFbwxyZnxYwBvf6e6jKdePHs0uIL4zyA+9zqod3Kl
9CK4FQ3cjzD3AfmHo9zSKoqvneqw1BXh3+jMXMRm9rNz2WfTGeA8ZhvUjDE3y0jSeBz8FjOUyy6R
Gb1AmhIPQcDJG/yyO1skEyvKlNrXB9gVRlrEneT9GpQKsNi7N8KQZZF7vj5FOluRh+YsPMgRTiFW
DzXcjb6dmG/af31POh7/MbgRNFRYGyHfrMb0Uq/mrcw+rMGrMJiUlqOP4NdTNtw9HhNSrO4pA8V3
OAlvd3ae2Ie4rtsGM5FPhsG59X4BOJJfd6i8hLjLlGnXdkDTzWVPRUMXHdxpOs8QjdUWv3H48gb3
F0E+tKiruQQyGuhE8TLuIggSLJUAXSoXObxYvkliMt24BGvIyZDWYCJQho8nHO39uNcN699cOccg
BehbPPuw+Yvnaf/jUAjrTgYiguv3gmptUSusrn8xS2jt6A6aFvU9KqT4XZVPWTnud4oB0EBWiLGq
qHYfJx1SMnOXlM5RXrOUHmeQu6oNIjZfjpw5JV31fr8tzRaYni93NQ/XV2MCXkAe1gG/aTCraxb2
SXFYTqceJ6kxyXa6SU06nVS2K75lDwcQM0KPbDbEou1hibhYkw/8V9rbjSMw0CLvfFUoQ+hM/S5D
25TrO45/157+uk6+aX6I2qxT6VdJ9cCtEg8jt2dJfgHKEXFRPAi2aHGX4XTVPXnGhQqkivwT+LpQ
0cuG4AHs5TiIfSHLYJHC5Aqp5BcpvgQmiupBb1V7sh4KeiAWExpuHculdVG3WfjgKGQkE6iiT8KG
SQNilCf0UFMJADdtYskApHT8UV+Az7UqP1m/I270REFwwP4gHgwVGzlD6oO3JjJxYXEGOsUS67QU
WsWxbKQqOMOvDsNKBm2+fgLIny4F8gV65IAvmyrG9fcXjAMP7a2sqqQMU0F6Q9MeoQRnQWBa/wh2
qDCUoDnXf9fdwxnhJ8PGwWdaTXLXALwKFxfTK0K1gUfQApFq1J+0HlgIwGIvgsgQ0LNHsvpqaOLr
p1P4EPV3kV2maGnZq+DM2gExX4zXT/m2DCbYMzdq0RC1Dn9rWrWBKh//LQIDpGiWKEl47hzhmB07
zDoC7U1qT4pMaQM577l+gafMyVCeoZHO0Pqpa1Hw0WXbM5/NExUpNbIHn/hIs0MHcz00wuU9C/uK
0SdQtgkWNZtSF7pZ61Pyt8vhFLevSu6N57NZSyKuDY7LcZbsZ6vExFawvuvWaIDHZkJ3pBFJBcEW
J/+4SDpR78bcvvOEUt+elN2GLEFZRduqFab/SV/9mVTc2h15R9PuA1AEoCSKDS17+VDGHdnpph/F
yNlGI7SwTlBLucaRW2cj3ALx/S7Z8nhVPWHBrUJRyExQ1RYVwGtpemxR/XyrFJapDFvhh6nCNyf8
VLffiKtpQINGX1sTQkf8Jv4basW+SI3LSSee3LlwUXR9WR24tRS8FgbKA9U7sjJ8kzdgchfr/cAW
3GHJmjBczaeXhQIbxl8m6DpAvR4L6xhsvx4lzxe6dQukSu8cyON720TkTdjpXVUhln7v0XworxiG
0Gls5GbD7Yo7qQ9PbyD8K6QkG5TRaauyI+3/k98QKEDHXhYL6b7RCnvSle0c/GTi7c3IY0Bxk+hO
9WNGlgmnLyqBqnQDPt0AaQptoRAdVSOnvkqdqvrVspyhqdLIsqbZxdic8emBMM7b15zTQUro+lCL
VaYXJYaXEJMrWV0QG3WFetnR4Nrb9JHNO9wI/xfAnNsmXra/D7sz/aGggv2Lh1wxg7CykKK5inzF
mgSj60yhAnnqQUud9OIgfr/AtCOIXOYOvbzSq6UagEqo19+5cQbLsvOQE6E/owXosFZOrqNy/faa
G5jPgLpBoMbmXKs+V1GqSCaApUYfYhsxJPNrKUZeoKXkE2ElT+Ed/l2+vlxQSiPaaW05XIXhqF4Z
DsqarT3n3yP+qLQQjxwCVlkZzpaQtMnrGG4hMoBuo6wnaQFIfEJjorJpLx+8Z9K/RpYnaA6ZhZLG
OFzlOwgGTndNN1WEubDLFS2FN7GkFyTjpYi0tnONuSW4XhQxxbApcMzL4uQr/D75+hjLLuHLCFUE
XqTG8qZ1yOAdUQtKVbvO3bajA+f04p/rKN4xTuCw6tqoPNm6hMqW2Ilb428AdwJChgWi9D3rfsqz
uCd2plqXcGvGC8Pzhps6zGubLDgcvr/40PMXXvLbSCvCe6vgCnKBw4UR2mds1wztCQQnFfbufiSB
cfoCd7lJhn4alm3VcnE3eiR2sh8hL9pCa8Nz82ply2mZEThwq8354BhjUUDNpuGmJtg7ttry4ObQ
1mTNmw76FdFYlWAvhvr1mgCi5Wzn+fAaP5epS0Vv9r12YOk2MLbsrXu2xdPGHEw94fMfltXet+HI
hipJTE2Aigeia1aIiyBfGBvVJ4cfA2OwxKLfG+/4QPPhmKuOpQF4sW6XDrBBH3V5dDQ6IoDZZ7iv
/oIoueM0fQX2NoMvStVntk0LtLfe6JDA1Gk1a3jkprHOsKFGDA9o4QM3fw/fiz64+oBYFzjtloy8
52SLy0ksr0aYJU1BYpCMcXbwSnbcwDvo2onK0StO6z2ZrZ8AQm3kixerPOq8uN5yqv9OpCuSubgn
A1AsqdpPXgubKc9/zRNYzqH7vPChuXwvhHJaW/4/OZ2hOe4nWQRMIJlGJkI6NiSrVk1wLrhkFYbb
gpqRfOit7/BA5oE1EiTYKDTzE24aldLOjihUPjTc1tCef/fhNil6HFM/wNnu2XRcQ2ga3UtvrzAG
1J5ReZV+1e4EUzC2fIFwk1CxpXY/evka/g4TZ/h69TQHBrHR4FfRESdlCq7/qpwtPbkS0stnPlbp
z8CvcfeqByW77+59fvtd9p4av0ax1zZJvhi15PHPxsZnkUfWe4YxG19Rkvjomugrl8e0G7XXLI4t
GVoWm5YW90hlrSerzByirKRYHWnp3n3nxLHOXE0HDz/UBBWQM8BBBSX3kcpBKtoSLp6RUMekJSlJ
4mHrsba2uxzknEbgzfPsqwE15BcGx+GD6ypY4a87vDlsUa+eIkbK9QG3PBqQU07QTCgI7BiCdbi1
SeWw4W73ktzApl9+CzAGIIQypndYwk7Q1GNjH20qnlzmZAPNXYXa9/YAzDfL8z9LQw8+lEKnTZXM
m/Zx4zcseDm0gMQHm05+dgoCS9k8ketT7DZE6wq4+0XRdzDHTlsCeRC/SQiJSHu7Tl6OAoK7tzlX
NoHS0YwhT7HUKvnSmfHWEU/71Gvb7fGYx1sMRIYOfhQjba97i3RPAQ4WT6DwaojSeNoEaY3U7cyX
l7iyaeYayrHa76opY4QogNAYHq9qAAx5fU710OzBHl0ZRAjQZFSZk5ggCOzijjFZ/r4jmTEDKH9u
HRLqfrbEYj+J4bxq3XUJ0xlK3P2HDNiMksAuolvraBbeUiCB6yKQrsmTxFBmJxXY5E3zbq3mzfUz
L6rkWgK8FISYgFxVaJhBJBWLylcjXuCzv0r49CQyGFuJbEahQCgHzdi/iv3tLuBeL7plOJfwLTHo
XruzITxDjL2CKoWmCSY3lerV3JIT8LRlHufAzRuQQzhgKTf3BnfNrPezs3NXlojevo/U9iFYhYM8
ZF76Mqcaf55eErczgu5HbXUGfXh4m4qiJdvwPRHdQ5ZzgLG1lJHtMiA/21eZeWl7GhuJjyLyu2VA
kUSPoCA39gVLRESAVQx79MLRN0ZACaiHassXNpslXPWjKCfRFpRHRMHS1/8mZ9+sULQ/0xqbaDkK
QsVTrnUc8aRjrZEcGMg9ARi/pwZ3VOxSRfPXwJjstqs/BkBQ/cM5HE56aIXd4YesfHgYDcNosgV+
MoyadgW57MpSaGcZbWK4GRioTzOxBj+ueiDnPMwVE5lrRLk3HdLLnsLz4I2RppGNSckax1SuaPMl
E7dYH78NQgUBv19uJsJQySzC5WhpKheZFZhlovi2mmEGXMVR+le3wBd6EOTQjy1/KGlmwC/UQxkm
E0kQjlnk6hi0TByzesXeHD6PRzJi7eF/MyuofF5cDR5YujV84yaDGlphYJMd69Wg8HvhzFJYzHV/
8VcZiSaJDQMSb4MXtFKgG3eJQPMjljAisSdE3gWb3SaMXk9JhtAkqhXo9plKmdMHe3oLWrWcxqKL
2f0tCI82CU0ZN21RMnCUmiXs9Nboc9PNmTfHFjrr0zZ5+0k+J6mXklZAni96Zot892pHT1UIFh1T
fexRYXYrb49c3L9HGBA0r9JEWbHbi6EK6IiIjVyo2kCMzIRCX5uVvgIzT/OqpA+lqCVM4AJ7ngHW
q5iInzkWIOMsCXBAIuDVdG5uzsXzzdTJ4qh0hAemfzkkYa6B2cdIl43gdhAcqApY89zZhLG5/aWj
qGem3b860KhQXcwPeXyHXt18pYnVVg7auhSB0tiLKlVLfS05B0Qn+sJAkMviUCu3HLgunjtANgTB
YVSN0X7P8NvrFSMXRAcUCz5kOaDaL/bACH0KcRIPvpz/mTzzLFLSgf9o81eCy+nVB9H1Sq88JNQa
5RfqcuZUuwzAgC4mIEc5Rb1f9VH92+Ox1Xqzrc5W/eVpfYi3Bef4xw1ASDSs+34vcoOD/y1bYXCx
xR7OfaliyM+HZdGveiJ2pTezD0R3k6/WXDrUIJ96BIZpb9mEqD97gQSAcQ9T3Dhvn6JfxublIIx7
qFDSg32I3RU9RtojKQFPI1O27RYzJ6z0r+rkDOgu+sLA1k0ZMEoc4m/R5KeUKik+9ky5Vk8azMZE
RGC1iQxasRzaf4jive0MGBNqmnecvg9kjlwcUZkWud6oLYGt56EaUrrC0PeUkQEcGRdfJ2Y7Tiga
f5v5hBOyhyx7kVvARqrCn0mWevBXFSjQFhZXj29yqEWjMf9fqrnNodtxKybf01PwkdTj5ciopH9a
61NLgz33K59C3T7Iv6Aa4oWny2H6f0GiFdGOBKLIM30pt7kDZnI6D3EwfnG9P20Y4ujRyJWVPITq
/A+bzs/qlc84fWqIqU252Aab++kBgtWjGIA/PTsdCE+xJZAQeICuTx1JmpY3urlsQfthBVG/robi
fAZKEmBrTa+U+h3aJfGrKk5UjJYdNiW2MGSIQJI9+uvz3K+969QYTjud9y6w+/1t/SF5+Z3c92/G
PqkDSqQNgBpfWfBCIBrPko+lSq4vHvvjIhLf7xjYXufLxbT9doYVAulgaraPu1Mj9t9mbXiuw5gK
+scPJadmNzwb9G8prUpPpblTKdqiHajQoqGSRtav4RixXbIvVXFfv7i3vw20MsTZxHS99SlioC/s
uknLkJox5Wosri54eyhcvU/BJDYqtyx3aP7L64I/+nCm23JqY+GvIUtejI8PL5Iz2O6AbJnYjR2D
ge2/b5QmFWMWeH7JQr8C3uEMr9M8ML1vR1hihBkqv5Lgj4Lb127vBuJBZRHhilDHBjaGsoyxaHDK
9dsGEXQakQXgEihYGTqgZtYO88vy0Pghwn5YKQWi8QrxLLlZG9/+AmS7TcpvJK05Ak0IG6/ecKtq
jO0+IntFqpmej6MQsRMzVvIIIqvdcRaHNGuIoluL/DXu7kECQrABGWb4GOJTay1Z1usRAN9MhHiZ
AyxH7xk9FaBXczvFXOBsend8BtvFHMn8GwdI02MJzC8ouKtm+TIc7ReZNSLS6bwzSVb2kHTYdeRw
ECeTzr6yk4hLuw6gffIcGSARP6urTTDp9b+DF1HDWZL4HMmGAqNUOoFjGBZHJldN0YpYwWYncp3V
ktxaMH1/OOoS/NoSG4uel6D7VrUmqMi/Tcn3WHRJneiRkRnOpY+wlyDRsR1lJnKy13zKcBUJN7be
hBKEYJ3zgMs+7r0+8HK69tDBmgMjIsWE6CVPALBp3LjWyY45pFUsY/c11Dom8XCOm5bfbVMA9Frc
6ghLjE0VNhWm77qgSFR3ddoNTwRKFJ/omx7aOkYbWPOxqUeydRikKNKTGLCu0nurAY0b9TB+sbpj
tZS+HxqJiM57NUJp3XPBF820CqgvyK0MTpgb49LsAwT/zBuZNTCBJYDJM0u8ZbEMflgL2nAj1br3
fcvDFHWZq1pQ1mL6a4QxhbsnSkZf2Y6r3IZqBJeGDwp+/Ra/D1lOnYM13tVKX3uqIYGQs70tuOwX
uRFBisgOBwAZoUkwl7wzL39HXxEvX5iZk30K54sw68nAFHk9nEnun3Qh7cuahlROxP9n7kfUyFcf
M9IhXnfy8j/ES5SkUxoe9dZNR4yAe5XW1Ga11EAAGbZ6oXtJs4AxbOHWhG4eGfxwP1Gut3z4Owvv
f8vkLO4sQNsbv7rwmsndQ57ITZLz8ThGMrACeCh9CWdFlWLoClEsJLIK5O84QUpQNxDpEwSquFfi
NS+Y1VR7t7iwYyGt+gdQrx8lVEMh7i5adqE6GDgnsmZWIz3FLX+VZyy3RGa6NXPvzYOunZdjMNd6
gAVthK+d7AiHWLuLYATrNCk8u6vHc/0JIqIUi2eYQ5d8hc2TfOgM1NArUTIpQa9U/3LaWISpa3oN
T40bxGbK+nygp5LtgcPwyN1rc9o52d9qkxb20Y4ZgcdZ44CbSDBiLYJ8GA+if47iQopOdyQiqGW4
0JPSFPPJ+MPcUFgisaOLxhA9DMec5wE3a9q6XVckPOvpGJiafvP1VxdfncrgSrHScb9Biwb0Cfy7
IR1RtSoA9a4Y4X10arbOzQlkhDS2KB8q8BFL43iwyx6SoLxX47IR70RtdGZllY1WF0i95M2LcEco
wUB5t3uX5rTLjFjzsbQ9sLgoF/7uuFHqDR5XE9ZUOaUDg4JuLDNkEw2wJpSIcDXondfkjl6+VJk4
yyVTp7LrBSTky6bfQd1oPlXpnaJGhBLzE/8eYHykQBUjQrw4Dmo53sf05gxGADJghleRrEInZzPV
G4IQsPtyht3t2OSOnznm82PN3hW6J/7NYT3D4QuO9KS0xV0HKxyaOJ6KLY9Sn9DCQPlL0nRiPC/6
oQSd2maq4XPepjiYVHa2LBuG4EOAvIhDd7mWWmDV/dP4SF5PHFiocbnQwAIAp/3Pq26Ab9bzyCAL
oXKh7JmhO5ypKcFmhou+7s6cq9SZ3YRyRIT9qUTek6rNNLkYm1IxmfEYgDZBykUW5eOR9kM4ASBJ
8FbWFxyAza4n2FmLCevxAtfCpEcBTXoYC6v4b9UXY1VD8v4rQFxQXBef2QKMGNzE0Jb5e2UtGCtC
CLYaYss2s13nhUrzuSfJA9YbIm6UbDe6aYpVUWOcgUPpi1Hn7rAscqJ7ycId0UjUqHvb5ctsXWJo
tK9aYn5NF8tK9FHdANXuQ3cOSNvcR1cZR6Ovn0hzUJGHnNfVc+1yxU+MeQP3FumjYSaPkkCHvcYz
E2Ezlt6upSd/6erxNMHlIOspyA4du3HGXryrtfaFFcaErjhaGgkmh0GOvW1ffhcOv/alcpi8bqdA
57/b7l4kZa4Nf/Vuugei+g9iC0r0C4R0N7lb1Lqs4gn4F1rJwE8jNsoUHProY2bhwraDFBr5HEKT
pvUbv5eEscsC1iI8zmDPenjE8gIYs8G5lOsEL+N4ev73GNcGKeNlNaQ0oLpUOOJxsz0Ud9hPlcNR
ZeVyYCuuk0YyRt6fPR5+M48X2Nq3uiz8OOiN920VbGro9J+j+ZC4iY+1ukVkDCPmvvPtv/Qho3n9
x1WDftsfHj/KrfYh3d+wP84qjaJyXje8ynuOh47n0Sm2qWya2QE0HmKJROCX3sn6Po0Womg6BH0e
ZKln++bXUPC/U49phtN1kMnA5qAu0dhXLIIX++uy2ISdJT72JPQV3CKKaoPXZK/rAHhmsm4JxKU9
lAt7NqvOWO9hWdK4oGz6FRIQZtocX+GFfMhQ2WgYSEMFY3Fe8VuGgMKV44npVOPEH5ID7DJ8M9l9
l9GFvJ0gnabpyRckew6T+YjihYAb5YYMxgAJiNRud/2NA7C8zseNTCN1fwTWfbgmloz4x7TLvYbO
i9vVRBCa0fEk9Z7nIgPoRZC0a/Dn2lP7BB+GC2w/UKujqYUsyLkz1FOT4OLQTKSsIwjrdlCE4beX
UDNbT2WAnU43UNWcWhLKGyOESKgXgn5XZpDcsmzLQV8Q/MZHQVZ3qsm3nDvGP5k/RpIqUmhUaDc2
BN3pDHOfpLDvsUpLU5OpIGfKYtizQkai4P7FsQE9beuYj4rFa2hTXR5odqMQYUmMUQYjhVz/16Qi
xSA4QoWzmKRswz3nNkZzGhQ+r1h6GRCYUaLjvxRzqpFaTueyPik2PiewHyXrRMM0rNvKiQouvN5b
L8L/LhDDR1zXdOqEjnH5zXZ85RSHnvnibOLJK1s3d/54RL0GwoCFIozVLGjPEFKZ5SMwoi4V11XU
UYsSrszlTGnUvBzAUBTp4k8QCWrtZGGp4AIA5eblGTvxMr8bDY8wiMt6Qp/AGQ3Bgq6A29GKcZrp
j2JpWs12DMTDpzL+vJdcEnbcn1iPfCIYpWrRPk3PVT34XwaF8iotSz47azLjplA5azFed9pVtsif
zmWJpJj5FFi0P2ljaS1xXiuUmuHJ+6wIahd1YX6r1Bi0vAqgV48ewzpLo6p5EFc2oc+xKmXcyeLn
5XPw9BMN2ulclnTZ4YektovZxhK8ifLdPWLyqwjBCupL8k91n2W4nWJ8N11iVZpoC7DWLiD3Via9
aP10alZiT10hUxnJYnt/Qr0td7W79STkMrZr96VjG2pTwlZdyHA9UPHKbIb3nbJJrOW76nCewREj
v4TqCrXqvnnTSxIdB6utP4X+/OPvK4OEDLUjQh+guYRDKZy/gJI3Wrc5Njhbwx0gtsHqoOKo7r6o
IIkpLvplpR1hQ/e/GJQpvrpf+4CNWfQhEzUBDOyv1JBRKi2HGMIeRgTByTDFX5XTnt0yoKp/9K4o
4GaAVmpYAYPLXOeBPyvO+w5CXtErWebwJBfz3e7oRkTXCqbqbLLVs7hy7/RurFnapWsp7zY7dpjD
y9mkC64J/p6K8Bgq12t+bydau0Y+ZCWicegzeuhEjOloxJ4Zfb+B9utTwP55bjOfS+MI/NcjfQPh
MvruWa0RUMk3el8tdv62r76h3hT9W5GeWlQi55fNatlVagkPyD6daCpfRGlNmKL9vwcvZpvgfEzp
pLuPXwZv+6rSogr5icDbnd6bnflgx35ZJnbcNpV1BYOolJImGdjIJbmx3IV4CEpk8/0HWnhhaYaE
5tavwb3rOt1lA/VcyuwyrP5b9K0qPpsgVHScoDflkHbqBecS6M7oNqNzuKuJMRRDOdLJE1nKUKml
DjOGjGJdLIITg/P+/t74VVPXQLbRKZuEIRD90y/Eoa0D7z11V6HYweupOhMInpAU2igeg54Cbkma
/+BoEjeBSMR/End6m1Fh/fj7dqTqYnxBKghIKxywLHUZ9LI2JW5m4/GY9E63cu/SweSDah73lCUW
VR+JafPP2lvGfbGkukjGEW1xpLSil8QWIXaMxzewSvXHIoPOTJRGIU3hDW4daraH0f1RXThBYmag
KjDlO2MzWszcFgoP+8kViAKqB8rQKQIsvPeC3sWTk5ykCGe3KWdGnRtTJ8WVIMnItf10t7jVcX9y
D30NPP21Pgeqc9NzDpErreWjUwTYcYWUfenez0R+IIoR/zpPAGWEePhb/Nxq5T0cDLyEqaQIf73W
OYYlXemN9s/cjZZP6jr0ChOsiVLoyUA1M5nn3yGApJBXOm/f0XqVHQgXzl9gR0fohk/fHlNNPl1K
M7fgC5vcTpTFsxwMi84gEz1+IlrRQdTAspQojxU3Nqk3P1ef9CDybllb6TvViUZdAY6ApuawV/II
Y+W+JUPH82l494BZsbbulCsAZIDHtWQHNVgcHplHHEcZ0K8GOojZ/0HzybwZTHLdnhmwfnHlVtfz
LaImYQs46XEbYYjRHvjaKHiIMpbE28yJtWSJRFVz7oOg3BM2DDdqnL9J8YM2U9yFSGs35khueDXn
HZm8WYWFMSJ83kMibu1orz2UGrh7mc0apqhJ+Mh8MDsEA++FVKp9QXl5UW9+3RLCidDbe8sASBT+
YI9s7vAFuccZY3mS0TQ97q2uDgUnmLSNg9FH4lY4ngr8Jmuoic/K90PDxmy3Lxg7K7SkZyVHmErv
byGLm2g50z+eTIAeGI5C3T0GDIjpnieUHLl5pt4ZGDyW1sgm66s22ixUSdB7y1ySrG13eewsTzdY
Gb643QbV5JfPR1EV6GETpdZBw7sB9vj5KJxQkNXkk3o82C+V7oStlxh8RN7jwFe+RUCMJGeDwxRG
QlZhdsHtgeQ0yOPV8XmuizIa5ZDdf3UoafA+rO1fRKFbdE4LknwzNiUqO04YAZJRnDxmOfylwR0S
WzzvFJ/9FZALQWOBWqIkIfTx+qD2PLjbB3/Ufy9nlkTh2DkJTXC06diXBYlcYuQjzLSJjXH0Bppd
iC79eoDAMQN2Xlw2NQ6diXR1mpr91l8wE5YnrckDRGhzkyDPquSsFwCpgpTsHkdgpR2Z2j2dqHJc
53YS8dNOH7HidTZC5wCJatv0u/GVZDqmzw3vH+99JUrBCSR8+/6ngU90Y/NTUtmH7fTr1/eLmYyT
lb2QyP1HQDBuE8exIPJ//z+USsq1AtjiQNx0hmz8aAkHHw2MNjdMz7jF5KoA0d7TGxKCknnzMrZ6
fIlMwsFwX1dDeyKKBlJP4UWG2p7Qm0znhEG1hgY6AjDAhmWtYYb/PayJQsOFYRQfKj3/iSnYHefI
7sBXiYoEjS56wZpceMWjwGtYDU2xELo+lkUXXprmiPHYWAeD4HcfWnEbQZqcePMHvwZgPBEaw1/B
uAI8/qX26V0/PlEtH+tMdBHE2ZFiomS1aW+CYgd9094nhkd0ko3a1yIbljN/OG2LSPERLwB5AGT8
8XXH02jjGKHWa1IzOAHLBVKQpN16XtOXgzS6+JOg6wtUlioXsxarUZFOh2D+X2/vQe0nU2x+nh54
EGJtCYNMVXMPqOx1Pq8q7Z02zQ1+feXTNkbZytGGj+PEslVVcwDdre4G2L1ni+gTguB/ZWDg8bMP
sNQtwNE+lH6DAYWgWJeOWocJC+3orZlhJg7Ukc/BeoKFSHsc8VEn0kff473jOtCniA8FZevV79wO
BDzsjKE6EI9WA7bKhMDNGJ7De5hppxkpRZe4vK8RdHOK+/8A2TUaIZ/FwUtCpDS3h3TFbHfktURk
EcTUBpCbaAk1BWNIBrbLQytoL1XO+XedC1si4jCOT/9DVG+i1c+v8Cw+tL5HP2MKHQlMKWnQ8d9a
Q4fvZlDhHYt20QySX+LDWSYa2ldln5qtaUXCZOZuCjBPMQRtnFAWtT8aW0XxX9leLeSBL2f1JWGD
ND5ETnzN7xD+u8I5wqHGygh4dS3qemKTYvqJCcyPoeu4fn6TRuMDvXfVICn3oVVuug2VnGen4OvX
SuARRMVdQh0qfjqwsWGMdHybqCPXb6uv81sIOae1bfL8DFzYHIYVewvia2VuLsxRqnjUk3ChGGAB
XbEg8ws66nkkwm8qkzcwPdnbA4xl5A3vkjUXnWDz6w2FyH9QrP0VeFKZ/oALFjxa1Ql4DEHCj3jF
siHgcTWL9hFLnLzEf+gASTHWP0fMqmOiNt/IILIA5rFEtLf5VUyz3mDSeVYsUM6bUH6gqQfCVuxs
G0mjdqYI1br9QahVf47fGl7YzGEOT5E33xJAgndrjVjdKBOS/5vjf5UBxtZTb0sGwJWN8ujovrP8
jJI4XPt1otQW5y3RnSiCw6NL8L+azRk0Bwgxi5s2oQpfwFwhcJh2zS0fC8L+3Z2xWridBUKyYAdW
4MXCfq2ACPx+/THAQJI1foteV0SlB1H31f1so6YtfrW15BrxngwAbBF6FfB8Kil2JBEElT5MxIQf
cNCkPf8dE26/wccFZBSYuefkwcHb8SgcqgCRS+dh6fGL159eertZ7XzrR5cSQkXUoPwfI6v6nL/a
YHjd6rSw+rzxvb9wQg3EN5ZIShMSpFCBAgBEXj98E/hYQCQyrPQCQNP07gakK9fe4vIkrMgKU1aU
3FGyj3LOdXkhGcnrCeEp0+MC/jHtc/e0TYHl8Iab9Nk5VO/6Ryq9RNO3K/vN4NHsRULa6pexNRJs
+a7ljWl3OvKmDILlBk28FKKObTqqoqeUKTIv0hTQkUOBXcM1jYMfXwb2V+nbq1/OHlTa66jI8lRI
dnRJp50O4fhyvjHU2M2X3tapsBz2wAGXslplGVYfsQsZbuU+ketVHMy5otjq6oSGxU4Ib7ZE8AjD
xzoWbjWZS6N96sCMrjztV52DBTvKENxwR270KD2R6G/dmrPkKXRF7mKbTzfDWK1Oq0o3in3x0z61
A992uqd5EuSS2mSWniQB49r0uHRwNWhz0KEbUWNmxxeNOv6kKDD0coSF8Lm2nJ/5Yvv/8VFSz6qK
JENDBuUR/veEauKcYs+NKPEWn2fyFPBFEU1zRBWNGw2/37/MNwKWCGUR+WV9JZhbWLFABUVOLjvE
tiN81WrbH0bW6+04UJAHDUM2YNJKA3AhkvE1Ak6ywQ4wZSrLcO7tFqD5eQBgxbOiZcNysRAGvHV0
IzyJE5ms393gVLtMP3LP89xC5zSknX570y+8Zd0f4JJGHSVsj18RFPc7lxiigFQD32TImaEVVLjZ
TMGZT1mzH4nCn8IikUYdRF3b9r60ohjFoazPvHmoVPpA3QuzuBaUhOWp/DLkBJHWCMt2H0oObElr
qbe1qZHsnSG0HnWE+MxCoSAj1phgpt1N/LXGCO0rM/TWhpoCipBDrPkgZhIGgcfE3ALmwSaKN7MM
TiDaqZJ3bq49YcQIJLm/9ZxbMIG2I4eBqKegDkYa6Puz/3XHYPwp078SXDG8QQwbsbzOmMKmfu8T
ceKf8Bpbvvd9a5bn08qEaf7popXju4slkwFma/VUO5m3N93cUdZQmYVRTLZ+HbyjEsp/oaV6L4vW
vHxkjfNz6W7sSJI2Y8qrhD3gNmqQRizwSmfZjQ/swiWtc2GAuw99cdUZ8BRsAL7U3lK+X49scLXL
o6Npf/6zwFOic+4kWNgBGhAUafPPkbO5k5sCc00Qma6lh0UNQX5MRnMKbGaBDSBn7u1Wt8OHlY2/
A3kvAW9I1S6z1xXo/StzMUHkqg5ITIhAbTHfRjhWEuyPUY1Q7ATGGhAo8vTUozxrMhkFsdaQww4S
Ek6vE8jxOXPj8dvXR/YkdAAIDC2+1uO3++VfugFWYwYsa9gPkcA/X2rPfK49KsBQ3KDvXQtZzAkW
UX/4fou7F2aJy7tAtT1HcAAsbORiThDkz+W8cDJYiGZVNGKYNdUnMFI+LWENiDTYbrElooo32i2z
uRhAgSbhQBWLteB8uAQl5eM45Z8JHrty5kkirsKJ+PMbsRkgBnwTd6EIDTMxEzEL644OMsTs73ps
bB9943Lo0aAbXeZEPCDT0UZm4fHE4kmrh7fMM5zDOjfBVtAuQ0QbpN771CguVc0fBoaoUKQi7bdZ
qyNWDqtxXcnnjoAUBpal/yG1vd6/1nOZIaz6tzk6mNDTsCmfXVR/D0sJlwuj//1Mnj4OVD2g5sSr
RJGQiJXSy96RT70f6toIQxBBPFBaWRnD/gmAhpUreC38mc8w0cFNU9H0jFTfokrmA7mLyzVzPk+p
aM073+1NPU6LrZ2RLaz6X1a+rBuAmW38K8uHsVpUIj8ayPSX6wDKsS2s/VmhBFuaCUpscWwqr+bj
sCVYvCLc2/awIgtktU2oXXXoUTNCidlJivH2COd9ZRlCmcmONiTUUio6DGK4KIhUpWo++d0Ky2eS
P7Vzwss6NxRF/9Y2zKJSRL1hgYFMRpM9Bczdp9FTA8VpNb9XUfkEClSFNZn2Rp5PxPKKKvffZsnU
HhbGmg5O2lJQfCeOLYrjxrZiUhq6JsoQ4zfukYvUiCu4cOUj9sYtNtwV0rRqvN/n2IMz6knv+g+O
Iwnr3yzYwHeN2jzXJOBRwiS7jHxNqfefk1nUqsuiX+66Cd/+IcwkxcCzZS4ep9VDgFyNXQu1G0BE
qRcwCjuxfgAhDMNWSh/Sqi3kkmbJy2rNQg7YimfhDzVyhjyqvdg7wo0Ow/CXLhYV0LFV7tgWPSlt
fQ6YlmBkqwXvRkhYNT2CU6+kzBzB0XzPqFJHResoSHf1KPqguymUi9qeimbhQtOVXJrPH3s6Vrs6
DzHuSqnM4QakPfh6GYgQMfvnR0QnzkGl1uhIkLa/jm7fdLs5Ll0mWlvPnBFF2dMyjDW5wDStyUNQ
/DQ8/nXZvVf/VbgLyKHW7vpwLIbrNoc5sSAy+gWuH+R5ek5fl85oKqIlfswZV8nbn8vyzbZaYHag
Abwg2gOcn/0l60LgJH5Eav2gPECq5xMC1num67iC5XS6SkrtlZDTtnUtK34A0jGbJGu5Do3Kjd4C
kI8dXGDS65Qb+GIdTY29ecp5xX1/Zcb9l7HqdKF2eT4R0Nii7JcIL/IfisbZsUR/b8hM+cAtPHmq
DsM7JhFTH6hUFb3QrjDOROHBREUZ0Jk9xXlLxN5CV57NBiNANp6fOBwpRX2/9pvSgcIPZ0eEdjXG
XRVOUXFQl9Ch+vEnDo1VOMOZm/XwFNNXsIIOln00JPdNVwewl7uXduVNwIPb7+wPTXnL+Ie6LzcV
f9SPyuPSomSJqhoj0Rzm9amTGV5L5YhBHa0Z5/twn4bsvuyL6KbxoXtgkoV5WwduuM8f1DuU217/
NFNzZGM+MGWP6n+vuq6Aas57EGca5cDl/5ehpN7PZGK+gfvwPMdm4n8+hmIkymDwht/AJvtgH+Vf
y5Ou4I+RsvjKsCr4l0fvBvHqI79vuK/jeIFFCt4aKICjcnxDsf+NRAJ1QlYhjc6mnWHLeR1bAdLy
e9ZdM/RGryslxlg54nC8jumVMeoBoNoTwZaJFZsi4pJLUY7SA2aGSsm5xIb84QW0hQAnJeNXYSSV
zy6PVigoT9rxDg8FNwffoFlyDmJ/FAtyyJa3lwteLu3kH7XzFoWBbw8jJsl6Bxig7WgVj9or4mFI
h7lyt96iNe/WI9KoFGp/i0OWHdpqPhkAeNdxeDPDzjU/3HEPjkoIARkntMOZVbNTDPCQFMY8cbNi
3i/lpTWZL191K8hMXsR6Sbktemnuj8d/6XHf7109PN5M2LwFOl43QbVpqz1zuSLsVnju7ZcTdEEQ
KDgYHorwbBgk3SXeo6jeBEAEKehKwGlo3neJNVoHiiXHYXGqcNqVHxUrX65i5I/KWcK7y9o4NHrH
MJVR5HWmOcWOUuhnMa9fqpq5oelHesdu+J08ywVNGYZ1oklL47rRW6YB+IkhyraZgTUgOF+3vQ0N
h2ZlfDScMVOPzXoKQvYz53B7/h1MPpb7mAq02V92Up0QEVa5toIpQLu7tlwVP+PHfkEF4n4QOTIP
hlOyo9bBQ0ec2+c7ANMIHlslNV8Sx5IECGzDN5xkSpwm8xvM2qV6DaRin7tvUv+vv+u0kSwAS8lX
F3GxiYS8GjBipZaCYBKmeAh1caBKx3CfvJMmulu+DQBfgAxycGQyHvERZU7o7BJ57Pnmqjwn1vV2
+1Vc/89a7MaB80JV7hm0Zn9iOnpPgDCNAPX3S0QulJKvP2QLDm4OManBTE/59E00iLMDehRIwGEz
CWXRG10hahNkYjqtaK+QNzh+a6TiRmzHqptSS6kajdedVIQS7a5MCfW6K5kJzu0Kx7Ez2PxrAMYM
2ginZiolaQ7/5lLDGkDA4wVZGfEVRFmtEvZEfxpDbfWboU8xUOKMSIxjqakXrD4suLAp90afRNyk
ee4KvhsggpzRZrW7hec27fnot5eL2tT/TYKtLMpOyzTR4STUbUzBnYtXBd7SYcOKGI7cJqQCgVwm
32P2dBdTbSiVLPL1cJDOAbAW12ljWvUnzvP8DnSiq9huFQQRDQW8IRMChXEcL+EpXg4XkeJ8w7SA
zqo3Ai6aOCxkjn6xKbzwOU/LLdzFAU1dwfDv0dqGMT5rV9LVzEfdWVWy3FoxRtOqxHypTRKCXyCi
pCS6A4g9b3oOW2V4h0rGutjJFMx0qS9c8grS8O2IsVt0BpmpzX4NDje4ct+iI6y+JyNYj6IFoy4Y
jyb70nnmD4pFrYNwpwkNZFn3Q+c3w+UHTkbwlPtNC/BEt7xv55acYdPpsy+t0uWTXJwgKs9pH+D9
oD4tIg3aOtHfX5hACw/eA/0P/02PX1dWPMCIXtCkOcnVXFaFaHbz1ilg3b2Gi+CsByLgOB0H13Qz
mJDFfGJMnZyYoCF/JySP24o09xzF1RHc35l81u3KFH6rOUc7yAcYoj162ooojxCPZCGOUPq2F6l2
YsS8C4ae9hiBZRoHJn++xNI1BPPWX8/D3dXj9G34xLYu4DxVrMFWWuG5pWLEMus9lDj9XS6XKueO
1a58xK4ais77D6f84dYWoiNM0OveT4n0Vl/1L8cHIaOVr4UaN3VTkhdAkQeuGThp+rkDTWVQBX7i
Xw7YdH+T5VnlPA3n0tU8yDEJe+cL3cw0Gl029fqU8ZwCqtuwphB5iX9WReJanE3Jk1ZW1DNYkmWi
EzqfkQ6NMMKZuXe0TEDswwoZRjJqmEpdWrt6WhxlLnpKvJLB8aStPX5rOCviEOKdO7YudTEfrnfj
7/EslhMrpcKil7hc7JF2vbqpztvVY+DCVcrFmb2HHRbsAsCtjE7voKO3kcKd+yFCB7rM0k0NDU/e
d+RxyV55XG42MiBGgjen3nMMJrIlrDgpEPeRx7wav6ru+0HFZUzFrPbkvkc8PgM+Ak/W+O05TfTm
oNO/VGgYjt6wt8N6u3eaRrjWnEdh+Vfo7JqdEDInTmV7a1aBImm/eWvWX3rjEYKd1FaVSCTflqSy
Da6X2UzJ7ZS1Qdg76864Zw4XIxRq2/LJg69/TuA7+R4l5J5vAF9EnYIwNVLWxrMTvl4ez9WjkyMi
ANHq38E/sUf5CZfiF7TEK/2xCvlAarCIUJYnKRSOk66UqeRPtxue+KwTwgLoy4A5sZTKvaCUsq+H
nfNdhS2l8+JVzrr7zVvkJWbNe+YHgUGAzgCO3PSD0x6G58lF6sjxXEgtFrlGlBqr/zw5Sb2VBTC/
ZTIqiqZHT8F72AxrmEqvaROqYMtOsMv7PTjupdRPT3wGS3bm89SOD1zoQA+Yl8R83K/0822LBxYT
Nd8zduy8iodxGU0uDVZwiKrfDRK35ay7+2cXPC38MntMhisQbuu438Wb3vDgufgBNwXyPOWRTg2J
EGJuYaOQ9KYl+oZGYt2kO5PbZSSLqunHCE8cSDUjUJyGmgUG0Hx5wrk/Vx56ii2ZTn6F7yrI8z0f
Gb6XS4l8JkLJ3Muw8VsSZpxvK+xF8FfZWWCRTFW/L0Yn2lXx6XfQmnDGUmnLZZmjsVc6jTJ2jnA8
fzpzi9pBB7Gxns+/Yig1xARn7N7C2qxtcH5VJHwr7GwWZW2bD9DXs/fs0CRbKthF09e/qGKapTeN
1FTnI4CGtf8sAHgdOonemBlpJ8hvJf7k0HqT/FjLd4RQozjNcO7kom7/jCe/guGlji0ml1CAUTO9
nfcUycPaSpOZi0tmZetO43KbWVQKrVOE/g5U57l6BcB5nLwFxmpPZkM2K9W+ApiYObCjh7dj9CRC
H9apZivh/XOQ0E7CzeN+GoFsWPr5DlaYQr4K45mdKPZUXx8ifjpyuiFjw77HWcoYTti+0wkU1yq7
bbanit4jSx+Q8sdiEVbk7RrLpRWr+G4kW/GhdUUQh7mbqiHz2qc45yzJwAyfjSQ+41U45KLCaHZA
fTfbCKExq+DKzR7MIMnpFrdx/KMhufm+AdP1k4YbdfouIpIuazJ0SRCg48uSJMCzppAr4CGJGf4S
E2ckHjliXZRsPObBWAbmCfWgSeXnx5tZ6uWmdhcxoVCetAGx0LCSYtXCyX4DypvNheNgZG9e3Gh5
MaXDdyHyiOxu4ZbcXjgN7IN0LS3T9M2t7M1DfbZJLBWIVX7fEJoRrqBOKKEjYKbcXavw49+AyFG3
6d+PAKIHcMqdJhc7/ihYhc8CsCEYxNgWl8hPovrkvDIFFcqPZJaSYUtGIwi3uQQvBftLeZ0uKP5J
iyWQ6H/kw80/YHUEuHOROXEa9BMPRjSTPgnpDJGjRdRpyukhUfdfjP9aXPNzw6F7WbMXIIDAzbW1
4c6o9mXFoNCWkW2y1+88Ysg4tpIeiQq2lAJpZ5K1yqzjtnuVV9OuZt1SGtDw9ImqetSN2K9cMYF7
CIRm1E+nWkRyDbH1y5uhe/AcQy6XYzKWxmkaue+5RCD5hzoevhwAKurlIxEWQ5QZ3PVZnjXuV6cA
KfbBpKNWwjPbAFt4sxiNlTrGP2zLOHxRCodT9T/eMwZbWe3qCHj2f7ruilJl8E/kKpX55uFIS7rG
QHsl05rJxGjvEURym6Fvi385mcoejj3JOfAb87aQLuHFbrgWSl+YHamER51Q5D9gmD+0f2VDHhSg
ycJG+rhOZJW3cFM0YSh51pAr6g6e832XsXOBEtlPJnolfMjsAki0dYMnMHLIJWe62j5KkhSrNI5t
uiZ+SqVRUvuMnDPl9gqznbAuszHrSAC5s/x9/tc3TGV2VqGwb/u+klXvQNn4t3DHkHzSbif9o1D9
zn80VbR/jsVKTj5xhuiP0+ClQsIsU9wugxGzrIzG4aEs2FTxVhUk5ng1HC4p0QPVLJRKqv3ju4Ht
wsOnirQzBwKdsgXA6xdu+2+xOY9eQb5DO9l9/Ktedwh2OhYsDQYqIT/WTWQqeAD7xvXOk5rQ3TTu
ugl3G2wikFpxvZeyVuNAXF0yvGnR3Ti/zrtQ78ywpGZS9ugc2RsmB9A/ZLzb4yc/WPOSckExLfmG
rpNq5rOviKTpFYnyheeqLJLQmPv34zzpXcC6PPC+fmwBfF5Jlm82jG6F34VRXL9sZj0e+aofojBd
eSMO3Qv2lxMBQmsnRgLsH4NUjq3sVYrdJeolQShN40CShp0xovOWzuYwHvXTpvuVbNwSaF0WfJ83
pSwPJZv4YahGl/oM5VuWxR4Qj7Q1O1+nlEjUk2oPbLzbarw9TDegpWtIaDdGxCp62mjFmfx7vu/b
1Q4vRjyfKWWUVGKcjnIgDIXqpfMwVDkg4ZO+AswieuyqPZgQW4UMslKGbacIGcfxYD2LIIOM0kEu
m0Q7t+DGZN7mdh1l0f/QiAF+mVxlCK8efQCXJUgCyzfFabL2wtNrWJFrubjpaSolS7XHPkZD37/M
euCVQqspwow9YihTgT+On8Pwqqg1FTiJhD+BLslHqtqdLcbIX2o7spWX7BvUtaBy3oiWDcEVloFo
37Upx4iS8UwqqB1BKej+Uaz1HUpBGwdlOypFPxydmHBY2rXFwy4aC+ayYLDJYTGsHneL0C3SMtid
BvSQ7+aoIqWKxWZFjmh+bWo1e7slMLciJa1A8VFHs0OR80aGhsRoT40yZjie7+NNm+DH7jJuwIg9
XUqT9IKf9w4DYryiioKZVjWYDIfvA7pzLddH/ppGjCP0rfibBdrAZWBj6YH6GkW0mGh6I7xQu125
N234Tct/6zLzVeT1RUzpj7f+X1NaIoE1F+2Wr32L9AXP7Xw6A36xiVB4uexTPY+Mv0fDXi4XFO/H
tlkHJm/ULh6/VvwQH43ABVncTs9SNHcLFViebuiM+vgarM4zJLsuPQw3PWNd4/eXwe00Mw1blJME
lTEmlqFTk2ivSbjhwHtCXwvVwIh30gjB3OPKQCHiv/Os2N0Rp+FwO95VJEiqrnYhD9bbC5p+anwT
LjEmb9n6VC7rGlyWYrPmqUGkcrdNCxF2Tjsb5vqGSh2Mxua0ypk3UpEUpv9Pl78ZHFslAMq/oQeR
zgbtu6iAQlfl8lL4t9JPDsNdFZQJ0G6F8ctnx+0mrKq4RM+kAg+RB81nFQ3X+f1K6N4D6GzC49Cl
dThP5Y5ZlOKxSNoTzx5CW0goCBHhJnMzIW3gp8YhJ+Qh7E2CbZ2kWIAgdMJ4o7DOm7d0e1oRZSLe
1eIh8Gz1JnT0dCU1sA8kQ+inZ/B82a4GDYjwhLg4jZnb0syJPbZlitLuaAdulSPHzrAwiGasbJsM
alBl4Mn0StxcMwkIZ63DlkZx2SpgSmSSqkJfzkmpw3LPON9y4G7C6rPe3ojBv5MCRbwuAynDT1WV
bHTa1niC8yoVH8EQ+OiZjTRuEVJQqqbmT00LgMTklmBCOppMWpQF16nKb0BFRHrklYEIVH3IaGUe
6rMAUusNMvM6OCU8df9DspoKsV7MCHoSpefBHNZkO3hXk4Fw4o3m2rjmB06wLpOmIkHFuGdcKU6Y
xcGYD7eKDUJ8ey7peOsMjTM65THj57M7ndz5Pi2PJ9jLJST6Wdkyc5IgHO2C0l+I+xS5+XlgDJqy
JIr2LvRP/FckZoE8oGncL+hOjVlzX2GuHs8JW4HQW80L6Ovw4cfbt3TtkafjNxvfPytl7QKiiLYG
Fu0NaKuR8NY5iOBSFackWw3jU+d+3AIf/D67zaGGmf9aqDmnCo59DFEeT2q9P+W3bqyHmYf8PUG1
GKJ+hJ9tzss0edKhAQImrB5gE56Yy/qESmEYk4TvDuDYSkzt/kTiT+unt4kLuNWrB2T3OOXvHQqX
GxO2d3yzkyk3zQSjAk2BY1wR0Oy7QJwhHrtzp0s1795QnavZd9fnC26kbsp2G4VyjtQ+MErjyMZX
Z3A+mpms2Ch932i6efkLwkk30FlS1jjbNIuJRTHgr9lAziMvNo2lPf4Q3wGNHf+wONC0E6/XSdvT
loiIkP/vZs0Iuhk0rA6f6DoSVSvjbkr85SuhCbhc5mhFbHlu997AoIQcGnhdbW4daQhAuQju71Ll
BEwCpjVszlZpCEMCehp11TE0r1Oeo0RG1QrhlOWq/EqlNka4OEIeHvT6HGh07XR/jWWSeKBcPbbb
gAUe3D3dpLrUHKE03bWcUj3PLJ+U/7WwOdusHnKvqFWbSEyG0c40JhKipxmY/Qf8Io0WvSCwgsh1
i/UMqd1Snq/IBfZD6iiJHbriIGTyNyFz9lKzq0BOPGsd7KmtaRnwl8jldLnEAHh5WR473Ggbs/If
o08Tgg9rn99RgCVVLpjS6hYFFPm6EwnwlbfobtZORcjy2UyzOG+LGA2RHvwDxYsWe8Ey/sRvCpsb
jJjGsdM7koZwG2pkh4vGIHIX8wm+6n8zBPJoUHHRNCekde1orHGQPgUFUEhZiawZCTfacB8eIw3A
h/j9MRvTGnBEZV2c19M2agxoaHuVPR8I/tcF0z9O0k+WxVHKdEYmLxljtUeTS+l2DKXl3BOMUgmL
P8LXP7+hnhqtWGCSMtUWKYOVU/ebvm6GF3s6MvGQ8smoJiFlYEBWzfW+P9Bvy9TA0ZJ0Miy5uR6F
VirLfGrorYBgmwlj/8CG0NaXpvQU75CpSRNKbHSTYBvVtI+ZnCASh7bFJAFRVqwq+B1xV9YZCvGa
OAOlltZxbDE2ZteQ4TjlyCz8xWfOlEgS2eOIOwwwjUNqpvpxzvMPPnE/RzHh+QcuE5n/kv2T2QQQ
17nUulkhSnBOO49XJw3VlWRssCf11mwOj+2/AF8zMfqwCo6Cf2EQpRnJ8rD7Lk3lRjibEtSZpEn0
VuY6ESSV8Gx7Oa6FAC0mR4X7gFkyiC6YSpYzfWK9ApqavNgXUfgRlWdDnf4wSXKY3OMyO0KproJl
SLSHb7Gpjtc0xar5wJI0U66TI1nY1A0/5MDxL5BKa5jt1tfVyOHTokvV1CEaXJCjM0hIik0FsDre
9mBO0uGQ+3q+UI1MxRYgftFXvZEbygNWO/k1dnm/0JaPypkvDuqi2mc7YB8Agat9Hwj0SYTTmpk9
Qbb9uNlD3Y4lsVaaV7E6YqlIWaMIy7HOCAlWQrsYnZlzbnV9TiarFpxwLCLKbbu5ixThWs6deqsE
DkJDzF+k7Z3gUdzcyWX49OWt01+0qEPvCYt4UqLtwrZrcxDPap/xCtOvl2OdDXdL3EEThwdFHr6v
xmZA4JiY4p/tqVDGVNRgXlw5T014OkMD0tA4PBvhKqLhuMZMIKKmo8BmYdOg+/G+DmNUP0WezyN5
vYCodCMJ7f5cmF4NtmYPAAIvQr4ime2lAh+jfMr9dXLao80KRvIC3CMQu+JfKp5bAG1tJ7NgF3W6
CFtMz0iCvWuoIdjd0jMeuG29msinvlWM4NzjZL8hks9LmHDGvQZXDxpD4MIFmbMHPPfwc1T29r4G
ToANETjrXs0QhgAlMvTOOEYNAsE+93E0A8T/q4LkhToj75SLoLmwTW8JF7LGWHRqegTz4tV0XC4Y
X8KojPup8bkEUfsrzWmFU9rIGWQ8q7UYzdyTX00qqNp83Ja/WmjcImYWvNBOn1z+cQM3rd3xAhCf
1ArJFCacouZdLEHa/ibwWvZVW1HIinz/To6pywfEnOGQcJetFo05/GKJeZw96JGOgXIo21mBfW3c
2AgNafoKrNBQ2fgqde1RdYKhxNWGsE8tULEU2MrEVfjMvB+zJswH3GnO+sZ1hMiYg7tQY/sD3PqV
rDleunImZ6YgepCPR0I5IGzAviuPGammC9+wt61V4UIcy97k9uG92+ZCGc72c+D44/N2TOWJFHoj
T+pam5/lTAh6ODyZeOC52OgF9SbH4A25PHQ6r2fqSUrMzKFZzE8cmNAyi4XEoDAg56qUrvwvGQHo
QBZopWWGzra3tgYq/mkA69rG6L95drhAYGw/fX6EzQRK6+i7t1tN+9QIwgJGHYY9cJYQRuI44lty
tFtKoIrwKEq/xjmsVJ+/Sf/zT6m5p4/6OaMfWqJ5PnlFzyeNNrXoM516hvcNFg8Nxx8gbvyeDK9H
s43y4YJWL3qBPx2wkLcDLeatwKOO+EmxIs+tW4R7XOLF51fgbJKoyhcYHQR8CLPc0G2pOJu7rRou
zj0WTTq9aW3MSNkh3Aaw2CiyfY5IYugqb8pvClRwHyTH7UEdjhGtazChKeGFR+Kxn8e0wBHy9Vy8
u6sVZ9Ke39Oui/2c1OkMXBMWscOwGbMsGgZrQUwG2iTB45c4GfWOWjOx9qT3f3485l4XZ/oQ32ha
dFNah5f5deqTgplXe15AcaVl1XtI0eIbGtvDW9yfSIb1ktrNVYFTHMsgV7igpMhRnGQzHJrzDJZo
5T2WCzmC9e6iwzV74TMZQYR2EhoXYYEjrm29acCLlcU3Db3WH1oBXlYov/ZNMuqdjTzxDjkbHT7a
aK4EYFc+lbyy+5HLVT//CQ2fdAXs65Yp8sKM+RaPmW20d/nfCJJi+++qD7PJ8+nvC8uv+yjdC6mk
9uUNCQUKDWvk1d1p9TJ4pNIxpdGA9aKIjkEW4ieeD7NBLm93Xj6Hd6WeAbsuMtI7qgSYG7EC/S50
bEdPme0f9Y7L6k/IxdxBjFijSTN0RWbNibVgpx28tHKDFPGIUJw9ZQxlyzWsh7SuHlwTmiIKZn9p
g0kv/Ui1w+s9AbiIIlRWPv9MdS/uZNDCaLk1mnD6UxK0UaJxdUjYc18vF8pVSoWboNAGOnkxcbAr
9UBTyaSCqvNY8gcM9owcwcjej/4Bfh2rE70DnLt7aT2RrkuowWLTtGzcZpAq5aw2Gbqg+mmi+Nyw
PlmwDublPUyH99M9NJ/m0wpsW+9al4vHHo+GvOsi1HKv1aoFSboKLepwOgsv3NCnMxjsdNPe/oIC
wful9Tl2gm36zT3H6MYoXeJSopeuUR410WLnVLsWs/lsH6ISAd8pBPQfvjmPPB07AFBK5RP7frw6
2O1onm6bvKyBGqFw53U1T30dGeMi9ia56SPnINzyta0MsKD3nIiMJrFHpMeA2KkNsfbDDBl1wDu9
czKlLbo//OcUa/E/xnj8sMmNPAiqIkzY0oW0INFOjVVjw2SYRL6Mh+yQajL+tnDyF4jBQDHlbV5n
Isfbo6kIrgvYjYlpWldZKRaqXp3exF7hZdqdDF3r12EM0iRJcGZKifjmPG/ndDcizB6WMXCFqHkH
1IZXSCcfB2lWyFu+xSYzOUtjTXgvID0R7bGyM9QMopQHXbl8rLuOfnLIXlDOYwV82BhCjEy2g95/
Bl/Nwv8ltvy1XB2E70aomWJ438j/l+8gEEZSO0x0QWvY26kGqc2wTzA1oDufzOjCQb1TYsen5wS2
tkfXrPxPqSU0o7UzefWKanYla5Blc31WOSYXs8gEo3Itf0maDEz9rQj8Bd71akj+rg6qsDSzvA4k
ExGdkfV7OVJ286B6bi1VPoIfzyeb7/JOUYSz0iY+0tW5ndHc5hTdoyfTKZUC+et5Uj9SKjEO8kBO
a2xsGY5QbGPTH2MprjZLsQNnVLtNB8qZ8S+fSM0k+64UTrsfyCxIGbvPzWxzrWd0R1XXLSFxWd8K
xSFODfUJpJjPQPcQiXkv8/BXCipeVazcIkHSplliSKZB1J3iFsfeE9YZwuvBafOBxHcaiJUfW3Vi
dTepR5SMjn2n9yX9Po2gMehFzVfIYLzX37hlpNAMZX8w+xTqO3ZqYIJWuVL6qA4HWY3m/dcLRWoC
gjItR8nsaVshLQRZPg+ylT5qFiEepFB5R5LT+HsLVgChvLKITyIClwjv0Bp9GUwhn6559Ie+7tgK
3JU3pyXBS3RPtNnzRE5Lqg0WMnJY/wUeh/Vb3OMm1dYlEAVjwuyJTf8UqUtn5fVV99yK4k70oIVP
qqwdF3lZzsazOLtxAh1H9x9/6UYqLoyIgqLl5C9JafjJucfNLkp0ORT/dVtHdfw0DJoRPeyrQMFQ
EGmf8JJ5WTH0oKSVU+GJVC7l/5G92eu0GDtqCvYep2/S1WCbcY15ufE/YwThBkDuzDKRDAxCeTnO
ndDa6jPqG/v2FR/vB9kgYfY8FElQD6v7ucF6VkILVU9sDPp4V3slGsyaCaYdC+Cb5Jljz2uAL5KB
zS57FgqjeHgPx8Qzr5xGKBz74qjwG++OwmJ3tXms380NzIapEOklbzhoEumHyGa+01MozKAtCagu
s9V3thDE4Q7ZAog+I1IHQPVBO5Y7u1UGfRyP+PzxM9haAUrQhi6lA6GOiSSgK8obGz2ziY3J5XZG
P1IN7D3bJBWF56Q1OkOtG+y8sxEQRZggUalFw9D6WzykmKY5sKpsRkxqoCmWdNCjbRDw+oJjYjrT
jUA55hfxvmI0pYw2eN6YLBVG37PicoygAx+1e0Q4Xks45wR4rMFEeY4iTvQI82WKLCvACfl1F6Cr
XHC/BeJt2YIFSuVyvoLT1U1jyvduQun+1ti7PTyep4mk3SDKGvcITzQlYOEvBtDg+4aapV8fukBz
xGSgrvkNWyILQ0kayA3lGa+ppyI9ZgwFiDZBN7bkVj8fcYAjf8gTjq2EiE2rMJ0tSv1Q44fPwpHF
gcbGaDn1azqH5LD50Q+bG+SoAXOirGxyhtRZZo3wXRco0aTi/aiS8NTxkE1Qd92dcPw/pZDKBiy2
NFuXlXADH6o5xE4JmhvC8+b1G0W6kZWvoys/vvTprBQrw+jM7l3Mo5EIXRggFImVlimDSLPlSMEN
P41n4S+9MCTSvk4d56Ch7fEizRtS/keGk3XizJIoGC0aDHT0YihZXmpcjzEMWPWBMUWHAJFJ0dmA
pb7CmCahPaajd2epI5W1z3+Q4acyRx+0QL510K/m+cVtPVSNlxERCT/BYKr9GBBkWAzkfr8tDOmO
A7NYWC6HL9h1CtLr359Yk9Fye76UNt3FPr9dUSihpLhgHUu17BQDDdFxhCCLsOfovSGHOjWONdtb
qMwrpnRK+9TN/jzBFUxLch1yZ8M5UoZ09MV3EoqhVC0QIF7R4eFdsgaSKOtLETuyaOugqpfIR32k
bZuWdqdw+j3gS9p9uMlSF4JR3M8kDG5REvrjlpDh/7G4xfc/yEWDgNtirmuXwSwkXMREo57HwXVt
bLEyl57CNsTYoxYSUmYOhgosohjH0JHj2lKqvGSki8iuSEn8gxtXKE/lfM3/LSxk5ECLoB7+Co8c
TlSIzXqKUFoYtWx/yLp/7qrNnq/pqEmKCcCP/uCdJJ6p4nayuDXh9s68Tiv6K7+C2MmWrc2jkF1r
Gof9PrfPrOU5UNrJ00nSZ+MR/oHktRw/ZzsgiMtatzOuusEY13F/V9cpPPY08iEly2qP9Zjrpc2c
bW7ja2c8xJfLs8DHC4bmUyiwfQWh0Fi4R47NXsjYhuiwbgT2ngu78LmFYHAntGHfkd9VC6G1vGox
K1Pte2aW/G2lT7HEaCQftZB8XYOlIfbLtEmLexExEBQm85Juet/RnUbNVNaXKr3NBWHiSCz4JVqu
cJ2UIYK3es0I6LgYu5RyrsSJ9sb44zvJQhVBQQcKUkKArIEdmrhi1srdLgyQaUVGcRc+mturTLgE
8tVz/8kA6W/kjz0HxnxP2OrW99addOBG0OGDbID9CYQwzmmizKKIznHPYOdekJFS2GZNXgvuzdom
Hhe5qA0vBKmij513NvwGPH0EW/NNwUPUMIVf8Dkliuo31c/RRDhMJRztM3OQQEG97qf/AUwoKMLD
WgskSV+zE3JjY1huzqEN94hNqxeFOEiwkJgppKXIbr8GMG07FTmnxC2PJ7iMI0p5Rjtg1UPG8m3Q
KrudKkbMDZVYokStMifIgCtD5kr6D6DEpM297fHgQs1JUoh7igl8mDiUf0OR4lIlV9L6d5O+IWas
j+pQiz9PYTDmEmSf4mH8CRQZN3L5ddwrNfU4fYM88HCRrsbDLIZlvmodEGEcb9sgtkhNVRU2j+wv
+kSq/FuOrXgPbHboJkBq7xsChPYml9udKA8RuUc2veoQcnmBjazF4Kl4lVtPzpWkMxHOMHLRySmi
XOnGQupPNcz7l81Tl42aDRJbLsf6rYEhrjnpnBh1bJnKGNuVCALcm8F25H1se+V7mpG47zhFHcTA
LQ8qmn3TcmqTB/rIezqA091Z3QNZ5hYQoC0V8xsvOop83JqF8e6xi8vvH/cbZhgUwZFyy/77H7gw
fAhKwC+uwBf5cshlyqHC2x6F1ou/Q/nKuX1cetJzwjjS519azfLzvCM1H3TxOqPY1lr98TFQiuq6
uRg8sxpNEG/om6yNUOKG7w79rgiVZfXpYeHfo2pieXgeBT1JZ+Vx5ZoW4OWYzy9sZ8l2iGja5kFC
fFJA4lQMTgD8WebmfFuBgY31pOqpUpj7J4t6w7ML3Vz1ZZR8YLvQX2HfIb44eoLOFh6+4e3cvIaN
13ad2/8ESKiNwUD74/aAUwLiSg/x/CbBrhdQV1cZ84hhUJJ+oSwTmsV6cl60fJUDOkbEe4N+DkrD
znYXg9L9Wq1mG8Bk/ZSk4cBIb2UHtUetC9PuTJgdAGwI+mDQz9HfAQfmB9m3RH44J9vp9/AAUrnc
YhnvNuRfToWBwNSwfyfo8codNrq2wyoblh4682ywFnA+Jkb3/WKpXQFwiHFRSc1UpsfobgRIuApv
bnpTshExb/4UxeI/J7ZNz5no3zhvDHVjBGI1JVsZK/CIVe5SsbipDu+d/QgC3C1a4712IoA9U39E
+DB1Q9N2YtEUjfVmC3EMrJypY1lMmoodyCw8535U5MfOJauHA1bUgeoAlbOBU7omuKIUwCNsDN7q
rEBzHxXfDs3ghl3PQMWsXzpzQWFmwxAN3q8k0hsT23SUPi3bWDoruceG0oc9WAHGrvrKAMyot0gy
RmJbGmiJHv9b913lM77yEJBdapESCO2bfv4o3n0jwJ6BF4Qs5TmMyKKJA8na9hav8kyRS4WoGk1z
5izCvZDE0kpEC5TXUjiPjMeGljFsW7ZQGBfIzM88FK/IDwh/0aNylHmmyL5kZkvoWtUCy/7YB6jx
P6dFgI+odhYBbd3rDVwi/jEOx5UJ/tZXDPYXwMP9AHH1fuyBra3WunvN04sRbcfsdRoUl7nG0KuV
utOEJd0hwZILn/jaBsnTjVqRNGr9rnxSsn6Kf5Xvm3YT7H3tSgSu1yJFqqAOuZg8CDqJcyF4+jJh
evq7Q8J/M1LkCMD909gIYD/sVHwsw2e5QAedpbb2ss1bf66xAvEiXXl1UAjX/LLe27Lni3hSEnaR
qPiDH5gOfj56XKhAKM7qk4Lf1tPJzyGPq/pJTBVyiC6CDmT/qHHsKocddZsrCy6dwpLTLNINytg0
wzdIR5ufqmehxbRw8YBei0kCXEQs+SBJhiPieN2WYa3gg+9RyFqni+xhe/tsBhD/+OIFygB7mlbj
6aE08G2ZODa/2NhX5THFdVchPPwZZ6Trbhe1eP16UvKiylg1K372yiyXeWgcaJabmtdBPp/xgQTb
A46f9IAYIIG7YhGiaRIKXbqQneNBS5P8wHrCUPKHk9hWMqehRzWIejte9c5pfQ5u4eo/OhXPAoo4
2yR2QuOWVGkC5ozT9xyil29sVEBs1avLLMsjP/LP5SF3P+vVeE3bvbT31yquxby7OqQu7rk2gAFp
DW7vHAq1RiCj4IZp+x2YgW7Y2w/IyJlvfADoobC3zSh9KByfkqH4mkhqd4IyEb3loxCpG8rYJ0TB
SfY9U17cn4VlCwa9TakfeNqo08d73YsPjPV4yPuBdYM9eafZhdUWfeqvnjePrEoLD10qXCRFX2y2
6BdSstIObCh6ygYW/5yKt0hZutsnKC5ZImc98Nsq+FigF+dD4nG2shuQXKgQUIWCpl+9iIEALWX0
wkXcIGpiWCZXPzX7GCgZnBJI+bpazDLEfWMa0rO4w7e8ru7X38yvOFcfFupixS1H4hrYPe82oZuf
QMPUsxQD1cdyAtdxIqIjc3uYU5Gt1p2bpmBxGKRqovdUGJg3ottbqTr8LJ9XY4cMwPs2mizE56sq
/2NdFvM6n3lAmh304nb8JnRFhA8wcvI+IFwGlV+jdt1fttEsIziPLCzM3lnWb92UiNWikBT7DksR
bOdLcN+3rukTfEHC7LuZ5MIOhmuEmVunugn6SOOcVUP9GrLGKF7dTx0BB8+3bUWEEs67eVsfokWA
a9hWRcvDBGas06FLg+P7ReuGul/Q/a6C9aKTh6XU8hodXiWAZbRFtvaGcm6uBntXnWSIlB4Pmo/H
vvxI4HTZCx6V27hbl6uxFuAgw8d+dKPf+KkATpmDarIo7dKzauFiOVrdjXbDcxYDNUWoq5wjUQJE
TptuVy+lU3uCbL4NM9jomnzfGvxc8Qx7v1cbqBwGLmPcn6BNXi5vLXDzE/Pd6CILOD20c5vV4mWP
2tCQDuKf77aTTSO/W+/dKiiLfEzTbFvtdSOa//R46Zc9Ppn0s7LcpU8G3U20T6FGocwGV/44L7lN
tmq78CFUi652SmZhYQE0+FybZyuwRqzIrLAHRcC9X/T8rKthJYW/LcRuqH+VfDTBnR/je91XKYDJ
T9omTuZ0lXoreebkOJvOBRD2rot0WHAH3YDQDcDCRCrfwA/7QhhgL6g/BtLOLv9ynN4XCehb+8YR
v2di0kRJmlM68wuevILTI9PPhxhEjgl8B6aK1U00y4Bx+NoXUGbe0AOeHCIQV/rnbKoi6OLj0nOD
p1tG7zbPU6okQtZ73x+MCITGGrG9iorxfi/ct1OsWCZahoYt8l6hVfPPs6R2KRAskeS5nBhS8Vid
HnXVx1pA9yglN1osynppe3OaB1d24i/RKpjg7RSYBeBIf1nUdJAe4zka3mIawdQItfzyvfNVkgiG
Vh2uuyJ7WKDGMbA7JYthtX5AXS3aiSB5AI2ualBAi3KVZ8SG9eZYU1dBAtEGxmW9lu3+n6u5qI6j
lemQqjTMFYE7A0WZqaPOjJ0aJxTXThlLtrRql2NSuwICO6k3m30U/+/R37SxeNCCfEp8hjbxD6Zi
aXT8LtCKwU4W1QIkxJAPoQSJG/2yHsnzzs52iTFrRW02pdta+2BOr3dH9bfsWNKMeO9yftZNNAbe
nrSqTXOzlwVZQlKrC756SAkprZgRKMEa5WB2FC6NUYH+OehzBhZWzrjNItRSqCal4AkahGNlwcp5
bXRtBrcdIhibkmgyYFuqWeBBVm+VN809+uU7BQ10nNLTeaRj0ID2PRGirwW9zYg+CRVbrPOO7BgH
sD0YzsSqDsEhPCRDAlLpJUqsKOh2jg5TaWqft1JKancHx7+DYf2Nlcm6dF3OSVN6pTjqv/A+j0yY
8aMIclNZDO0qI1o+hAeAzlKw/Y1Agrja7atmPW734UXSkp2rQYm3cSTaanP+t1L/KmidKUkJAh/B
SOQNfm/B96jgz1sL4VzpZzuxfHyjI0jTNA/HNoUiVhMFDtNCMJgIpvvmnKqz/wLqBoYSvvrS6tFQ
0byhAwEsg0U99V/D0owWGtWYVXZeoQeawyTLS2bSlPeiMIH4JEfArfGZ7Ma1E43QoTDYADJEebZX
uSDZGxA1s52qdlwu+KO2Fk8tu7dbIDXuhUvgrGIk5SyRSwoyCGi/bScIoG2Pre0BnfNr5AFHbvOY
SFP2hzF8tu71W90RRpScUlyrz0eqAvbOmlVxYsQCZKuHydJTDUwT1WRydR4ekDQBRIxgsv2Euoga
hbFIvq8AurgDMHyb+stHHFyVKFuRmv7U5NIbSHCUVTuQKhfX/CbKcI6larq+gkPBWIOCcQNXI0fI
3W1xk2beklW7a2Ui84co4vXHqgWGKHDlHUSD3CJN91hb1+yMO1JS77SqhkZ5bJKRTqjyv4H/W1cd
xm36TOpHM/DltelXIoErOWoWbamWgZa3t5sLQayB+rVDAeKMEDap69ObjIr+zSquh4gX3zZjBBiZ
uerUeqo2ZBv0i/b6JXud0tFhGB0RyMNbkp9pAX1bIbRSgeHy+K0/rGKCFIlFaxkO4vY8HBcJU9WA
A3B2BIk15J61rjKnEQceoypMlMbN1Z9NGTF1BDXPLLUSaoN6bKLfGLTqC/eT9OhyAohwR/4RcKNv
rqZHSPlCZWkbbQhR0GZwJmgyOJyWckWJQDQ6pts9S1Raif25EY2LTHsbzNgudxnq9D8r8IcB28H2
Elf5zmfF3iWchYoqNI749puCLyTuLk74BDgUV3JgAVktUA0nM/hJO2prub2Xhb8zlhrwEzU/XELt
TRYkoR5eho+NgnK/THXeLoSHKxcjtLv0LM5OXjG+h/888+VzjFNjOoSeiqws2OJlD+wTxkGp4zxk
jxQbbvM6qG4a3xAiHwOazQ7eAN1oo/gvVSSLOKpdkeAnDHl0ksb0Db2wylEfVLeDbEsYHOCkAs4z
qG3R+MSWGo1zT4TO4i1ONIRDz0v6/jqOG+amd9K7oQZXO7MgfwwLhVN3V/N5FvQuQR1zaP7Zl7Xw
kBcndVNiuvgRQj6B29mOqGxwV3gQeDg9H34lMyXQELOaNGXW/GtnXFw1lXeP0bd1NpHpDa7dshll
OdGYA9//jpFyDZjttycIQYjtdeLXLfKM4nO7KGxiagWd6nJt6LnWRJJbc04yZ++JY5cgDICzVVpK
vgrXmhqeFN+6REf4ksiyHXZ5GgcTH5gvXeYGRoFyGwVWKuciP1ePzKXVRFoGeblRhhdk0d0hP+n1
uaZmiI+0npgictAZdKwmKlBxJu726L/UgFqecwrLPnvvOgB1W3Fd2VpymqzQepab9auIR881ZfFN
hWDvS5Pr8jrVCZc+0q8QMoQGFhzuOqN3Wp1SQCMd/floNuBbyqo9pXeBBKPkcsl05ErxO365bxmX
+lRz3e8rpegY1pYscisyw1xtmNimM5Jfz5ovHf0DQf7ooj3hG9+tiFaC7rFuKxl1TuvynS3QjRfL
Xx1k1WyotzRzpVHA8E7wJEEimCK+9vZx+6QTSEwPht7c8zQB2O9Zqf0LrJl9t9BUhB2c+L8h871E
DB+N+K4HJy0fToAVOJpa9J/5NtFGaOihXjZWk3uUjCOuN1zigGXqo2HuSH7lJtNVM72MxipkNH5M
7Vo4xLGz0vPhTvM0IhiQQRbt33cq+SbUmmT9U6Mbzii5TpfKArnhKjl9bBPGCk93UpbSUZiB9UGz
euGTl4BnD86bELwyq12W18r+PVP0MQ2oVSgknvLcjDJE5K5vqcFPpu0Vw0FogxPaG9U23T2lviPV
OSyZhZO/pfOBxDnV8DI2BQADHl6YKkBJxkXiZIuFORLp7vslAKsr5NyvverQVnvODIILNaI7TwKn
cbhbvWszjZLjfS45XKS1IvkDNG5XN8h/0GqP8OkPe5GezE+punvHbtcuU25GSjVEt0yDFqZVHe7k
jyVG54rTheMGIbhsB9cj+h/bSj2t4ywVlfybNi7tiU9Co6gUJWOf624+VEZCAUYzbY+kyQdOoWto
LPmHdFVMDGO3F8GFHYt0iKnRvAyWDLTKnaZPZen8eLYbIbiAfL0LwzOTEf/vIqTpMlaehCbH4VaN
23VxCPMnAeiaEnMnODJn9tqy/4nKsq85eBrTSXYvI24bXQV9W8XtFbLBmwESUxT7/XRMWOphz/eO
c9ygaJU4vXEUzctPpI2lS9a+nesJsOm8temYnc2l2ZwYi7vcAH1JRwNfEIt7L0IMritMULeLaIOi
e00/mkTo3uXrj2zmlCXRk0/JadaudTW5NJ39eZWn1c/RS7kqLmBXmgXYFhX+RH3/pRz3id6Rv+we
T6EQCYB3Q74JNhVP3SAfpCUL6OwEFy+qZplDRHFh0M6RbFcpnkrXVW79vXI0dl9VdshllQfXWLhD
m4wEPtF2PXV0hqsthP/D/BtUB8/9/lmlJKNXTQfGIWVtq/YzIv7JELIZlFd/AaX1XX1UxQr0lPS5
1NEaUykKGkeZ4e5cNqkfyjSBHYFNLT4BxjyjxC9Zt7c/g+tnncm/6R7SLdyPQLl2QUP+9A3vmyAx
MhlnXIvlnlNnii2/4+8axnZv4vCPd21QZxY2nZifk1r3hyu3FTViLwzQSu6x5LEcJ4zSKs0fIW1Q
U6jCIsfP8PHTDUovgH+FP8OPbc+t+EdrTrhCY9fswMW2N8z1COFtvZWt/hkRzWmk78IbNoo1DR+x
gtO2u5xNByG76/XILr/4E0MwU46xpk9cBhcW9nVEbMVzuEwy+Pv2OFEWbCWWo7dTW37lP8dYOWqf
h14AEd3VDEJiWSyIUg2zxhc6XJ/b4pD3L89ST52c+fHSNBoMaj3ehBUZ5ejvDy7fXCKHjBNKIp1a
8Li+7xc+WDXQfQS4zn9rOetacoaXs5d4WQDo73yFI9aqpH0KSTjhUh2ul5jOnPm/bnqQQr13Frcz
Sz+7cf9q1Ft9LJ/JYEyrCIRMkYI07G2llCJdLTif5UFQuw9+e3G+pjQAUY8nu9EJaWQ41x496lL3
exnypJ9hKvjElMxked7te8KKZbxepgJPWSvl5S7iYH0mUjsAR/Fa6+dhBpCdMvy8h3Yy0i+wl0mr
QxMxL7s6ce3i/J6kQMEormdnep0Umnk4oAVGYsQDLpU5FlLlv6Yf0h4yi+PkesW+xoExZRfc5+2V
TU+kuMcZFeam1ggL/NbNKThf5UMEEbdC+1S8izy+8LlETdfNnnv2jlRzHNJY8dZLpDuTWmEJbwX3
6XT4aLIFO/qkl4/WaV/8sbkFHZy5KrEP77Khbxe9AySVLpVqmslxf9XcKYyoGr76rNXNnxLEL0rW
ba5pl6354dP+Vymd3kq1lRzjCzb8XkpyKtxG1Tfi5LI5weuwFLa4Jk2Bf1X7TSd0VnIBTcb9DpJA
0DeU5uohWz8WWMS8NRzWFtRk8FC2B2g4Ipski9PhR0ciwAUfXxaGgiDNXXewmU2sSZWhDLy/OuHt
fwQC385rQrKw4ainUuD89HHPCAIr9erwhvffo0+WMfpEgJwx0jA2aR0NJ+LpmmcG9RB3CZcCNVrA
MK7muaiG9btQ7eNqz6p0gwXLyv9fE+XgRtKomEitfEPFv+rFmR2v/2WmZ7hJ2q3vgXfFLiAje1n0
Cf0EGOwUNPhm6ie0ECnNckz+ZqqcdTGJRDBbfMGUhXBBD7RamobxsTRfWc2p5dIW3p1F6kl6kTcc
FCvXxT2gETyFZ+VTn5U/Al8XWRLDNubgsSm2V7eGqdKxP8DN7k21CTRTkJPy8SyASTIKJA6Zey/z
o590mxknV7EAAkSU6xLtjFSbXIXp1bLq0Mno5cXK7gNEK2NdtIeDwCQHzqcO4rVNkOzOl6qBra71
VD7zxE3eMAMgPmXlNXxM8HuLyK9IkJ6pbpPecyaOUyjGbN8t3G9jl+dkqECvg/sfLAIISIvm8xA7
foeMymL+FgnytBjcOSrEc8Grd1Ipc9zS5gKCZXvs2qnMQNhGCcUFDwTIZozjTrcI7kI8b0iO/8t6
ayAPtUJ/gY8yr5ib23pEbgDIqjLKNj+OXBfN74bZ7LTTMjjg9+bhKp3ycRMJNAzPtwnst0WSFs8h
oSdZTrUqyRHzJef+77NFPgFmrfZf0uVQ8YC67cBTkuLYj1YC4ae88EmLPfUpNzKI6ngY31oFMrDn
NwKp1ZuipqNHedyLot2jn9n3ZwXFFZxIp0doo1M6pICwA2PAA0qGwMP2Vy5iN7Gs3FCwnxaToU2+
FmLnIXx6UX9c2lf7MXZmgwSJ8+OVLiQ+75go7uNs8oHweiAd2hnHXdD8MZZlEKudTHalnMHmNmO1
HNRfx/25ju2i1gKD9GUhQ+RaohWGG5z4MUgnpR08dEeMRnm4/U8i/Iny68uOedWFnrxmj76mnfqc
vlXH/UyU5lxSdH6SaneEBEYnZEiucer4TsBgNV2Y5Tn47/Wibk76r0iV92p5n/zFCu5kBtM0YWLX
cX5Q45orMgD0FVPvaDvQzeoDKiPndgB7b3h4UDI15yT+CMrAa5JKvcefu+7G6fOZC20IJPDRScIB
PdmMYzhtCfsOPs/TPyrLt4qR6Ff5tzoAVbdk4YrNo7tx7RW00RGEANR3ofg/U0gRGj4nmFyzD3oa
2zDX3Hu3GFL88ExdCVeHzlLIFJJKosQ5pBIW/1fbBupBl1fQ+jfR6DDVNfxrODdX87IulGVDxM6X
qp6qy52JXi+QpwE9XTt16ah9LejZj/15kUIFny8SAc9uZtEs2H5fkgnVQt+9COio6JRYnQ+Pwqdc
eX7TEtX7c5Iy31R0g5TnsqvP680g05SQubSPGXTi0JlAWwaz32ZWZIF8D9EXlGyLeYC26mXSGrHY
FkhDhsTiB4qxBEDTtm6ImnOratq1caRk2f5VN8Ob20rTCMcFZG/WSnCRkbdONj73fIVx2gSJXgvn
UIHW+HgSy3sccIv/PfvTJ/yLph7AT4fCoJSvXsQalniznZrf/MEAAX2YlPsdrRR60+jXPHFN7UOz
MHoFSuke6hzAC06IOup6eUxRsVVNLFoNQm6Mnfah0ER7q3WSac179U4g3qWd4crt2AEuuz4q8TsW
U/qxeUtvNEaKLJYjQT1IQKCng2YfMuTFo89R4esg0rCqqzV2YiX1vxtzH8roWrtKicnrrZkEZP73
mAIBa6cOlbskV3qwDm7ZNZOOvkR1mTedfqyNNuIpkNTagzBHGHY0RXEGnO4UI2bDKIzhKpu7JLpd
KRx583BR95h/P5z6jUhpIXWiZ5VVF71rkOigTD2AA+9u91aF0L/V6KVCfi43oLzLgZ1tUj2uvOsv
IsRdC+PMdvmzMfL2xnhlSqqwFj3Uru6BOhPyvwoblsT5EBrgZCoRdcDJjO/Ph6vV0SLdSsucs8yx
JkELZroMtUkwBMBJ4kC05EKCoCAW5bpAjq3SWtfKIZzAGv9ILlOUVkt8eBtsu2IRobRDYhzsukkM
n+XQuunNBIZ52Io5ME+lJyeRlJhBEV24RlrauLpvx87wR6D9p2vvyem9vmI2TWjyDbwLQViYvYAy
5Jx4G0GgB9Sv2BiIA6n9JTPI3VNsCxYdnA1pPeQGvFsr+V8+KHngqYsYUIs0XiyejV/LYuxX+LZy
xaRBcDezKlqgY7/17XARnk/SqyOVJ6cx1xTGfadAvnA9aqD85H846jOzicx0KVFYtZddv7VmX6tE
o+Oyp4meAkBwy5vdKS3ldYWKaPgqjkJUvaKr4enXsnkJN6gDPD+BxacIn10BXDNjnmCGeNr70lWY
lO6sZo64E91ZJpOg93AjmI7MRwAfCFSITtHz4KS7fJi0Nyzt38DHbTGmQ1fHezTo/vb/CKXnjDRI
af+YXOndFAnuaYCwu+JbrUZ8s8oe8uNJfbn2Drm9+OINw6eRoq2ykbALTs810dPuk7j93Wry8U1s
8oX2c4fKLLl8tHdmtHGyTbplYPzROp5vHeItVkNzf17JNXnHLfaY4MyC/lItR8+Q6+UofQQpJ3OT
SjhJao+Dsub0MH55tfsG9Ec6whpdd8O82u+5LgzKWHLpyY+fd0pQti65ELfCpASP0L4uMPUAgUL6
oRrTBnFVtI3XKiTjjIxfWP4UqwU69U8Up2yEJxlNZL7f3T3iPm94XoZgiBxDFL+PTqLdW3ZkkXUH
Q4jmN79MvYc67dgQt5NfOnF+WR9w1d/2hciWFt+qxeYCMlQoDOjpD5BbAFRnclnz4WisTs9L5Wxw
W/gmRXH1TBfgGE3rn//FY4U6sSRzN5ndtiHHK4RiP8LShH7UI/e7h1eQw8XpJfWQI15Q5Pg5rKPw
lXpO/xOwqYZxxwSQz4v178f/f3nQlYm6AJXR1rTNVIPdP5Op7g8f82JRacN+EWPWulYQv+JCuc1e
qS/qIQa61+Q3Yvkrz3viDU3GH7IaSZlNBxgOPB+dTPz8sUaCqCSKoJ++HkCQPOMTiVpASt1GeEJk
Mm4UE0sRrqONY3vAAlolXzrno4Jmt+XlEZEhICEnxJs5ASdwV1EqSiC1NfC5pdO6TBsGBIsh0LBq
LcbQ038RvYKUaYJvnAAVgRxCQMHIwVPtA+jUedIO5i3M5XwIQQf9odjyOPIA7/QdevbfkqfLoFP5
+vaMdl88oVbMg037sUolHgcs4fwN8QuGz1DTipTsEBeu1cbWg9K5/PewLDAy+cgqlRrvln27BtVE
btrDk3LtievhrV+vBAS6G19REBN23FIXIOzQDvQo/TvU7ktbYhxSjOOj8jlUJv+th63WgrJ/QK2c
1t8Rxvgq8mcFWB0mVhPFCj/KYUwcyJd/flixZxzYkro4h2J3xcXtBrv1D2menQEeIb60xGz2lkG/
YOcoEhT056FHYXql2VL7m0mHBPCtltutWsygDjORv6KkW6jcXa2EnGLyGxA9nkzrGo5/kHk/8r9q
eoCKfYy5YHMRZVbYiNIKD3FAEvKf0BHktJ2gY78gKNcPYrHjPUIvuGvnpoeDnhMiMxD73dLT+8uw
WqTE1zspD1eZpmu3EOzhCeihsrBJj4DQJeY+vWq+nQrLIuv/zl5txS4MSuvFmrWDpRHI8+KNPSmZ
10kM5J+FrKXW5B8ePU0WNqqngI4g3FKBbYz//PgtlDGUDuW14QBNnxhAIRlwtx/uUHmbs3ep7dhp
ytU2jqgKX/+S26H+wHwFkq7ZdNI/BFPsVT+xck0XqObgxGEw2rlmjJgvdJ3FuXdDqv6HD4n9CCwY
mprzpbyevZ/YInVqcxyvF+ZdivJGTv1f2ctDsGYBwJQLIbv0y/IpbTYtcdRHEN6lRgwv/jfFRBm5
i5sm1vxucQgvC4LdJeQlHzPDSlzBNSQp6xwvpZ+fHp1lH66IffKEOiL59pHGcfB3vh1iddRaTahc
5xXspr7GdOBIkKVgNhmFt+L0DO1b7IGZ3JF0PgqEC6Kw//t05JC07Luz3DKi2lXNaSNYeywtl0yz
16WV4yiom1nJt8TwU7FG316JvZXUX4TYREoVZQeZLasDZ4+H/YjQwYB0FpuBZuHRA2PHhEV8k5V9
ju4jxJ3lju0Xjaz9Gz+zCALwFfmra5WBSCnx18/zjeuY9nHlC8E+0N7FJZ3BphaPe9h4hZIvOxqU
/N1g4qEpr5RN+3J6z5/+vk1Wj3m8NDMaPXJ2g+Nxv1/gqO3jSfHOhXReIyw71j0N49i+dfYUX7Hn
TUwPCOmKax/y1kT/EHPgT6AcU2/tak7ZqvK5yQ9MZmN4p09Ixru+MKGjiQbj31di+IKkEOots3ct
0/q18jNcM08PQOzkxIigr5yBhrv6nvS3pruGVHaXLCXm84RcfdWG0baSoC/UlXdWY+u00uTymfuI
YvdSe+2zbUpGw4MO2/gtIx9gSvAKzfuINA2ux24EKj13hOBoLTqRQiilBLCecwOKO1NgsR32ny/p
TzXtTL/voUf9jauax2b4LAwHPT+dAnvf2UCcR4QqHCc1vkF0FqaQuMhuFxAsGbWEkEW3Zyd1wQTu
FaeTP1I4nFrh9Tr6oV9YEH0+zu0CNiJBumKs6RxdufZICY6e0X2Ow3hpsGhLVOtH5YnUfJ/cotbi
kxFWlpQI0e/3/Ed/5junB72OPWz3wQkaDscHN8LiKzLxJGieu2HWsks9Ri7wuFGVMRTsKsH9nuC7
ctXD3xef4Yv47NfJG/FDe4I5hxGM1sGHSL8t7TcEydr48EWwowInJu+jmc1PX4d2HJYSzZ2AtLOo
7gIczJ74howZSkXxknaR6y8FYwsT+p8ZZLtoInrlkul4o5xEn1P1xmVlWqkHLljUJAp381Aj0YPj
FJOC8nrUlvn/iX/vJFCc9uo6oJIO9HL4tk3XHP825QIC+A0Jb6Ijm3LOlIA8hqBJlMaHBiTvxAIT
m17j6rTM8b5r6msDQHuMklIoc9FhjfH1s8zIE7jiw/8VELI3tscxrTIV1W0CCOA+pH10G+2V+IV5
HLrD+WQXDLuAZuIDw2sJo+X5VshyGWdZsyVu7Y07tCtGj5KyvvymdCM768v2KNlx699K6Kq3pwMS
/MlpiN3JotEfl1dHhoQRwaLxXB06Gc5E/pglV/VZ041ZmHccte9O0PvOVZBehuD0ttk3GTq7x1bq
wDzfBu/6e4mhohDzQ/RFp3zHYH6hOzuPkeB13kavFYqHbgcdIiMuWb2+LY5cE+WX8p6QWwVI0Jc7
n6HE6u/xmK5Lss5NOXZqaDdgtfa3S6cssU0BX4+MH8oSgvCTBefcfnkHGYKEGjDfxIaT4Phu/iRB
R8BwoNNP4Ir8Zx65sYOny3CpJqrugo6NSSOM+rUrzHl/zp6ZkRAkP4QD5dFleAEOnhdtTPZicHgv
cKCgwU7obvyBRV5M92mS7d8aMezn075+AFqW8/1hM/GQoONt+TM+VVkVIeySHgfZqxD/QN4UW9pi
2a8DGE2W4d6GSW7grwFrZc42Uec3/Fh0uEkyQ7+aoQvGaM7kqTBlmPEz8bItE6wre8mfv0ALRPkF
iNrqZGzcM8DssT5DtRA1SqjBlLlFngZHUs7J0bAd9Owt7xqDWoYtijWA0xd4TR91AXC0Rx0IGAq1
fuku0UYeM6yYCMeCbJ0LcTVPQ+CGSx5+TPolM3CvZBayAc4kdrteMt5K0ct27qEbUyxBS08Pffxs
zmWUZvLfjXttrYQNpuapRzmnxhyHd+cUoAVDvOZww3RapMX0w9uD6wqMcIDF03pUx6YxAap2FBlH
GB0eZ1b4LLLrTlQ6E1tU32ZFtKTZHeYoeD1KoI/KIOtIyKiKLDAnjbLkQ443o6v3oryRUwfDTFa4
9dKjLUkNc38DK7Xk7lHRVLcrxT581knMs5gjhzxdC/vFqfWTrh2ZPZx7lM47eFIHxhX6u2+wygdH
07CN/h6cB2ijA3Ra06fwDSvY7wkga9dLZVR1JwIQ6x0JPmo1wgejbTHqd+y85M63h8Vn6vvqfuwL
PltmIfVUtdRiWLxjmDYnQS0xXkKb6yJ4qm81LTm77xXJN2arjzXD42UjPwtD8CIo+PmYqG1jgmJz
wR2NYljVW/Yd2I6LNWrN8oAiDrEsOvl/b5qhCvEJjiBszw6vFP3nKWEeYzvqxuaIzx0SUl/qDgLO
a41xUR9F1tGQQXyPYb9FENh1r/lfA/Sc35A4Awyi73rWfEstZ3cz2OlF1L+ABMRCcSvy7/uXee4i
Za/TVvnxG3xva0sh1RCq1Ma2o4Ta5gHpgKaD4PpB7KsH0XS+KBgwGiPp79DR2mPA1B1PmHMi/6JI
2o3zOagrBh5B7y6W+VEvy6JAslj5ZDRmCZWCXXM5mI9h2fXRWgGiP4wirnZ/BKUx7BBZean6GkmO
0WyCi2+wOcQfTA5oi8m8zX/y6Ursw4DvX5OqDLHTaAK58Le6lzoOlBlwfTtUyCvHUBzp8kuuiO+u
kSrtEyopKP5aLqFkhllsOzOXRQlxPux6wSs+GGBkMuSyZDhUeQMpOhJ4QskmPjNb2AkYKeW8UfiD
mGBatBiPqwUnKoQ+EvPpwTGaqKjcQ6g9K5XEdeKWDIUXyjy7iLXf3qDn11QAZBTorUP0KMcLGf04
zRQhZtlAP+Xbv7YXI2pM51etougiKTJdkrKaf5Z3wvu+OALTqkggGnm3wh9l80N6AAuG4eZXwfw7
Gdp5LG9ZSVlIE/n3AqJA5kNnsek2H0V3RFpDXJrPkmkdXqRTjtZWWDIElZ5Z0m7biVSrK/wKmhbP
9xzj2lA+Ou08TXaDY3XcZR2FpYca7arCjQL4cQug9ihCpxeMDjkNvt2vJ/gu3B9lUtQPe9dqZNBi
8msTSlCHvBipI6uIXhJUyZ3USihm4n9RET2wOq1Lz1HdiUJYGnSUOjI7KL8mL3i/FvdBq0AUMJpD
Mcc0JI4YL8IClpeSL1khqc8+IMKmkvkMu97S5nXeWY7SFqvG6ueYlq56n5U4kkJQVZ42bpTn+M+7
5oMZix9QmDWXVhF5UTg8s/RGwxJ4MqXoyIHlbLn0LCltIiThO+uHu525gOI3T8orVxI52ouy6JZW
EGuh2swrPqhxjwUvD8MYjXq5ioK+ECYrVaNfcFGcc32SYi6yGlTb0XEevDWL3da3EdtObxweSb0g
dbEhYMSEIGKWN3u7SMsqKvnjYPO5uwxBjil5lQGXu4OxMz0q3TIwJMSWlNBamLpI0ie4qMEpV+eH
DwdBtRkCfySeaqw2ZzLJjzMOedtfJHM2piP0OjcQDnB8ss0hzGwcXJFpNoPvcbpmcyuyPO4MsMvs
nRV13W51W400NnOd4ZAMIjreenfp/z+F+TetsfHH3ebV5Qd8yg8E1u9XBOLirONiZ4lGA+d43cNy
mpVoxwwDlsSQaZt0Szw6aBPscrWD5ukl5a590zSGxaRoM+glde+y0dqmx0gBlHWdFXu+wMNa1QEP
vZvWn7l/lUEbspmBd1hVwQaJ8VzzdgkKFaBv0ax8DcCAP2eL68DeLNBgdnCtmfIjYOVBladWghDG
KLXTMoodvVR3Qe7pYeSCXjjD5eBPOqpLjSORSt3vygY7SlDrqZYA1xI5aqf9WzSb1t8VZoNBANSd
h8sCh/HuK+lXTWsZcvf1eTCjQLO6lDUEsPXNp5j3tJO/xa+W5jrBarru5Yc8/YKV4FSZytfgSAzv
CiCUAGkJD87j4CYIh3IM8S+fFX0DBJUDZWa+N76yXB16XM3J/bpPaRusTiKRDG2WY5nUK+ozaWkk
w7qjnaoKQnS4675iA9tnB5hj6AoM6F74V0UVppIJz4wLbWJHbqPMTLQKhu02VLSkYr44MHQ/hEHk
b7TJcRnhmzjZupn27+Fcy3KOohqCcXN9Jops59/5e9C4b+4B0Oq1pCpWyyZhHAmZVrwZaYCPTiHj
mdPLUClwBMfWVNNL9jYujkNdtYs8VL1cYHtydlpt9d/jPNeGVszOAjLlcTlRmObaVE/jLW2k5opj
60Q3B6IjtdqQxKmKREes1pzn7pBAJLvZKSg09Ej9ZYuSOKT65dSBOdGktiBAyXdP5m0FBI+XLfyS
scQwXheMgEXTm4h4z394qgMlwM1B2msu2bKXnzWe5fq6gWri2xLhrwgLFponyi065Caj0Es18UcO
JcnZXTfvIvi6///OmVjQpanM06hyK9s2mU9iVVQq0TrmzE2DRjpPtCKQZ10WLjU3vF3AP4Ho6oWi
SNty9/87HNfV7wD/yyN1gNI/mIpcVMsaJBoGYr8Mfpp3NJivrOyZAzPyhqaBXrooR3Vd7NlTwZvt
mPC6dZ+NI7Oo7l5LU7/ZQKeiPzBSxIMb5nranPPHdcYS2OoWfvK+6aUs036QH9VLbLmBmBG4ayXz
uLTsIoCwMjVskuvBiZgOR3ipSvjlh/85JWzcBJBeOgIfEQlhz9pTrb/vTOyUnsCmHJ1BDNcwVB1A
OAg1QL5v4+lWp6exbsxnlWMH131C4IaVa8N47O+OmhH4pwOPDatKgw/kzl8BQr1rnij4diJLg+Xy
81YFxz0X0MbVqtqMTI65nvivtjtqlkhKFmujQxXBCnzo0ErLSKOn8TbJsD5gVh/nmvfX9hJmTAcQ
FR92QWKtJRaV0jk+SWv1QlZswZRN1IeKrjq4ntcVJ6c94m7oNm6BQ18+lbPI8+Pu4JGSmKJWSpvH
0MNRdRhPbNN0Hxd8hcasC2fHtv+QOWc2zv6ZtJCozQBS4PhCFeVudfNaXkcovMZmwUVPEtsOudHq
s5pVYB1/Du+UErlwQexBB1xzy4ud8V76EM+r58BfzMJWHVC4aHILPLa2Yq4rE67xPQWqaAFUUmNw
05aocVgaqocc6/6fK7BmlnU+dCIYNxintfKF0g1DTcyPF12+7A5HthH0sJEEVOoaZmjYez1JPoIT
afDt+fM41AqiEc2TG7wVlhLXJetwBeQfEiCbwXhnF8z4fGd4F8/RF5cxkAjoDzN2JxALXecKW5qA
bgxUm12JEMplHwjqnU6RsdQ92GFkbzSQjUqu/vrGKZS3Oi9wdV2pvde/o0N/7E6LCdJn25QhpIST
Qjal5c2VatdcMtGlK7RoyVwTdLWzLbvCzQfqiMqAkx93lx8+p6gjXHrSCdP5TLjeRNR0INpzUBy6
gQ5VpKU/+bSVckRcaqvSch8ZK0t+1tCns5KrEUtmWpwUhciJ0/HnIKecCnjkj9krmuJn3BsqmTfG
ZEvL7zvGTuJH9ZxTq06TXPU2NAyCa2a08DcwZWA6IALSBbVM6F+TeF2Vgbsw5q8DBWPeb0TENCvo
lgDbXqPDlN2AP/ax7F82vD9LjkhyPN3W+rkc9esPeq0zhS8fUzbHvw2vgElvA6ZusQ94FCqi+Vxp
ABNK/h7afTNIJTq4Nyfkqq+/AmoMVHAjSW/yz23tYbvjPM94io48KwWRdiNvzEIaoJgzcX91Cq1J
DQs554IQRnoY46Atsu+3SuCXE1/RMGliM//nGka6uL3cBgQr+aQ8LwHevUf3//DIyIloBnIkUvpS
wp8jLpNCQPitKG2MJw+k9jJYnjNMqVJXA+RQ0nEMBMCSdnGJWX53UiUXXeS2FSEOHrOVHvWMQy2T
GBBc5W/aGjz2X8450DjyKOMPKRyq/Jn6BwLMQY6zRnQqFmDASlxtqRBAC6N9rPjBQ40Aenrgd8W/
ySQwKaNYHzvaHVeOlyvXEBFhNunaHpugEnfwr0cz7LglPcK+0MoCQ3xKlXhDYFMF/DnPJGikydHb
ccUhA1k0DU9BtTcq0QQun/925ZAYwRJPCmhnmaGI5PDG9rDlDi0mztx9muyjFTcpr47X5rLJ4HUp
dYqU/vz+HczyImC09Pg72tOnGyqnvCb9ZOZ773ftmWelhK7kwp6KLu9H2au6VtAlgWqiGi9eBofP
1KSBG++OEU/gpCsykmo4JV6rg5Vbu3NRHNqj/nNP9cF3mjUOD8VtsOAVx7FN/9UAS+dr6Z+SUwi+
tIJCocMw1HGtI7KSVgbCdkdy2cwYZ10x7FZqJEKoWO0fPKMxB/aENRDqPgUeStv1JN+l1ebpqL0l
LEOcEStDR8Cny2zhlyFvZN194cr+0dJvgLIB+zpBEl26gZ+yxHRz9WxnFaQUruX6X40HFKhzMBvz
9lRbBq/7DeCZVk01EgwFHzKXLUuFPk1nUDlUCOhtV1bRFYSL8uFfQkB9y0lKSJaGoeMFQPgZWQSp
naGCwclt/PhyevHsbJ70fCoQibkVqZWprslsxSkhF50vuFwJmSyhpYTB5ovp3HMOVS7I27sftIOV
FrWqnTOKDmM5MbQKC5cYs5axIIcNdg46/MCb3siL1zO6XE6lNaeu6VW6VN0LtBCC9cuaMbawqiG3
3iFoMzCGdI97icaqYFfm1xUSDBsHmw3NekSdv6Ps7FWXCA7Px5X76/tzWcu1VtGIAonTKBskw+Rp
uPH9GXNgi2gCLUZnV1gYywu1WKp/KGtpkLMSpZ04/9LGCcXIt/ufhvajF0zkJNRWPJ8Nq5CKK1M9
9RUIBnkyqz3osCvf7qymv+g5j6UdPdK2k4wVDmzEaFNloUaWrq5qslBsbB+uMOCQViURKK9bkaCi
Rxi8kIhhs6RtQgwSrNB5lLfDSFQUqYxQJxrIqPtzl45Swwm02oyBxSH1zckxEOk933crbuSlGpLq
lDUYLWZOyVqTPwgDox6TUOPRLWj9UR8wb5XyJtMXDcZ+no7aKfTcF9Ylm1BnHPymU3wSR6X/retw
chyvK8sV+/wxTH2+GrKJSlwiMRCobbqn4KxR6KE0CUZlcVx8s7CYW1hQa2lgB7LO3vXX3Pcn2+2B
PlXf+y6ju+Xht8mLhKkyp9Ao70+4CYmmNROFtNsQ2N2uDdebdlACBCxiu7ytkrMLKE3oMCMEKmAf
7x1/167aqgvi9mQ8KrN4UFXZUhBVQTz7v2bUOqykwfNcmt9qx5sxRYNMAaJQc/pyurLqiGiQu9ka
oq3vdIhhGbCwLl+oRp/vgd17HE/G/Hq+RlLex3qTI7PVDhZ5hV7LTK/j57dnXPBJghyML6+A7vtf
jiV0UHQ2Oqt3/SxuVp0Li94wtDxvvzjKO0sS78rIMoXguRDuI+pXDhHZS23WePyPGHO04j9dUnpE
ahK8nVRf+Fc1rf70Q0mx/t9hKCLtfhRKRAn+J7ldMFyXj6XadXC19mA5+LE4+/o0xOgYYP/h1wZt
BfIKKWlDT2+8qVbNBUnuediGCyCxYWxlvjgd12kO5o0ZxIIl5FwFsvXz3rbFeQTziNS6TjdDD2jd
LEv89OtcQlbCvDr2OFqvuvvjnF3tol2HqBtAPNyoUOr0nxIhnYiygk3pe/MlOKSPloLJtGVH3st/
ifmny/YA+dRyWSgE2Z6ZjCNHCYcCdtlKxf6/T3R7fQGaqb7V9+r45ng5HU4rfgg/6Yry3HGDM9lD
XzuZXfk+M2PJhl3i32WMV9jPtTdxCp6HaOs409cFpsmTuA8i6ExJgNoSSXRjjtpOPbeIL35hpZfK
dH2f6I+mRpgV8s2SQnmiOdh9Jbl93H5/wx1UBCywA7xdV51c2gz3rr4P7e+O9lRBYnHciD0jmadM
wk03qmOeOsYi9Kgo2h/Gft8JP1635VdZQZJKnM1Exu1rjQ6FH0IFO0wvnPP+x4abWGAsaDCJhjja
bKJdxpZ3X/Gfa1ldX17kEEvMLF9ThO5bodUqcyU8AQB0wFWPRcNPLX63QLebRYq0P6Lf5inHYgkx
NiUdIMHRBYGKhoI4RNH7xmXs/C76l3+0PL1vRWMZ8+e64Ir3GsSdVz83dcaqQ/pXlp2rC3/Sz3ex
ryXEGbwgtq8MOdghhxvSsJlN5LNOOU7MGFMvfBkensuT8d+2/tK5laUYVDX+YW2avqHYaJ0cfCFs
1q0UfKEcBpLCoiRduhBLy9XXYaGtoEpXd57DmORHi+xUpOrAV++FUoGvSSTq9G9/iRu6kjDNM59k
au11Kq8G6q66nVB6Xsysr0Q+WeyEskdm+FmLunQbqVtTsOnBFbsL6cHOJMfG8frRtHufCYFfhdJo
qV26uxtjpcfZkQBvIdEHzb6volnWEltNDyM/PGnuAZPms44TlDu+3N2LXiwVige8Isj06I3+ZIWK
6DHBp+/WzpS4k8gAKPxM1VJVtio5ErFADPjyqcVqUWPFVKhEjYg5JwhLwFSpg5lU+jwk+3BFFgKI
1m01Om2bQW2mGmSJwhDuZAn2QTdJNNYewFMTwoALk+XlffCdNJwBUDO0S5Rrii/5ZsVcG4rS+LNi
m8C7fb/6RcD2QNJKntA4xqbY5MTJ7ely1kcakGQbx3K+3q8Pnk3V/FdJ0ZKIvneTV8R21Z6zJtOV
ine+X19L5LE7Bro0JF53XHmH6VyOXTw65qCg8oSWrzD9jAFKmk7zxB4hpH+TJOCqwX//GpIFZaHG
knZpQU3Q1+YkMDCbtbDJDqHKcxkH2RHhNPCWBpv+6B6OycY2b/IVGGqY/qWZ64NmzKBZ4NJe+/TE
7dIrzMXQLKQFeqDNWuV/wWioHr3qDugSfF2sh0KUDlAOzYVnyvvTUI8J2nTopYQ7SlrnvPr6MLko
dqXMESvvakACwDGA8wOcXxDCxbpwBYxtQEaxbTJiN1qoW6YqK1aZ8JCNEqLE3TPiHXGBiE5Ruh24
qNXt9FsxV6Ser51dkYtw8Ko5Bqd1FQ7h05UuHo/FILFIqjJQbK615sZUfe3ofVKMdhtFaMDQCcF/
I5Xh7pd3Xb6zhuzP7FHC2WfBdRHt9saI6jKkM5d18ePZI5XDSEGvMq95bes9iIC7QjY6vI6yCxu5
5jCADP2Kq8emftz34Fl8sq7qFWIaxaL4NF9LNJG3f9gEZqeFsdS9JzfbaS0D7S3zXfUDkf6Ftb6C
QClCCMXOYSxUp0rMXI7Kb85p+GUnSbrySLBmfOhOfEamDzOV1uBxgpRksW9+3xi+LTSrIRjxBSDo
Y6oWDJ9LC+Jcc4gJjPgWD040lP9MuZY5KLL+Rh2HNU1E6skRaITwZ24E3AbaXtX6EMTvKobWzs+J
sRmdfMn+HKF+4jDHM1vbE3PCdzk8FCR5Bhdk9bwG21bNuF60K3ONlXL07ytPs+LvlZHuAq9cdj6i
iUYxUgIfZFviiV+szgSCu0ZTiYY7FYc803/smEerStKNYXvLC4ar/yzuTOLgM2Q1nZONKZ0I+tC7
anML+7cpuveVAsyr1kszXQcds0gz8aXf3qWVWdGg1+q1bOhj7Bn86vHrFSUmWo//s3iKWgOx/g4a
UNtyQmR6qwHsVde16RnBYHaErt+wuxn+7q/4xE1Y/VRyxKFxWKR6Yq2mcn/ZhspoS9maO/jmqcXe
y7eCXJIz39o2vMOFnH1MMb6KbUZ4kq931v8290mf4AhjiI63Wi2BCRhQIb2zVgp9IFxiRFKWFRg6
ysVgIIi1x5/WLrpotbVpJ/NGCHmAa9wSCn39tzj5dwJXYai/PuO074KVcOE70Ns0sGkqdLauU+Yc
AfC9CS5Pd5GKSD/zxeUaCOT5vC/AfwL/C8Gi6Jvo9x+1CqiBwx/+JF9JZFK7PUglwL1WxneBUVnY
n1m67X7ptKzZwFOpiZWGxK/oajy6muCqm1qOmX8g8YFjh4VKtqn9WFGSY/Xf/N9EyVSDpWI1uczP
zaGO4d3dSi2ZrGHK0Bl8jy0FcdfU8yPbydXwntLyilsENS7ezNBjb4oSiSmmmlb/pvSbjhM7aUug
PRHnzihPIihuLm1BUpeorG33QtcuJue+CnxIgLy4uibCa+bbWIawUkp/Qdq9ZY0zWL620Sougvrz
hUigGC1S5C+Mzgq+1aj0McxiUbajfCzdjRt3Jg0CIK8UIVAvfloOHixOYEyKlRNazzlcTxKTuHAk
vlxIGSb1T1ZqMFP8exuQziO1P6nt7r+BiHCFQTo5uLp1eG9Yeu8hiVfBYs3K2y+1qTFephabbSe2
3XlWjzrmF58JRgUS5dj7FWqNmKyMILFCmaTscNJUCeQPm6guWls9uAzPwOLpXAw6YxGJZPe6kSbh
iS3Ab9o5tRzfkRtO89rvZ720lvQs5F/Ca9qDFlZzlqDNxs/ktzEihToQGli2BTe5vnCjyxitRsVh
nRYUitDbTxnPN1mChZnhkqlnIxxbF7okLEonwio+Yt/iADchBkMCghmkf/LO7xMKKPJkDTmyqy67
K+abkhH5dbgbG2lrjF9465nguiV4g9GdJ324+updRCtCHSVfNucxWZeJTr0VYBqdt69Em6N8aQje
XapwAk+boElDhMamdj0+iuFaxZn/Jq/IVezLjVfvv++UUn3zQC8vtOBs7NYoTT5+oCRFfhtBpvKz
kf1EUbtX4c1ooBlKv1ngYsbbSAto1yps6iJTyjH5jVlETN+ph3Wx0Xgrdr1BiYdGclwmfJUdugJW
GAsnqNxwbTYe600sbaeMpzAOUrQ/4U2caFk82RSfBDMvPmh5Z/XBPmipwcZ6cwOHmEUHOG1FtWz6
nmuRrYXVXUVxW4ACipvtBX+JXmxV0euN5Z3tvo7+okE4+MijqqyXsVNMooRzPm5zWfHuLkWlLc6q
aaB1Mokn2c2KrnEBYuvQDE7mMtYpumpZb/FzbM329cdem4Tok/J/LhjEwvvRQ1BJr0jFqq6y9OI+
ayeMOMrfZH0twXQa1RW0TbsIbM3TUJtL/8TU0qn7aUv9lonLGCv4Pj9qnAt1ULu3SsYm7bNGAqIg
P2+6FRj11JQ4Y3ZrPKHuGAmXAViAZ/TfYa/nEI2P3bQVZSPEV+44sGFoymvMHnMVSvNItlWOZMoJ
y1eWxSAvYKGo8Sjzg06Tnduym3M9dj/N4VYn8Up8ftWO1UPzeoLwO419HO49uMCD8mbuw1dD29Ii
sI4J9DeTiy2Kp/wXoiMLwV5c/4xupWcj8VlxGDku2UzP5+L8aCbYvfiuvVqLlu/QcjHXn/YvYWBF
UgN3v1TgEmURug70S/OVPYhXqgIzAGKejq3VMmy3+fgj/m7XUQmNgrIdEb+Ikw6cPDn0xO4+NWoF
zf3Z31ULRtEhLuZEXLUkddKM6GJq1FnuN5ppyqkRvuDeoR8I7VoGo95I5fYXJ9Gx3n1E+K3qYIp8
Z2xExPnGyCK7ppGvRyBpVZDQvRiDlUCKoeXYJQhDjF5i3wxsQAP3x/2qEggacfjaf5Jm6tj/xeyv
lF5nFwa4EpQUC18x3FbfkxfDFcLEzcAPtjby84hwB94Z0ArO2c9TR8j3jLbUciBLKxPt1GJp/fxi
F9V8VeOSsYB24JFzrYXyy5HzBQq6fYFnllmYLkFMl6wrYGti280zJwN9xJnLsBNh+s0TgXvgo+SK
u/atOIJLK2baAL5vUpfhXNFV8yDN0V8WAK9+g1SstMTcBsRpGUrveWAYbqalTQ01OgKVRF7I1qAV
akmxHqDtNvSxa0TJo2FboseEQsXMAm2Bm0XEphOZRe4OsilWAT0Xxs2wyYrK5hyJln2NOkppahv/
+PI2tmARaLCvB7FDeYhe373pGxc0Z3/a9Y3VF5NZy8Vao6yHyKPH3v/fKWpurJ3vV70B3avlhnVv
jOOW5+JtijfCG54rh/xqNDYMm0r3lFnk9aXkWkTWZGiLcg19RYHhSRNpgkarr/m2AQeiQwBfE4ac
U1BrIA2WWEeMMs7FYD76QX/CfzBoKXFpSlaLmaLjjTJLB4TwUfDVY67EzXwtVd7Z2m0g44KzxzSh
j0lZo09AfOk8Ggsz7Wvdle6EGOEDLiyJzmlfkLqQMxOB6sFrPNVtP7A1F44+4Ce4bksAduew3TJa
ihaLJd5qqh9g1I8R5eAP9jN8TFkuU5TuUksxD3qLoqNUMtS+Pdzca7lRzy7jAqDh9Y7zlNm/eu/D
9E11OaXOmS6WexNskuLpb76rOmA2Cu2YFOVerFUOFKhBYWtuH6BuRSZGIEjNlJTg0oiOHCvGbQJU
Ddsh/EvGb97vHfPPZIrco9lHRHHSW2eVJvxVLQKdUN/BzVqMVZruPeCyXZJW2M/exkI8SKEPq73T
RtE+A9FjIGdXpqq+msy5Qqa1/oiOmGy3P8q3V031MzOadnWrLlOMnBSckV6BacOVEzUru2uF0ory
cabQBWnIE236KieNty1kAxki2LW77hkdVtBp77j1ykDnSqWtwPfZbLdYJkHwlTA9zCNzoFeRkUfz
6HkGYCgBUbSpFuyhxhJysiOg7AghMUczTuYQW/EXsweYKxuJIyuVsaipQmTthprl5o12GXcIhfsE
AS2GVXkzahHQf+OTc4dPeQPpPT3BkYX8JI453c6tL8rtf+jl479ogC66p5ENR3qTENxz9BXET7Ez
mG9JGhDk3JCeNZzEY7eM7oFQ1kZwtXgdIAGqjE0+nw7u7170our/s021b6YTYKkTpDuo0giDT2Qc
ucQjLv7Um3zJKvqenX/1wD3KWF1L/Qf1FBqa0ZbAzl+/+QH/ZmJDRMmRJJ7J7OjFUncIGT8rO1KI
HDdOA/O+AlFj/a4WxidrLfcWYqs8wcBc3nFVdY0TVY16UznHthb/gGH4yNgHIN1SIhcdx8FXivDI
E677+h501lBQyaoA9ny2PkrgN3avXeYjz0+TnDCXlx8cQ5xf1fhpiVttizv8iA0ZGvqZjfm6ggWG
tQ71HMg/x2kkcNoEUl3G4RVuddVNOx3HQwy1PwgsJ2o28ml59lmJV1swOKuPmSrU/wjv2y9T3rNZ
khfxi41588Mw3xTgV/VgYDLJ+a0OPgeHeuWQW0Sf6o+MLpRgPnK12IHs2yOaU84LUYilvZWJMEhf
ukkYQcJHgXFj7n7yTQY1o2iXxnnFZnSo9zSBDiN8pBfqvbY+0nJrKTivvKg66Y5s1/SYS8WxmyWa
dKndkLx3BEI7RVPqoGTkEyu23siZRJTznApZqOQdP6ms03LbtMC3VuZQkb1x9q3t2An6/Hh0wyP7
x0Cz9QObBk3sGAaaZwHM1ElRyqSR8UveCfPEphUqN8cyXIJ+2QWnDBq6YQ8L2erqUMc3I+JjlDhI
POWMJMT9jY0vdKMQkJI/jz+HJMJDdTiBnsdYRLmX4e3g0VsYCwxT+ZD/heU7+OMVRidfKD1e2wFO
8kZVt8brutuZN+h9ybIOmpZdelDLFuqHkkxOhjO+WjDSBphp9wIf+eD1YyHzGAMrHPJFZ0tQCy2S
TncD6SdvgPTHE8yDJQyo9s+ia4Z6YMuxe2554DQrY45qf01l8ZbOuRu2rff7Hpy3iImrY9vTDtYQ
HUoEuN2ebUEnErjN7AsYFJtsjjzteKVTQ2Arndi2ivKopw4K0WSn2mtSX9znblfeJMwHUe52VDr8
EObj0lLabo8AWtOtrkL+qIQab1Rb8UsUMdVKD+DYvsuXmx1Q1YjRSxHiPUjvk4SpM6jjOIuhAMrA
/zEY72k59T+N8mt5an9pTdI0yPy0AH3ZATxVTteIaF8t1Hviht5d9ZaHCDKsopT9Sw47BVVU1HhD
PMoTVHwSA4tpAxKMRvWSGo8Jo0YiwcWkZQIZvodkJHkhBbi5iL4GvzEhQMDWqzC0oKgUscDvcqP5
5viJTIPIbGHxy+9NQ+gq2MZ+MEgaTX8vKthTTXGYROSiR3Q9hk/O34Gte4q93ofUHlfAmPGgy58W
rPQeVfvEObMTVUW3zNka8tmVDYg2nEKgD34+bkR1C/M06ABnsibBHhafXk20PdbZP8o7Mchca2q1
1qbzjM8ziISf+Ijpvxz3oBqPpNtf2hZdOXRlC47MWBCXIM4ZhAC5EPsQZp3dbd8fii14tUm5V+Eg
dDWvSOwTFue4M2G6b5QVFPqXr7gL4griBy6P0u/pXei1EyX5/Lmniz2j+bxV8QyxL7tCCEv5uA+9
jRXmaP5c3kKrVCVIpmWtwYhqOoqPOx7A4skE2Z5Zg3BySg7peoi6LqI9JFppKsScOXx6iXZxp2FX
lg6kfa1PTRP5mjQN99Znk3nwP7ChMeHougPiAyR/MpNznrxSCBnq2FrUNx7vQzwYPD0BeqJXZ8Yu
gJKMZzn2ORTGtQckaL5UXeCV1hHpmODH6RfXSpYMc5yT2u63HcSJWDBIca96JHzGHFTvB21uvYZ5
88SAbcsxU0t1IGUWeNleorxZg75qzKD2JIy9ozvNEuDYDZWwNjzLTUP1wKtQsC+SCoOW/OV1qKgl
Tuf5Mcw/sbSgbMQ54b/dR+JDFlNP+fDA33UZDaz5LoFPbC0yWdQiKKzat6kQy/7PuTrGS8k0bma3
gUf3iJguyGjQohBAx33JMKvn7dgt8vjFD5FfsfJgYHjJ01n9Z/8KIymPIttP9cRQq4RXfX2DKIyZ
lXlHHrbZcTzioWg7o57Vugu4RYKeGtO7KYhmiVM0WLpvExSIwwwC5xeYEYBPrcVdny4CtYG7oCik
m+QSq8HpKsBDIq1OHeSEdRb7AG3slUqn5ED7HfdxJCcKmoIqBlcvxfChWHp6DVWdA0vWBqzkppSq
HLMuZDtoaWBIWH87uB8MIDwTbb13rnCa/SUMVvePrlduFAnXU6LAy/YM+WC/riXgxkCbgGkdxj9z
b5wUQ8aacnPHZO520xdzCo33gYL9Vz9u6hcJ/CzoN8ENhNPrJhXXODbW4ATSjOFv9qIXnuJDGSpD
RXFnK4ghnXBQpGzsp+oMcqP6TxogFkUJBFT8pF4tray6Sw6ymPEDNmdUZjGp6M4u2wckExSY7VBG
CVZRt14D2+jEmwz2XfwP5K/jJhsjW7ziEEESA0C73dgI3miTZaV9C/RXLqrqhNtYZ1m+AHE+HAvT
+41mjzxopIbvtjFAQ46q6aJX0S1l/ix7262qx+LWLyajtseNl05EOWZvINnsk8QXAy8y15mzABnf
vLpEMnNfqVQFIK0/v21Jsdhh9MkjRASvlLc66OiB348TnTr87udMZMK07Xsv1y5zrb04FV6RV46w
GYrZWZE5cSiy6gffcVmXeX0Bj6Te4JDygIQApmwwC1bTeYL2CLHOhJz819Dwnv6Qw079/7C6Y8rH
jxP3V5GiBkfJ4ZRWv19jak+Q4/DJT3DgolJqoV4VcpS75rz62m+HyQVDW1xSshFoEWYjs4opIrGR
rcgjjvfOihTZ/RP2CN2/0Nh6uTcUBmBDPZeHUN1zCcfoOJgjhjoToRdRCqYcqR9zXoIkE75jBaPi
tn9cXi1IUh+wart0iKk86sM1wvInocHAG4gA80YE2wM8gHxEa3lwlOhHku0JK7/GDgjRwTHE9W94
WZTBSqOS5qWeuRbn0yYQpOFqL2hK7XJunZFEMONJ54UsghuqkdQfxLklGSrgeh0ukC7DgeCH9ZYk
yH2iPmRwMCajgoFEAfA2yCpOj63caQElE3G+aBT5ehGxXFKjUydk+BA+YMcxUuoPcP9c0hNdBFIp
j7jok6g4/ewqyvh6HFZNaDVu7pAj6lFfAQX74ZD0WRAMhNQfbqhwEXwyEACvFn5OvqB/9Y4IMeIw
B4vkFHlKRAhoAubY7m8Yqqt7IwD8BYiGCK6hrhhXDjNwrzE7TIn+nDrdakzb9IeYrWNNzNS/cO4i
FmoKwG+WInggivSYVFLvPUVuURS8BMvjyBzWcG/OKObFidvbbGfbP5FzkEEXprZ90TS+yggHfGuM
xIK9Wlzm8itab65QZWily52Nj1V7UqagLfgEDHLrx1FlE+gSBd/E//mLBrvwo0u4PFFondM1vXPd
9vQQUxV69+2yYEjNgv8D8xrcmU6tjRsKM4x0jgu9ngO9Y7z6yh0YHGIy9+BABNBXTZ0t7rwbgce0
9anuTGp/MPy2aOTs2MWntwDZJ8CMxCGs3VO9fxny5PXbKUz0Z+xykq/5MfOQcHZb7jUH/rTHBZVj
yHJS6H8D7eoQ/JErATgI6BSALjx3drlYek+ZwXktVwLnrRogMEjmTIov1IYKyzKLtdthXQFZaAuq
u5XjsIVeDU2gqlhmupXI/OYG+lp0Y7acRvCX2hE8PF/pUQw8nmLPfIcTO27AilSmTCS+zfFVV/PN
QBSNWs1YEXPmbK/79cA/V7g4yi/rGvdrbBLLB7Qr5/KwDVehUULrOc07SWC+IZ9RLsSUeJC9Tghv
yCU59hXtWGpNzsB0Vl9EHt3UFu0G+RsUDI7qDfV+WCUW2OLEUSmhimnLoRj1cUIqn7GPhf8e5EGl
/6b7udzAO/qDLZUxA+8mJG5MDouSdpMXSxw4fuoRFsoZp27cqLu2+fpWO2jfDNZrB6DWFAgzvb/k
UyJui0liY7qatcbT25tBj2yJv0B5DB/9LnysVLj+wl3+hAtVEXmkad1qKODvgUsQupGH6fGihR18
R36nPyNhF97nHpudSGCYqBXOv9iPy28XS6AVJhMCU5vP7wtELFhGLnh0L0XwNmXFs35BC1MTohMB
DxZD93YpK+yMmpm1oIfhBUyGzkmGgT6c1X/uJksj0wEafAPFyRzPFcy5VAIh//1T4tRTeqIdCBBi
A+PXsFQl4I3JEb3oJIi9urpeTG5qp6AT2JEEAZAMGKg6fZwn2nq029IfW1O0740zS2rJDCSrh4SX
vx41K+5bVOBXbSdmF1XbixaUYWnnaspQuR1hn6KcTmHuFeoMsy/NYOXCBsk90o1C6a6cGe4qOK1V
Jc6dy35YXFWlANe85hOiQjWzdHPVArHz68wlhu5/DEQ53m0pGFR96qeqGuK0+Pji06c+G3xc+6wY
e4nyZhgU684nEeVjY0LSz0QNNnG2mI41OSQ4+fkeiFK8+ZrhQzygYrHe7c9NplcB244R2Tx1hdyC
bbG/SGPTYK/lnYzzRYb4O9Vbxx5UmHSYxejfQ/VlYbpWA7VNfyRSL4AZNOtK9ivS5gQQZXU04L3m
LKnKHx2HbWSOkjftjRPSkijKjx6lTARwp0y21tWsLlTcLPyB+ybglwjczeQnppKtx8jdf86Rb51A
yFiXGDrrrQPv6WoUuvhEK2Rue0gUNkO04M828/4dS+Cfxa2zu3kuKO5eQbpW9jJO812lDhrDhrd7
E/gXNuKMoX8eRF/g/4j9KlGAn9MtXQaKi3CrbKekBm3Aq7GB00SyyatqjIA5Qp7bwvusFcCp4gdm
OYICmi7iz2wwf17lPQwUTTg9J3eRcUuKUMCNLpxYrKSgBUJgTWSWb+3f9fhHOlCbasAdeDsVKsbu
5GPF+whKKd1Nr6RIDHWJQyefIhRBX7Me8tnbjz5unet2rFR4Ev5VEzZFEyaLmg92XXR3KR7NaEqG
mXJ478ox4DLMD1Qob8/nwkTAONhIKoLif9a5Q5F+OfycjGtnIW4F50Q4kMIr8f/Khbl5u6knalWW
5w8v2R8yF+6eHIvZC1P8J61VoyMt6C08qWKeiphAFSimUqT5JRW7SlGW1z9CNCDGbTLiZ3bMAbIu
s1NBDcm2mTH4FLwrYtQifM2cHHhLCmiYlUWaNvc3XUldUaJJbPApFpCSOkwImHwRZVl8XiQJm22H
eeB3QvNSrZdp+7Jyxn5N2BGj8l2BOC1mqK60E3XEEVkBNrUZ+HFT3KuZ5kd1KrzdiMYquvBA6RH3
6FfI+z+WWcjTYl2SIVlxaVcXYFjDgGnt3VN05cxcFhAeGd931jpFl7aYUFfErV8nC2df+4QzD3qW
xX5/BQFFj8C9X9doykdoXfeybQhVBy72alSb+8i0YkO/UsmlAP0UTN1fxsFsd2YYI8aG56tkEcmO
VwlvUOEvesXUpUXqCd9DdPNTusO6vCB9r0Vlsk/rOW3r5ugMAzpaOXkVGOqDqehdRO9p1YRDFR1u
eFYGq1U09VqGkDImg2BQO14WxagGLW0RWhpiU0nRYsjnSA1IsclD9/Bp0wDQobAVff6dzLjboEuV
h4NzUINJrEP9huRFKIXE2ESs5XFPiRT2XPqPv0S/1Jgmgezf/bjy2Immgh161Vi5MMWS6NAeDVvb
7rffhUoHKXm5nASX30omL7NbRWBeu1LE9vOvCW4/Y2nWzh9ZjE/ez57ufvpW5KHKqKzFlykHf95P
4/zDkcDLCGFUkCdKJFe4F+QJsYYJs/ooJHt6PUnckVtbHvI9Wmwu8eeoifktu2GMLUYNfFQ66exY
a4SIb0jpRTBaTxSBhY6xlv61UCGbpJK0toT0QgqS0uypkLETp6Xl2Sa60w7WBCCe8aS1BPSGFp9K
YrKCT06Gf3zl73JfpJBgImAy67CEDEZEHe5Xigxrn8F/cQjS+7NCGFAV9ChDv2uFrFvJs7R0BF+v
+EeQuIm+0DFgM1G1dSoKvwUJ3XhdeBIB7NwyphikbSxFPeBdv42Qo4cES3RIE07/YjrNdCntvp9D
btgE146yUPZuydWsFexb1nY1xK7XE/lgXrc7+x8QH4PSFZ3HHviy/bcQYvWeYgwOnRV6+vU+5wR1
4n/j5Fd9yqWxQPnDuUNuLVOxGXrj2OWwBN8l7ya8BfZdMsfQM3ulg6QzM61gyaUTEOW2eBmPDt9C
iodO2rk4BrU43GIoD/kFR9iX8Ql28aGF9rUK9fBgFloQMeFW1FGoveMZai8piarpyJhkM+q46YX/
yoVQYf7QeqBQ1Hfz7L2YrNmrg8vWZUiUm8a7Gj4vkgNQH/hAfK4JobGwrr4xo74UBhoRT3KfLQ/f
rf0ZxMn/62Ayxf6J96NYxAgZktQy5UwUG0i1n42PVgijz5YMKIGtiGsPNRKxGzQMnCJEXTj+NCTj
1XlpRsgKk/5fotZegf+bWae9C/8LQbQMj3iUvEnVlN0fR6bZ+jecZjMW6Inm1qdXNrPUMv8O84sS
hkuCscvXnovZu0gt0Mvx0QuMWjm5ubb10AerzNKEU/SHDe51V/xsaOwMCnobl0u31/LKdSMjwpqK
FYSzkXLXO6xQptFJBT9Up+TCeLseHz5A33yETKkCAjDHIlJw7XDy7WmAt8zdWPpwlBAyo/PavZ/M
DaE1CIEYISJG9UMtZ6Uf//R1l+w6lM4AT7Jf1GpqBkEKVaVAJjA+85+HRdnB+97rEIaEqJVBMrFE
SmK1SXYqyKFxVcnQOmmrQwvV5nx0PdbqttBqGXPaSKjg/XBTIEoEW02rDY5vo7RKlCBRpsAOF60T
rsetw//rpF9cKLbF9Vt+LcGtfKUAxWD7nWPxRRpYIBydadmEDM9JluWKAPO9qonOaHhwpLzcvonx
EuKVzD3FZj5xGYld56ApZcbzwM0BSpfGeYQTlSoFy4CU/W12Sn6R4MkiNpKM9mu81wLd44igI3SA
3hJM2eAaV5CLGzObpOrWv+b5tBTRPE/jyB9SlbAKFmc9Q5BTbxWpc4ldt1OsArj5ztr9Xfj0lv8/
EVaCVXkT69LlrD/Y2/aXmznC52Eyy5VcRBFdGtz4baQwwh2nISA81rG4UxGlocNLdlYPYngsNSlM
kB1fYcEmRwTFQPa+9WNupu6IE0aFS+W9f3ZbBYhm7dP8yrgXFN6yadTDaFvM8zyhbPzU1Nkuxt9A
H11niXLaDjiMjqSvnbey/ICAJtCHxtja9eN2NgFSlOhcLo91APpn+aKIRi5jfzaWI2R4902zhqAm
n0SjR3Vp7J38gilfdwfQz9ncnhhTvJbNgBIon9xz1aong0VAOtaYaTyWOYwh45IBDJvMmw//jHjn
hv4pRd3BKSKMcl3PvaqVgsDP8lziZByPDCXQVYFYoHi9lXvxcZo/hzzkhCLuvReaME60hs2hFSCA
DxHJOQW9fzBRg6hGY2GFeBhoWlV59i69prZ1wCrTXEqh/R/lkFXAu+61A6ahzfA9zm19gsCC9ZOu
uAbtNTwTA0qGy/iMw4CG46kiXuejgyXokU3uhUxoYt3um2u5ms6asFrpKbNefEKKR51E3TRgJSxQ
Soper7084S3R1jgHd411qqGv1F0KjT9AOf3XlL7Yj2ZtHBII2yAc/TicYQggjAumCx+i6qLox7nK
ovrbt2MvYD5lbWKeidT29SAD947HIdmVo72Lop/eg+qEMTgydv6Cq1OuH8WQbjjscsHCkKWsUiCp
0Z7EQTTDBeF2+yE/VyID5CF7MSRgVpo8xiyB8fobEBd95pYnvfZ6DU183GrAr1ujpW3VqVreF9EL
gfYpmiq+K5QIHNs4EiL6jpmE8PWXqRXcnUlAAsR1GEkAlbch5O7WbcTKlWXc9SLvL0xnQHbPxMp0
hykBf/D+GClOIMTuAyrLWFu2rH4Sp0vp5SLyHoedaOiNsi2ROJWuCUVVxyonrLAL2FJv+mOZghMj
fKB5qYrg4PnB60/1ZVvVSoX+gbwy/vxQdbYrtskxR5j7ATLYf04v1qRXAcMQAOY/NV7DHAHDIsIW
qkxC2ndCIMcl1IbKfy5WHFno5Aza0oHakd1M4sieD3yRvDM1z9nYPAZURYuxUNVFYyVguSjeRjRz
Hhj7w0InpcBfM/6VvlYaOgKh8pO98uqCOZo/Zn+fTBdVCovdrsU8791LWiQpUExP0fyjrqKInLJP
Jj1NQSXGnIxgYCeactdey+gXuYxMga6f/fXQKf5WTT5X2efEK1HttWTl1NmOWp8BQuGJ504673fD
bXK8AIi9lP8HKUT86JlHp2XvX5sTZiOFw1YXCXWeGmGRstPze8mBMv3ugW3JyXmsqYlvub7e6UbM
6N5qTqnBMEQ3W7gptfVDcVJ5/wjlhJ/9n9aNZUkgb7rD9uFWwlmJwB/TCMF6ZFT2zfK2O8ZgMPBu
YgIjLNzC99lHSQS6XgqRyXvfVnAlqX8s8q5vpN2bYiw+F/BLiyhSNsiL0uQiVhxAOdcu/vpw1VUM
GfNQurS0tbtyEv9Gu1Q6tccY0Fr8vgSDrz7tDZgQODEAxfpYpysTuRJK4cX3swlhV/tD7zUgd5EZ
VCXJLi3/n/r1o4gSQOpI9rICYhGNuH+sVAfA1jzZr46bCZdNOAD3H+nDnMPPZpkkBy0N737iKcRV
a7DXOQzXFF79WeUjDq+BULsvckbviAT0sC+2EvxszdQBQu3pyCzWWTx/sbZuQ0VKyNREtrr2+mKR
o8qNOF659Ho7Yo1tmXULNOALINa44M/ZUUnDoEKgo/JZQ6aFgBFWTNieYmA0KYSBHQwJF0MLjcNs
USqZ29l4efOTpxwPY1ZGkL+9V4rNEq0LmCaUyzBxOYpap81InVcCK11BUmPvGkkw2QARhnhEPvcv
KFM/2FiQfqxgG/325lh0o0s9RZe+IPP0KG25aD7tyOC0RvVGSJxQsHmh9BXHrxMstP6UCllWwBvB
ODJ4enlXMcMafCLviHdRMMfxJBbiB0+481phqtnL5FzsQkkC2AdShmpEWjPePuhdoGO29ZwS0HbL
2VE64UKUV8n6R8XGvZQuU596mujJyi07mUDp0wTvgdA2bVaKQaaLcUfi4Xre1ZDe0twgIeFmIctC
kKcqhjk1xUizLcOaZwPsgfYY5sZtVAmLUmfTsQRR4tCvDLfQ0Jx9/wgIPkdsf19IwW05G521NUCp
S8bBnRyoYEzkzy4ttCsOIFb7hjwYajygJ8V8JZBMqIlZQYVUWhFQDtuTEINhra4TBOH6D9VIRB2Y
/lKeENtJNyNHJoK+ZNtBOTKSaJv7LZ17q5mZjN7h32gK1D/wIPplLncSjfvGO2fdja75yv8ziSHm
jewBUCaHzXsMi/Pl1lNVm6xh79XQpxc+N331D6ZhM/2pCtleajVAsp5RE5PhdKcyvbpoU0MTEapE
DmcoXJiEqqG2DFN+EG7C/1H5Zce8ICPCDYUW5kuUxBM6srhN/FaVunhEMGzhVNU0JT767rU8AGpD
K7Vyn8Gegv3XjwMcWh1171g3B0O3QCOMsOPQRxZu5V7gIg26CdVXjLPNPraJUyZis9JQT8QFJLXb
Lnq5p5krhnajh/LKTDIVg+NLPdKRi0pRZmqx8PpHIvx2A1P7NHGKMlfwswuH5wv9g9V2sr7kvP9y
nsUEdspNSVmMZNdKkrmKFmk6p2sUGTat4Qnf/IdUeewHK49JjUW6E4ud46LRVlZIBtFlTwcIpxac
KXtjzdrCpAdWF4X7WxP5um+56I7PYg5Nc2S7OB6bsXwstxtJsS0Nrfmlokqfn5wOEGAZ4+wUh4wA
pEstxqnqpnUHfTt9iQ7L53rB01Kr9RAqZa2DRVBgHLzpkvy7DYmWBSnyuZ0vUF9CcbIJQ18IYBiw
P03fhafjajhOsSDMbxGfr5oB+J4x5tYHQSq1E/68CL4T1S6pNRjvOIMCmzf64Kkgbw5b+GmJQWWr
ft1Pluhdhwkf9WjrYiKj/pTeiNheBNL7rVYsYBvoXrQDp8SThLEbU0vFsthKcNUbToNFw2xdy/1w
TcrWQYI/4ZsGpc3CF+/QTW8Bwihd1Mz71h6xZ3WBj3XEKItsC9oaJK+vsQgucBcPcw6r/OW+hpoB
hLyFoLA7cOwN/KqT+b+Ssu6CWZMaFa8Bbitk5SbwV6NS4iHJ63SS+KRPMDrv/+Os1MYz8gwkxOMw
WUTcq+AIk7rPLp+92VPlFGB2XXjFL4YpNHVIpge7aBElOZQA9kNQSfQ4l+sPqYvyJLSUgR86YcwB
SPQCjLGAdxcEiWZqq29v9FPrKWnxtKIP/ncC37RDUKKV1E0j315I276pmJKqZkD4chfaMBMUwvUW
eMz7kd2sFNJ5iPzZDvyExQD7rLtzxECJs1965LwzM8hGkKtk5pVsAyXOW4JQI91DCFcBRVXr5nqE
HwUgZywopO1l8QQN/m2ePNvOf/Mf5TBUrXi6sFED0UIFyUiQJkq/m1koxKXCHqDXALxERbM8drNe
biXh3qDvM6R+IiYmFv+ZG5W5d+EUqHhOlBwtav9ktyJhiYEH7V7Y3esARkn2wnC4mzZiuQOpC2bV
T45nQOkmfRpo89CRVwI6Eehl1hH0uvSQ3Q97a6/UwaXIpmoNbt8EMmPZH1EFqp46toFwXp1fF5JB
Xr1U2Wv7v2rNExZgLl1UX5mInJu9e7Yt2jNROwR2UsvX5AKucpPLv6rg9ww3WeJ+0wfQAWEIYL9N
rfmFcTlZg3b8Ztz9JUQUl6D04MwHYjDvENy1ZEAd0TvayI895EZ2Ja9g1cLW8Wzdai48oW2l2JXb
c4AIMSZCXcbyC1UP+b7JK5ygY4hEV9O+XPbar3u0Pk8EazFs4bjyWBt4dAYVFFnAFXpB74wz5hnQ
/XVHRO9J7W3vM8RQyWwUXfIMsnGJQ4MPCGGo/ORR4deZkBQawsKT1J9Eire1HPnq1oEUI0kxVX3H
/KB9/2up1kazoN+w+D+Tp1n/qx7VNnYYq/Wf0k+yIpFJmBeGL0NPQJLyGKYDIZ6m6uuKsu+2njMu
mW1bdadmiE2mnziQ93eXok70/WwfqWZcFXCodjGof9Ru0SwooHJzlsAN1kLy4qvfR6aU57EkxZcR
K2MsKwJEus7ZPL64vnZWU5S+W4/egpdoBLaXtL7g84pfjBauMNZCE81gCYqao19y2gYwQVkVDVlS
jOG84Cy1gRAocXrXL1s8ERcx42vAkKeH69I1JjCGPPKG1qVeSVnzSGfkHgCBnK2PaVwTGcKUOzee
XDoOefFzTEtRWBms2MAf8sEe12nijhAG+VGrqFd4Nb4OVTj/k0+rDv7YXlFqKsaJwNbJHC3eJxI8
N3eHGs9npEp4kMWycvU7W7TTn5w3MuNZFmAqsYbwJ8/b/+9pv1TpApfTu+FoHHZmPval1RVjifVK
IhCGv9IWO5LuyP61JkVzfHbDDApHOAZYW73WyUvav1rA65lCdszu+XxnzJ9eqngpDZyQNG70LZNa
J2hmzjpQTIlezgXql6NpEXo9nS/cEImzTvT/JoHjUq2tMnawWUHNKbyC+nfz8ttHqOOf9DbK6opV
CunFz2JH6L44UBgXwYpb7Gy3zFRFbOgab8j+3x36rPDL4A0+XWyb6KL2XoOLJpKi3VifbUR1pZpM
tr8wD7jOoqhs5B0uZ5VtCFK2XexA4430F/xoC4TQWQNUjO8Unh6E+qp2QthkzFYosp+d+Bt5OcjJ
McmCoh7hZKceB/h1zXFS6ok76S7J19ht+7+HF2xK8phiIV7abC5s2jmc0zaPu1NW5oFjtTivhA1G
pP35p0fTkNxgyZlb3ih7H8+mTki4Cb/wwRiRK0je0CUakv/ZdryIc6N5aNr8k5439umHEdESxa4k
t8T14BwUxIYtofqNMitkE6Jnv11Xx5CDX6Yo6o1U4yzDaF2kKLxgcU/5AzGcD1UXCXjxE4a7o4Uu
fGY6bpB6RnxSeSLLMjXdhAG5W0dJAr+bTkkE/cdla9tMXwpyiV/07bZ9eAm+i89Z7Pya23skXSiD
9Oq2DA4EA/aTJLoNfvxAD7sShoxjZhrT81apqzCbOiXlPSwak8926VVb3x2MS+EzSwnOyZ8MpY28
yT27wyGdp9FlxdT273q9YblktpA2fU8PN4Rxcta7zzLBpxufLjNyhTlGIEbvniAOuuX1aRDBjS8b
jnyYe4UnKa9X18CB3JqQpb6mcAvPvyjUwH34CP2KjZAhLqAi2kx+wPZd3ntjRxWGJ2pmMtVl4WHQ
pe3w6aunzqhDDMYv5PMg9oVq/IaCZ/ZrYGKHfGY6cxYtQy2Zx3EC++udvk6F2vXo8TOTncLHDlVK
4VZRSoSBGABFvGp3buKXctTGIoFfoErbVNXOA8TkpD5N6zeeaepG2KStV7TmBcFUwML2Oamj0aho
dYFP3frx4yUxjrFz5AUGlKRgwyMUtzWYohwtJqg61ByBrRHIF06s7kcKa2gLA9Buwxi0ka5i9ipn
ww4WK8WTbNmVon59h9L0JrGSD3cdpw/htfPZGqG9XLbwrR9uS+0f1PcuK+PON2jOQm8WAMJhee2n
G6418uzo8IoKueR48mR6Fgt4FRwH71AqPUdU/QVBpbMOQFJsKXyYD7knTm4t1UK8o2sOJYBeb6lw
vjMxP85scqBB6vNoUI709oDaXR8AlqERfK1Ts6THuikYQdvz2VVXPsRCRucMdmyTTtM3ohvu7eCs
XUGmv6ojHxca+d6D84iSQhBALT5caQAVP2pK5SLGLpAmFYynOb2CBFm02WVpi5CfJDxQash6bqFe
xy2oZRGpbgE4vT3pqaxpJ0CiRCr6xcD/engIjhmLXgqnfLP2D89eP6eVB6uH6l1ymStcVww1p7pY
pIghZ4zTBnk1OTpt0AsjVPZf/YYAd8LemhtNrWCpP5uAPsBDOYW4wU0sdf1o5uVZHmXtyOlZd6q7
xSavHwyuUIUKoxCmD4hn357AwGoQOGtbAvwBXRjgdpXqHJ4ckfw1HIWMnPWOD6mcCLTAfkl43OBg
K14CRrWCwHYuXRIpX18NXaoeTp/wJtLOqCpBpgpPGnB1wfbP7ZhSy7CWiT7LfnvfASnUwVDwBSY4
pcrCVhVEp+5NRjr1bnBBQGv63/7x7j9QHtjYwdLXbZy1yGE/r8rvZZlKJvPNBu7tfbu4B9tXLNKd
R0WRMHzdNKtvlmnhPdyFt+8BNV2MdWSyTYP831koZpSklkHt96Z4kuqqoe+lzPwlpluoexESTWB+
fLXVbVBrx1QjY0OzzUbUyWN7/i7R7tf5IqDVKXlZZ/DPyfXSQbk2Vnleisvbc+2ezRedHfraoTbO
lY3uMzNGQrmkXFrZ4GPcYw3MSE+NiwSFTUWoxgo8NG8R7aNmEApU/LwLvhK+kcUAbJiALiaIzl1k
EvGYyEcQ9P6IqXkbbaYxjWtR1vHYBt4RT6O/Xrr/zK20zougx2PLiVtcl98++hwvTnguj1oK1sEC
6CvENm7zHYTSf72wq048Lzs06SMotX3SaxLweFqrCcM+uJNaUJHS27XlOs+ZT+09UE+xY7BBK+wi
uZKDqRRjB/on1x0a4wq+v2PtgSk4cYFS/DrEsRuxfu2jyxnquFteeA91YEXs/Rbp4QOZK+ac2Pcj
b51zdrw1gGBEyLg+q8FiWEQed/nrOdEYItQ+aW+DYpESLzXmXG5TUfbqDMi8nHguBTxA+XM/9XrJ
ucyS3G+SCKIkIedcUte9AhsM7v1b4xObtDOI1vQb6DQCirOSXPHP5bqXCobI6w7W/s1HkzdEBD0q
HS2Hh1BBcjn2l+asupOIiiZKftK//fVaQ7E6Ub5Gs58zgiquMsBi9BPJhU/B/Nxuslx6+cicwXm0
Ch9sI24cTIDWW+eok3dDw/z41bLGpfcp6D/NqPiCVEqJmZU4zoOG5eK7+fY9Y6tIymGtBxTYPsIw
RUe2r2iyS6lUmv9Is/HnYxXPhKIp1Q1TZHCZV+lrG3cyKH1hGK0+6yO23tIto5BIP6sHA5583yxi
yhnHhaEiG+6diCiADRUbIYCRl1ArenX7I+W01gkqksmKzROzcvrZzssIeEJklBS+NW2tgrwjj2o9
+qqLuEiuBNzdO9hWAbViggwFs7CarBc7mlpZ5cdSvNir4liEbZkBGizKgtjIEkG4XedxOYLG7rtr
kC/jEoV0hTkeZYLJ49Z60kv1HFpoAHmlMnuVaWzabrI0CSA26zvF245CQNi2YBpr90C4ONabOdqK
WOMf3szzHo7VnA3yYkMpSWt1fQ7XZqqUradAYMruA4RvuSBQNthQiEuVbBGEnzpSXqxQjkfB7BzV
6vhSRvPhGXzinpCGU1vTVfsN+83srJdmIpicedDTYb2PzB4BNPcl06j8xYYy3bYWjh4HUfdwrQ8p
DajPZj2YgMb+CSSqeEWRNc6Ml72VKmrOxNZPOYw7iPji41ezRqPdVcmZvtsOZkaPR/Bi/zfXSg7S
P8Tjlj5mD403zI2CgJSx+LLpPoXa/HeyeqmvYY1csWHNAHthgVkQXdUHTo0puGX0Tv7vEGH90qyO
z4VupnxQCvE9yahGY+GKC3bXLr6VXziSROmJA2QwH2groLLBSjrTPyKbeLMCHR/E9bqTaKvldAGj
BRpP4BG3j3Pil5hlX8JAYzIDgNZ+aalMSib9KYDzWKOIqinApQtX74mm/YQuv43fTUshG4fO2zoG
J+e5ntPKOWWdghXTWYpfsrF9SuJ9tbsraxzs8sCbcHYGAKqV3ksAnn+QluueedHl5P3n5LrgeuHr
wvq1RvhqP9rxLPYMhAoCaosoMCyFGI9HCR2XvRMWpGroqJY57ePRxuiR9yFpnDiFSB3/mb7hQsAQ
JXVrlQzOSRSOqXhkNjwrly422GL53hlGqknzc7mvQ0RE2m2TDgwa5xWd0j4wWF3XOtPMDcbCx/yM
B5iSmhyGYWYs9l4u+FQUnw3zV1LQFSY5Z4m+HQZNWMEAQtNXa+lie+IId1fBh6RCk9beg5kJ6QXm
4NBmCTZMTh4YrGw+dcfaDRqMCOuuqhYoAyv9fxoKljvc3AKiiFRyxgYC64slZybV/qzGyEw4bV1j
LuBKkudajQjJae38yJjkamZbEDThsO+X4BoA9Ke6tbeJWqrp1nva0pBgS4T/UJBh62CIEX2TbEYE
mJc1zKDZV17UlQAc7U57W14HIdKtutFxl+PmhkxuvXuIGxiaXtGIEz/dmDfg+DkEjfHoCurbP0xE
A5h2pl21FaL+VsLHYdRgxwL79DWB9s00Fd1tyKnamRdswVNEwKyPk/cWVBi8xtDo2nm0fJNljETc
RNlTA6ukWQIxn5XGJiSX0an+Couhsoz2/eF+aAA9DHOcYXlM+yD0+TGFAW1Bn95ZG336ar1BvVkr
cAlOmDFTyrOPpJH7JsLCjOKj3jfbmg5BkC3BDmdxJjNASzzPgrjawYOiosLg7HZySdr2q2vtP2If
Mw+rxEpBZ1b0Goe7UPxDA173DPPeALKs1wocNHO7361EbesSm+476MbUetjdU+E21NHwG/5UqkV8
nIPOGajRGwyogbThu6pLpI8lb4r5ubdLXjGrRipyE8G9vh/VhAlO2wRMDh2rUbyl6dUeNBiBKD3A
Us+uDupkVlGsk0bH6kltOIKUXLOQepFbwWccKt5Q4fMjGRshr/cK483+6msJGr4ENOp4ti9PkEi2
Ls6tiZWdJE+nCQ4LTpLfCIsWnxTaBd+7DQXcaeIWk1AV6qe2xPcdjM1vlwSsARN8l0hYFxpCVI9z
qLxWZxQSP9BnEceeWkBGiZFVECCOS2CItgi6aYCfqRrKfhNijR0iUOvFN9TPWRlu2MBQyHnahDQA
YeNiJhp5YT9BW7PkCWcDi/WKuNFjHsOya6awVHNMQMXfhplKsr7jL4Yvl4JZYcAyVHvP5NgB02IT
yaiuZaMHz/3x8EOgl1cP7Q/peelCaSSv5rCp+hL5mVmF8WaSn2E4nohQJDo6k5sECJz8dpSRRW1X
PJk00qI2kc52Oc0gXKUu3CkzlNbQWQarqqoBqe91tJ1JPeK7m6GV3eC6jrOExNV7lmnu19FDubgT
/AgxoJRu19UsV7sU1jHEYl0kAssDafuK2UnOi0kMIZjj07vrBIVfryz4b+cEoHC6FgASE9ItvWyj
x58roVGbI3q5swSiaWgwg2RSNsc0kXk0S47jIp1n56ARPiMn3pPMHLrFbmnnXKhS0JUC1v7MxYtK
ZHDZlhC3QKLihMSe34Krjfr3BepgDDEZoP8f05sG7jolkB0ADj+iwTjhO8eRE+g5P1YDUCnABcyu
DyRRwAS8uBIAmxwDfWA8YnOyAq6KPRIa02skoQmdED+nsWCteLJcwO/6WdlaQ8iH26ThFxUYAyqL
uWz7Ina3/qiepRVr1s42wMpuFbq7zXhNSzdpz9xDzoSHtapsdj4ivfKIJuptDw5DmJhToRCVmdF2
t+ujyQFQ5WmXsIOhthYFhFPRf54gPv1CohGmpXOADgTXtLq+f1+F2ahhmIyz2gyehOuWb+uflyh/
R1iG5R0/KqY9b4nNSKv2m/M2G0cjfknaIYxsfyXvwgooSFlbxjnMkp+xmQYT/jif2DgFsFSMQh48
M7hR2RGXRybK/UCPZal7tz4uSTbFiM2mk9vfNmAlN67535hGBGcdOciVKjAXt7x8ZZ4MAvYI7wwa
ug/h1jPhDYyyvLeQHaSNBS4KmDWWoRm+8nudz4EVxf/U+juOfUsKSvzWQbkUYon/skj0wB53Z6KB
WgmJNWLAftEGgmldZ+MOHtuuK+eWfkUbOXx8kErXXfhtsWmhBd8poTKltFDgGeK8OC8Npuekprge
iQZDwm1/QF8GDww0evP+T7OgU16KtK5QYgaaA2HFFZma/RTHTqSKtC0761pX+2lMNHfQLkqOQSNp
mO5Yd4E+t+pVh6guqrguG0ipjlDImTEOjjfEFM746hmDfCpYNPnmpNM1+4GxzurHsCZ6RpbilbfQ
f3uAgX+s7tPl2X4T5kx3tRG93/K4Yux2Ow/ezXlglhl3zwHhxyQtnD6qmrFt/40huD3hItimXONY
4UJbznXJg8DVICMLRpPbzE8ndyH1oZAX0hcS0mZ5jC9i5benjJK6OyeDhXyylhsaGLTWHHp5I9o5
0x68gbbi89Af+x7CZb7Jbvf8ds0Nhszd4S6h5o9RsI7LL0KKT2ofN3K36Q9Y5XwdPbcwFiXaI7tG
ju40aFwmZhn0mvAEV34wGfp+fm/Rt4TtAFuxXoI0rzz6paQCbPLieP4jWYkHZymGjqLiGs8ziUaT
2b4W7i3dOXWqUceFiv9B537K5/Zgjua2sbofAA4idZsZ628iRpF/+JVLe4ICsZ2tB7C0MORCu7vr
MUCYZ/0iUAt6C8BhG04PwBjKpJRKB0rgHJ4Qnm/UrWR3m/JqNylhmj1Pq9B7qkgUQdKP/XVoEC8j
U4EdYgV8yoWCEtjy/c5+ABGbt70qy9XD/gpMN31KSL5EKnH904/Ao/0Axe2yYv2QtpeTdYJe3ZjB
vOwP/OMS3hD4MYYLArIktJHP3A804qTrwH9j7x/bXylMxfVKgGspH5o965S47xbmKzT9kZY3Zh+O
20fmvCj+QV1mK9bZaCj7iOdR8CeftBm+pPsZQrKIdpe2SJpvtKWvUxKUYmaDbBntV+j09XDFeSEJ
DS3h1MHUncZ7AIU2TjlQ8BQE83ijYEzfi+0TwmpjZVJXFTeX4HM3CoN+AQXaNZbnGGtQgoYLfjxG
UsSdTf9+EMTpL206kEZ82GU+LXlPWiFO0BZXQH/6eXjbYh5XlL2uiIcoAF5U2iN7pTrRsl8ICIFW
lEtkD0E/5qytnyNBTrv3XM+4HIDPXSe/DWoflm6HxDGityDRWfG1auyzLHFjMlQNJ1oekiUOLiAO
djYup60AvySetM8qy1VqQ+MlO2qjPGfwYCUTRijhgIp8pRk/TPYQ+gTZxwIlrf9BBvc+4ubVczMX
NmGBPHqBByfBtqShhk2MjUFWx0soIuMn+wMCDdo7iezj3IswaoUINX2xCZXwPYnWAEEbqIAUyoEa
a6/MbicdTaZf2rLDMKsxr041HN4f8xKaAl3GPR527T2embbB9/MhD3U7I24mPdooHabhzfb3/REM
ZJUrhI1BuZBGddkav6nNhFo5+uCpeJ5Xx9dKOIcHvh4bt2ByntQrHm4TepewVku7GZQFClxYZ1Bz
I4NgaYWaXnep86u3sMExEMKNtigeyAAZ/tGjsZ36dY5laSZ6S+BczJa3g0VPHfmfQEvu1SMf5QfP
P3XWHe7EFPd+QA48zNGZSgDZqLH81/JApq66hRvNQym5JuRn4M5+enTQBtBz2qZxV14Jsl1ZDcpn
jDjXsC+9SqrDwFMnO0LPlxPZGfFkMc4gK5xtguNSMtm45mLw049JXNOWjgh4JSwDWweRwBgd/HrE
DI/AqD9zc8dd5q5vnWnwrHmX/9t6rUt1dyp+UDgj+W/htcI9b9GqxiASh2/GL6dOFjqFWv24ot9R
SHZCffO99205Wnb0Wflgi0jjIBm3EUkJThSlzQBbR1+QrUzoPGNGhZ2fSoxWV4PMW3n9UTgecxet
/k8jw1Dc5VbnPncCJaMyG4hjuoqGyqQJfzYn9U2ZKjFcA479ZmOQYRCIlqWuBFPiUSTAUlO6W+o9
I0VlsUBsNM7LG3aO0CX+sY5qfX7Eb6G8X1moVBjsLuAL2rmVdw/XHWZA6JQIqY4M3zAzQms7sls5
gxUDYhCuZ4BifAj3vyWFAHuvSItyLFYU6mdjVC38Uuqw7xS9GYVF6josh9kETgK8uwbmsUPBlcbN
vP2YXmrdqkEh/u2gUJ1EeTjzxV2cEIgky/8IXLZkr7spzIiyhYILiC66eXNhtPMpC7j6F8H7ejAP
QqfqsOmp7bRYcMrAPj5zIrCN68dboc8ffgRTPylj3QnBfTsFQbRj/LnuuwK/B7B02l1kgqMMB2OX
Gt3GkePpqK19o2LcoSG9vlXMDFUoITvAPTrhS6pRs08FiWZUrE3JjI8Yr3lNDmeP4SDYR9fkE+Wh
wPRfLW3hvrHRWQBszvQoOmeOdt8x74GOKdxY7H16tzjrFJJXnOBpnikpSvgQCYzSG4ixGDob3oHD
+ZqmlLnicO6MM8kkPyu/nNLnbYpeEa5kftxveHiX/qW8B4iREnGiGl8rwTA3lZTcrR4uaUZyfKQF
yOmNijhOlORf4Zax9e2HEhElUeZlFhohuBmqFSPvu4fI36ibkKzUgJKAcIW9gQPClDfhWeH+oivJ
4kn2zoUc4LGlX3AqBTwo3G+c7oBFvdUPer1OTaiQoOqv2DIl5WLH1mG5ay4aSb2oEmAdf1WDdk0k
zjPuJb5ruShWQ24EuPvxvx+g42dqRb3f9rarjlcEoYXRGoQbknBFscustOdbDwRimUr9yO/KO0m1
UaWQLEguxlKQIoYr9N/RCv5Nf7UivyMAOXahenFQH4ABIDBEskb4RAhV0w4QhcFI1aESHMYIKlVx
/lzK0M3+A2QgZ6hKBdTD1GnmAmnOt8zOTSBUXW65v2p9/j/8JKbOqfDVAz9JQx/GneQjcim50/EJ
loIazoBmn/AOPTmq5rLbjOin2jubRntgBO4TKTKt/yJasphHI0JABGWrVqtmsC1tZRQVA5mcqzwJ
4+g4mrdYK1BUikXLgy2466LLsVl7Kg/Q91SbSL/UWV+PiYRrYhmcCTeJRVTp1i4gjJhDcleL9Nw0
RAsrox9maRTS6IPRlY+kypMtugBJQhAxuTt2TMzM4NZg9s+3xdrJWYrp3Lk03oJQuAOuD2sREmMG
x3EBuDrncpDNw8Z3eWgjPEhrqCLQP9lKrVNPjNlpcWWTsX4qqgbyfLFzxZ8lOGJ/4e+eIp8MtQdw
weAUonJcwfQfmgWDO2FQG88KBX5pP9zHY5CNa4J2ecP0lSZTZoyBGBsN26RRQglrAMPcShAOOgNH
kDn95BH7hL0uyyWTlKeefKfL83dqSU0+GE1O7oFiGwN1UrgWlAztbtrSU40HgDd997Qh0SmsvwWC
1J3lULbepkvWvPmkM3HwEGm07BSKcrmOJL8/Jm3fzaDdWpEtpXnTzUdi9V8RFt+aJvDLp0APS5wH
XiKG1Pv5zvkODo3VA8lgpNkyvCidMBvWD4j2aXTJaz8zwWViY3vrWD2CUnoE+pL9Zq/WR1DqyDA+
OHnvl1MVLZXumkWsSi1Fm49SzGWL8i6TfWbEMbvqGHE/QnajiEhhVldw5ukqoINuMh1w0LKg1Rsz
ZatXiKRK/+iLLaPosCsyXQlEsirTqaOY80QT9N/oC0cMd+jPBO7OymTO/pLvv6cdLvd51rXMa7vS
Pzy+iLezyrjFlogVuv8+TuGSzjJIpLtljG2lKY7OaXj7Bdbk4W1jhl2hAe35PT1Sce+gy9VZnsFw
Im6+ZBLjdlyrGj9tku9IcJFCfAZjfokWSnXNBSnjKOXG9uN0izMtTLLkb9XCd8pf/Wio684cqoKS
kcgawszX/p7elDANJJIJynz/Xg1kR9YAJAqnuLheDfNrv6Y26C0s7eqXnwDkMocnaBj+lu0dS4/b
Vep7RujRfHN7mTNFIjayycgYTIGgN4BfJhZTU1WV26LvIyp7h/ZysWw7v4XhCIm778BySSKzwUs8
+wgUI2u7DW0Sc68Ak54w+nkvTcr8ivD5B6FZ8t2NFluNdzFgxWU6X8NbXFrNuqSawCLGCqHgv4Mn
juojok1/1PloT2fWIzwhlttv7jXwStWZgAnSmwVJhd+K4tNwD2KKBihjpBMOmNuYM8+R9tQ7ZUZJ
tiLvdgWpI0hP1310jZgwQxMJOR83qpoTm6OsOdaKvbnxOpi3zwVtbLLJXAaZw5qQkR+bFTzLBYY9
he06MZMsGVb2w1EdmjT+JcxdrRuUXaB+mk3Vo37Yxu5CR/ZjxhJXrTQQJrQmBYvjKeSUSDoHWqK3
a32H9z/E9+xEhtXO94dgXVsBE374dyVx4bidtmFDY/9dijg/2TLSAFLBZgzDZSj4qZpZbcb0d1f1
QsUc1MEwaWPDYkxQ+HFkf8TI959MXzkjMHXrHamrP5UsdIQ5yO1nfu35J2xeBE6DiWLARm75dRlv
y8dGUhCJStMp95sDiuk04o1mwdNCJqyEOQGk+q7CTLupRq4rOb1L/+oX9zwWyETK8mfEE9JXEWwM
0nYANMF743/6OjqWSk9cLdb55AM9Sn2f/8Ttm9qv9XkNjQRIYhwIb/ONSfX4pNXlSHPrefhnSlEm
ivEhxxQ/DjLl3rp/uDBT32D4+ng06e6Qc5WWOlkaKvYH+ZwEs1NQgQcaC3amvfHDSWrZIyB6oIc5
82heHFLGgzyGQ5P4YN7aQ1Cql5oYCODZV8Qi68NpsnZL8pzeBV0o0WYEzBP7B9/H5XvJGYMN3Sux
ZfWCqLx0nXVtAbSfHLJ3lQVAH0Jmr64b8cWDqmdR+wWK24jxtSEQlfmUFrER4eubdL7QjMokj1WK
Cfue07SCEUFLp3O0CRFRo11Gf6pRzKOH5FSXRw/3OjSAXlrFcuxP9TO+iA5fSK21Flh3l65vkpKf
4YbEWM8m4+BVJ4xKdwIFegnMQbpxYtBv9H3prVp2yaRi1UDbLUe0LCKIk2Uef7fxBvijF4TVfoxW
/hR4FCbJGGzEwMWj+ml09Cs+gYQg+3QnVznr48lPzf5WrdFqvFZ5xpptizZ/GCDS+V4QmkrkQF8H
UKcZZvbz+jyqAe/WlMSOkmkkK25qr6E95n3EFPU2NEReJ7X3FTPi/AFSxBIJoWmDPmJzk2StvkkR
2FdakMyP8fwIdZ9zxPs8lmMcVJYEd6GcW5kCwQep8sdPEJaBvYnpV0X2p2UBCku1pKLB8JVLd1Ub
+xsnnCD0y67dIay83GgNBfe8vPVwYDEF3MgX66bpMaYZVGBM6C1/plwVm4LgQy/YvkN9YHR3530X
gnLkOzUGfUkhcieLR8Reyl+hzBI1stcbXqB7EzqKOW7XCG9QS105ksuKjrR6EYSjjbKFbltYHJj3
ZspuotFkrjwZyb3LRwTI6X6iuRWXdt+zuTB3y3GtiVrowL89cuPzcYdjZhu4CkBL4XtWN+kVM/VO
aQTBUgaR/uS44Ep2z7TBBonuk/XUEyPbXEkxZ8RFZTmLUjBj65cns15R5nWEzkFP1yerCUnQ8vDw
oPGAmbqX/TeYyX/BAnokqGPnLPmIpo26cf4kBhYzgW0/yzd2OnAI8SbTLSAmbbDhXNcowLjxLnDI
UE0ydtQgRj2WkCcxWjihfv1t/Z0wzCRrIoxWkOtWjaZtQOGACo14+4eOuD3vtiwHLMhd9oT6F5n1
58jmwG53+yzJu0l4aZ6C/oTKZAoYyNMjCuSNgoOXHIUBXiigtEr8clAGgU5XEYuaDWRSVEgg7W8R
D2zWRlU55gcN+iyDbiubYAHzfNJY6Oegh3/rm9YV1iooKDh33KU9Ii2LKHuzjEQu/F8Rm8fx4Ac/
uU3Aw2+6rqYjWwiG5kbrxJxaS6v0XETBKuJGLH4btUm9C8a5GmK4x56DA/SDAKYDNkbtpkX4we8T
DFoVgIwAmNdK33K7oCuFw+4YWKSZxAKCyDsXj3PmFoJa9OmTSdRNnr4M83gp7GEM0hqY2FE4xjBJ
STVZjttbW7NYyaICAPI0JsbX2Mby9Qr2QtEFUKvC8v41zRDolfHw4bC7nfbSqB3YSlssM0nsq60K
MYhbjqm0OpNidmh7X+EBKphhyeFxuBhRCdwSYDoTPuIPO1LAjEPXy4gUqfZmBw62aMUptlSYSxu5
IZ9fwggZgipiVKgeF0Y+fSH5qXFSQMcl3YE3xOIXFTxxQiS00x8hCUwjbXZcoDLYipzkfVwapAUQ
2PmRY98WTPgw80jdrCtkUc2+WT0il7zLXG7N89G+0nM5hwIceswQZw/Z/X9gBXN+6VhX2Mhrzmfu
CGL66uWL+C6O06YnbEfVSbYp3Kn/bs7AZVUY6UI1mEsLEqlMVqtao/r2A4lS1oRxOj3zcVSPRxLt
J3M9QGqGkUTpmMvSTFx2rF1uvnK/gbvyvQhH9gdtotFN4QXR59OEo7bX5YVXs/rcq6+DP/G3QPL0
o11ZvgLXBMfNV6zEoi9GxucOUknfX8chERc9PRfPimnd68CYu2LMT8NSflX9cCVY324aNoDZB5xW
sm8xNsDZZaGgNS8UE0LfOFSKuSJBmc2Cq6sGBrok+3S8J383BAZL+ucyXwp3XuMjlnNFRpQ/t/0t
ful6WsjfUzLOJsr7pQZN8CXKI4iHJHe29kz6CeFW9XPpvGywZW4PGM7rLGl8VX1OXEENdnLxy/hL
FAWypb9wsJ8mqbPDzNVyMJI1RMQ5BGWUwGo+FQpfhzJWOFT3xtnb1Pld/xWUng5oO6QBrt+gK1ha
VDsidbKu2Oc8IrCz5oy17HGGwAkvsU8DrnVZrJZlaEFMipYIRNuxEP2eQORLk34b3DwoGW/X45qY
SpuycV3oOgo3IyVjkpv+L2EZ6vDrWFAO+Dmzsfy4UYFmdDbPKxlQEqNruN02OPjA1XDJN1jm9DT4
eGWNur26c25jtgvuFkSEMspJSUr8lrne6yL0kmL253r2uSBnA6rsNKmcmPaeQLRetHGfwIMJy68Q
KsNsdBzilSOetP0mIup0578s9tJwExjVW2HqYFF5yk/8lt6Oi8eTGv2x7rqj+xZ7Icwo+cM/qr/p
KAHZBNdEF5SDCI0sL0NJ8+xO4WNyba0r29a05q5iq/JbHWoVGNs6UmeQDCftYbczwo6NHw5e1H5e
hr7+WvqemAAv5190OoYXeJe2E+L2Okfl27IkEqlTEcfZ+V6qJ1qN1B9voYo/gOqJ+eQqgsNKmzb4
Cxfd8vxSvoZUjAF9IwBLu2nWjd4O400L7K2ebiOkGmZ5NHkFhqdqKM3r9YQbcrrb86JnEGsj0abA
dPSrjjjBCrXCSfezXTnYsBC4KdnaC27OHlKS8+9JRGK8c6RQWh7b6aOSXq02kBELhLgk72CUPYQf
StzPcPVWytGXNepn3NUNkDbk4KpqiETc5TvNtJw63EiSltgXi8Rcu4+Hv95APBr5afIoVm4uhcZF
tIYjRuhsbNBaD3yQe5Hzce+SnSc2z/tLL7nUCrEOZs0uOyMVQXFe+DsPSJ6ssSjKoSrF1/uK/r+U
Nk/g1edakgB3EJE3KKUssGCAf5OznpkTX7PB3JeRhHHzndgpVb1lcKoqebaR9igLxzHKge4aufYg
3eLLe0hqXuEC2clbBBmKl/MxlnAtusI5PNh9R4Gpqy9zPW/HUzrpxkTiXFolpKIBIHrCLVgLrEXJ
hLsUm5n2w8815xlCHVc1Ns/XNR1iQlK70wXelB657nx2eFZD2w6i/0SpKd+iSvWGQ616aQKOSvoV
Kd74dJSbtuqY5extao0sA+eXHsBXSrGlhxAxBl3RGNmXR7UiSvFKxhpP/UORVNXyqQoYErFmRL5t
B021DmB98gseyk9FgfM1GumecRlZ55RWfOIRTSsA5IAaum/zPlXsdfvRW58BoAFxTes71Bcaxtyx
WWl2OqqpG1zAhq/gG7QkTlqLOhX6EfXWN7t+4hXQK73plrrTXG8oIoZvji1Ef6dk2Yey7+my9EDh
5WxDr58qKv+5pd/0zHP0Pi8u3iKdEtHxTiT+YYitCvdB8/mvHOFNZJMOunGA+2nibL36DBagzd/g
pVyAhBKe0g7Yz6mie3rylytKEx15LhsfYts6Ui9JrK551vXl9geNFFm1I/8CnH5wf+KZegStuqpj
FMTe++7DTTfP5L2pQJuIyaW1Cujk+Hv1QlqYtVIHFDCjBtDJFsMuov2EYdBGwDZUDmSxVBgxM8Tw
RBIWkUbH+wKY71TK/pNasEehXOS6+cOODPwBDyQIOFnj1IIt9xax5cjMcZdbO9swDLLNjWus2LMN
MTdU1vRdxkxxDCAbGvQDkGTxCpzor9eRChiUIMF+pR3SrsJfoYMDsl+/d+gmUSnaWW4FQYAd00a9
FHY7n3iDA1X9DR+C4s+UQe6mcqkRTHmqVxCIFd173nAeLrcyQSEf8Yz3u4ptMgqry3zoZo3W2Gg5
0WprTKrAbTJ3aLDeYKPKaylxN++zpxkzYuJLJtv9OODgsYIA4EdRMMSCqHMJkfKa3v3C3dDPKxKm
8igC8EgDXwISZuI1yNjDctr9h/sAwG2dUKL0NEXBmCGQCFKJE9oRL/AcPw9/E4A0jGrQHTy0nJ8O
YvQSgPm8aOg0AQugpT6jRch1AY2Pv6anrlz+FUhiABi764JUlvjiZVysihxd6uChPCxQ7nixVIFA
K1MBOpy+SFTXm+JL8HYJS2HKWmV92Oms/V0o6ZwYtZpOQV1Wz+L8BFCAJW9SQ+6yrtry+AtK2Nv5
JUUo6UPWkhOpNjHNC+XISnjRBVwl6rdcQuDy7kXeSQQTjNKrXtTDuG6RuKnyPIlmUYOLde75+2pO
oR62jjYApM5c+tqZg3ZnDf9WJlU46ZRqos/cwq6YRia06USK8vH5GVhejQ1wNt72KYNDYuKxPY6o
2wLA9dZ1FLsTsom0Yjg/L8IfnvG2dclYSIS3FqJ0DfEaKhHwp+WKIAbFnIgTDlmAeRue8KlIsc0D
GipMmKTtmwtmbQRzMbmhRAWutEBVCrdGsun+TikzqW4QqRpRw/azQeYBSs4OEfLNYJH17o6yQ+SC
ruP3o0TwfefKO9XayROHvjH1jcw0XKHIUVJg17ouCmmBg72mHYn/FVJRF7pfsqb91wOXitAQG4gw
54LPdvFK+BWRM0YIVtRLUQjo32fVW0HndQ8gSM0+JIkJ89tcHnaczZY9JD6PvnebCg1Y5px1RZjR
TFd5SkRDc5iSYnY6iluID4TBv6xl900Rq3Y+En4aHg6NxjE487QyPqJLOPJf1LaJhaiUNTU1tpLT
CU14O5QgAu2klVrbKxDqDAglhDd1ncXSwuJPj0KMmEEOnttxZWqR/57A4q6yTna0IAht2fJInmsz
JodetVl+av5nedu/nWVKmnTMbMvXBF2Mea3DRPlZpd9mVdis4Kr9A5Wv4IUg3AmTljLuKffUhLOn
RC6yThrTOkDK0xTd+bvsi/i/LkY5F7kxaXYUrwyaOsIe625/C76qjNI1nZaFpOTCZi5TPKPtIQk+
cQNbUJ3RjZL1TcwkAmUQIj7nCk1l/2yL0QYrr7+wJTlBbSO/WC5TZ3B32mWYcBJ/5ibrI9CcIY8X
Uf4fw0ZmP+jwbfmku0asAplbqQEN3iwh/0DnvWJ9qUfi0Cl3m9nGwHzYfZDkmy7ff+zaIe2pzDbV
qw+5B8jfIXXIvq8AGXsOJWuHPpl30NrFVvxrLRxD5hbmMSK/7jRq/B707Uh/Ja/wDXBUqUDU4u9h
SXm02gQIGxhzOhObvliYm2IgDNYc0C7LMUdOhmyQjsxEADCrMqtMHPNsjlrr75jVJuQuBJZJPGOB
OqlCUu/e7SIaSp2hzqZQJt45ebGcFYYL+MHOiMtWzbaB5IyRXauSflFsudr/ddxXCZnVePjRxu5g
Bhj8jIx6gl9+dvMjF2e+F/xox01FHBrTTeZhRBrpI+J55O+PqdiAdmEVc7McALsPshbbvGNCcKRk
ZGwqPo7aAImBmjmaLDd+ERUJlIU1wTsLXYpMRseQM1oPOiS73GK+hTI38GoDCclzzXyt4DRm9gUe
psAJ4S87GLHxvIlZjQ9v+vd1hG0COn+I1W04Z58IEHM/bltg9g2WMIBb9WSvxL8C0tjOh+u64WwM
H2gyFFPDYDXVwuiYkLQu4NNITv4lErhmzP/gi6vebDmTL0mXVhDjzIPl+AS388BrtQJqghNItnz9
50lIRDEwW36rpMxcTd/0HJpX9En4j/AY8fCkK/CuaD6sRyvtFSlvQIoQA8uVVwtnTO+kYLP3rZ5U
tYZqe8yXVA+e312Hbo3aQC2kDL0Hwd5rcAtuHNslu4QZAD27tomiy2qwD/xocl+IVXK/1zkzSnxR
XcmQcs8GQswweEk50ol+cojzCxvgzVoRVJaxI3ItUmTYqi8vY6clH8oJAPSnUEO/AuQujFhbDVGI
n6OFutZculHtMlKGLh8a65tDDOYGN2auB1gvqZo6YLCwxemyvwwkdB3Nu0HMtwx0V2ti7uDwbJKY
ITJlRsvV+c9Txhd7frfmeMX2l4aA3BP2An7aJpzHcN3aleo9lsB4WhKH+MdsCi7JjpCH0L6CROYh
MRycnwEaIdkqSV36zN4Tv0JJXjLTBLIYblBdIsaHkSLlt+XJuxBSRyvIMpDq+/gXhVJAGsbJ9wgh
UYK6z/kzUZA6vmQgAYssCMOE/svzcULw4TI2BmohFEzNQZa3dSKpjfjz41PW0TbWlRlXKf/OU28b
EHhQzJOG3RzeJ+HnbNu4r/Qc/wyAX+sUhnc+K5hy3vTiH+j55XTqociBOawpYEE8AUKH3J5g0AI/
3DSg5zXlkG2Se/DLGc0zzkOXyNUdIaCJSa0xDnPX2qMEt2dZWjQzWnlXEKurAzqIYoicRCzMmOT+
shGqod0Y2T6UTgJVjTifq+Jf+OdcTUYQhkcJHaQNOYkhFXDUPckgRMbh7uWwge/KWa0mbcFYohtf
gLIgFsk01J51zQijkf+xZIEKDnK84BQE1zuWVPcmllNcsgUsTQ6fZSqZuxS4Vism1q2Or06wH5vY
G4G6hoiwnn9mMhberFyJ27ptIin3KMY/ETQyI0tXlGAUAwYfqLSCXv9w0J/q985TweXxgZTWXcDD
SAAZqn4lyn8S7kdJ9r20bxFc8hlNn4E2qljIIeRl8eyU6OICJ7a6W9NNe1RYJSA28jdg4VCAOsQG
fAjox8cMB4RzPH+MiwcGlnRmJgxY/IYiTkj5nw4/egVVJctEHuyVwOfkk+hUxbrtlwmNMoeb65QT
Josc5uGG3BsiVRtxOzE0hr4w5P5l4kqqCxGz7yFg4CZkbqEMCv4Xpm9nHpAjpMtJUP9LvDmw2WD3
b6mEzABaa+KD+xg1MOqZzl2kSgg/hRWSTr1H/pzj3F9RfApzwXBxB8gdVDscO8RqK+GEeRfEw7Hg
aFFsEhaVRpo/nwBayy96i62Wd5Q/JDh3qt2sJ8p/mtUt/T+34Tv1r3NMv+bkK1ZC9nbN3rlm47KJ
2PtdjYOrw7LJs5nLpsuow7g5JMhAAxVQ7s0BNyKyWg6CFK1QkKrZkWtQ8gPVC1pZXUGCbzz3YqYw
r87caZYUhyIuXzuV7eKf3lglSlgLeEGG/tIzWxjBvTmAs6RV92VLbKWiAxClOPbdFLZuDtwUL3I+
KRaX9SZfxVPuxpk7vrzBetauID43sI64e5VyqWtGxWJ0nAIJRwBKXgzrkIKM8TJsFlaic/+fu4bt
dT6Y0D0KEwHc+ZokU7AFKF1dG2IZaEXXXJTq+dRrC1Xpwmukre4FP1p5hcFlDH/cQPvb/mEDN27b
QwvbdeNF7r2EULvoaHeY8989ITQ82wxIJZ1DRPULXtc8blGuuLKNCAL6nWeUU9xIjQL0zEsoqurY
RQO24f/am+Jg0Ob0YIgg2hM/1IJ+bgtBqRPGDKHhup4Vmhtd9VCk1U42Sm1cyp1ZKcbfV3snlm6w
o/20u7s203ccd1Etn4ULqyHelABVQSQeV9TyqNrfpE52j7c+RbVlhd7PUcBPaTbEWHPx5SH5ST0y
U443xv5EXkNMIfPxNHVZUD5DpilTBlcyfe5g5s5mGndftOSJ1eVFTWVfRipKKgAHrR3uqWpZJO4b
2ue1Z286HYtI6HK3d6yU4lZnza33F62MtbeJR1O3furRWsZNRy/e0SgG8T6v+AWmvr9jEb7Yd7Ij
sG4qKomVM6ufUKASoRbAJA8nXPabdJOWvEsAMQ+PlOaEovYWU7ulrsyzxKQIHZ5BU/k/+LJXAxTb
+1D/Fr9OnMEcuON7PmT0uN0332ON2bzYVAHKCcopRZLuYk+JGgFeZhG/G9bEKA+OWwGuwelqeLVB
kBPxbwuduNYmSfpG4bUr1X8hfMoo8waZk3fffqFYJizW/k1A2ApN1knuZqftIVmofbWMoyuwXAy2
ziPSAD7+keTwsBxnk2TR+YU34K6Xf9WBUXYwQ2K/6tJM6lwRX++6sn3HDxS5rMG4dqzdbspcgE3U
ysVJrZZeV0Q9UDGqOlvYp7LwOwu+RFPdFv4hpvZOgA/hae0JXLz4F4SULJ+gJjKiOJLjRE11qSel
3QQbkvoyGVKVYN4Pld0ARKq2JN7QLKxqV2Nq4DFcMdQimCrj8abIYjH/2mUA20L15v2UijKm8owV
e+FhWtHYmdqk3rjNuQy4hE9cYgvBT25NmcvktS+rGgWeuIhwEVe7+FbfkE7ulgIJsqXQ+rpd9NzB
p9t4DqWHn9oVQ4BnhnAFvp0UF9Vk7776u0u8f/3LGcBt2s7o5WyhpWKr5LwjPtZKqiduw9twznwg
K5+gsfdZHQHmkmr39LjskdnoZmyqAMHwTzICxuK4GHfj4/s5qKjO+tlLRM2Q9ai89IEHG8GD9K2E
Spn85DARLlYgJJ975hgvgQK5SEnqMI3P5OWb03LnG7gbSZalf6VjtiJpAPbdgYbJQrcjd68mVjOs
0VHxQfGizA3t0K/nmxE21wwGkvZtTRw2u9WH16CEgY+z747ia2rXjkabJomaYUVcEaFC39+Y6DVR
2nKXXSF3ZlTFAcuRRpLdOPbUiJVyApc/eA1EWr240XpkccITsFbCICoyjceT92uf4gB4sBAMQlLK
WKe4C8/sc3V/CQ6lm08rrRuUcKGRRtHXqk34UWrBdzDjuBTibNmyuUfKmZ3loL90+pzquUI6uOPo
zwYRzv6QX2ass0IOHBBTvJf/nJ0fGfuLPP5XZdOhU5h4Qzn8IGzWu76W5kt1gC2RT7lBWrgsvj8J
K4+HDSBDdAxUKGzHdEOUdZ714iNXoXs442h3ihCWC/A/O9LVQZ3pPrW3O0FSckzyaoh1yErIuzky
GJ7GMfx2ZZ70to42Q1Ff1jYS/wkxxOqx8udp0Tc+1+ZjxLqrqBgRgJ6E2hewSIp4P+L0cJskga0a
F1H9rjg01INQN1w3CQqqyI/o9xF/blAPK9CsvUMJYtLGBMNgKTkc5/BuyffA3lJMd3vp5nyFNhSs
xjG/v21GJAKeJvg9G90l+l/wpYV7ZrVRqzezXvCTMw6DJtB8EVVhvsMd66xNcY5gQdXjKuSMaShP
rtbcLFRmnZwR9KTHYl5//bzHaYlkgedRaLChekc+3j9+xXQXwcRJa7OEAw2xYkVm8h6gF3P6N7TX
6wjigguGj4X6n7XU429QoyPGTfr4IaqSDyH2kLBsEeiNKdEUirJKBkY4qFrk0UhX9UO1rQn+U867
fpC94XP0GOtoPDoR7WiFqayCQOEdrsO7UraG3YPD97h3QA+xXzHvld93IweDSvLOTmj1OVM12TRs
YW46p8/9+FRp098RTvVGZH/yEwQQcm5Np+6Hc/2HxmB73z1TtbIksT+slXO1nwFJVjfMPKFUXCr8
DBrKrkfrR7hAUUpv5BEmDzOu0bGC0JkCYfYotemBPcm/kcbbwce88Na5DF2qvz+yKy84peTSc9SL
8giVdPn5xJqEjODZFQEvzbJqVm1xIKsM70p51CN2YIc/jHUcGM2JU/hRPYFrPijZmfKbyxfD05dJ
GXKGVj0Z6f2yffu+nuY871/KmDgNIZljAflaj3ZgHDgO80fb5pkM9u9eOiwuI3CsFbRYBQgTh7nx
wYNjY7m9pMKU+WCoNTzEu9uGeV2yQxba6C3S2rN4IDkXNYSj+wxBuS01nv4azkCoukQaG9xa9XZ6
avJYni7yWsde6rfuCelgbsgVQBqtbECPUPE4ml/sD7+XAw8wM3P/xZZU5zHABKuuFAzlgiHAbvNl
u3cYhDpUOzyqF3AauhmU7DOswRtePoN7Xgae/mOG0Bl5+eth1EldYRhqaoqDXLyjcAGv0jCr9O5p
WeoKmcb0qpVfKpf6mi82KUh7sRF0J459SFhXsHc68J6O6GQ0xaHBQUzMg+a3WkRqkY9OfK+62b5m
yo/Fb2xaXSymg83aWvU9W6HzRA8A5Pbb4mwzAqOU1oYZeYsZyQ7rvwv+lhCQc5xAsmljMX1cm5YB
AJgHf9bx1u0kbCrjr85TQN8/mFLQh9/BU2vJpfG2qD1fRoIFQ6D9cZe5aJQbnvkp/hTLevKK0fLZ
amJeJ0CzTLJz/eNGgSd4ezREMSauo+fcf8sujRCdANNtwCwb924kunfucNiOrtEAfn+9rXmHXe6E
n2YvqtlFPJBmdp6kV9VRdXueTy3gP/TvSiWr13Q9E0+gbpn7m/9fKi0O3Mq7xqj7KYnFF2zjNPMV
xLMyHKwiESmjk697WaNLRF5El43fgwDe4aPH3q324QwX7pV6Amn3SP1xxB4vhTYoqRPjMuQm2CGl
VN3ZUPO989BM37gSEalEn2oTNVXbAKodLjQm8OO+/FhX3ArjcRQX280Jo65DOEQlfB3GFAgDOnRo
BXV4Aig2cqGye4BmZr5HpdT4u9OkNWWdwY73lUzaUScQR/xZfMKdPe+pvnRIFEJMDtoTo93MZ1bL
WINcFnxTrquUyokGp8W6VaSAfCjGa1BXSfYegoeVSLwgsrxfxt1Wg3DQrDDT98t/C/a9Ivza0R5E
suW9l6GzApbIpUlpS2DXEAycu5UjTGDoQpobx2mM8UxBj/N+zIildOKNV4J7DRvp93fIU4rzueTg
IcM6p2zSL8w+WOWVlPTd9Qfr6vF8Ny0tydUF7Ex6ibUJkGwmf8v35HIaxp7X2l5c9XLaSdwj4gxe
iyccejr8YN2fOi/U7kNBP6zI3cEsp4Dz8GiiSLaerTzfvZWDck0krbddjU6Acg01a/NeqSElUZA0
2dHWUCgdYdR2k8tkCd0UitgLNDopw5mLc+j1hiKI2e9kD1Xp8SwRV27Iba1f0Pk9lMV9sr6NoKii
cVfISn/VEv5QYcNMNOIfLRd+CMomOW1UfWKxbz9Qs18o3Hlh/OWzacigocfiGyXn4o4HwMR6zpQX
za3c4eNpt15fdkoRthXeQVdUl/3nGnuQHUhETRsF+s689k1qVrSWwzQ2z7ldW74og4UrDLiJ1WcN
zt8rRi+byPu3bhvX7PcUM7Dt40PUMsmPgls7nvQUCkEZ28F0rAo8ZjkcDMRLxwvOzHuOKGbwfVZ/
OyfnR+CqR3RWFdOm2nyrG4LGpj8gHCEuA3u3ZCCzPiPANLbNAZV0D+etVgS/I3fKukpySlWr6ty5
xXWJNqwq2ZuAp5jGhHk96BZrlZnRdlPSrfrLUEe0BZwm2OjZR9BfsPNeHQfBo4iIU62yx2gFToUx
rdxHopjzsLxVC0zzIJlJiMLMt2xpIJVR5TDblv+0fMEnL68MlZI1ZAhdzcTb9Uz9c6omiseYtcrC
9oNOoi19RBIH1hZ12NN4qIMKfDywbHXFzTyTETa6gNg9AM7bddQu4k+zoidaR7xS5J+CgXEqjGNh
N696hpirFp3scf+wP68gNh2p92dbnUoUIZnpxEGhuw3GfehxObxHC+8VP9arrsmIKWTRo0GNdUi8
p/kKIP96wsNn4oolARDG5oFdyyi4ejCn21Jf9vRYxIJVf4apagX72KWXyN9AX7o9D3Z77sGB10rq
YIadMwcG8Rq19DEmHvC+WJ4/lPMl4a4qzw4Jz2kZnJlQLjhztAO+1lmWJ3117VAks0cLJXC76Axb
qgPkPqmHP1V0+Lfp1bOev9LDwGszzcagG1WJ27xy2E/heE9BhCQvegFLh57jyvVxWizzE3XiOqQ1
5S65wiH2tcHoo4J2sd4bBhC+pwVrFxN+3KxCFAb7hF4pd44sTHCvKXOkGeNOGyJmpJtNrVIaAjJT
MSnE8oXhlquSDH+J9w7bOoHrFESzw/QH2dinC0KMJfW5az4jg+EIFoPjpPoty632NsnTOuWlsFM/
2e1nT1s5H1kARN2t8oIWsnTcU4h1QGVj6Ysi832iLEal2QZcOVoAF0x5UY2X7Z1zf892lWSocP26
yfBKt+I7rv5dbRmZi3HIRY8sTsfntqWF17DCqbi6PYWPx62fixfR8T+hhgaOYz4nsojG5mHHoiFs
I+8ncNIVTgFE6UC8YRe/4ZjJKFbw309H8I2mVCJe+aaV3rh+8Yr4VKeJbMe7yMQv9QsXOv3VhRTh
XTJ7mSR+uRy94ZAqMBUFePIs+7TdMirARA8oT5FjeovcqfYDOZVdL+qnt/XJWzh2hQpLhuzNRcU3
Uq36vo79uIqU67bUhbVQtfNSGDm67PO98jOAMgk+vJyq2HdUn29gG2WEhVPwUpaSslTDmRZ7O9HI
/L+hca3HL0I4wEYRsMRv3BxTwh6ClnxSaCERQIivUdieP/EWWNffsUwGE5qNeM0rWaGcw5a/aA9O
3fWXIrjzOSRmiwrwUeAieJLT62LAXLSxYOw43KE7N9nRG7+co2+RvneuSd6wmK7N+5L/xwGS8Z7r
a0vHXUACMomc5jTOrRyE/TpAZtSlAaOb9gj53JsTDxLvX0NZAP1WWu3sBP+8CV2I4ekabc5mb/4S
uXVVrqCMJ96M27znJjIdxbgkhKlUHfSYpTykVhQHwuuh1hj0TwRexbXQ09rQOO9vYFFK/aIGl9fn
rhtGZlmIXWCU7sCJQ2xGItus9a0pHpAogrGDInJtz2pgKNn+Hryw+JpceTShQW1OfBVyfsqE1uiC
22XfSOqaRSmu2EGPUHKNH4b/PKoysgm+FTpmHuOa0B43DOTHSN8PD37GShhV8WqV/Z7gj1Vvjmx7
11J5XVtyiKLoh4F/4chO5lCUjUVackUK/HVAaOtk0t3iXhKROZvKAJtHsPuY2av/eyiLJAvtNhxb
fPyYrGq0oF3Sl/sh+HkeYLAX4ZbhNjPSebYEjAqrIkw++DD/yWYYUVu3R3234uJ0clFO0ReSY5vL
D1BnAXGxLnTs2Wby8acP0RqhCPXoZUYmdevpdFCD0Ft8NEUHtiJzc5ghTlifOdzzhLB0eiiQXDYh
XwVVRdEdZwSFx5dOJGSbpXqQKkNQEWZ9GJSrC8dBz69N9lWJQhQFox/p36NEGePgJ+cliU87m59B
qOutqJsVjVDLfnDu4i7JNo7ICEy/m5NELYvwyKjj67Guhym5wT3eylgy8sewbR5/UysdvLXa0joO
VYCEkbbehe1iSx/i2W3B0bNulBlUk1cgIkmbhs6WzRgjTHlbur7ubWJrlfblYE75RpreFr1jc+Ik
s3NMClX1ZL/Oumt4Tbw8oZL/Uq2N+HeRAgejnSn6OCAqGCSqGd51aK07FKS3+qIIkoTPw9OkEl7U
UFKfw3q9ByztcoqZrmHtSDMaSW+DO9nInNZ3EUgSVvKkqBTtP+ZH4vHBFgWe10L5+PVDrLP2DJ7B
keQGD+1pfL4H08F0XdLXy9zQ673nKdTNtJEB69fssxP7CuKddNKL6AdTR/3Hte3yCagFhOjWNaKG
yLGVyWpu5sQk5vUrj7Qfezngp/6ObnbQgE66VzuSbcCB6MTW+ANey1FXQb1pBZCHOyvuZTa+ngdm
7dihOR3c+YwczmdOmW5zv9QNdojgBxHCo90FY4IJ1CoW7lVe0wOfv9QGV6fxg7bVT4Ic1fXDR38o
YVwZ05aOGANNKh0SFmcULtv4jhJ1Ed+bBTju3Q7ATdY+Dk6FyOCqergtxDNTN/cfAi3ch1m3OD3C
0ECFQOsX9cJsqYzwUapPNcmY03YTqEFCbVwC9RAypdZzOtXgaFfcywwZRyC9CMXmoTcIzbXYj4Lg
gRR1d6oC6T6fEi+n7JrNBvZVLNWiuAiT5bGu7U6GII42dVcCkKn0rLG9f5dKiSDJBX5ACCWGQMWo
+ZZ6WxSSU8mz9UsFCBN5wmspIj8Z7ismLVZKh4iSyxOir8SwG4w27sg81rrUbdS6DDebFVLzJVX4
/3JOZFCxYu+XtstvJlxL18tDRW0GfZpfB/JvyO7c9RtZ8JGMr2tZxNDDhtfAsqz69aBcH1r1zJbZ
4eUF54Zq5DsPF/DlLVkUST3kP1KNYeIpyD8AG2xAhlRJYhnwjac67B4TY05/M4qrPckormljdKnZ
bo4dsEfFajARghwrsXCXOM04Grhk9e6M5p1m4kagUE4ere3T1mXeC7YpSUoEJXSDxTshaMUEEgBi
5cGNtlqLCgpbXcXHxPUdS1rTCryxm5ble502GR03gWlpNjjP+kG0yT4N4G4QgxNV5uPcbO92ZfMH
s+TS5ul4kfXdp9gSPtongs8CKbesMPjRuYQphCFAQdxoaTqNU+IiRZxznAV59WIzX8c3/rVNjKxm
8ghINqOFEQ6GpxDPBCX+TRyvbhfcozAtfyBP7sw3Ez5I+NXq7C5PZJEN9Rzhz7rrghTywNYLkJGQ
5U1SHmalUk870aynQuV+0guvHkyI1SNZWjK5vN0mFgXfg70Zzo8hbqzzKv+aYZQdHhNcXPXn3Gkn
73CjoS6xdmFJxXwaFbz+S+odi+nlvI6wavk4wb+pSyb5/YJZJ3Em1xRFSf54EfiAbYmwhAUuWFoo
k2XNjjnTSW4qW+xoA28IvNN1UlMCgOGv+KI+QImJHu+2Rv8fP52UGq1/qSU3s2EuZ6evD6qjWbD3
FwH1XG7z6g3CDOhpRD2p8IZMG1wlOI4yMfYQEvN3X52T8pcV2OEPvMRNzH3r67DYjRhYMD8wR8vG
qz8BjYqbxQ84iamvpNF9VS8vTV5mS+j42jtsBvbK2rkJI7Lgz0cSeJFCa7YUbw+8zpe3u9Ix4zzt
j7CE9v9uEa2rCNbYXK9FKd+t4wyDTUEm94TQ4aLslXjIViHOkDwBbI1Eo0NVUg91NV50SeQ2kXMA
1snHxvfXE9SJoALH0XyBCxOPMPDfv6x1UORNXkIVksEuRNkx6dX87KaDQVW+AmxaYp2vTpn4ItP+
jLg3KLcmS07T9kV/+EQ5XQ7hfDA0wc2I9M8041AMpVwjZd6h+TnPe4r7v5WPrTrpVHcrh05q2dSY
TLGW3X6EQBNQTA21Yl70zUcDxqIKOOc8/+gLH6rvBYYeW2fd9Is9IUFKFiG4q+/SyElFVTFQ2A9y
fFHE/FKDGhiCMY0J6+hxgaufab4H3nc8cVyDczk94Gaz3GGQ0MCu7iZ/LGCN1omzIJDPKfrElXLv
UKAvH3BYwahzwKpAwFsTtka66YeVbdI9dH23Xo40fba6GBZIMiRWJlIA7KqfZQa/EQn/LjftyTAF
UJkeClmBtH0OSvZwk+3Ku37OhjLV3dDfTV4Mke1Jj+TAumv1BM/ZMFUB6eT3eyhI2QLw4XCpi51/
SPSEZCNpRWtyqPb0bWo0gghiouHCqt1cIxHbaabdu+ivjX+EwNwnGLx4fxLb6r7gaA8WBuIenNVv
icNHC8Q/xcrL3eu3it6qNWqJdohTJyYY8n95hmg9I2e+8hZx4SQ11hyKn+Tz9dX2JAs92LbYYp0t
81o9TxWshF9S6MEBYe5JS8kwigbDjva5nbzNYzfoL+8Z7JFabaQNsbqc2FbzzjUHQXQC8Jus2B5X
qbrqeJPSkv/BSI6FKw3jCISVCMlahHRfTVqB3mQud5eOUhFqIB34+m8kIUkaL+GW+cWN3Ujz5II/
9+MisT1ocmdkhAFyvoIWC3ZY4GRdUPF9IG2GUtw8S5Rz+qMmDA56KRjCBOg8NhH2SSL8Fc0+TkoR
Y2xUtnOBT9c+7cb5WdY34gUV7MUrODjPYE+o99WMV4NWn8c/aY/pXuSkf4iv6HvS9ysVvcyN1YmY
2+T0dOPUp0UG3QFi+y8aTHsST5XZgltTiRgrVyfafeg+q0qXhNXQScos9Y8Vld9oGUpH4sg1KWl5
z3aOx31BTvBWARgjsL3JfKYJwWeuvf+0sVZSTzFZjPYsOYfiE8v46VbN7xmSKbIHB8WV872UTMYz
lCkweMzgqUDcjQWiPnCHvQ6JA/l7ZrF2wRvsR4aGDRwtMczpszssF5N5Mwzab4+h0/LenZnxBtqX
gVkIUwr1rjtA5IiIuHGOlksWS/nHrQvHSoye3uFTcYxYYsOFOSo8fdRXw7EvxyYcVo+GIyi8t7xL
mMqOCDsfi5AiNzWWoUvAO+ukNVhPAaZD1mIxdYzoviuEBflukLu4egYWbPwbZ1SYlh+WGKFN92nI
TdRR2I1L7I2/74M8o93wb12BO2WM/qMe1HF7rdnKVpHRAHSlmP2z7hgUJ7Vb1QL5g04fsJ0sPcCE
CzetStJnYwhAYUPrVeWCPJhBFjxkAzCIOrS0VGFS4D4PifCgqnKZcgl4gPOOZtNkyaKpZnitgXPf
xzjGgzC99osl9MFNWeD2bNWbCmS4WJASK4ONQUD+kpzpQ9yjI5pJo7yGL+x0pNsfVGpcOR69IeEX
uGL4AKsGJou8/fTHXdXFcXDP4UjkSLNaa2NLVPFlEtPzffYZmNu6y+sNxD70WvUXXLxEfg+YtzPg
aT58ZhWZmOFe0w4DsjnFJ6Os49Ghzzlfi1nqm14sD2dm7WUpXmSjkvNAgPXHNujzR9YFPWxExaAg
x2NF2rCd6VjFFwQbYoTj9o07AEvHe4E2VFombRk7BTBDwiTVz5lUoFqJIN4yZ8u/9f0/AuPUt2+f
CxSUnYbKQ6+XO7m5tbL0uo0ONJuWIiEUVNQ4vp9B9QzdIExfwgGaGC3s9z5CLIzHAFEQlJ8q0dd/
/Gg2S4XmEPZzSzYGEW1PkIG+Ua/sTA7r7KaBnMSuvWnR1Tu5ihWytLpPBWcSZk+oL2ztaK4+gJ9e
We2+hJxpuN23FvBojmzCrSRfrb9glHAdkpi4gn92frx/9CzpAVTZrLtQcdRAQEfSiLpKEICvG5AS
+E8C1vvtCApTmJLCV1zEEiq+NwTtA4zLYYtlkhuIqceVMMEXIoBE1MIDMk4qICJmw+XIoApUIMXv
7GgAh7dxGQNl5lvfm6vLBJiJd257ipLaCari63TZ4VKZJc2VfVMEV2XI3DSV989ERISM8SCNoUsH
sG3HXCD7nhIQsr+12L9Y8d8djeN6Z1TEUrNfTghnWidSkOCmUfoJzwzN7kYX+ZSHd46q4B/ewqjb
FSUbXia2/nZmJOnKeAFz/ywwLhZEJ+8pUafCFS0YBb32kXnTSsW7id2h5QsdyqJYMlULUf0+VmX/
gI9LBZEA00Dic+FbtCq968pp3/wroJfwsaemYxEmDXNGVukeXCH54eCyM6udixdI9O6nhN1FL2mO
Xai8dn6FuNIQ2JvA630tMj+7glwjsFq88bov+XM9a6t13mE+7mUfWBsEbN21V7Wj71MUhGn/iaJ/
KJsp24UXsvpS0mJ/N4yE104C0NPYgo82VgIKMGDioyZ8yK5YueAuLxicAEN2axvhLLtvRyIpkQ41
t1N8ziRTqO1JDW5bMXZ1gDYMeQuyJIvmMZ/tfh8duyxd97CZMoNPvCK6KGEfOF2D4SmU4BtUhiBz
ZzRh1RkHyuRr6jINs8i8AH4+YOogn68Rsksn/S+72BBae1rcM+Yc7eVeBw3cyyGejEPFVb+1z/zL
pkB0Vc/rWS3kZmqnkQCbAUHsdI/WPMm7ntpoJTHATc75t0GI8EuTIMJvSa5v1FLsDGLv/KkbdWyU
5HyoAKpeetiY4DdxvmGT4kveaOqR6tCQxuOKlEovZFxFO0kmvya8iJOXXstMQo98goG+xfkSBhVP
he59OBdX1cwtkPTa4jeQkMeTIud1Jd6qK33OefRvtjHVoEzhugesU2jv6m2Ix86tjtXYoWM4lQB5
RTazzzQQLixm9/b/DTH5c0sDggdMuGjzz94mrqkkfFQhL8LXACay2GwE9Z/lH8o2LB3wprrfNOQK
iF0KwNoqTQQ5hyqpYuv2f8Q7d/mgK5z9FAaXOqxYlokiHUgu9VkR+ZPsK/V74tIDgx94qknaKeMC
Eor02Zp9dPkSBcnBCISktH2OzsY2QfRMV2vZ+jo5Oc29uFX5HGutNCN8QfJtxqpeqzVsLDpvzB7B
Icr8DJVoC3fBWOnQoCaj7/I5A9M+vMrAFkmOpfcfMjKTP7cL0nD+wragXaSU95hHqMHaaMRHBkOq
AhdIjawp8z5uBrT/zQIL7SCmoTN6qRGfH/w1s71wRfWiiirLdEs5O+ehmSpnN2e2UBo6Ix5sr3Ho
0CkVW+xcClxwtYBvjBfe5hmEqGClesBuNIpEXMgtZ2tmYBMcGtW/easHLG0hR+uyVo0dOAXek+sq
s6EgjkLbJ5HioHU2/ZoWOo/Wt7qHQU0OEg8tooJSqAS8Ojbk+DI2Wrr7g6c2R7+7n5SzUvWHFoxW
rmoh5V1aeIz8LTvqgss1lTrm+kagclGUB0VSby/ZdqM8nt55vI8JCLIXfl3UxdJbk1ibhXiaGNkt
p0VO1rGf1pqmgOeURfMLjRrnzdk99Kq8a7oFsrIenhZeq2an+cPd0BI5MTIZ5UqRqouMw/8rgigA
F9SWYyLDmokEvXGAUXXVDf8ZAi8lFxFmwNmUKUVfrTqkZL2u0KHoWMthEE0YJfrdJILrC1eEBOuY
FrD/3uIcd0HuMQl9mp82M4rEu7gbHiWldEgooiaV/dXCiz7Y6OgNxHmrpWlhZw/3dPeXG0LR8RSJ
SZASiZbXUyMQxr1yQ0+ikiCqMFLuUgaQBpBeKEWAG8rT9vua8YoQq5EhJyhzhj0NPH99jEimAz3l
n5fflT6pCrdV0oIye1PRZAXwMhWVw9wjRmpbPcFjDRTWTnwJ88zLpUgBxNxrGt1YI3nhAEe8mgV2
jirtQHM0rc1sU52F+1Ejkub9hORzTRbHndUVmIYbqVXJ/DTnm3Zk1UBNK+z0ICdNg63Q/xrpM01V
IXLmL1c9tevFSbi60LToYFUe39ppBmT4O9qEYl808CzGhdOex4yGr2uq7alMb7pZL0+Bg7DbOmiW
MvPAWPudhjRchwp1daR0Q/vRBF+8GrGdYUN8D/jNiBoUS7FCAPFk8LJq1pbLkTXPxRq4uTvpgcXv
aA/Sq/Q32niCRcJ/InSsikBnumUkqKADDAmQpkApcWmBcbB3s5LWl44RQcRm268vckojkK/p8V4q
PYIsN//6L287iHxFuzqKamcw4fJ+GutbC39yA5+k/B/d+gFDSeV4iXZwiediqKjLQIlHO65f10vT
+xledGtiDDaIl7FXGJMzXD+S0YMP3pHpH4XZV9dqbFzK7JVqsgOvoHK4m9/Eq4ZHoja8ExPAgGrF
3LIQ2nxZVGevdrGM/OA9ohduCtTi5SLLZWUPOv/x0n8MejQzGQIrSXLxH+/fqbft09CqUwD4SHJ5
+cBkvMCdulH2FVp9BT5uwEr0mlpfqlMiwwOQFI/XwygqQ6rBEJwVr/NaJzbE80GfB7LblAzAYmZ9
4tlPF78nhglTdzpCxDaoinJ+PP+CHlXRrMEXiU2ToSc3nJyK54vgiMkI+Pgu8n84v31k/ExJpVuL
XtgBSTOGsAnrBFTKGC9sodlGy6bT1aHoyaSnght0kXftHCgHpazZ1NG4bFbF4q6qdA/8BbAiU9NW
WyjaB6MlOUUlOsRE8uivCkJbRrD+qApgwXyRRvJ4hGntJfdobFTwSsQi/2J40mMqYJThFFNhOYOp
U20DTBYw/PEWAHvmZ0p437IiWNjpVnGuvJfmjSbJr4lUyDy2DqFTdfr0FAShiqI5CUM45oI6wL4S
qzsFTdf4hFCF+7O2d5S9RpQr2qTI/s1fyCAjUJKw1yJjWTPr1yTqiJ26TM9D2KguTfiZstQOXTUL
zrRoXv9W3agm+bAqKxgt9phUMrjbb0ozylhSrahWTylgnmJPP1eP/AsZS7IvkPt2UXMLDn0PEH06
xPy35ExHD5iXERgmigFUl9cjisePwWyjBk7uJO9EfY6hzuWzFTNjKq7SYjGJ3V5gd3i2mYZL0YOi
28ExyLrxTtxSC4CR3EVdxyunL5hjN6TMH0XYXlChRY3l/9nXSjGoW2A6e3iUUd2LvLPFyotr6Q5l
q3Ry0i/Hvp1xs6Pvf3LG/VgzzY2FgCfOa6xUb4HTllwQK9aZlytOxbASok8E3m8GNEBAI4kU+2wJ
/gg7wi4JIKffn30cKK7e3jSKKePnRKN+2TSXzYY3waxSKYdLNqjAKdicF2O7XMuRCqOSUXTVc3xD
Jcu6osoIRHyYFvQVh3iZAE8P35xZ6OZt8KadvXIUNfA3wDtHVI13Kw5/DSBARXvp29jYVaaPri/A
oiZCDtsmCpTwr8osbdXJeS7/m+ZaL/vH+BU8RBh22QQck83d+Wq8jWTQcsKDDmDdkpiz0PrLZU52
jbEjKe/Hyeq4KHhN1MTxUCvi/xeYuc5l7+S1ms6Nfsq0tWf6KRp6TBdSNt1i+NKKlwaQ+ljfTmUt
Cx33OgtdSXYFkyQA49pZp7nhHXCEfIF/Ne5ZLz0/d7qOeYVMAlVm9wStD+aiM8caKuwAjW3k315G
eXxbVNGMk9M6+dWc3jmsO96Ai7tZ+4/rMo7Qd6ihbxUgsh/RGKJH9UJvsqz6kcKkixF62GpEBlMZ
GheEKUOQgA5lPNT2yqSQcGZNVJ/R66odOV4Sd2X0zGo9zwTZoeW85QvgAhKLvks3r8ymJCIi984l
OsvItkBHTorQfO88xD0Xz4dRI4cynz2VsLlIdPgo+O1LZVL8HYBa/6GKZwVFZcyonn9VxsoCfHru
b5ITHWpVAojojCB228O+xf/v3OkOiDiarqutRI7CBqe0wdoflgLccgwtLykzR5BCxhqLYveABTP1
YRKqN3wwkiycR/el22k/Zbdm4HsPwqGxx5FvsGc3rQiab52bODykvJtQ/h0zz3iKUZCOV5R47LiH
ScWolpxMGpZxfozwxD0TqomLQdN7JSwaEKy+ZMPeqs8lD+XqQNSGBvFhYMKra1JvbUtPO3PauHlv
KyQXjsMUo3rO9pR3b3bHJ7OdNE4OBYMiPsFupSg7YXUZT5Uu4e4f0+cwyBokEBUwgudtgZmLzs4W
7mu6UhwJz3XJOXmh01fYhvPd2TgW/DlQ1A7oX5Rc2simqvWa71RkA9+SvyNCJ1bN3qAfWxSgEqpx
3Z4WRcaC+MHCFDqz8CCOWR+m5Sj8q5ayOnT7PHgwBCzYvb50RsDrnAxcMYFn7ic7d0Djw7Ykd4xr
zReAAFeAtDuqDQAsbiPMK/AR4whZMfPNLH4J7LAcQcQ7BIpI8sKbMP4+N0EI0RUnQVv0880T4t5K
aeBqckKFGfA6gIMNFz9aKGZo2unlVsUCb6vSWV5UkoMlH114GlCacTDbjTw2ettCA2+dMIgk+Ak7
GjFzGI37ClwtRUS6S753T1PPIKr5MK7LnbTs98ki3wP61SAq9EIYat96RQapJxAfhd+ltnNK3hmP
mrHYQsHLBmWxBZ+kVTYZkS7me6u6WxqFmbTEJDCT/+dYAcT4HB14E657QzjWXktWmRO4Ec8ohjLX
CMlVvVSbG8oCRT5725lIBjh4yyiFNn6eqRD71zA/+QIGAQ9nDWLfgdjT/KlURQrxMBJSZMYg0uue
3xE28mIQ48Z9LxElrnhx/b5i2Tm7YNvJu2FE4+S4Js7eer6Qma1ipwb3OsUROU3D3E5yq/FDboS/
UH3VWeXOl0ABs1fcm+LLIMXyQD6uljOmoMBbXeMFCtv0bSsZnOY+JasFznt3W9SI/aZN6lcLkGHh
udDvmyapiUbV+DpfhlhnHPwTcJZX2YVOSFX0pwPjpiTvjFlNgg3nLyljUTL7Gy30bLoehk/yfvmt
11hYNIgeYvS9Bm4hAymsHgIuKPthbPAGSyCzhvvM437ByCeEARLABpTKdKQI3ZWccEevbII30Qch
K9Jr8gFpWP1K5N6jyfnhtkBz/2FXJYDTd/I+lGJuoahQ9rEMrEUfSKEopB/X4qkx6iT5YHDwPh/9
yCRbS6Xo4meSWPRSj5029Xr8m1+yyvMXMAB87tucGEHnxCK4PwWRXiJ3VFDzBpBAG3lL6AoqLewk
//QXIyrU1nsWbi+iK2XprRPi/+f497FUzcLZbH305+STx4RFrgRNtSTEcudPfQk4WPekg130MZaa
91BJO/F5hDev/oHhr03qvVd9QONl02iFxprRgL0ogVOlHHli0/ya7CSRY3PrYkL3XijDyfOSXmJ8
xTFHTeAl+oSKqlyCEM2WoSa85x3goIgn8zkY9wHIxRS+rxjtUxCmyN/D/T51+I7yQY845NSgRMpX
IHzvHrjx/7GFSJ+YMr9FG68WBGPlgvXFdJO+VSmEu2MLC6TwbaIx7vKpkW5FBuK3rkVs3iudQrFK
RJf4HfkF7kv82UTXbCwGLrjeZJeOLLUk5+dxdHA60t123xlilQb4yG8vWLC61a50jxnUe+Oua6IT
nrM12CRMDsOVxNbhhiieCEfhQt2AgruDPZQdlomUTEEIyAwqxNok4fyy2Ow4BvMUjZ8XTbcS/eiq
q4yE1mXRVmr6IZrmMzCF5PKIY/ORTadaJ9WLa6EPCzVzyxT11uIJZG+djslWO4Ll1ETNFLYgiuPQ
+KdkaV53t4XIckCZZ/YDZg6geNk7k3FJzUyguzwvaM9u6ZXqf63wa6ESnliTmQuYsfx+h/QVmMu8
FbCAC2Qyvhuj2GEfwo1/bzMTMUC2nL1FYQ9hKoS77+qy6Ij2fQpC5PoLdnMRFEoR60EUGjcWig/C
6pGjdVCYal+pyS34pm+bZRXu311Hxs+vf11djMPQgnkbKbpQD2ZP6sE5BFxpNYUWE5GwR2vWzwcK
n7YS/P1Z85ymBrphk0BnfW6q2zpVVoFQqVar/nM02YZOXQqbwnvrCFftpJtlc5Ri0WFddQDeQSa8
m9GpoBaIEslQS02XlN4T8uwFe+hdiEc5WLnCvLtyG+suC0ffwj0M4aYuIADSHwPQ0p6UVhOJC5uF
0C15qfyLcsqvSYrGfZ/GeDC+Q8qBW7LtIIHPIylOflxyJb+fOnhpNF6Zj2wGViXMUEzXC33+xxB0
IUEO3ZZX/k3pjpsuP5ZRg4tK4QIMNPdt3X9K1Evi5uJHZrmeyO7skU4ZGfNiB+T/sgcarQOcCuMK
yu6db19q0esPc6m22vF2Q0VlsU+Mp4JF8pOaszoGi93UmMH0SZux3pO6ysACB3/zMv6dpaadcR/o
tvbkLCLKlkqLfN1T2Th9rBvjjh1PcMhhRygNwk63gbXSnVvIsjtgVTOW3aTiftx629O0Yl8V3yrz
a+4uC3lPVnQVqBkduEb7s+WkS0PI38tAureqQndwdLJoez24+XMM6vAEJZ2uKUSeJJbVWr2Wn2zM
ueiSmneK6Dq+1JXnHul//W5SfE8SqRM+XadmLiv8NffITCqN1gZ2z6LzEVgetfqfDDyV6QrKcEGw
2D1ClAD5SsrusdLG1JkDakcnB52chvoQPri7MIYNMIsSWM83Xk3DOF9iWupVdL3KsYGGisGyVYeB
06G+Tyvfv4d9VBSpkTHIiffyqHWoeFaPFGFjeyKeufKDEwwDzKuKr82lhlvFKuNGM0o52iLJ1soh
pTSBBFO3kbx7HeVT34lCeYZO/hiks1XDEQe+SSph9p3JG+wARmqAfi8m+PJOAFtXg3FBs8k8IBFJ
4vKWUjlLL1wL7pNk3iKv7zcB7paTrY1SvSAlROIy5wbr3aaUVAtlLrRd/zhYRvS4PGE2aK/FR8Vx
XwaF+RUiS5g2mjXA54peDvSDskkRw+WmOHlM01U7LhDTQm23zyspYQBmqhtAsdObHWGPmzFYrYy6
p4Q7msMp5jR0sxu32heboV76GpoHBeaz2SsN9317WCcDTQxNxvmhXhwlvgWCf2RXzrzmsFssWvSh
n9Gcc2rrQUnmEfdfH3Gsnh0FzIwELY5S5So1Y4868PLH485efd1Qf1V2DbV0A6gRrsri3Vmn3Huy
rzzmJwYD4ZjFlKAp7pgiuLrVfROai+w1NXjQ1dWTZICa1NNXZRoMMObCE4j1iNc81Y2HLm9t/vHF
EWWcCJiNvA7olpp272N2rIsEeYFY0NYmQj0LNd3OgF6Y4wkESY5kgV7QTCZZI7m1RkEKM+Laz5ST
+hGwph8/xsUP5GNPdMOvu1M2bMrB3OWdwX+F2xRdnIg6wRWTazub6YVwtyk87yjuir2NryrhEp9O
z7FCkCulHe0asGwTIjZNVt2HCrL2yvWnrwOnkjQBWL2Co870mBe3VIQe2chytt9zln5npkADWH9P
Y8Hii0lGYstKgI/yHWerQ4nBECCq0z6HT1pPplshI8i3IVER1J8+EIJjRXGR0HFG5X6622VGQyOf
4QIrt3aBVGBjP+NdE7F4J4H736kXhmxNUf0iPNg/NfArN2JpYJwNIp81iMjDSiILoTirRMwQc91g
DpK2cHP1ttAdYBHgaR8EF6/A5VI6Xa8mQ4ippkH+86mYuM3KZw5HryrVWORJTRUtz32rgn2g2bkQ
PMI3pRKpfHw6bY/QvOE/+06xQc3vZHSiUksqECEP12uwBx/6AfdrANlp2JWENu6KYNSjn7gtw8rs
QGC8v8WuIbw5osI7TM+pJlGghDPAQgKifVVd4PWr4HV4srScxwlXPsZEkCv1s5mAutusvOsrl4rr
dsEVXxK7AUsRq+kEzuqHJylTBQUVR4re1NDvByQR8sPHEkcRXeUzY8gm/8Id8ahtViMfZemVg9yS
LiRr6/2a193+tmEUGfsY4nLSiFLgoCC0Bsp0O9ZkOG54+VEHVMYoxzpaNEYIQ8uop20sjJekGt5k
QR4+ndP/RVuHpmutr1v9XRcdQ3xEeJc//nHXhQNlrTsK9Zj9tMn3TZHY5Neyj70U+4fEch1L6MQ7
ZYNrMcjP+v2FCuYR5cLKqG7CAvnb8jkKpa3OpVF5sLGwXykuMwaaRUQOVCLRfOkV3fmoa49CPBI9
K4BtkVx32ewL1sjkIEr07rwbliGQZHqvF2LY+tGg5cN4bX62Bfk9Ilqeu2iS0FT2LxfgNipR5hCw
98GWevv0pBBlO8Mt8qEPJW1ETdPP4kwzxaMyNEWc4k4UgYhl+XvdVCCLad7Zhf431NhrL9P3z55m
1W49Vykxwa+ca30i+7Js2A6aMVGXa7b4TSQ6MTvapg4o2wNBxZJA0LoCPZ8c4hmtJPX213brGgEW
f8pQyR7Ku+sMJsRCILJPbc3IiO16fMwfmVHr1uqLB6dWW6HaTOezQxZFh5X/t4meODJrNDVy5xuR
0ePRkxvbbgJmgvJpSzcnCdfbQxytdOfWS8vxO5/zqQTjOQEfpDWVbtf7KBX98QMDB/I3ijNpudGK
mWKDRiH/fy4FzlJeU9ON6Ao7PIwAkmFTq0VSmQUm3DasSXurBadhcdV3s4ez/vAAmRYzZm2h+mqF
YLyadwSWXYYvdfpfYTe6AAQN5qE1yLmnCW3x7WJPlH5/IQzXUHAbVd9KkHuEHMreBzG2iKtZs4W+
Bw6hfypAn9morwx9l4KjUnAOsfdQFnwPxjlchx0LXPVZhV6jn9t+vdpSnhPprnKYIbdnpqlyQB3V
07zUls4t9qLE+gUqOTH7FPuiPwbGNy6SX+ztvzFUSCzmxUqIdv9CXnHEexuA+ccatm+cI5G8eV40
bnLHKfgdpESzSh/Fz4GCehiDlGkD4nlxy6O40KD57aHvvF2qo+9ZUm0DBdfZEpxc6VxYWS/fzV2Q
acgoJClcOWO1uXCOZX/J9iv9iaklHYWx1HH0w96Qh/eL+2EINx7PmFUZXWu4En6PRghhSD3bvr9J
RAAJ2AvRN54PUoIzsuYD3dQqgLenRJJjwkrleU8ep1W1Fpnx5psHQcd/UqfSL6Errfu5DHJDHAcV
eMyJxNKviYS7z70IB9NA3bMtmxa8C6OLAdLX98kRG787tF40Uk+157F0SPRaXLUFZVPBMT/mB2hI
QNaii98G9SG/b4C5pygGxFbcTPKhlMrK5w9HPJUSf3K40oCwWBJwkYiTEATrwNCLf4z3gijCFb63
5hVSaOnG+eOOkOGvD9SPKX12rM9r37quuyjYmDwk71MXAN7D8jl5Q0I1K3hn1BJA50A5KbuDFpn1
wyiYiACXL4cjhgfmWB6JzxuYO6AdSaEnfbats+QIZb8PW8CsL8QqV+wXXpTWZFrVl+ATqIk1Z0s/
9fcF0/Xbt+Bgx4xCF/6dwYe0btpqRNB2NHa7+UREDtgrhZvDtWhxaDv2YsrVz+PpW+hab87DMtpR
OgSjHWGeUTxPN+6M4SSjETinUvp3GZE9j1JybaAFyXtlUKnkTYqbgiJSPc+DWCjdcUsEmaLuO4q3
yeOCwuduHz8D7clto/CPB+rO/8DJ0nvyzxLnwEYGPO7SkT3ojII8dWFVigcg7rBvQ8AtwaeRso3S
sSENLXHsyMPzBsEuXWRBOFfOYrZcT88hTJO3antDiZXgAs2zz2nuIA+KN5ZhbsLrgcBgk59dHeq2
rMH2likh+hjQe5ILVEsgD0jt0TXHzHWv8guqce3HtsE8OqPPZOt1BEVxUNxmBXn0XL8i8cMaCbKk
Qqa/zvb8HQvvZczMYJ4B90ab+dfVUySYG+B6OPdLqzpjwW7AbhZTfK3Z9ZfXu/Uibt2khFTWd0pe
S2Cy3RiPM08OK17tO0EidAPtf6tTXEE9LG21QYaph1Uv2STI17qvTo0PfUI7EiDZjRxShg6FKLPu
nhjjcGg3QT/BaT7QW2+1CdVSkTDAtkJs93CJ516icgUc1UYneve7WJCLbD8zUnw+IDqlZ2lA3lYp
fYLp6Kg9M5lHoLxX9LtZHXTvmh8jULjo00z2SM04lWwlfH9AwDsSQfXw9HW0n+Zgrs6iwc4WITuj
+z6n4UTViAxaedNqeZIcWEyaU6BL911n7orIqZsmutcGY+fMibdJLktI0P2Bpj9Gi678kBcfywB2
/PQ9bvL9rRQuy0ZoWmBZUKC8h8zylKqsz8GHl+HQRfL7GpwwO0OOjb3tzxSzhw5yJe332OjqoCr5
NhvnuALrAEDIditCZ9zxeqJN+PllTF5CJn5QQNsinLaDLbERIwm1FGE3QB/ZPmczYaHS9c5mpnn9
Ja8pEVoik2zJ1/Ah+EaMuxlHSe7avS3/zOwoW5DifPNgbNEYLRSCFlhZgCCe3rUnDD6zffbwrGTk
/XVfwfY7xpCXN1dlEP+OgQbrzSqEiS/LdlJdYJaNTNZ01coZYXfj19WeqlYIE+392gxfw0+WNled
Xxg0BYhnYJGv1BrRl7iBXyAR3TDKRxN/TneqW8fGPDq5eNtBAI6pg3DSP3dTf7Z6jUILDeT0+082
yk9qiIKm8X5oco18OyL49Ezgw9xSVlNkuKwqbuvVyU6gDqNWeYuvgz7awdp1WTPxVUBb836eLlpv
hbzOKNmZ8zivYM2xkzZd/9SXy470qznbzyw3BY6wPeVUU3gXH9vAd7mXXLVMo+o4kemud/0dqbjh
FSidodROQJcduMV2lMqGXoo3H0B9rhnzmZh5oHw1zq0v/kcxA87CminD2MKMlYwdpXV05G1mBaKM
FsCFCiq+LuxmYX3nzt2Ma8JgwyVdBb3EPkQ8PJ5hvlzR2uDvFZ3C9QrUykyHdz90lSAnUuPQ1Yhv
X0FaOXN0NVEH7xTyHr1In5G+ED5dEr5oX0aAty07uAuein8rZitK8fcIM5DCErWvAusDlbkZ006R
dUXXBVEYSMbTO1PvKHI2XWgVvXPPE+URjGam9JfaaXVlvz6DaoLawnrBTyiBkM1QGMIbgqUIMK02
x9dh29vh9XtkpAc+fnRYs40sq+LKLETBZtaFIbSf9GoNGEXvnvN8W4GQdWskR/UOBUUok+IHpm/I
7fvakCkJ6WwwnkC32J1BWA5VTRLpsQRG5u5uPc0vwGOlRK0DU/Oiy+3RytE5Brw9VipvoiuO47t2
4ojXZ26kAWu3+GyrgXKj6+x0ejBVFIf0j53FP+vT0OneoYSp7x4LVLmqFTLfJ3HiZRlNnJwbV4SL
MiVphkj+zRnXqz5ngUJ8pbQTKskn7GpEG6ljdj7MSRFfPyAqj1NpstK3A1kfZjImFQI7nRHPhn4d
6ZZ7x5gCjdH7OrR2IHLSyLb4MRG5qZu2kXd14IQtHdSSCnkmweZxQt6BDJHlF7Fve+4G32m+J4EW
A2odWkUvuIrFv/KMK0X+KamKzNdWkpqOjEEHCCsh5bZM97fB2VWd6L3Hd0wfHeZdRnT9CJFC6fS6
IdrzWs1dxFaSClV9hC9IOR5zZO4M6552LAOqOs5c0S9eMRJqvXkgEqQvbbox0QOXyNePptFnUh4a
RjfDODFFGVPnzf/IgeHEMnFcGtuO9ea7I5Rh/9S9KHGQ19qKzFnVOziSUWs08itGxmQzoxkgtDpm
0Rt7N19ZTkqjqqkmBWozwCkLQWgenh4wSshQMnnbCQD2uxF3gcMVRPeBUVmQKUyQ9GLNjV7hrRIz
wogcn68PCYHAmgYQ/YWiYkvITKHDE4KgbwBD5PWArqQgqg9gYPU3xo5OZWNx/l5kCntn5VOCdTCR
m5rcNT7dJD4HuUYfgM0NzjDC1y1AbQ5fAUpOgjVLiyN4WKRZAHRyTzDWqNDN6X30nw7R3c7SiZxe
3ds+6FqLfhsmT8E3ENJ5Eg/i+rvnY+bmsHx5xNRZEFEZ6wMmh54qUlFtKCYvnx9dmI/0QzlQo+L5
StnljuavkkHDAxnoh22DHMCddzWwgThSENZsikK/qvI1PdzuAk7hyowRC3bCXnxIiLOUSmVqpbJ/
L9ZdaBsLpRa0tRssKSe8e9j9qQsI219DkkWt4wVpki+3iDKX3jM+/2qMFhVG7eJuq43OpF9tSvdl
sgr1ioCp+Td3xQQ0jPr+WYmt/l1PQkZCS/okeTOyRRzRLI2/tIVzjJx0H2oKfQZB4UFbowSB0e9n
OdlToEDPb8wMb9Xt6ZgMd3GMi6LFASczq7e3A+hYjkYT/5YrDZAAUA6YEuLiBtd9Z4XUXXZqh9lT
efxCa/eSlB5U9YpKxR9HXuMDZnVQKBSqD7a4gVLtmzLEUELf6Y2I2MBp0aqXVcAXyyuKzlPBW1Tu
qkDzcpXNsHOCZF++tRjo5zS3LGGHgWEEVbnhrnK+hE0mnmc/Fs/6ZLhwv89a105pbAlC4LjS1f4X
oM/HUPxiN4YR3eqUgr08J5sM+Fq2p0UZWhufs+njvZq/YkFNgL/5rkWKpS/M2CzK97PKiFhGDmAy
VrStMZ9d04MO8z1extPYs/NnAsyRmZQT0hOpJ5KlumGrqOvlOtZwQJWPCzrtlmk5wCjU5nF0nV82
T4Wh4j+Z5z8PdzscQq/kI3LIoM/+JIbBrkNal3cXIxRgJI97S2Vhb4qdAN+KkH9saJLp4ooUqc/S
V0eXbZD5KNkHbRoibpX0fYu+gl1db49wGQm6p0GD48i/OzHZPP3fUA4tZ9/5ivlaxZY0CWewv5dz
oXd7fMwJp+1NkjowF3XdzTaeiXu9ZwxyA/g34TNGpT4E7W0XvCt+mDcKR3+aRlGKo5nSvD2bOKny
W+Ae5e3sAWHbV7junUG6XJDHIWKv6p8g4iWQ6D5tGec6pj/pmuEp0QxS0SNRrqqGn2a9hGDnOgDr
YE1I5U9+PWMriUQ2hlSfD0FcQC0oVbbAAKwgqEtqVQ1LpxrjGP6SP6WcDX88Z5QzNdGNPEXQPHBr
xnW6BRwbO4tjpkE5QXUiU7MATSoNszlT8M6dV0perrS53MV7+nUqeNbr5FG4qnHyERcEj0+WqtC1
WQ7lkMI/OXtkqe04eqgDcrMm5S/F6oHhs2uUWv1n91fSJM6CGscxnwR0wr8WPIDA8rsuYFXo/N02
4fimtbazLf+Zmqzu9sLtbRdvY1jCJfUB69Ng18gwEohyItJ3RBMkMFgqCpxfV2WAvZpbtNBJOxWg
7sk4LbN4qCJolk2hqUS97xHzI0hJJ9z7Y+NYyBtZuFPDgvORymG7Z7HZWl9F+pAPDOsT+dZv3SaL
IS8mp8+536zqN2kAGSA7+GITVUIw+DVK9i+2NwHNGSWC+gh80MSyqcVpHPsajJFkfPuMOl7jXGrA
nCOcqPCrRLeUq83S0r/AJTbaQm6LXed/tgX6da2WIg3Oj2SHPk1jMEAlnhSKRCIGc0E5unkGeR6k
jg0IJzN1296/EZYquUT1XDAFEIN2q2kodOOsgVI1gqKhluTqVuT8/zpdvHBKNJvA0YbmYsMAOWuS
rudE+OxsIjtC8JMRJi2seBfdrssbHi6lRphyg5A6UFtQ08mVSo4EZMs0BneL96zqwxz22169EPTw
icxCZqYW1f8pqKWP2ur1Ys0rDfB7z/fza5oBeI5CEe7Zyb6cTgemBNdYtQo4H2G6FHW7VYIUssUL
HfxoN3Dh5PFGgb59gszP7Wu2auuDL95rRBNliEvG3u43onKcHlknbmBLThS+0EtWjmPKNOmFLOHE
g6TSCTq0NwDjEtFouPV8s5j5RuTDoBjxqeCaggjcV85t43VEHo0NuWVfwFZW/YDAD9b8DdsXoseH
Uto2M2PfFtx+6l3pD0ytUzufE6BDc707abRQkNo5VJRskENxZGxw7EwYS7I45qeQ41Qrah/5Q+YA
QHcmxLCwMeOPKh3b7d/28F+ECUStMVVw7pq4e5VGGfAU2aVlPfRnBHQi/kMB/qcothWhqn+qdXBO
gIDU6CXN477zxndg1tU5pUIfbN6CuCg1iGUe39hNrNZDf05XamgxERldz4Yq8aYea67bwRSBOx3k
WEoo/hUd5WRLwrjNX5r5PK4u3zx/5w90F0wNvV5h+Q7iS2sSoYj2tl7s7kKCcvjo5FqA7FFQnggc
vY2AhvmOYgcLuln+rwxV+Ec5cbxefeD4Lt+g8AirzGWI/yCYMkkWFQM6ur83sjvwyXOBlgejfpEO
r/IZ9/PVOgdeDZ2FwBvkJ/3Eww+MFHmHE8GzMG61qe4MUxHdic/f+ZW+4L7fRQSSxr+9cuTCPuQA
2b3a8U6T06s4dwH26wNNCN/iuFdjn6Ws1uyWUWzEw0vq0R5FluclicVAsIGV4J0Fy6e2J98nF43s
SCQLvtiwhFAaCx5VOGTlgs5MzjlStp7bb0QeEycqINbq5XWE4Q6mJ8sXzqQ5jXA2fDRjFFr/y9Ne
9hTXH9wfPODS0BFzfv91ZOvvTPRWZn/hz6chhzZ6+o39wfnvITiguwlFMZGeAH96fTOOyhye1TRy
pCzzL76Z/caXPcLe79YmnNcJfH81Ux0xbsl7cOobl0PBSZlj8dt4nlhRcbs7FwclLrrS866RkO7R
kJ9Wh2+RXgQyYUMaTMg30F17e0XdVwNnOVyU/Csj1YxzIpd4JB8u8S2DIDSVBKrPoLNIm8+DQcem
hPPyrfcSRyfxiHhiMm6pR5drpcNy+NKPw2h4wO4+VikgevD9HWewzD1zP8PDBWbR/O/QlENQZRZh
hrrcvR3fYbmTfYnxIRR2zRo/KhyMzzofxElDeQYUvSxL4kELL383bhPaFHP0nX4Qc1MiYVZnMm1L
cO9wkXDicpSoz/39/k2IgyMtuJJgtGWG4U5UifH3YDWsO2oj8kd7Y0as3HXfI67lWG5cGNStxbQf
Nv7N7CLoJSGpQqcAeeG06m7p70XbDnQxODbJdpbdPiC+DnPvjyGUqYSkSBkKOfsCr/GMG3mI5cVp
9xUn3pM17EBS0MFwfPsjqUqRM83rRDLYZjpjOIvKPQLSwj56JicrsJjuUuO8504sCJfVnNS+jtow
biNBVWpy5LUKtT0uoaucbDyIKIVU0cLuORIUd8C0ZkelkrQKLYaA7FG28+R7gmCaug901rukOD9i
7Atc/ddc3UmHMfFYQ7UojazCIkFrj7zz3UjA/0S7UaU23aBsCXjrv1J0O4la3RvrOQO+IxcRbxIi
KeEO8ts9m6U0MactNCPEcHxwkLSjxUQeYBDxA+5xYDBnTroLy99sJTRBeXHGt6nKUcP8Yd5LBwWm
oR3AtmiTNs1L9rGXM+dS16bW0QKN/+5nCPsSdevVCPqnWJqqHvYsbpafp//47B0aPKwLdTWkzyyj
XcXjlVnWPZjATOn3YlEMYQ5XjaNBSyC38verQUwe5iROQy2u/16tuz7btIyUynQ6QXZ8SMF8iXsl
x9k1Kmt9qRatQeeV0Dvnoj5JNuAtwXcpQV86Wg1wFdYjzuLEcnixLJKlI+JfZ1pTFvx5BaAQyH7F
Vg2hBrF/9Zl8f4biF1Gdi3mAn3alMAEjYt0CV0SsPWpCwxALqdnyAL/IjI2SaoYBotqc5GI3Gkno
cJuRTB0Oy0+5zxG4rcMg+mVLbwPMuQn1cYOInk2v3wJ2IZ7rYHcWsorinISv/UNR99GZxc0BMARX
mL4ObWS7UeuKyEjQoY01v95iT6Ilt+/X6wWP5SpCpI7wFEdhWzxkuShTNK6LMBu1lj6U9tYc8Ny0
DTjsu/4u6C7CBRNxqjoi0Ejd1lV0SjOkMGGWff5pfs/3+IMgQVDpdfmsPzez6Pv0M+Hzx6b7Oc18
PugJveX05gWQo6R0tfKaRbeS/WjDuCa+CgcWfuZGe+3UMa8BRKXhcK0NpO3D+dD94NVOjC663ZkQ
rqIoJj5oD30H8/zb3uFAMs6kkJ4pu9BUKB9iYCteL045e/Tx4pKU2dIkbaz/gKAuvk5eIvvwiA72
+fqUvXGti+kLBAWp4kIiqxZC+08y6o8u9awT8gmdnY0hCnI5PqbzsgLeAxo0nxqCmcEI9CRQuIqg
NH8XSb5QbVF0nJeADzRNPpNBlkeHBRA0r3ydtf6a/RC0EIbCNvrk3akhozjXmY8Lijv1dhtRyR3O
wyMOJ8yJGvUX9JoAEI8Cy7+mMVku/U+JcaYXZr4Ezm9uusUxJLcKHcbJbJCejPJjsR/stwYLiuI1
WGxalIYAFXZ1SNh0WkIKOPM6nlreVmWYg+blgHC06jaKXIT4vZiRLkalY4PmB5YXA2vRf1zzGZUD
R9wMKKLlaCKyc211KNqBOzBq/+1qaoAOeEu/Iu2GEx/h44LPlyvRIT1DUCvj+qBtHTDkDrZXV8ao
p24vAhZjBNH0azdl/sv6bPhs2fLp2OvgdNq5AIPeo1WasltO0C7mxrIWkSPYMRLdxjdLK7DtyFgd
VqUGWb+4fQqu340BZpChfnCRRF3a76C5UmbBil6h5XFjggnioGG4vFlZgaS/hBHVZgcjXA+Bf2kC
vmIDpPr/Be57njLXBI4CP1g9UOWZi2YZ0HzLRT9+LvmFx1lhMfTlTibpDEMglFkXzyn1/uXjFDc8
HAFHOmRaQqvdpc5ZYrZOJZ0rZMIlJl2ysa3W5x+FWoj+CBKMU4DnFLfU4gj5RlEEmBBPcrXAhJU0
wapMP9tivP6nE83JDtjH8Z7RnwMQHDGpXdlK8GOwuKs4jije52tZYxg1V+3n4/gnSxi2mvgY3Yl3
L0UUX7op/Z/KFIMvy4UI4B+T9HGgMxJI5w9Nwou4lclCqQFhnWvJLQ9LHGGDPDyld2MkGZqLhkJS
+QbvOlt9PirmD5dIsVQZIvjFAFIkRSk4U6G0mjaX2uOHyN7k1T4D30T3MRl0wWFdxCQB1iabMT0x
VFny0/QIGAy9wTRrDJe1D+BG3IQBMZxHQDwdICmyBCIy+2NATZB/GjofIGH0tIfV73Xw9D6x2EJj
tdF0dixzn50YbFpUKdEUzqaaCx7dBQL2CcKgWJJ6lMDU/nEgm0ATLf2hXb3TKHzTZRZxyheexmhb
u2kYNg6EdxB7xHpa2rx8EiB5R9PRI86DG1Hmf8RJ+5X5LdXGOofEA7IT4lG+cZ/YnNe1TyK2ukYr
S8CaMUIuFO7t4WxJ5f8l/1PZHOj+Sqi/8mhu/BftGqlkWCFgd86zayqV3DMnqi/pdoh54uN1gltq
h0RmN9F2p6OFugYiq6J+vL7JQFFLqFyXYpb0kV0sRRiRA27n6Lq/BXy/nvuXdAfHSY0GvKl5r7A6
SNId4ZKiTOBZZFDhl0AbaHzFqLWI9znrdF4QN50HZyhKY0Hlu9F0M7LbYVo995lEWgF1X78iZ3GV
sUH4sbu0L5o1ULz0Wypvnnym0I5ON06b/JEMgmxyzi//GdGoHpTZkuhh/8rI6uGGyni9c9f+QTfa
oF0ShvQJ/JwS0nOHRjk20olJrqvNYUe7JKrEWTkEmZggYseW+CPJiwQq1tK/dOA4RJvTf6EQiEFd
7k0SfszmGNDBMB+sLheuVFbE6wMV8fXbG8riMacxDaioHo+figp1fnk55TOp9VkSHplEfyqRqBQB
Ddc350qe2IYIVq2Vuw6Y4OYbBUDyIlRin6xYzTUQXuD00gm5cyepk0VTD2YbpcEMZFR/3Ml5+DYR
icVd8boDWT5oBzlZnFNFb4bQJCxeN9RlOa6Pg96vQRf4cbI3UXF6JQRtksf4oH9Hss3vR/y5BLnl
1EGDIgyIw9LUFXWtzv1lhispSQyN2sXQqwRSg1crld1evjjvkhdNt5KnG0ADuNbRJj19iIVwCp0p
jhLrsNe2gIMWNr/ghJCF2zeJFBb5p+3sXPtwCsNcPRpQhz4WOLFFgJImzNiU0fAmZDNn8zGvzA1y
4jZ5e/busHLGhQR7fvySYZSe9wMTi0Bi/MejNAsF9T73LUlajhfvnBP8EJjATk+gG1mEzrbIlhwQ
lWnOFk6CtE6CkQClOT3vJPef2qJOZ56y3cuzkfoFKSNAKEKPfwuJdyJBlxPlQJKww0J9IpJyc0qc
hC9vREEG/+1A7viORxD334mP0X1cB1blPeDh8IRjODVTk6JI9D6LDhRcOC2rZF1dMemjG/GlmRQ9
toJZmb4zCwME8/pbg1Ik8KQQOoc7Kfl4qv2v8iXGljpNVnNB+Yb7T6AbY8VKi9Zr3rzvO/MhVpek
0EEL4YsdVPKR0ba+JWkE8dBLrkDrAwBSMCWEA3pGvzXA0R9hL9rACiRrTbnpO4utjbCP3wvhL2vO
FwBhquXQL7WpnFH8tXoyvIMrp+8c2KGtfwyrWV2QQCcxZU5kImBT9+T1FeolX4yPSalYfizIrops
KMo2QgugSrFxexzrlYX1wQmNy5o5AKlnFc88wLw9YEaSDst6mNlcpevK7ssYJnLHBkA7bPc2l8Oi
tOpD8XuXOetGWmFx8xpNcf1+v47Gk5rNAMQGTYE/gpYFioSGgluoJXLpOBWbF307Xf0DQF28RaRp
KbTNG/MhLqrAPJY9CiE6h7mc77O2zypBYD0dheAOF8qK+VxaBvJCW8/q3TBNov2YrXbKXlnitmk3
3dfW4AeGHpFIoY3fduj4+r/j82+Xz6AqPlJJfF148+gT1gaevdRQxwX/Tfuh8dpe6I48HhS5YopQ
R/zF89diztRzYr+UngSwIQ62TpzuyxWd6YPaVUR52cSV4tS8ULafkjsMFGNfdV8sIXOnGmvSTEFr
iEiQxiG8AfjqiXD4mzTlSgn/d27BDEgRfroULRNrWq35WLHGy2/AdH4SrmnXByy9rDthmZLvDVkL
jxmMLahvBOua3Xu+nuu+WSDqw5AEuZkwGZeX2WamnFYkwVDzX9H43szOdoEw4iGo9rG+5XLUdCEl
iKG/Lb2L1ZOyDi6//qFTRcmW05u0VQOxNQapmHggQObOoU17kpED2vkUT1EV//uQvnm7HVrUHpRu
cbcmeZws9prYpVSl+CQRAKQyj3rwDQCFg9Y4FX479fYuQfbMd3IOrbDQsyUNd35W3qh2mDnDZeBS
ueylhIcSLHDRn7fNA0msQr/tJ8GineuukDbECNTLvdDGPTwo9HxmfpZuzdTxj2F5LI7mbZGAXwrd
n+Q6bj6Dkj1GZZYcknpSWBE70/s9mRoUtxIlWxWcZxy/RVYAVXTsQf3GBcpXt0gImuvxBUwQHMY2
knXJmfycyM8uwsaf9pUDnbJUgFWH9BJBqp8zczuDnFjD4wW1hU3/FqFiD+DAM9ZF++gtjyemABus
vj+iYC+XFR5R5OyC5rfWqX3bEGKpuEdscAaM9SKIQFZtBbGxtbZSgb8Fjm14gAqL3iyk7pZEaV4N
d0mCd+SZFvlKFeSs9Sd8/Fu7ML8LCsWtF4s+XxhmMy7xsksILWo/IFf8SBU/GrWUvXCVLf2cBZZR
mswiMcX61O1YOJWm8gFxViUqxcxI0uG/HGWBa1nffGd5elhsBRD8pPNwwU0G+AgJqJXBVrr3ZYLc
eEHRmPKhng6vhVGK1Sz0CNfe0ryhxV6wFuUIbZzHjycLZGnLfnRJhJC1wJ7Od3pZO6Lp16VY4cvM
cXPKJcWHZAtRs9v+b+EXunefZ+2TjXa/Ty8KEthGPHWC0azYOe6eLHzFugGccjlu/eLhv/mbH5my
XL2cFP7gd9mGi3a62ypq8gSu3ZfhwGXc1pwDyXkvSkVeww9UHLzPk5rvnBFkhBJ4kwJBz1KDMjDq
j5NJC6uzvC+pKrQek0RwqWNF9KP1rwexo8HJBSY2sDmXxkldzAsU21DvK3wEMqildy/CZfDC+PzD
+k6gxyZ62h/mHXNaH5Yn00C++rzaVQrY0n2G0fGIlv6JqGJM19yoSlZxPn52wJjnrsNI3KPHmXuq
3zJaZeUU+r1gmZ1UMSYCO/dQgpNeAcAMLLwrymcP9Grg59thNvvP7E8V/mi/2HyHwnx1Wte5Td3v
+XEYk18R1Fp5AaETP3+/U2kmmLJInra5g/2563HsTNOZPtzRwWSLtImxNqSwaWRnowtz9DpEFTqv
Pu8px1yT04f4RqVfqW19hUupKH/zeSFG2RBSdbuIrdor5w6bYsNJ4ON7br2WVsXRwoStGiLlUAL8
GPpK+RKUBDgHGYGVxDtnTTO9EMn5vi7+G5K4jYFpB+93nUrlhbr2leUUJnr6wYsGmtLbD9wLUiIM
N6TjD3TJok32ZHU0gvkNqiAydhglLbFDBUrMtnizPzRh16PPLHkzSmAkiaDUhrIT4RX0A8UQ+2SB
92suf8LPK/EmBO6NLQLiexAdiXVv/f+6h7UbO3AgW1hRZ/exBFYtWobFHNI6qfqk7uXCVkX8WYzi
YK70dStQxZaubM/Mdq5xYzVZxw+0jiV4ikIASvmLTZNrZOisp3zI34K0mmF+Cd1JUWKAnu00XFz6
1oSkLHwNgpvs+Vap02IiL2u2XxCfn64R/LAwxZZ91xKUoxul4NeJryqRQ1D5ytkKJrjAxgknJDA4
Dl4lMc0hzTp+vxMHrfdoF+4c+keHNuY5XZdlnRhxj0PAz0O+RbYs8zz2OiAcue+HphWKhePKxApC
nzXXvTTJ59Rg83WOpy+xG9Y4oAgkWmG1kGDZr34b7KfGotOGomO3DMhU81ye0xEJAdp+Eq+4qpxQ
+poEl45UsTFRh7pwtSFw0saS6kwPe58UmX3QryVWFNzxkxTozG6OZhAXslGVf0iHn9mnXs/PWVBx
nwgtywTtztAl7ju3hugP+ZkZU0fy4VGPb08wRji+2iquJqhyDxB81Qe5XgIjmegZR+u+rDeq9yd5
T0tUaXexsPefYggpZknyQDCinZgvBMWFjCq4jysemCG4fe0wHEuRuDcge6mKG0dq3W1puf9N2pmU
ZEWqf++U1ewNu4Lmhy+G0sVAX3/CilOyKVYcPH+2qp/1yzj54yqrBOo1sUA+SFnsbHl21S4GDrqI
FADEHGbZsgrnw6wf5XxP3iSWDN/y1AJ95otOl30ttdn5cvR3zHXWYzP1SyVOgPX8zZUMxL8nqQGz
B9oFaNduWX8njBuhq4WvnhPS8ann50KwbQPmsQcrypvduGrSrC043MWzHz+rxgbE7BK9p1udo/3M
mE5mR02xNPnKbGMivhe7SAjL9VqTGReAmr+FgNdyCtnTr+rRlPnid7SlHCAMuTu4HgAGd2h33u/U
6PgyPTlN0fkdNhU0Um9OWsUi6GVCAcmv+Y9D9h5+pzAsHWffKp8D5dFjxFrvCvp/bmQnaMxVe3k8
5H5viN/hoAbiRp8fvXLjdS0kaBwb9aPbliSTKpxWBiWgPXTjU35LjMC/3yNnBRZzxqnzNpa1IQrC
gyg5DxflhuoHPGCOc40PgtGreTZQ7AI1nVBIbbQUkvuTZrHP9Rdxrh9fhC+3GrU/yy7NYxOr7dRM
TSP5zeri/iSKZ7ExlRznxVUVDjcV2b4meQ81iygx1O7A0I3I0tKYI7jP647GNlP7TqkUV/DWvM7W
n7DCPC0yAG0SuRBxLbuexUovqygezxjBVQCYJwRGH9hVB3Fsj8mqCTw1wHjSAv5rEQjVfNXqfysG
FnybfZmXAH68oo7Fm6Gr7N8oagJcMifmPqaPPNvJieWPYnSMPod/mileiCR20mhB7OR3PW6aV5Bh
TciBJseMil5jKDPw2ZI06N+EqQBfKheKF3VDQhxf5QhP0eefqXlvbj6jpukWr/6avF9/4PCgOUTU
bGscgNHnk4D9Rf2B3HCPiFl+zlvm3hOBwlc+ZDwPywD7pcOTpTrJFOlzn03OsWV1lyL8hfco/Zvx
y5XedPVZ5RwlPO1YbtPVbSh+H9ao7/TA6bpW9tLF7n+hEYzqPT1nR5biON1gJ3wp3qiZbg8QqWta
RQdoAcC+S/SjzArYY5pMykAo18eMGHCryS2R+sshMkCIZqs8rEn/wywSqj7TH6UjmuUJuT9J04ZV
gjU8EqhlPrwhEKZJATWWjof1yPhg1eyQecTddtvTdlpVNSJUPSwTVQkS1bRiY5VFnkI+Bo5Pk+IO
//hGTMAJGSzsMFxdc2b5KNcVDIMrZzkS7G2ITyZcZrddfo6tNX9SUerp9SvM/IxWGpgpUeYnFZYm
uUKCMcMBWW2egLsmK7z//o5R/4g+B5A29JVb6HtuYhv4Tobb0UMMwJfkGlGU2aM9Dyfnl+Ye3q7i
iyZkQyLZ+UueVdffbZFQxeAuRgcswd2r3enjFQ1b+ee4DoZ71wH+GJQd7LFzqSudWAXpf2P4D5tY
OZJIrXiPonfoEWGhnRedPxhagcggdHttURVd7X9FEMap3SWnEXTv0wtgt7pkCX554zz4wa6FjT7a
AyXoG3Ii5gRi2iybiE5FCCVqS0Cw2YbQzD8aBxsvtxDrH0HwoMiJbtDFkXA9OVjiFVmjfZgBF8Ut
Ja4f8OrjgNNzpy1TfMklYZ/j3ltuM8pbJR+BJbWMOyrbmD4KVw0g8/fDC1g0hGsKO2Q+jITEnt/j
P8EptWdygoi/Nfx7qWddDEG9AaPxg2W3nSfxSs5CrldtVoQ3Y/7zRtVcwSwK3s99zIPRB4meBjjd
5ZuhvjKNqy30+S24NcD6ceb/JBCp4iA04VQUTc0vhFxDoUpP9d8wS/XVLIgG3rRZvP6cGw+WcW+D
yMHuFkVfVWniyLqU0r//v8OcSeMKqwTb6cXN3WN0+vmANKLZA6ABjY5nbmFnWby47ZFljz2oGcHh
uXnvHuOdw0/t/FM3/MhF3O8NyqsK5wj/bdqqCB4oG3fRlrhLBB6OraKG3vHAP25Z9CFoBocRrHvs
uAiStwfoYEYor6itD6c9dxdEbZNlU5xauwXcVQMv/uy/MSR7vn5qs7j2zTUhBOdKkKXOuZpJS+uM
As6h6KteSYt0HUmOR39Mlmz+cuS83Ow9Ju3+kGJV7O7yzq3oQlzblI/emxB4r8lHyoD1Cky04E3Y
ig8Ob906kKm1W8miNHkRlgpQWGcOypV0s5aSrVu+fb0mZ2MRErXa3C7hVt8ablS3DyAOAVXVfgY/
3rfl1lBJVwuIb3DtYCnmB2yunAlNK8DZPIs2LJ4umiJPvYzFKJFVixUher8IYFV2hOZbmMTSDXKu
ZTTFWC9Qwxzoy+rW2+/kAYECWmnkV56iJBNUXlDPh3WKaHZ9rhuHzYbN2BLvboaDPSnkXWd+MBHg
KwvDqwNtqXVsROuX53CRRJqArh957rUqowakspJTXmfochNm3BYwKB05GSx3/dOBrUcYTrjAXUkT
lC4EHNKrRoWoKDfnyDntOWTSHAg8MYJG3jCxttln4FksG1rfsGCO98MzyOyog8WjLeRtvE4lKbXt
2QS9RV9gN9mfKHj8a6L6vdx1KuE9oLR58kRE79x3hadX6ecHZzRqu6+FFLs5Qsl2n1oIVFPyE038
ezMT6bfFgdr6itrYH1lx3HW8uXoObJZkkbjqKS4RzJPZNLOOUpiOHb8D8BLelpAT1qfvg8uav5k6
oN8uj8Tsq2D1BAiL7EkPTl8o6BXeAcrKUqu2aFFBZytg3RbHBdaqVaTFXOYIumJSrZwxQFXLLH50
hOcyDB8hujWSdFnITk5Kj5bXqDi7xZF5vk/6wPjzzjvHX3W1zJCxNzEoY6KgIcWpbIaeN4bhJq9b
6PxAvNZahEVFG4q3s6G66jKUJxEPNcyVfbzCFDfa6Q5zqbR62LRK2uYGv0YQ2CQKjvgxJXvmTvQH
CjY9q8KMUm3hHrMyEnh4/6Rh+Qgrf7UGq14tE4ooXe7EeF39tShZm0YTwIdSfRuq/doWyUF3nXR7
MkRjY++8d3I8ISPYbs3UvZe7vgJQjqc3gw5o1PQ5d6wF1fkfDxJx/MXiRFoc8EgC2tNLZ1PGmpfg
h2YsyaZnw/VXnOW78kJYmOkv5BCOdxnMSIaV2mTtKcI8jh/1CCG41Dq0BmGUbZN24oou0l2oY5OT
z+q0rKeeMzCZMFXjKqKRxC2kSpEJ9afism9PYJkRCgEAbNahEnpb+mo2gcp1lrugGGRChoO4I2ao
lqkDttet/eiov8g5CcnxJz2cQIeRl0hto76FsA2S6V6jFIj60lXjlhJQzgUtbuUc6MxAWKxe1PqV
QzeE5Uu2vIS5PKPYXzjGG/JHG2NwuDAqtcm/mn5yY95EbTMIAzjrSFLvjF44D8v6u80fi6qqDSj2
Zmm01me1yisTnID8RXYtjnh4+luxmwHNzL2zeaQQ7HPBkayNWrEEmWGVGf2bS+VKGl0o+8nkepUV
w68dCB+mMj3UnN7SN4We78HJPYbpFa3CNlhS6DyigAnq8or9Zz8pANmxJq23vc6oDM7rAV4nbBwJ
iNNHHvo1Ns43gutDgLoko6m2tiU7vLvDlaBMbpjv1N8PWVPDaTu9YFVhgQTDdDYkp16VU4misTmV
00j5AHNhHIWjNxUg23XIny1LXXw21A/G3XoK+0plABDN51Uc9dTi9lHg7HiuZDf9Z5zsOCNmZ51k
VM30X40BXwcD18/9EaaZygPekFp+10hCPxM6hihdy6oAezYTXPVKjiTcu3eTCLlYq+8VQ/72PX5O
xgVHZ6BAkaxOXCBr5Ajw+BWsltZUwC0M6eDteqS12JTxkPoB5oq/u3jX+sIwsFUXfPqTxGHuT1Wb
pmfbE+1+eHc7zEmRIBi/x5dWOdKycCXMOx5UwSHJSQeFnMkrcbhM3BtOn00I3PR7TcMgXWzjwABg
L9oalG3Q+vO5eNhH3SRuXSUq8TWvATQ/GDnnfnOnx2IpM8hTAyH/i+SLukhgTOAuWbo3augsrArT
cuJYE2xc9IYmhHUAE7ewK4B4d50v85UaQ1/7qOQiZZrSTI23CPlCdErSCML0xbPtryVUTfJN89QI
N+QT1kX10T4hZx37l2pdMsF2mASo/ScSPTBftA6G1oPWgrYq5JejxQubG/BS4bOZSEab6+RcSa68
hhqV9uEGbW3WlXhF+plNJmkKjlRZPqHgXudMbXZgu/vBV1I3DVx5ohEsk8rQpTwG9mQk2wKeu4VF
k2hwwuMNoWDOj6hmYaArkxSQ/jv9Wt/InjAypti0atsetI43kolfGlWay60XpvNeXqSbr49Rm3AQ
VUt19i7n0W15zN9EGuZb3GyCsUhMmn70xUlci3uo1v8DlnocvLNxYIuD+FH7jUolT1MV+PxoroMD
Xuqq/OecYvYjxZQjN2nr7EOGxe+BiU9xZRnZkVhcImvQfNzjzPdGIHAeVWBeYp24cnmj61fzINp3
V60qVK6flEvnL0fY5BdF/FOXEZyQdMVYj2h/95dTg0r87CaaGFcQM0aB0vqVbXX/XtByJle5r6Pz
ljQgwMvwlu78MMiWQUbcWV9fwwjdsW3jAgfkeyu2DGYMH1SEnjvtKSzi7cFCOyTzbrGR78cyVK0V
0va4K686vHT/cvIyjacPe9Dd4Q6rrq6WgL3ffOS02SufdIIhm2b5Tw4yn4yv9vnxyzn61+1n8qL6
fwadBPTqUF8w1k657/N7wm9fu3Q2gMKOF5ZgdaI2e5T1Kz2BxAWZpfohpqIPjZ+bdMUqsdUfFgEN
RIKeZTMlo5iHXg6xNP5x2Y/x+Nl/FGGpzAbGat+2cSE/HUC9aAotNMsjaEpvCMlz5gC0OMcxrsdg
FuwGHUkL7zyDbv44IddX8O9rxUy9RCvkrWorIJDgYji+RibS8ZVhyRx/jpNdFrxBVSclW7BCsyDI
FuKiY6rhM+Xe7U8rKIXmUjyk/UxJOnieoO/NqD5iMg/OYdLn4GwhdlBcMgB0zG28b66wAP3bttkk
a/6vJLEIM1R0oyEvfTMaKNnoKsPf3O84o9R7N2j18YoDiBwJEHxtwECmBv7IacMt0JiDWFqNsZFj
CLZ1Ul8RUMQ2QI44+eh3+EkqcQeAE4Gj0tTpkIhvWwapULv1Sty6JGvHsd9laRvM1/RhNM4XXEGH
Ajz7KbqgUeZpHUlk1h/kBPSMdkCKyH5uzweabv924RyLD1x6kFTW4oQkspJXpChxHK+EJg1N76S7
KCM6/kLS2IaoLsNiMi+FlLG9i014nE0IeJOXyQkYyv1z4pYHBQpJgvN+MjHxhRj6DEm6u+2bNELe
9cO8kNZDi+p6Hxpu8DnwBSOwle436c5vKArIiAOnWRig2Xq7Jvkw3WTxAZtxo7A2yXhFbWRc3QZh
Rv/bXZAydGWeFTDTKSOS0fBtfb73gHCJMRGd07xvrilovaLJyrSkpFhJpnJPYpZ3aSHKpU4JbSWX
4JzgXjIhODzr1NkBVMaJm5XsTws1C33jJU93VyPg5eW70aje3OwqiWmdjJF4XnkFIsCwC3JVGDN+
adrwXNHGrcVnyiMwTZLa8SoUDLkoUVaQ3L+nWscYyluJY83rUGBdiwh2PqpCeEYUAEe5Z969ma2m
7bMiyiOZ/8mOJP1C6o6RXbFaT6OwQKU2c5faZATB0TXKvZZNJwmzwCwmOQj17Mh2x8vfmThwiEoR
OfHFIAvXq60XXu4TbiT+n97Oj8CbWi5cbUGv8UeSk/3RDQzpWCxecKU9dxJ5skcPu1PBso8y19JY
9RdBxdBZxO32irNrF3VyH5LzTM7r/nQmEAa9rMnFuIpD6WozKEfplv/v3M/vWsbl6qyWU9PcrTeK
643MYM2jFL5peSEdSgx0x7FeoYjWmcRCecx0FcU0bYCMjY0WiJ2SHOlAgN7F1fbE2tXBimd8KopV
Z42kB858sN+YnGovFNqJLmxhRrpNyrF0MR6B29+9hMK9QqzMviBi1feyioJLhdloRcILMK9pzHGB
gSKMyJEhWbcKYaqj+B+2Y26NfwKsZwwNxHQGby0XDRArSjsBkUO25FFmUGcayDcGIU3SQzfT7xGd
Xz4R6BpqOGimT7VlJPxmV2f/mPhun+sDadBm04yFPJ2fZXRUfmgZkpJ+MM2XIbVo/6Be8zu89dyo
Weom2Cw/fIoSGWmYuq2qDWxSqUYw1mWmezhvWmITtYm5f30T/WT9s1iaDt+DvLf8+0QzYk3wHsbL
HnYdFKjU1JkJS+g82woBNcmLOPUNvU/3CLx3cCE5+g7GWDAAYRus4s0d7lOWmLC6ootfT1AZkSuh
4deyBiuEDJEfeiPj55b3tNhptYU35xnpmx/H0DSXSKdJf8LtQ/q/YQA2VfgeQ07KySTOg5Xx5xsd
ze5fnesVSJ6tZr7YnBlSTLEqWHRNNTlRZlICZ6YI5KIuqhOy7PBUD/iQzkgGtOQvoE4LPqKadLBE
YGX/JB8ov/+CgmCPhKuK1NGRYs1V3ipd/wrcIlu5BvJUKlmsWtrJ0fTs0AFYnNiIxDPwL6S+Y5b+
ofg7kgoC17tjEF+EDFkxlp2FZxfGb0xbJO3hGpdiStx0AWlejZTw87JXSyWijaW5lZXe4BMzZvAc
A1355+A1UGGJVMKAs+ZoosI37RHLv7EFviCMQHoaMFbUUGyrDeFIX09/h395VeI9nWMplsSAnaoW
XLHekeNr2zazxZBVd/W9E+td9dzL9RhFB0b9zUPaEkcWP/IB4IHqSeJwlTzi5AfTfDpG68zyiShs
uOiWgwqrNYpiMwBYQilCyVIWhcusm5n9f8nPu2etscIJOVWW9Ph2iO35N4bnoJiaN1oZKemjWUH4
c3oDZBt7Fnj3DVXQIstTZF9uqJDvQCCyTM9swhRgCCoTR57TT8rIfxEjF0vd9TAq4kRi+KIkrIwR
WEQxtAFyAxzGVhKGhSoWp7MH5rFYHCePc0MvWl6AFd3T80h7n/uPSWMYbImuRZ9WmcFVZz3tQ/cA
s+QIldsd5hrjMsFrVwxtk5aIymVVKjDavaYfN/KUIL/2Mj9hUnyMB7CnO7xm0Gr/rru5mjG/liwW
fMbzvIesZVHviv3sNwR3KmEHwlJDzDWFqFyLM9iasLzlIvImQEcUDhsF5QUkPhQPpjPN3s2tKUDL
QbuuNWPff1G9VvfMxtq8PLPClhdxQUU1ePG/taoHN3/HdTc04yZzAffWzmfUgb+x5Y+EIDv6lFQY
765V919JrGhWDUcOlFZeoJ1MIoLscmqz/NKcC70/9OKJ5dTHQGOf5AuDOguu1KpMgj3q0icAW8Qs
mPcvPhP3kfbew9Bpa1Vk5qnseF2JLoaM9Cx4nyLd4T7jP0jipWceVoMg43LaFRIyRVHF3rzHe8Ia
1ELjQf73M7QFcybQo4dWpUKZYRO6JPIVg1foD+keCdnUBjOLCEhaHmhckDYHrIcg+ksHP8Vr1Pmz
/pqjqDphDdBNsCU7gWG3LfPkW9VGsEKCqHcf8lvoYR+BblNsNZVTzh3IJYuoogDwixn847XNb+sr
WhzIb1wkWAC3+bD1L6Ituh6KDpi/7U6FzqDljohApIZ4OuA6eD9Oi6nNt4wEObeF7ZPX6MIDGXtt
xhjf5oaUc2sMTo7p0jwwH3uYHimFym3AgKzEu0P/8J2c9OgoIAdSr4rEY8lWwZO46x9xcdgfYw9N
kJqYaaIGfbcRKTxVQ5yYu6iaOqyh6gZgK+0uqExNUYb7wTLvDOK0NPzSP+CwiCK7ZobT+t8sR+xY
zNg7WgV5uP6n5iyM/mFeQNUMxQOJKAyM8QMqAf00fVlwkQnNnqLdKuO2Xr24qFiTQO9hm21vKaWZ
peCFVgNQr2qvqjJEGDeYdezLw9lGnQop7GpICTnGF7BVFFc0FXrOVnCnpiDt7DAO0IWWUjDWrVg4
kQVpQnqxMw5mQrU8HsxOpydxQDqupAG/EGce1e4/3dm9PZvEE97c48pDg+YECUEO9xqDrRU75zQ7
FmxvEMFJrgMD9V2BFWS7aMIW7skwMgDbDXAa0lI+g/LMsx8KwdBDBRMYf4zRpHUY3F0uvRgtaIuW
dCN9xnA3goZsE5xI/piHIjUDpZCtA4z4ABLEltQ5Kb3vrDktneAKIwvyzspBXhU5XhTpKvm3QpKy
L0K6PjrgeYLo8dciH94luV/CUZ6LvR+drwpVWkng95gKT3zZ/090S8nJ8qIVAyt3jpyLwDipGcBF
JJsh0ciokf9S/lyc5rS3JJJBc9SSNHY9/kqi7nY0cxpW24RJgE/hfHurYYIqNfUCLOoDxm3WYDn/
MBUThiaNKP+hOvgtjioKVdABknO7+puTHrgSJLrwX/eQx14bATGS8gNiX8hr8iy3q6bIBMcO4E4K
mh9dqHfGI+apvNn41ksPzG8QmvnAVUUQ4nQmVA95peJBVAZYrxF0Yp1BoyDhc0kJ6Jde5q/QnI7R
Y4nSz2WlwFm/Om0a99yg0jVR6l4KehOPb2Secd4Ah061Rs/0lgbnF4MEYI16/132eVRLP43fztv9
gvlJ82QdRa1TFD22CWZeg+8UrzpLw+g6HK+wHk6VE7akfIjqXyq7GcEMPwWEQy25l3GjPWWJ8ZLq
zz1WvvtHYi/XSf0HNlSNSIthnt5qJ9LzPzp+cFcI46A4XmGtKwe9ytju8YKQ5Nfzy/bF/iP5rjG0
qMbN7lFOhDF1MwsOMrH/WnxowVKd4c55GsXhoSfrII5iSyvVLZ6L2a/V6XvitD9xiS2aUUNr0J4f
7HfyL6RoQeeHKzrlFBKh3iIFhFL0hfa74W0ht4KYghGYbH1gNQi5naFcwGChFkLkXTdGXmabhjlS
UP5D8n0wApqQXB67DdF/Mm8LCsnSFz8Y0aW8xAYbo75YxBPF7D8ShpcuSBuOl6uBZq67SU3Y6WlI
TaZrtUTbrBAVuOcNxPta9JRaL560kZQKFZyQ9P0F4dfFg9wGTJev56CpTwCUx36g9Z1pzkzE3wEJ
Ajs4fIFX7FfpuraJC0SYwuxe3ojJgCDin/7myiw3GR8yNc6MsicCF4KVgPRlFXypAgylx4vmAfPu
ohYNr0pzVuv/wiFCb5rA+leEZ7eSK1HlP3whI7GqRk1yZscAylSIjaayW8WblQ6+pUAupy/DchXx
WAwU6h2EiGfxb6FvKfTtSvI9Y6q9u4uNoeQzpkwHsk2jDwjreM9y0v8fUclklNkrFKRWeUHYLWiF
zLZHX+tZJlu3xFTuSgEezvMyW/RY6DGnW9KDnVyDETUJoCWcNQroNMXKB+PNDrn+JK7tnxgeFBtS
yXIVRzsbWbRAy1GUlp2LQgBia4xiNNGeOSQNmEY6LS7r4QD71NKpwngU3/JMiiExL6srJcj8eGna
50w5dXI8CWhOkbqWYZpxrjoRPKliA1GP4L0KcTXajwbsjRrxsCLbIxBWHqGVhMlfpMmbHn+TqYea
TUtRw4ZXWZTMhXnACMKmM6/OV+kTCTxBqF+wMOrjh9vee0UnGTobsN4pF95Lrp+0bm9cwNO5uF8c
o4b4Ihm+CKfsd5HgK2cxNr0lWh19Cxulv993BBD6w/gmTVSeGQPdPgGavDNlIZ6tcdZsovDGpquY
IJzDaVPAxiwxMhpvg76IzXv6XqAJVa8xcod2oV11V+c3xIu3d8ghSoPVoGRUBU/rL+ZPn8+lfHaV
VSpsI5xZHBY03DzvvMWFjHFs/+38wdPX3ax05L+MHxZ5ykJ7C2ojVVDkWqz8sOMBxHdCIvMjucqp
evgLxAihkuGOEKKXLCBsovhYTYb1bDfEG5M1igXwuWPPz3Z9WarbZyVk1xjapW6bQpikfMYluYaJ
8LMpo4ZoRd+7xcNgW5j+l+JW5RvaJ5mdfVkHoBj2240MX4zD8r4J1O1/8OXHyOfvNxTLzTX7WdFG
zD8Vvwe+06AQhAHAbemqz4zXAZu5U3DWZoPf1vRwNooHe2nPFomuRxr3etkp++8/IVxqosvb5/FD
KhJMP5KsSCaX7h5kE09PAyccza+tg2bA8r+RAfyHCUDOtPZ2OJYWmIlZ3DfnBzYhYQ+0I9VgsazY
rkgqyGDzQsLTSFGSsrXs8mQjpnJUdK6qp0F/CxMEaWyBwFR1a84RaqL6uWiot4btH6ZwQpzaXU14
8mhfVSX5Z1XebhBipm84k8oTSpN3dHJFeWdelKFY0zZohBNl2KfKZn5EjXRGsvBOXj7vBnpZWpIw
P5hnV9xGc/tY/e25V7oMUekUCSRPf7UD1JOmmpqpDkz+21trX6VQLXjnOUbl7M0Gx93EgHYO1Qlc
b9hbRjHiNoqdmjTAfxMOQsexd80NRBssXSwxLGPWAhxmZObe9bKTBGReX/1eMex9wfYafj8Bl8r6
GdQ8cmKgJNMmaxdviBBJ80VXKcsUsQTIe5lNUfLUDUQT6jRrYMCMg5hn8VVpGrxPisqDOwdV69em
5d4rbctaWzuS+W03iRwoKraVRC29EO1ozJ7roHUp1JQjB0n1frj35PfzH3MqWs1qNDmQ2ICThbOJ
d/QYChWMWhKzrOE53Jjlbhl0Ba0ApaGwERBuZWln5eD1KMnqfTjq+HMb0OjIXrRGznP0xc9a+iCc
s/OK/XzJPrcj8B+Jou+eQdcZmC9YiEnaONEcfz7MhglalngEfjbh5sf2LEvdzRv4MwdDMDnHEXUR
CqREqRUHtfDkvrNFEKS12pXexxRfG7r41GdjQnYosseMEucVF3Tnak04J6IRDUtR0NSZ29mJy4rU
KfQAerXWbDpH2R3DxVio5Eg9vxOa0WAmbGVIo8dXWoowdS9aQRTz501GrgF0zneUOEIKmUWPfrcl
9b3ENtOH5cNYZCKwhfw0sYcrG1kJUOeuvMFY+MLTV+cpkRlH5T2HG8V1DOmMZqGcKL0vWGWoXxcu
Vmy9uPWoy1Ljv82nMcawr1lYWyZ5zqy4zga6HDDs4xJ/+CJ5xCDGaT1N6UCaAcwpc1wwGYwJRH1J
3GrWB9xWAJ1i7roPMS4bENVXgsn2zjoEqe4+dnCT9VLvpxelYutccUdaVzUQzdZdXW8+KwAvC/S0
EY30E2HjqzoI+vy0erdzoXbMJvXG3Mts4wwfMTvMMeY1vdxVGkirX/8YxHO6lNGgiXnrCasQ3JZm
ic/dlC/17Fi87nC3ZH0+WpvML3mIpb+gNoaqinN2ba0mXkBkdu6Uie0u8LJxFbWcD5bct3d3Egqy
ch3upN8LTnDv4SFBuYxEL/WtBkRy8wVmdDRx51UouvCxf20Vb9gfiFbe4h+myF5/BNu7G+lcE/Mk
DhbhEaKB5kFza3GYsqDSMEBnEKnGSrLtZXHsZXEKM9g99W5IInQmTDlHzXneXv7vFqdf39lBsmGW
xa7dfeBBhrhzLMFsnLHCyAd3KzUPBi8x/4cFdEIWokoJuWajMyAY3fbO/TVNG6me/rjFKrj6dFxG
O0K8swrIuJeZpz/jI6menFncz4epGZD1w4T4vz1UfX/P5XXZCXrUZcdsgSh0zNYZZm4wW131CvAl
ipsM3UxKZteJVZQfe4RiS9efRYsN2+QeYEPqsjmowbrtE0jTfWsRtHsBsWfy8LPSRq3g0pALOF8z
TMuKrP0k7AG6LQ79M+WnDQ5Ezf4SYR7NH1Bc/OXY73U/Nfut91EiBRH7p513vPlRtz4UIFn8LuiK
O2/HypA5kwhCEy591xPmz8SLP6dW4+tWzo9/7SJ+iiSWW8nxydrc7F8JakBp0PHxgixwnnoF0E0a
Hv41E2eKQQYhJ8gIzMhmOQB2XYmko5Z0GhkzZrzbYJwu3LW+LiEIOEopwQ0eFBBbkrHbBUbBaJKP
WifHnscGPHRKnzsz4/2HVjN1JJkIy2F+ryQGuZvDwJ4jfCzjB0k5aJtaKIZW7vLfzCsNgt+wI1vW
EIQuEKsS3vY0LE01xVW74Q0oCDM81+LTnAf4fdwWtCRR+C8nGJxmE7AleCM/5/sYp1LtsTUDURW7
9hSuAzGX+GkcdM9eSw68URGjqNSl0vtl9+LV6xMgdTb54utBnuLR2+eqfQyQgAOFQTHoT+zNUvGC
nK8cSc23qHQzB3AS9nfgLtEvZgzeP4g2HOdnCiJppZ291l/Y3a8+GeP0EXJDUL23br6D1G0WD5lH
/mk722/seMiEK+L2WLZ9qa6WViN7Ec5NlVJuWT94DP83iWbosV0sZdSOqFvyUr67+u861GgdF/nO
7AT5X3fj/aST7JpfQym9SLWC0QshrKxV2X0IxyIJDIOKrE/0Vl/RvpX8GjyYyeeKLEB7XOGagfde
/aBkxMBsJ5LLpBq67CYYAb8JK/2xksJXNr0/8G023xgVtsamtH/DfaNuzA7daOCE2FWRdPmsiQmh
PS4DUblF0f0o5IL8Qb9jEQ30HAVA75n/hDndEHC9iSaIdy+M/gO1TBhh5HWK7EnfSIrNSup7PvwC
3JfaWU/GK5s2AYvADkROngceiwSI47RQDsol9LrI74CxSidik5QNTTV/i3rMgxXTsPSUJaksEt6j
sa6DSUnti9EZTMLkhxCUBhf6LFbeCcdKlD7OGhiMj6oRXUKBbv8fnNdg79+jj8NkzgXZxrxCHYqM
XQ8drLjpgDFc5oXzssBcDawcN2gk0Uz5A+y9mO260xSxujlHs/Qh6DvdRpxRyPgkOIqmYr6IiIZI
8djaXGLsnXk6P/abJ5X3m4Q1/Z8sVklCEJxRRjzb+xDLmILTxt+SeoBwvGVnMh5kw7WRth4XQ0RO
gxDn6BD1p8IPmYgF1JhNrLEAtZh6d0vzUrbDndPgVWzgb4rBTvVwrUhEkYuxEGfF9QcUBJbT3TJ/
+LItxFw/hs3krr+/BJJZEJUA8j23d5PrbWBxeAojtS5b4jkqgdtoZ/LTfxXtAiBXM5x/BOAnnVaA
3M28gkhWVo8QBRwAuTIlxaLXUCqmHVLXkdq9Fp5lWx+QnEwe5F2I/mm+/VIXhWKBBcJNgHaZ8rYC
pSLZb385CMlUF+7g4EGSyfqhas1udx6sz0hOkPWAOOkoVjsGBO3V7pw3Tu1uyPP7NHwmn5KGShf8
n94Th3TEbh0yg4F584t0BJqOzazKxrWxl8EXbdD7t/ob/Zh9uaM74RbMu7TKlBZ9PbQJIsdiBgby
Z8GsFYqIyBwJPpLq3i0Kj7ta0ENiyOJqGCWHgqVz5jZ8blZqyWSE6xl+XWNKAy5DbTLpOzofydSy
QOeafm1qoEA7o5Iyjgymwir867QGAQYETiJ5VmLShoWGSdQS12bcxBmcZQtkMUOpncSzQEzczurn
mj13WTGcwU4Kc9wr+PPLHH6OowsNJDGWMYdMIelvTk24TJ7w7kpnkQiWmTopGIY1vLB0GPPf4x2w
L2dyD5jTaBru6py+3ZkijAFRGGK8GTHiDxDNAUpwi0IRyaHkpc4juQQ3P69C9UgVQlY1CbJmoNbC
tvaodYjvwvVBPYDlM/73etyCz16dNGa1gVxf7NZ2Zm7jSQV+9GQrOJ8MwOCt7FWCUehGRrZta9Eg
CmpoLNoM2nUmpg6jIPJiE92QdE0C0+ofP7Hzj3BJrrc7/fwvtdBXuShf9lmSFjcYDOZ8WsUzDLOf
bJ2xxF2Aw4XvriJbNml3NVtvsic9Yj8iKCqBY5rrK0fw9/ZuADoe96vx0SRecm7xlsL5/GwF5UeT
ak8uDk5NGmjjjmXSTyTOSiv8JqH2M95TTo+WT9/C8OA53/2ZoSwPaRxwXmMecgS+vvFSEwvdobZD
ST9Tzf3u9twEVTRo1nJFHFk6SFPqCeVZwsQzcLNlfzZw65XAMRgPIiPc68jVdJEtsZaD8a0NziR1
qPCR5MfL12Et6/N0DzQm1I/NdlLe/iRRSGOySMHQKYm+hIvC3q/HRGZgukc/OP4rILqdo/jqZhXn
VOh7Ey0mwL1RxjZzZejaVFXheJTNQ/IBiTNKRKNH02w/ThIAyawMz9mVAyW4wnPAD0Bqu/xKcdEI
6RIMFWdbLq1c0n77oHZ35xVZ1znE+54NvxiTltIYdKKn6S7xWwTXgW92E7FDzKHpFJUykwIbQBG3
W/u+UJDEnSrc0NWuC2O4cgNdWXI/hbawAFVVb6BvQc6S7UAnWOIsDTf5KIHrRhDToMiKZgNMNYtU
l4ZHSoamdoSvJzIPrAFsI0eL2bT3Z35PIZNVaVHp83dvGQFzOSffbWFg1LJlzWmQRrZb4zqRjNPS
VLNkl3fZtdmFtrL+Y49voI6hY8L1TBkkImcREQY0bjwTR7BNphpQKFZr/AosUiHpHYhCQNCh9iwZ
ZKkJ3S3AY3tIWjV7PPwx5FdYX+16Py5RHrR5eXbzEM0RMgdJ7PcT6L6fsApNf6MmJ8p99e4bKw8c
vkHuy+rrE+sF/5sy2iBqnpRnh/BjctirsnddJo/I3gWO4L1Yx8SqgC3o89BnsEA565VwB85QZGfZ
/NBHM20fxccZjhdzBIWT4DDYwKkcd25HWvigUb8WwCj3T0W0WQfdpT7c9ajB8ZRF7CHNfVz3NTcZ
gsB2MBsj3qmLod+VINiT2okv23tpkpOO0TpHNGVq7Tm+T5K3qsID/D6DvV0xwQyzI2DHAi/bgQnD
nyreZHvsnv2G+w6vuemYlFC48iHSwXp6bXgENjUmavNAlthsnol8Vypg5nBrdWkAqMBe4EQL5+OQ
3SV64QtB5pONNrDfeSaK7WFcvXK3FawIiJzcxmdARAFIFCDltLuUWUXdY4ev1H/3I6xr886sBo+G
ucgPQSNdDFszpaWWkVk/xYB7/48TzsQyHFL1B0mI1cd+eDrdsw9vuYVsyzmTkHz/+Z/9NjVgU6gi
USqgOQ0IeWwUUUbnX0d2FWR1wmyWmuo9kGPE0UtdSTNvKXXijThMpcZsXbWQ/v6dJQDaLKQbDakP
OQrnytyn9gE+9/Xlk+R+lsAiPsLWgSRmS4ZQSdI4K50V/hKLyVKT1dY78/xSgrKOyhyl9nor94tm
XMYkP2czmdV1ni2du+wPCyluDhIP/9wkeZ/ufE+8opYxkzl5nBn/58xCjeT/hX8Dj3IgWeXXvyPO
jf8RoMBroSwQZGZZpvlAFsy4kczFVShBlOcG0e7BAMQ+eaRbt5M3As+i+MnMwoIqPg4KouDt/0bg
AX0Mb28/kiCGNYWOraW7KGwLpJO1AUXqYcocnGPNTFMFNE/ASfox0ZkPaScLhvf+VjsPrbyJYJik
ZrBRBTXOvb5HJkiXtxJq734+MSbFZphoAqPzHQK2dN5vhnygV1n1ZbpNe7mQxtO8kP7K5l/P6AoA
f5HMcjMNPpxFHEKI7+MeNgxPNGm2Ubt2mgZaSGjAu0X//2LV078xL9vJMDdNTgxbdi+IaxDXU8Nc
eXXztNDeRoIZGIxo4ITeQb8+ND7e9LgTnoPSwztWCnCi8oVEHpI+jYfCD9R5YyKzZ7tHsV1oL2xZ
fMoNVqyxOGeCIbJRypAluPO0XGuuy+eaoBqNDCsFPlbCsNX2/82zRhTzyNK0g79Jh7QwaIUdG1Ha
gS3wfEqP5A7BMOmMLJU6DWznqjIQ4o8RcsiJPUvAETA5GkFn2Y5Vm2Ze4+FTPPc8h6kqpatOhxNM
yZyDabhYkAIP499ktlSmZ9i1NrTGatL5ZstOPYorvFd1NtxfDIA2MxAmgx4mt5RqDmDNj9Wn95hO
UL8mTWAnJSuZdBeXwTqgyXeHTzaykUp7cUeroIkFrd/rPOPuEkqH+SAZNCxnrwiV7hoMYx5jeKGn
8FBbSuBwX9faTtz98ZDIoHA9D7Ho9+A/aJENDSQ5fL75MslyW21swnQh1xx5dn6Ubm5EsD8hxFaj
MJRKpcopp9C23YhLfyKHezqib3F8xrCVsX48mAOJpU1J5VVQ0P5ktAr3cFgb5wKfmBtWQABgP7bx
eTMtKaBR2aMnFlsfWXJPbmGQvhA5bMI5yHEzAbk8q0TKwJ5ubVPNVhXW6BaR2t2X4CqDyhRBr8Kl
KLH/OqiasqVpOWx0T/d7q8cmsqr4ikpT1yWkRx2elZkIkifGfd/B2EIN55WPgwDFaXZq4whu+9DC
HcI6EBEbirFnFOSolvrM98H5crN2rSHp2DtTzuL1XLoGENY4UTl5d5K4nEfWHs+ANhfNhctTIz23
VYrbEVl1lCV+s6s3p+4MQoDux5aFLB47L7Y5fGz0ODhAnGcg613eoZh4fIxveL5rQaz05RF+pRx1
jU/oi8eoE2v86dgX92ViAq7ZOGw2Rmzwq+4zC2kuRkM4gvQnfT4iSh7ih1FdYyKCDWMj/Dyh3oqZ
vl6S1hsTTV6MQfAPZluzH6Cq8AENqkfTQWrl9pdSptS6M7DuCs6zqYJAo9invAjKeg/YlgE5EuHE
jJp1rDDYP2sD2Hu7cKzpxCYKHAJ8kn3eW1JEPAQmHOSdG1OfWbEoAQEuYzSfwdybuc3IWH74J59a
kaeY/mRPFgQOvcX7xqwQNsuOJhpHIrXDetEOTnsEoulGavyagIAer2htFD487Kz/ObwculhAoVn1
rQfXS3/HXewVXR0/ysJYy/nsvk5uGGAcY3zmZpoet7fJuXWFyij6ZU5dhe1oLXWsMuedAQ2SwmGL
mbXrZwRN2A4aen52akB0ttksr8WfRUba5SanNebBRnUpRcCfgpqgsiLUZpOk75oT1H04+q9Zjz1T
nIXNv4a+9e8OIxQ6+SDaLK7uEjaq85wbkG0ACusBnK4L9NehfrYUshCDFYZXwe6NnxzvVpCe0Yh5
pVPKvDkGG6UvQ0HPM2ah+ie21Ci0RfjoFXJY6KwIbTBAnp4jnA+6RGaF4wesBmyY40aoy/Bt13cS
vnSv/uGbf04dnoJVbKfD5sUH30xrcvQPG981eq9IkVeqEoq/RS29twDJnU62ZVVX5IxbqC/QBza1
wE+9lrOnEn+QglLFmW38K/YIn7qbFBz0S9bkPHqXiKZpcaApB0WbXtAfa0B5GW5neWirULsTj6JY
dNmn87ZsXxHiApl8XqCdlKJlte1cd5kjF+2WwBGDWkszi8Jtt1oLQXjVdTbsve7WIuOfs9Ywez4a
xH+EyiNYnUt4TfzaZqzdmgoTqDTbwLEUZEJugcBBP0RsQlMiR8xGYOkC+XE1tq/kf66Z9bEtPCaX
k+Y9ZJPWLBT43KwJ6fyG2+OrR/OAnQtH9z5j1pcQ7G309nXsjbrhdFipfTUydb+zCOCHmbDs/T2q
U3YDKneagUdnx3n7HOOdWE2Qn24//LUb44vPKx/e+QZ0b4XCZCQYyY/bwn9OQiRRYfkAnOagRGJh
+j15K9e+EjL/JtzVvD69kMHy7duQ2IDALJWkCFq8dKlcDBYpVz2lZZud719cLlhF7jgjDf88+ION
NCtFktPzpnufpAqIR/+cF1nuLfCIiGAe0jp2Ke3/gfJMcBwxfLsYoy8bKHT6rItAPfwIKPki+7+f
U8bP2dHAvc8J1uCKx34NqAkqEHJYPkv8943lh/vE+rD8w5yANN6VBC2oq4OatFdN7sMuB5xrHGDO
HxutldsQsPWWgNMz+s0d4Ynxpx4xiGNcoReef5cfjEs2yQuglv7cifL8rzmvMPTNiEfKIVAdMm8U
R2fwIaDKo4yM1Xda2u11aLVrBBty7spL7mFNPZfmm2/utdWFiBAduk5ZOMgTkR1rq441SuxU3BT1
bgrHT86Fm34Etig8bXDcU4x+mNvb2vz/TL99okMk/6bVLNKqWh9CAgIlE1BzcrtgNDD6uuZJPPK0
W3jaiyMm7evXshTjszYfrzfovTNFk/N010ZNTonjOGjF8GQ5lGEQL1Ev6KvdRra3ubvVl8ALV0To
F7ZzPH6LIcWkq38UdK8XXAS9iedo4aHVOm9gM0YqB6oZ1s4EcWdfM7TqlsMbnv7vApcwXBsCQcfs
D1+3lJOYGWLyjGbnVNOvOTiaEPj/MZrzDqyNL3gGht4py9ljmzwb8TtqRLStzCHeTNLJPf25vqh9
IEsIhQmNVf/p4TiNDqLqKmeKYSelPtlR/Kgfmj63eCLNyCzDCy6DO9JJMzr8Wh22bMguQa+WJnId
yhNipyFKAuH3B1qY4BHbRDuhfpiXH8KfMXx4nCiqlGKsKweTxglW3mroUJl0cMvDwL5iMx5HvsLL
oD43BbZis2jajiDtxG39JLbHFHwVGU/7GnQtP1GbLkOQ9aJc+ao62ab5Tn8MZifW73X6E1GrHQPv
CpMhJwwm1a5C92F1IznIlcwxSaDhEOWx5D1UVL3m+t5YOlRlmet419tPxNTg1Z/AUB8x3AHx3D6k
0H1cQoSxROBXzfAoLIcPjUyMQ60AShmVesEJnvJfhtnEMbf+SCFqK1RimZPoRn6KEcd606d6zt+w
0q4SxEP5jhxCGTxFGwArrkd8v18eZ4CMFqW3/F2KF2TXYa53nrr86GbyvrtPRP7MovDxhnrxAPJH
0VQj/qvmkKbxb5XGmyR6bPOkyJXak2Xk48x4E96PAZtf7QRZn4pCfwEPq6rd//cts9bHQU6a/CEH
MPkRQqyzUKsM1UGh2O7vSAO4bfE2qRd6sdX9Qe2edkhDVOWVfAcwkB6W8KOr8Ipp7f9diRm+uLSi
aM0ceilfMnnjd4qkU35LF+3j/IJLUXfNoARv+xs1MBqF0NFp9Eaden7RwaV5o1j8vAWLsrI0q9lO
y2uMVh41I5w6bmSu6pkOMWG1lFrbZGTnngC1U6wII+wn/JE+cY/SLEj/TK0QtieXMKCd9CH+eBew
1JHWgqD0VafJ9zDFa9cAGpwItPKNaBfDqtWLkCqvAyMq9wcbiY6bff1T5xppqkp3OKStorvTLyjI
UUdlIw39Pjk1JsI6406chbZOlkPKwSZvaR6VEREeE9hCYS9FErh5SrdtlsxiMcONBEzdJMfcGPkS
OXJbZPGx4oEuCSJ80xr2WFth46/qdWxx6GNzBXiI74GPdF/95GUQnp7FUYIgWoMJCeb20TMDce0Z
UBQbgKnFXTxYrueldFDaznfM4ouuJq2A1rhq2C7L1F/qOPrOTh9yzUUTT76PiO996+NPxjfMBb2W
WKY2KGPus0QOZbqokcbTVDQYhXdlvqD7dJFMjyv5ngx1RYY+nKI4F5pb5Y7/CxfejIE5FzeRIUxi
KPgBHNGCm3LUpxstUoHncJh4v+Ru6+51xbtc4MgaGbfJlkMpujKkkCusqUc0JuFfJObyUFr5yx/1
KQGwogMshfSgWewpOqY+Rvq/KTD+beT7Pga8TDizPNG0UVSNXkEBWVNTJak1DTDXvm6H0RaMNW5N
EZ93e3XSjfQfWFw1aJJyN89VwKWSo1RM44w3VyYx2jNJYrKiEGDxI77KfPzMunFWwxrHAzrN5GK0
ZXzpw7kYV7fKVLr0fJ7hM8DNkC+1EXquC4duccEeo1Tgsg4xzWkLiBDweLaDq4mkRpOgg0ZtdV4+
0qNfKn4BSRvzMibxAxCTT37UrfjDpVeSmcIR7g/7gDfNHD0PidB+aMPruHO2mTETrOMKBcjBPghj
9EPmmGZOIqhlqCJ3dN1xiOLeqgYlKuIL+4XfGPRyEdSeQ9g47eflZ6nkQqgvPgphRA9WHePkvmMy
UvPiqnBLX+dyVN0L0yvAy5TSnEzDo19gDcfWEerEFhn8etk+b1kDa63gRYCCzdC+56FVI5XHBMaQ
vs1uMLjycjZPJYjZeg7S6C7IrdexpBbkX/TF1UulotC2GOPbrLey0gBNYWOweBctGjzX14aX1AHm
yGXFvTBHUDswUHEYx5TjUbVGyKFmeChkcH26L+Zn92wKxr1RWo6z5LlJqy3M7x2tEvX9SWsvS3+j
JmU9vNC0cblC67JFW8AC1GYLYFzHv3e3Wd3RbgrOfAg21vmhq15GbeT4ApHrOLie6bozxntCZcDH
9OUtXYSowgXwNFgSCMYaB3MbJMDEMSw+/Lg/zWZJydUS+5A7Y3CRFVVMaOMGbLpKLMlBKif1hPO5
hDcUesUq4byl+OFRXxQN6VE+ZAFM5iZOK3eCGHOSibYXhnGGxyvwFSmZtIwAdObtubm+yuPrkc5T
PCfm49k7POSN33ftqr7rVX+yDufNTxhn6F6f//+l8TqAzJCxaDwfdvqG9XnRIOT2HcyAQaLuTP8K
8hnV6fomlsY+Hkbre6YPwhAS+LrR4S1/eSs9up0LGS7CsmWKquGfAAa6RJdu29qrbfd78w001t47
p6Q04GLKQLuECGSVs+6a7YNf0HE/o/kuhPJcPSMvRs8MiqD67ZFvjGv7HZp+0kRf8v3T2d2x+Se3
ly6tZe3B81sQe4a0db+dfifI1l/kZ81DkFPH0s67gHaO74T/laosNuBn5cMZNesb6ZshSSwSp3e3
d4qHjjQ+BeWcAqOOKBDO2fBCG0JANgyCdgvQKLhZ7zfnq90/K3BRHTfBcjshortAqD/yxay1kRf/
MshxraSJTEhRRxsUs6usdj8mpn1T+kT28xfV4kjn7yiStS6BzFO+qMsFMCR4H/qdoJWQnX9RA3G5
cOVFuIo88GB9OyCJYznyxUi4vIC+teJO5AElYKKj4eAxejEaL1e8TSUuHJD8xFD0Z76JdPrfT6Yb
HhSFGmlieUdkewOcotYsRaGdTM5OWWojLLC15aT66I2Ouzah8l+czqU7FYojNM8o3GgWBrM6GpEF
pdaeygWNuDRtWi4OmsBIv2xvPZGTScpLBWvyLpIFRg8ssO6fBsYa7ak3Q8FiKHqgxBcxvlds/mqC
2Eh/08PDIgw+NgB24I75M9zc2wsTerLGofECvAuu5poHtjYzf707/Gu8anfDGXCgovpRE02aFQ9x
uD9JiaC3Pj8zMRA2yZ/3/0Gyv6Tk25eMQA9RaeX3BD3O3uagEwvxbEEcw3rdqkWJDk4ZbkHZC09I
EblxV82TZ+B2OBb9KWD4s8SRbupsIFooNaKjfq8R4clc4+7pCKetZTH9vsMLY1mbrYbMTO5IgVNb
EHIepmA5xiUtxbmVEM1/FTfLOezSEOTiT9go/e7kZuoPOFRyrbTSrUw7BjcjjxAjtGvfRokDX/Fp
sJWyEuVIgY69rgMnnUrWBd0TigULLG6kUIWe9hnhnCTTsmLzKuoLqfhuEGE5kmgpaE9dMWsQbzVB
WvahNfVQTbKZrwyJqKKUfnT5XBRQw5yERIQjKbW4AjR+KJGmO3pj06neXkM179QURNQHTAFd533o
yN5rq+/2naRzaNa/AFZk37TcqRYmIZMoEw5qAVMgZVWDW93lCZ6EkyNsONphtM4eXxMZys5hXRuZ
pq1LzqjS0r0L5wupqsOrd5kWfvvqL8Uib8WeuC6MTuhJCWb8ZXpqWleheGSXm6M39xfU/l3+SJRk
K6JKl6Ei8v8eOyKWQ57+57MQwHyUe+eMkIy+eYnCV9yLX+jJpiOxMZYmn2ibe3lUd84J2Lg+JQuW
M0thEitR1/ZG8RP3VhkcjgLtEfa1mWQlMzqzmjs98golL9Rv19vsrvTa2W/Qb5HSEN+rNr6CHpDL
LSljD3S5lSta6Kpj+cDKlx41rWg2IAQ35pIZh7racmnS8FG+A9qiL8xYLNtZpPuIkCjZ39mNqm8n
VXg700IiwsdkhocR3MRiAmcH58AsCmyKQBnK2AZ4iimhPshC+fcNETa3cMaH5pBSz2Hz/kJfLdDw
rup+efdtfSVBSK3zSSKWtQgzj4PxbOhc1tVWuW1su0W+PJMwc1hkW2BnU+yqPHnNQhf9z/T0Yz/d
9TGtrl188O4KVuVf9G/2LTJRjY9Ez9FvSZ5Rf9wO5OaWBxIlVqU9JdBXEIbeAiM3BXNbQNaluGoo
m1YI7dCDa+l8aQa4juukFRj3rc+W1YRSJXabiw/OlGhBkMefcZNoOlXfDY64ms+AGyjrwXBOy874
TbrmSJscjEktq650XvYzYif5vmxIh1Q5Cp8zrVRvXP0mOAVFbrx/0nPOhI/D57u04luTv2w78amz
PkXUOy/viq/HtdoYGHZBAgmCE6H2EqtOwRZ/ZaeJ+UpHBl1Pmg2Uoss3tF+I7+Tois/HcU/dgMfL
BEMP+kunI6tF6WtKcDBqkd9QMT5b2c77G8TRWn2fL1bRlQFt0jNloNVsvKoHQh3QcglkGFICYDsk
UvZrTe0vBFM6LqMcep/azezCNkztWentY8+gH8pGM2kazFRsA0GM1sH7Mx8qu5XZlSTuNua9LtSC
Blo8toCQQeQ26yLGTfrPYDKAGaey3/6TND9r5+gQPgSQAzP5NKv/HbKvzKxFtI/OJjVpPq+pPHzl
+QySyOHDf5nowYPaCnfihB3+A8kKHFm4bpRbdF7znJO2twXjQ6ntazRp0QRBPfUp5Jm/AiGenv+N
4hhCTff8QRADpzpgYU8Nr3SoBtOBFET8xfebRr0S8UCUw+x6KutSi0RRw58Qx6tw9CdqaqPFyxTL
ZFlLZ6bCekDeX6LQBTvxVQE/7F38LV/1Wfuyz9Y4oh2KokH9Sgsnj0fAiqFf5wKqx3V6HSQjokUP
y3ttABWcWAkUAYR1UrQ/MY1wKPkvHW9Qy6mbZzgQPJs19SZd5n7TWMTFzDdBU7tmncm+dug8GSEH
fBvWvavH5CiclPle45pYtiyXHDIRAoOlcmzAUn/+Q45imNluYM7J6/jsTFJdTBnMIZvrlYHOafZF
pFprVBxuFDOvmWIcOGzXCjtYCQEWYOEzuXITYhyLeRK/UShS6p9wNa0SruPb4f4txkCGSHjj/jEF
1qcFTkq1SC8Eb/FXdBU6WjlqGgiKsbKaD4Po+zQNJot0BoNVxxExeRDl7VCpwu6J6DqC/LLDk60e
b9xvIoafO24tW736Q9D6xeAzrHxRJfXfKt/OMZi4XLKVz4pjg4pRIM3Hbolo434cQXl0ra0pTQ5S
i/CgSGI/z5LjptkNt1VeyI8Dhd97mwuGkBzlVMkAWfZtOFpJ8NfT/wJXxSAyO4X/4QEZ8PUPicPG
sJzudtQ36gP/JIrKUXy3lfYtpTRTSaGHK5sgZ8DSu3X62YbEU8knmGZd/W33UnmxJGHtX4PMhQzL
NqPZrVSHBL9q2NW+vp40LVSVzqThKuU38M4aFkTUzk+s5Z6khN679kssOjpeSlfK9GDbh0xbk1pU
gEd2BybMnuEBcu0psvrKK1DFHwuUHff4NJJs8SLBsjJa+uerq1pgRlyvVmW8BkiwGC7IYrGbqEEo
zpO0+CVP0UK66mOR4nFW9VFvS9PvI98Z2vSlz5SAd7Sj2HhMTnm1PpPphvg4yrm8QvOm4ZROdebE
fNwM1bNMb8bl/PIqVD7kYmMPNETnJqA1VYL2omj1yTQ4sYjr01lNfT1Ca1iuMy1+Cmv/U6wPO8GM
T22BtzzC/2fol5iZveBKlzVEKc61wbwQoHsQVB4ScrWylKJhBTljFaHQsLAsPr1t0TJMYCBoXFiL
aSa5wa9XtnRkZqhdOrXA9wGvfJMdTxjJdOeUHyoZIbBXGKGnArpzaeF9uh4djpGaOop12yyLQu/g
70ciJ48MhMTf48xOmFXkA9KEtj6UOvtYPXuKw+JCwRzxK83uqmYN5gj4wPWrh2tjNoHwgeyK5pQ0
XKm2priCfLz/cJBmECQd8C4u7AN+c8pugjN8GOwkEFlnrjt2MI+1zpzZXnjHcvV36g6LdK3Qv4ex
eYyLqRqKxvtVFHYVsM1SfGaORg32WpMMDT11aVRu/6arBOMXNie+Twzlka7oWvAYxZfHA42Y/uT7
Hwj1g8S07Yw3fPnt36UWYk68z6ge3uXDK101Yd/rdKTgHRxnENc6NF9MiX1imPl33DQklR5Po0/B
TToqBpVhPiNJTH30qthJV63T0sYRPfFQ8ADLcUoa9OycnJP3Ud5vrMqlO5XYi9ng9oINjqO4Dmam
fG7wHu2cfpIgIOlEV63GqsptYVFMUOouHujKbncjnoiFKSaaluAj70F3Xw9zQ7IJIXDJdIrihjAC
tQI4b0pEP30KedB5+l1lQlXdtteU9qGP4EfnbUcecp65Eq6Qcx9cKG+bw6UUTDmTaGNpUQuEf+z7
UgzjUBY6wH5qtG6IAp7/e/rzYgbyAa9f9a6Zr1IctgreyqQ6ZGm04gbshT6Hm8kLNaY5FXxV/0X7
3wCbsQ64k60vxiCplx89dQz1gwi7C+jkwQOuJAb0aiErUjkx1UXTm073xgtyMf9XMoq4UtHdkwOs
Ur0xuVpDbOv2zp0EWmI3IEy5U9qtJGaLiaJ0g/LTNmTehn3Ey3tJF1Wl8wBpiiafD/Hbxn7VnQCm
y+HJhqHmvXFIb88XhwOcC6YjDvTWMmQMZVpw/HtON8lQjoZNLzc0sPxdPwXgoai5ZCqffKIJhVZw
qVh0NHXgv/rOZRpX6BWflNuKR9Vy+g9tXh/DFwqZp827ANb4U+3yx8g7m1NeqfeQkMw4wEbX4Tzx
ScGp+Naq/1u8M6H/fBVvfsPjK+Q57HmJgUGbKNAbasXMEKmvFYviPNCAOtcXYVuQdaHleviLmtSj
MLBOIG1AdnHC3I5mfER1W+IBmu5NHTZBVxTWJaJbgIUc6vTzDfS7RBeigYcSVnvsQnoo1Opw58z4
lRfZk4fBdRJdYtofnwKG10U2Vsuu6vcc1yjx5NG2lfrpfZ1BBlrpGW/dwhsbVoqkU/Pm3E5wECT+
KPYjUDyt8gfr8OiYsOn90ibmoWdDZABV7D5+laQeBz43h5rJ7GTT5GHOQg7SGWa6eTDXfoVEvLDS
491Xg91SfbAPctPY61g4F12k3NUOt/j1cb+kvWNu76wDMCSCc7+SMTRX+H2Yy3YUG9uJOTKS3pfT
9W/Krw0IkNShtUvA4Kv84WfFz2xrYaa1g94tpF7Xb1N5RmiMGVYsKGJzHsjfQOvNAk66SXwnbhnw
JT8Ws/eUoTp/2NA6CvVNdzxOPdnCEQym0rVcm51p7pi8ptyjMT0IzrgE8GtTTM/+a5H5NcLsiOji
pcIuyICZQhjcyhkshlQjRkjZm5MBRuNFv78xx7bUpSAZ2mwBgyY1gT+WE+cfN01CFk+w80yKPNca
uXtZ3/CCxxuar5vgyZkFr5guKytr+GER4juoPW90qSJplk0h5diOsPkeX5hhQBMmJ3ttCF0l39Lg
sAglvIrLwmwUVNrGdtZEuexIUxptAcoy9XVA9F+PrX1qiH/PtjgNGS1jwuFugM5aJNcL6Zq3oSQV
JSEpD7Ox+lYF5S5tI3zgxcoiphXvTbetQmtfm5LOfHe0ns2nSN+CC1GG7lgT6gvMLxN/LaKbY/0Q
+0i5gjoXT0oWfpprV5AKDoqzE0mGs0pM7zh7r+WvIqZ1KQZak6eMenVyoLf7slrMZPubLZuyeT5D
24qzxOrF99hZexlfKny2WhZs5KIDTAX0aBGmvgy9V0q2z2HpB6q6ZWO+k7AabpFVbtyhgqFuCEyQ
s3lZTOTQO4Erij+7UgR2WwgHe78x0ryVIco/mgvFlqJMTBh0IARkC5GHnHJTO9ZormBYd9qJIS4x
AQDqNAuhGTFRj60LZlZxzsFkL8u+cvCe1nQIqrL/ysV1RxdVRyCsvm/nsEH82NYeQh5+QeMZJooB
OuCZL3ea66DLslqYYz370NYCpqK8zclJ6kWg1iVuHuJbttST0bDLMlF0TY7cFfTZycWnJz2Nti5i
jufVOC2s55Qk4r1fVf6FCsocMmp6aKVfvkDnwBiChlroynMkCkumnXC/c5f70eL/p3xD+cHSxSCI
2qyzeSKd+2fUQZakROTD8aA4TUPfTlpjhvEWlCbAZxnKVV60m+G09N54RjrMr0NFyjKxNX+dyyVj
P7bHGCfaLVudddiD1z/MPqS4ULJtVG4noUvRbEl+M4TSB6YgYLHFdDoNlJ8cmTnyD86eV6ZwCcWS
OB5IGtyTt5FL0XM3Lfs46oHgXBN/GdxjTa6vCFgTENSKkheXRlqVlwdoRHaxHXRjkfoYAKZ0+Ee7
eltbGh7pBQcJjFdGbra6k1v4IQbUAwkj5kMMZjfNFhCQ9dBCVqyHL/lCs5kwAhdSHroa+V/eEFHt
ovHW4OgwyKaPhOY3tST1FpO+iepYMM3Cm0M9a8Eptwiucsq4iUzP3HI7kst4ldbzXr5qQEdBZNSP
6uM8snSYlrT1a0KsWs6WJIGle00fzpQxHz0S/KDnkU1MVM2yvb+4ZF31ryRn5b6wUt9RmYlM7B8x
wuUxNfSCA4EwYLF/y1rdkluHhh2qAzwBM1SivfF7Tm21IM6WjS6TDT3tKwYwsOWa+K0uu6tV49n1
wB6aSE7Gj/8j9Y3rqmmOsuU8sLm3RYJ+waYGT5i1Qk2d2WQLkwtMxrdXCBzSWvbnV52/aT64Rd6b
Hhx3ZUYUqbl5o/XJFTKqXqIFsA95OBqPLGrNIkfH4tbQ7RnjQg1hGVysZwRpuqrz2TMaX9CElG9w
Nb2etA3qVUWvlyTCb7rWET/0xxTnITmi1HI7BNJ/+gZsKmarl8P4LxLoK1zR2ILV+4PSnajRvenN
XW9qvLTVx3YY7yvaZZjMxOfqUm4GPwpNBlJp7Pl7+JstVq2TEipXK6fCfXSvWeISqxi4E9fqlM+M
7xF5VXH7fTjvtw1ImGmUum8Ialp6/1eZaxLD31Z5sUX4AR3nrJf/cwP1lFK7Rux/2Ddw2mt5qrcK
n9u5nULgJh09GQQ3zkkmdKktmwHUXvhpT2bCt8BTBzYvnBfVT0LX6taDcSGMYn8TO8LMUSqGs1tw
znrjDzl1Cqn/Twk9Qdix8HuePX6T7BdsMNNbP0XzK4DQmU1RDMPeoj+VLPNz+rp96qq85/nLRCYb
OHXOOBjVO/pF2JY24bGg1ony8uhJ2DFosOB2e/3nkL4Iepwfg+Va4YroJueABlGH+EQEndMhUj7t
o6zTDqyJ0Jl4vYEWEucupCxB65J+dMjgkwBBXe4aJN++fzUy+RWhUb4a8TwtzndYhgcnsBic/NJL
BVb99FfwHHWIeaLPFtEmigwC/R0gLZi5tibY0Xhhn10AX0YycpcV4W9Yyf3ydEPvoT4sGITWc7ET
cskIDu0SoAdBcg8fhGFJJ25qAzNKtIcfIDbYc40QT0n5++9SF2uhFxvj0c6bw/u9JKfih+KxtULs
oZhF8w3S7SbzCA8S86I3JbtncUraYs63zeB2Xi5o/LbHsRtbdUDlVs9q1n5+lDsLn+T2zaDfvEQ7
BVsCrYZAYaimdtokpp13hyCv56GDdltBNftQiLs8RZ8rtcy6cx0tipaAxgbEM0V7OKa4lkWAQTwY
Rxtb3dNkdEbXMRzw9So5+uc28cVx1v6YV8k0fsg28y19c25snUNrjyOgY2TXfjUK3/0IxJRgd4hN
qRHRjzFxb/PVU5L7iVY3CXiMSGh9cH4NxonfmbNOTa7zTdz/pUluHPieNeiTYNzli3Q1hsCBY+mP
G+cQUYgXlfQ7OJlTAHvVQL7V58GEis6kMkle+48pA4NjI6OnEE/O/fV7A1eia0wI9iXzORS/2YTq
frtNMNG+mVyhMIkH9eFkrC+xpFNmWivmIdT22lgLlj9EBpbjYHAe8bOLFzlEKVQo8ZE0nzOb3kFf
WCu0cqCUHBpxdmG/G/E+UShXaZacD44QcaDCPTdFbrBdfQ4cBanLe9uBdCtGgfDRmG4eU3POWoJw
5PcR1Fw8yVxCdvbvOdQ/QYneNX6gKPiiGPqp1T0vVYlyZ/SsnD6swP2ShYFSlg1/KyH77bRIChFx
5NT4NE9uSokxMUT6tbKr4vJS/7PqNvwHWlqISRBpbmq9Hb1iCdyuxxTvDtIQxkggTxpBE0wsXDHZ
kTlxUmroJhyyVVBAGwtpJ3lV5MjonEBm8mHqv2j8JT0LcIrOc2ckYGL0wFiafBVEJVFBwHOuLk+c
AWYonfJEmRavTh6StHl9F3TR50yrh7MYpICJ+hohyxIxxQIE7ZfwFiNrFvekDZ02rwNvd//sRuv1
8bNE9X0Em5uUN1RsRgqEPsQAW+QzjXhMUu7luIqYQaVkgzS+z22aIEe91bmXL7YYMcq23xczVALS
KWQhAwWqrKy62nZed3DdZlRL7DF5v1y+wIv7BeUi9IosMmkEOmGtj73mo1AicuJyAVFOXSbr+WXQ
WGPYwg6D0WP2WIbECEFXZK2kHFV65fkoqca6i2yefqp6l6ysuIE7vbPHyEGi8RDGWBTiu2xHjf2q
RTjXE+nSSq1hsuiyz0wjS5DKeC5nfQgkcFRcS2eMbvJnDDtuNUEFfNDpFVVx2SKvhVnfHrdoifev
UjwYD5pPU8puMU0pPQMD/olOBXxq1d0Dwqr6lfvRq9+fEWmsVtqNYqMH9ZzzrIgnele/AVuZE1Ni
cqPM1ovbJB1JqBIu9wKhRlDadms2zeWlJJaMJ5OyBPYIBX5EoCr/BQogqHFLvX7jOQ4tbLYvgCIE
yGl/5N9JjYsB8AqXl+0o1MMUlOdqBC6vfpl7RAYNNiQm+blb+A71hVz2ci/sdeKFOII2YJb0nkJI
4K+QFfVV3P5ZlkvN57QdpgKbFhUNZqUKyzChYTSgiGkm/ZEe2W2LzThPOwl7pvuISSo0EWJjw02d
KUzonG9wMzNyQhYbsSusMQ/F53VhptfUxUNijyyVSAV/vx40Qii0kK2wHna6mddAxD2eYXDrBIxG
LL+lu7xFARPjYs2R+LV6nqrEL79piYNCwViGdhyHq6/PGY60fOD6Pip5saC3ukwZOXAN9A8yPO4g
ggOuftfzyIVraLPBILbdGdkhukNctW9BstEXeQWkJIGsKpzUmGk6z9tB3CfCvPT6zFq3MwwEI6ts
ITBAZpK7U6UDa4TbbBo8da7hFgH2Pov97lH8Dq1GMoFx41v74z4BX0CaoHvnk1Rj3V9CxDkG842E
nDA78bfDSBrXt/Oyp6ipMo5l0j7kMmlZqA7TMy49MXRo1OaFTgOV/1hFl8WFnSsrHJaK/77jxG87
xYRyB3HkcC6mpixN9OMBixPacRPLol5KahJzmuB1B8/RmaAPsHb0J5dPvOn68jzTGEPWwMLur6jj
47lK5Jou2SwzoZrGOQB7q/7be5lEjZptYz1HW3zhiYsUmWDsjUPTF4FmHhvn6xmkfmC4PtF6yZq6
/ZtZO1TOAqxnI0F8Gkyz+KAGu7mjm8K8nH/lJpbsG3IS0+8a/ixWn/AdEJXBohp3X50ThF1Radxa
c4UePoKOVgLsWVI/iX93KJH/GDedkZextSeLn6gjlf1/h+i9Rse99h7dZ+bsDyMY2RFX7va78rL8
+RFBxDWpudrlxGWNyk98IMJf45/ZCrSzKuWEQ8cYYHqAowORoZlD/RSt4I4jOuLOgbFl/dycq4Lv
siuwrJZYKAOiYnQ22Qlkf1No2nwa1yWUhxhbq6zTB2KPi6Rdwd+8uFvnA56lscecHHVfdRT/AzwU
/DVJjnRbxjydgUrZPLQ2CWtI1V20DPeLP5yqYBLId6LCYBDWF+NdfZhUdpHnct8D7/MYbfZcDK0c
KzLpcDQTmQfsPbYaf01cCDT6xmeuqEkzw7urcB+cbDWtejFTip+vORiECU2NzpAuC4rSUNXJaKJq
eFybrPockuHjH/1fW51mmWohr/a7eT+fZsikXdVWlbBVZMgCR/hLbY5fcGmR3eMk9Pe1J6eeJhb7
x8nwn6+RM3BomolfjGNEKDM4omO8EgvpUbeaDIyJ5eoOdaqET/hLS+kagtiiAPa3fDtckOj5RPqu
Ki7dOdm6BALOvS8NMx2/1+6fFI/uL5I/6GsghRoV9ajvnHp9Rzepg2rVJrTMgaK9wh6NGsvrTVRu
BKCTb9AY2RGXQj8VgWcJTz8fOEwxb5Q0e5puOn6w//X2ysAcfKG3yu1GUc67ZbfEtWuVRSZuT6tg
XQqmbTE72uv+Y36Uwl+JxJOEEHs9roMNPwF9hBChHtI8ld5TwOJ9zvVKuMGO8lESsjLKAdGTkriI
UtlhjkJzfhY4Pb5Ich/aChY+r/2/ldbT0zPWXVRKkUoASS6LJVkiNeSVr0f1nfyTL6sH/ij5N2x5
DKodTdUEOrulSmriOOUtfS2H1CHU2lSAtKjWiaDkLe5Gld1a0Bj/BR99P1FZTHMmXawFX5e1cA1Y
10ulppiaaq2bAKvGlUM1QHyUDFfa3+7+jwWIgRppm6eQ8w+rSeWY1wTl+9NpcfWJ9npiMfIW9fyC
Vn5/7v0CDt2QMheF+lEAblUWQqNHZpOns7EZoxivh8pzqiXdMdBm2R4WNXjGW/GBQcLjaAmRd1m5
POTeaYbQ1B/nX7CNgKKhNayqseaMiazaffxexGvKnhHrVjP3K4+bgVEzCBAiY+42dFcceiZ16HfX
dBIp8yyJ0eyXruQs6E4jixGspjBwzgZNotisGXfhscTWAX2/7EjAS3GaaVKLTOsDrs2KxWofxP0q
72ZBIzeebKIIzkNW+NtqiA68cHakY/rF8lTz9tBSb4li+DpSUh/ArxANZdyBOovEAmRMfIl9VdxH
pc51g8jF25pkOryzul+AOuxR0KDrGl6PbqTHgqKJPtZRmxpDu7GfMAyz0SncU9TiyqOIqxCPo5gG
75dpR//HQ4Y5gG0CpO5p2RQUJW4wuYhyVPA6jf4sm8fqyvTq/xuFp7V8EASexzoTo+cpspAVAFHo
oulp81esc2R6bfmdpGTzzBfbPPjNGhJJEqWMa0fcyRMSVsvbUy7T0mhIDT648goZ4B3fVKlyKUoT
MpPxcI5nf7GfKqIgO4TycGIJUyUc4Dd1n5h9QeSuWXca1whJE6VTLjtaeZ5foB7cRdgCnE9zyr7J
1LaxrO7t7smV3h0xF9x/5sPnNYcp6umwfPRlt8HbvkQ4IInClLLA+yXVEWvbdywMwbImO4DR9Uyv
aXcgdBgZyUK9nwk+FGL1ls93kIDFjDJJzWXoveuSHpDfKrN3leXMljNIORt6m8HpVxnQ94LvTytt
kkNUinlBiEofFA8ArLbvpgEWOj9iEzvO8mHar6rh2Wd6vzE0UExjnOLLu5oCDS1a3ljgRZXGUhuA
WPsdZ6yV6V4YHTHDxTh8OTdOZq75nPdbqirHZvgYzR5g3nXvM4JGzLgS2FNUMktrNlQtZCYbr9/v
aigLLhq5VuEgpajX1IV1hK7Mc2Vk3wh83okSOSxB3HmLvBjWIrf/bDDClEM4MkDl09h9iD/Ih8kD
DXP1zlA4C3+cnEmXV7c4K9XFOJrdKMsDre/G9bEFnhQjry6Rbe3+gviSRlnWb9qRgC6lYN0/v+Oo
V9oYjhLP8O1ZI8QBFLp/0ZlmElAXdSxm1KrEKE5+ORrW447YM3iMDw2RiQy+LPzWCsCHJ56Cr1Vp
yPiIEjTxTv+qjaygYFn5v5mtR+wtlonJqm8gBS7XD8/3zW13osUKgTaLkGgXWXR5J8bm1nyyaWo8
7vHVrA7F0l1qdzLJjdgkOIFvDC6+UXTKgx5qHfIwN3/6ObXKhQyN5gk8FiLexGqg07ZhQyqOfuKz
tp8gg2MIJnQeG4seB7/6vQQe7j2pZKtMACyVLeGvHNsq5X4k8i9PhLcXRdC0Tt6g1prlxMI0nHbZ
TSHTmbP0Gviy9Q54t0L5yXoXcF7e6VsBYDHWJ4JzME3vCVnHapbRCELSEYeqwpPQGvD6GHsiqo1T
C5L0e7ZXMnYVs3kLBRv+rni43Edwb6uoDnfbobdSrRDkEWkw6q4fkPBA3F0/J4lQSAvrWgrLV6vm
X+izelueNEnr3Of1KsKwGDLgp3zEBGHwZ1HKOp3LAwf7mDBU6n/Ii00QIAp5PYXVnQ0jIP6FUQ2G
3NZmszVmbNkCPxifmvDuyf1tzZHaUqKFAOkdN8pzYXJ4ioWTAdgoceMSXxWTGBcKZX5TMlpb5eY4
5bEtPyicv4kB5KlcBMdZRhucxe6GCNqkQSpgxj/df5Qefelq02Rj4Q02s0diXUGbqTomZaS2fex2
+qK9G3X+gBu+pA3rhIpTTkP40JKQizDm6giuXG7fRSudA7Jo1Iut7LJNYDNWb8vySBgAu/QS7YNu
6bDf6kGuZUbP59kSAB2cw9kBWyehTVy9Lwz/6aLZQhLtw5unBThN+gpOshkc+TCFqEVtKPwxc43z
ydkYGsZS/BrcKcAEfLNcJ0PvfIfEaH8p6qrfTyZs0ZQNNDsx9fg5AVzss5t/GI1iHq2MKoK6fW4K
njmtyr70uvD9yTHjmMh+3ZR3FxdxxpqwxL7YPX0NritYih/4WRcpGMM3R5ZGN0j9dUHWmRBrbH9Z
H/mk2xi8EcphnYs1dNZsJwOF4Ns4UHuc4WdpNRIlqZ20+b9R1MrY5MeWbmJjywOVATq2dVmHPiI/
jvaljvcRmmG1T8g/3fwhjh8CEpmjKLuaXdrgOOXApXwcOShIkyxAUCAWxLorpgMZCYZvUuEmxTIB
947SSwA/NIvOFzIIYWWV6WfPtp2cP41qbXJ/m8gcGpqYOdSgOk+05VdqUKvPZti0HnRjU40Bv9M/
EZ9vFUak45f2BSgMcDjzjtRNTvc3r0TGZeBxUtoVRgCOrNhGmLtW/gW8YXv7Wi1amISGlJxQt1sl
9xYXJhHqmI4pq8Uja7PFItZWSDt9ATrnE6pjblj7lpSjOtcW1prXicycOVvOFpbI90wC7OelNtWu
dyq/4fAZJeBVR4VnMI/F3dj/e6qB39zRNPbeqw7YKLAnRoD+qdSh+oWNOJEs6AWdawT6/NIz3ynT
En9Quf38coc7f1IYohVU2cYn+Fk0MY13NsSBJmEuEsOoXa1oY+o1rUXx4VYmwx9964xgGqkJp7T6
GgYqbDk2lvUQmpRsRH/N4Bvf2q+p2aHsrfBE19PxK/JGHdefbnVUJ2sNql9PfloSb1MoNPTpGvNO
a14bIJk5qdgOPtvRoAh8K+QeRG86hI9DS51uhc1NwNYlDDGSbeMCePN6j2P28dZalo0Mkyct7Sjs
5xeB3WfiycnQnTp/732EIkMRb5K9Zu6EFEUMxrRx0TLlwZhk9Zt3v69nW3i2DflYRq/RbjIeJZ29
Zl2+9LMWjp4VAsHbOqgJQnYTuOons346kw8Pdk32mVqi0pDSHbQVtHin0ml/LCdc3uspybnOtLLa
JmCfpvJhUpInT/1abq5bZc598PKuTAmGrC2Fbb+92x9rdxG8QeNdYdOPinQCb02kV4dSDrYKz+YS
9uJZu26VoXKtuKaoImnNpbcuXbeDrFtrLsSnkkHaKbDYbtENAC/ZRMf1J4ZU9m6YrXj8LtzcJhRl
TLVl8M2lI80PKTmskmdf2jS3Ekf//Qlzu1FZbFxNlEhT04GRXUvNje+Egs8ghTrlAOpzvULK/1yw
96fPON6mxV7K9493fL3jdXuzvGT/AaqN/3gQYNNO6St7YGXBzAlJDcmACwlTj0bgnUYzWljiD257
V5P8bxT3lKZl9e8uXTqQRx01OlQg3rb16wnLkdBQh1YQ7WVsP+sefF7vz71EYJgWX47LF7cOY2eZ
XTvTdxEFPtIVjX3l3ZJXSUK0FPysscYjQZ4ZgRZmUzo0cHUT4tDRFV+joCzqdJwiqm1uKj9ZTnHg
bCLRhXpYxy5B15HcSaT2we4cZZxGuc6RkHgpBCevVJbC++ofpi6/jBYVOIrX27wi7RekJJVDFi/3
OIQMgiYef1fdTM/Qd8LTAxKBxSY0gEO6Ga90jcT0xTa4RPjWjRh8TYS85UsPgjpg3YFlvIZuH4zl
HSb1cIZ4tNXvbgmN8JXXkpSD+/7wK+d/1bvzVbwUkbQmlZhDGgURZjFl8nbl2FxaNq52NAyeXU71
zUR92XgjG2N2ktNXMPx/5TnYqxU9K6dw2T6q7ovfCQTuhkvR0v1h9d/fEMPMeH0LsVvvOA5+cLr2
M2uOCir/KrdLPvpqKfzn91yQl62FuExZcu/DJYieHMg++2J2Uy/v9gIIgJAuMjdwLm8bHsBpz/dC
buUk6vaCaGIBrqiE0xFkUbOIs1ALG1ekf0PgHiUYdiEnZgsIuXqFzZTpDuGcbPfuNT/rNZm0ePSQ
phnXfYa9AKG/xCE1HZ9F07jT3FJKLHLzPk8DhNKIV4GAMFwxY1xNv57RV1TvaJQURXmyjj/kGCka
NqNCAe2qJMwA48IJnilkDrsaOmThsH2zl0MjvB52wjgIdKCknfaRY7vQAiNZoq0/fspA2OSvOyCl
P5M8H85OHxNxPLQxTPw63fLt0T6clrRIoOwcJGXaDk9Xe1LNBLCXrzEW4buzfvgXOJ8W5Z2G3h4L
gaXo4ocjy1VokljNons5xVv6/ibFdSPHc2CTTnpfWOpifxd5EYRgyp6To/pT8zcwT864suAGlFjv
hVqgAbrB+77MXMgFC6MQNDDaDGqiJzr1MzBAcyNwA+AGjHTpG20yImzhV5L0H1s6IYrk+VxUGz26
ROqed2WaendlCIKiopwHh9W3nH/4j0robgeKiip72hqPCuXyH+2TAj5dAyZR3bif+ROBkXq9ck5a
P7Y+GCr27i4+p2s2z+5Ceu4hzjw2o7SkvehS9pkyzXbza6Obxz/WgglN9a8xB76HLsDws9zzCID6
Sd8xmDaKCsq8TTwmx6goU89uNT0VWJ7u1k7eKnnrNJUJyPk0+J6z6ZHsNnXNdrabgE1FLHq755Om
Xc5mMwpdh6P3V+Y3YM/U3xvMBp15RxPHI7m2gIBnej4BXfOks/59bcL/mD6LaOCiOsdNIeTvcCpw
kQ+8Uk8Rl57B6smQOg4ZycazNLR4zQ44wt6RJ2HNgZwp1Zw5z1Wp9m8TNIBQZ3kVOHEDVuAWLoIt
sy+DkAdkMtMBGSdJZ8+e/ieRjoj0Biq+KC08oZGn5D5XvGWPCrDKcEAxZTPoamZqKv1BUaefbhBw
GqMUBivu4dF4mcabA4+1FbZxkbbizBO/mSofzA7xFbNLOfMN2XfNDtrB5vKAady5pD/RlfvyLumr
aoqFkWT6Hl7bVcBFZsKW3qJgzVw04lsVE1ruGUlR1pGcbDKmiEYbNL/h9y8gs+ZBu0PqRTo32SJM
UrNNXPsA7RmWEZ4SYrKiu4zDR0Yu+rtGW3gvt6tTFQGsSDwQM9ga1WcYQs94zsEpspIUNwjZv2oX
EBPdUIoRU7Tv8SLHgEGjNojhvSBCu8BLpeGezfcF9NtwMjFPw1AdarOYBXVN5qlJP3NK4UWAT+Ez
1srp5TAZHtOcjpQZTLBKvuLWs1O42jHYG0Ufo6pQ7MiDr254VXdY31JcKeI8/ddPLyIm+eEZp4L4
qXc9CIrWcvGR96hctcZld4ndMt33xPhlNEmgMSBpb2puwhMVC8eXFzHASLpCbpoIW+2T2LcMH5MI
f2fLEIDAIZsRduiBbvTMkXcjJ/M6GO8hQCGpSSV+sfgkQJY/xerWafy/9vigSe7aBUJYlg7v3T4Y
sDZ0U7ZkgxXtYRkvJpnS7WQ5mw3VwtGxOdBCEtGx902sBk/53xJf48/45LzrlOSjmor6JJCG9OoZ
lhYE0VSkN6RESKV96O2FHE1yedUinfgAdyLQjjlacKpnlE9fyIefi2bqmD0VGZwU8eJocpSj9beX
qT81S8Nvr+9dMP4tzU/38+oYLva0HiJBLDj+r6/jRdXPDmuKvo29AMLPBY+w0PwyVdOj0YrSp5Vn
ZVQGHSBRVnNUUQTeKk4FxYRXlbHzn+Af6uFTsDoZsXguJE4HOjARPWHCAc2Czeky9kAFUecjdUoC
RQLH0r+g2yUitLFFEmlfVP7Oz0Wqd05xCeBnwMwjvaGkL3I6X9GKi8JjJAb64EqOS2euxfDSTrhs
02ZcF5AE7+8dQ2R6a8BBdX+kRH2nNvGAqXvdGfHxmBcbJLmyl7sUADtjiYBep7hDM/oiWHwOQZjM
JwpB19ukZ1ZEX20WbVd6li8c10daDnVYBNM5qHZyI8OG78K3bxi8sfnkPowv7PA4bv8wNl50OizF
MQ/4PHkXdUR4sAo4Eo2KsIcLKnRJRpCZwgYS6IhM2jBCiu1HdAQPQdVKieIDHUvEeuFYJcYlVqaw
spICeEmxRhCkZdUO8IyTt2lHBigbIVGpOskl+BTw4lX2TguzZAXs/2uClGHz+jPpiJfaxeUkfSAJ
CCLdwLS5cS9rWmtYHPIHCdETtQHUYB9MwiZKrRL1YJt2I6UR5VC0mlaTeO49maoJsFtxkSwia+0M
jpF7BEdEv+Z/0kfuik+LWtoE6CA2uQARhgdOXee553FkWKbseFyyHVhKrZ7IC4mliMDwEv9XvfoN
iwn5FKukBO1Cxn/GuTodkkW8FCRdQ1iuycz9M7ToeAh1nsvo+UrezLP9Hz2VUs+E4LqeV8FeUTMF
1J/60px2t5LzQ+1jQbtLedwXh45J+kN860H+hDsBqpyJsdg18W63nrQv48d/5DN+P30Akhqis6F4
BzB4dQX+LB7pRTwQThamIkIDUEGbrJhH2N9j4mR0tWCyr9tw9efa3+zKSBmjniGd3RTC+U+i0bIE
4PP0zj43TV1wxrpTyVmZxPHAd1P3zzWmykmWxoWjrvKBDJLCV7lgtcojnqwouTOdf7cHb1dUqQiQ
asc6FoBZlQnVhmhV27bj/YTTPLoLpSqZEfdHrEesbvcUnlUrEcR8X9hNF6osYz34sf/KerlWeKEc
cull9+tyWPUn2fEKovA2ixMnokigEEAfu7LKz/TOh8F64Vw4Sj118ae6qJ+54Y6on7ntwcN9ByIk
ag8/TQ7ynYnICIo0KUSuwwNbks2OLIMjefEC1U1AvplpzIW/EKsQjYsV9k7RFaxkr8CXBIr4vu0R
tcYQq9kkemwTTBsSOHyHI8q1iIvsGNJJGqTZfFbWLBHx52bqXI8BV71QEcx6qqLHGbxj3DxRfaWK
F5bj/Y7GoXVBNY14PAb0mc6lZ/fDpaK1qz8rLwuorJS38y38XOOMdvbLp2ikgu+YDuevUR1+c9fS
FSau9vnQzkGG4DIUlDtzFghoMbVqBAQaviclBbnB1uRUJ8/Odefaq0cFDLWdHsk7x+DXBT+dNRya
vUdiUspR5Um/WfHTavf1cjfCwbkTju0YiaWtwsWD67NMB79YRE++jm/50JkvMdDILPi9InXnaaFk
c2e558Bd1fIy5dOgLKXQqW6xVSrffgPzg76IiRr1L5Cz3qnUlLRwfjIeAC7NtzEmE8o01WB7CwOr
m3TwKeQJSHkf6GTDMuhANzbiYtZFCFKoA87zAfx2qFf9ASo3ucc5+9fK3c5tTmCBFa8H0j6wll48
TI0UqqJ0X2PrdX40iSQHhlIeRUoQa4wp8hMLO33PITCfGV9+sRvmbduSJYN6IIm0uPtimrvdPV4p
HFlP9Gk6zaPwV6DK51x5g0xhdeSRxAODAj7aVWoSTihzEXOsyN/jTZKoZSvvvbX/IABGTa7AYH8z
8UT5qmc3Bhh4B1EFVgLRTxC9exmLBkPOUH1CTJ6GpybDfLruJCOKNxTVVwwMd4NFp3XcWGooN5OK
rbro7AskgCuokBqPIWomNZ2HJmxvi7IuAuAWz534IBjeuO+YdgTKp5gjcp++Pi/43fBgj3GnhCqG
UVi00koK3lN13E8rgIw3l8mrgGzVizc87PVr7jfWGqw71jK2nbjVVY3BxiNcMkFNbIHD5RX8mSY1
0W2JFcjM5MuQ6+jWrc1wignw10oPKrs1GaFola5OeP/ggFHR3jqqmS6fQ9oFS/6IQlbgTwXLjtYc
xhqAbwig3y6cVhfz0qIlvD3eK/vPHzfXWAQvi2QGpe3lbalV0dd1GskJKa7KACzL521a8r4Z4CrE
Mn1Od9qGVnD2FtduHKMnr+6Kzct3VFHPMTU+H50NrvWJqLN4gwPcz9y0oN9+PZwD6RTzU2vUTV3u
m8HX+jSc0MX4O6RoywnNv/1VNx0EGceyUCTKggG7LSW36c8xI1x5hyHjN34W6JKOmh1GE6bTpUP2
TrpxuUw91d6yJejMXg6Fi5fcAGvdaGGF9PrvdO69lT1BpxXnisNr7ddJWJCFUTfMIJlREQSjuc9H
exz23S3OXCRAOEDiOZmVREDz8Xrv/kyUZdUQV5R3DGyPWdtcskUJJkyF0gsH0gsFgL/+MkWQAGJt
3yumx/ePfyPlkXmE2YaWjwasGdr558HxDg2MPSR5wMWuPy1eAYKexcGJGPhLG3gEjdUu8/cA83jJ
d+EoFlRX4/J079iatSVtQdcSzjYlefcqoFQSKCHxi/i85gDJClLomHKyieScxx9C+DDQ4lO3r87T
vKx7LQtHyE0tRm8GzoiS6aUHXa4dxdlq5EjwkjH/Ja3eeLGUXg+xVt4FM4rNWau48NYoy8gGX5G9
wecdcz+CaY3u1k6Xq3Q6mbD81c+96M0BN/0mWoTBqGvog9rdVjD4YMh9ut9sbW+6pDySh1p0ifNv
iYODEkJ5BQkqHHgh5/htHrmEoepDmKgP/uDpe4njPPI/Fh0lON4DcN8dnG/UZiGlOSL1m1SC7RRL
fZt1bFnZFspXexvYVy42L/FWJWQT5KzU3uZnT5rbnArmrSTQ9vs6AtGNWHtrzzB/WBEg20jAwTNh
k9IzQf8X+HDqi/kIhBE7JZfq1ybPEGxOm8S3s6oR0tPiwbCji4+9nEJudYjfOxjQRQ7BSdByo0ew
CGTQMyr7JERCaxwzoz4H1VOcxmHB9CcjIyluhal26sPxMTqBmfZxc+ielf341o/iH/u0u7heMZE3
ybsDhqnwyoZimm+t1uatmMClOBVYrFUp70viCFajXb9Cv5inigtmfdekpoeb5n1p0DSlFj9l44nq
SNLTocugXJmkcCo2/A78GLGqa1utdsjHSpucbg6z9xaG5oXx1/IA+oQKUWPAEX/sWeomjjSy05kA
eJdPMyVfB2iYH+LX8E5mDWcC8mrpyWk4qcGXmT6RfiHB4WTC9F1R6Gtx0/DuOYDeK6L+NtSnM1/K
OP5rr82s2Z92F+zKrlRwNyobFr1WwdpRkytmkDx/ii4YYsJknuIm0VeP7smtzotJPBuQ0N1Knf1/
oT4l8kQB9W2U4yQ2k8xVXTX0cao5hCwTrCbIIJ3gDeOOY60jL2EbxJZdaaMSFTt4MXyHrlSujwD1
X5pdTIoud9mmIPmhwiTVhIQF6cjFdLPRfvEAAMaoNZ4MAzAFsRfxjsyGF5POhSWL/PgXpFnunSQq
ES3V6LjRW57PO0vXp/BW1o+4ml+BTl8CrIL2V5KXsLFjb6NVgf3AcMlt4p4ix2M4/VNjOxAF/GVW
w3/euVosOt5ZrooCGM1I9UX9cKFbaGgO19PeIXJeeD9CkKnlYg/Wvo+vwrS+wAPOeID9wrhMgQZ/
QGOQxIGK/Ecj2P2kdMVW9s7jKrVPqzGYqf4esW2iSX5ed887NlpMbAxnJ9vZ9Wage8xH4Gpgn7fI
e8ymWPjfgfb6zI4BQr/LnUG1NfLBXigRiIy2G12v684xN29pBHVGIx3xFGHGJ2/H8g+/I194akUm
Y/w4jdTlueD01gR+WfkNwSdfzCIvDmhZrBMedgOhjWcnfkUUjCau38Q59768CWkkaWllca9e7Ea6
z7u9FtjugDowrVfS9nFyVAIb0u3VoqjrVY3X1Rrc586whYUAFEFVn9/rBw5+wtmNKfFLMWM3jKRg
WtN5vUlRtcchpDcpUwLaDxZ+XJ6Pwe6k1GgV6Mlq51lIDnZBRqFhfjWD8glxNyHKMfxWgam4fOON
+OGHbgj9sxDdBXlJS7/1IKCrAGejSMKrnlDwevr++ezkLYW6+zEDNtJFsojPh9w7R8ZlpnmIx1s0
n+7OPxXvyISqcW2l6Eq+WcPt/DVyaCX0xMpQd5zEx+/VA0tMx+OyfAljOFUVQmKsakCRwtH6pFuN
kMJNUEQCeGbnbrRE/QVKZBXdTfdZi3SIZfHgxpGxH4telMGK/LB0ri21lLLVQfjmFvV8+87lS2m3
kEpQwWFroCDYJ4aSihzIXPtatPMbtwxrZkUUx7Cs6EPneeuUtO4UyPR0gJsX0tb/PDUAc+qPhZPN
AevuPyna+M4bD0peziULrnoatA8YCLHVQp4Y9Pmn/SY/Fmj7IGwG6JRIWjKPzG607DtSqKdIn1UR
dZW+I5hnsCqAjK7BsjcxTB2dmToPs/V7b1hGOVrS76+K6cYluv32XoOxTfbD9JNI2wmHUJQbL+TS
P8/t0mVigfUlR3fgElzgdwoyrPVbO1h09pvwlv7/+I5kYE6uItUWmrwgCc+guuRfofaKiwrQv4ca
PltrwO8v/ZGe1/2bHB4BO8jbDvEVL5WIJ2uLErFemnj1NwEK/K39lXGcVUKb0ELNirdVx6DV+bUR
nId5x7FWgL0Pl256urjqNXN5hPXQvVtFUv8WCKv9z7xdKzM/gEck/F5EhH2V8h07cY/dcCIASyc0
o0AuUrYXYzq5W8kRgHkxIBWvDg8uNcPa0S2zq5oPx1BaxSoN80dg/+qIrWldjRhyZ9YQ2d3si+ZS
PwCIbvK089Ft9Nb8iv8vEcbMc1rYxPddvXVItG1rUqtnVZ1gUzA14HzgqjNfZ70PMEjJ7no0RuRy
gcEuaMlwnbFJVSwjC2AOJG1AydIXlh4TmjeLePgkxL1w9OXCE5lkEuscb1Jd/pDRXukIIr4CJEdi
6FT+jI3H5uHV/G0/I3Z5hvk0Z55seq1K36M1aC8BwhQ+vjaI2xSLxMCgtolAdzLRhiYLFPQ1qdTh
SD3DIcLALvryhALUoqHfZdvciWkyI1B07KMNoFMRSVT/kDvk7XFmlOrTEQLD1T+Gv30qU/aiuOLN
l+qCBUSXkZ2mS0mSZTenDKkNx7PbydR/F/YVHAu9Jb6hY7fV0EZzSvcFAtjkdY5hJMj51v6Fajc8
L/xOFjwhUS4XZyLozW9XR1sUKA+pIPUrw0UM+QEHXparTKDbrIsHWGl0M893dC0yZzoqbWzfq/x6
MOIwU/ts9noO8NNhlSgfzVtBICWxTjQxeBytYNmJ7i21b+P92Xg6N5ByxWCYgCNzAESHk/pI4gQ0
/V/fuc7hsikLnc3Y8/dLvQZb5dQnFbGcZFjXq524c6r2XyQVpZvWUx0VI4uZeXefFKgMDx8HgMYR
VQbAnzugvka3DfYlzIvAn/QBhwp2FlGcTFYmKvWYjZtO4xd+1rLmy3VrTsGfu3jhvMw0eveqqvrq
dw+eXj3y3RAdhTso1AeHo7WI+4+T+MrHMcuw2j/PR1c54aLIPxCJIeBPqUdVZrVlqChhq3bANhMd
zahdBv5aP21zt+DU4xi0DQc7if449We05H2ZaBIK6IDOWYJKpkoyrkqhSXTHWnW6o2vm8jiu5/qc
NpmMWo1asl79+1xf0eltAR9IGArneAJ9jCA0pH6iUO27tIT4kD/bXqIKDn4RkO+hzdo4kaOsUkAn
+Gaul4vDtgfGpZFflego9b9Q99KjJ9DTgGL73jPtnXKvO+XI/T4YHaz8sRmnwO45YCMR9PxjrXJy
7EosXupt/dtp/ncDusgqGLp6RNhJxKZhTgt+MTZT/qccN4Ry9Q/S9l6G3fwdi5p1SuxsqFuUloK+
Zn6TzuKDfBhlBJJMbri2aCcpOCVInr8QTiEk8ORJ7Nq1luAa58ULm6jcOf/souyxFRT1H7St+7wm
ciT+OsgdG2oPdE5xfVvxstE/2nn8nWsKaHVcJfKXvhliGalz/dUBcVL9ZuG+t1+lizLSna/RBUNR
Uc4C8SUbQxwEJWo64PLydsDUIrYDP/3DNkseOx/l5K4Nbb+07S5m66g6r9k1Q4adMnz3mA6oTJkN
YdEnMI4gDQuAQ2T76lqZFTzImCPLRZFiRvOn91pNKaynC24NXgrJhQgy/+81vbc/Hinuy+mQe7ZH
aUKPlRKvhDfSiDNKLr3ZMjwROUH0uoIS6pNNId7hLcgyX+CEDr9hWNKkCzWlCV3W5y9M7Gaaw1up
VBecpsoKbHPmhahmn8u8js4P0Kmv4wYNxpC5hQ/CSOt7xo8ziWYW4fp7pXQ2AKGGj7HmA23+23Yt
PnzYzXEO9N5P5kIv408XOdeb6RuMObnBFMgPNR0TIzrpFDlqsUVebmW91+zjt5ZqK9wi0CbAu5yV
yXkOep6CJ6evxDETbO4o1it2AnAxVUPEIsiO6tDR89NaZB61bT+iPZmgLdZSiYcVLQQESVvSyvn7
v/IB4VikgNo8GrE68MRG1lm2WE2WfBP0/X6rg4NN3EvyOlGUa10ChJQPpbsCwuBxpOX2nL82sPv5
37obUmTJIDgg2ds5VMHH1Kdqv1s1mL19mcs6Zoejm54TExdV8jW6B8o1Q4zRKKkIuQlvkOTLmZD0
82AmasPx9v1Y9tznOwJGb8pXb96mojp3fCEzbu1GcenoaOhf9iUjuDxPfY1uAo2uhUjBn8KEVyvA
gzdSp5Nc2dCKcBYmLp7lYcpsTxZ6WmhI7Fe3bNMhnmXKGWX/CvSSvrH5czQwra3D35xrpw6HkfqU
eXlis7miPb6MSubbFOvT7k8m8pKN1ks2VlZX2VzE11kJ6ZEHVOve0iOEF0bjlLQwj/MTuaQqoc33
4nF4xsvPRv24inkol2+JLswapd18/3B7R4Q3GYv8R+Rj2CF+wYPw+Ur2S82JSpWu5bZK/7IHVKVm
mZISSPmSaCBVw9godYW2eDHozNihwY+Lpw3cYo/HFFnI9XcEvoIoetfWLb9D0yFMK0+GQp0Qnqmh
bGM4ku+2NZGx2iHaI759SVFHkv2m7H0STeS0Rg0fY1W7qw1aL37/y7bwpIirJuhAn7Cewu0ic6vY
8UZN5ukkTTUB8P9wH2UgzZX37Ku+vVA3nN1TDBgejdFy4FvufwkN3GWVnzTpyApYIi6BYLIciiXj
fMm7QdsTS0yZX5J1+hjN3QYUQBBtubYfYmnStlS6FZePD/2tM2p8XulnboNxnDDF7uSQhVhIdUKj
1iulYmzbvCjbhufrqKGuslT3eU03pOL9WVjU9uLjxeV++IHxQ2lwV+zdmccx7fZGLShHDkmiUV68
5tOrlUs0hsDKQMZbPqAuVzgpAeaKB8Qdj5bdausKvHUzDt2JUHw9oVoO6WicXBLgbwL5a8AiGDHw
Fnqfmgt5mYHVQSb7gzlrXLNj1jPpJQKCvt9zxA+lNWIjiCDVrS62Srd4/1g24BlqgQyDDPIcK7yo
qk+ocspqYZXNXl4yWCEeHfyMGNmOHn+ki0IKyRFWFZzMeIUSdw15A2Ckv21oa7uhP863g75pE7rK
mY1fwtAQGxdhTolDYxnL786usdnxkqSjCIwGcxmI1j7bfVCRvsFyyc/zHFv0bQyb/xarHMata63x
ZiO5rFWAU8E72uUFy088FyHE5yfBD8jOi5mu4+sjgJBzdVu2InIGH24dU/02QdlvBXWQSYLRN1RC
ovsO9kyjH/nzkLAp/uHlt2x54izUqUrTD+afqZHSHwYrCdYp9Kh513jKg5ZQopGv2hGheYzzSK1G
5XupXwe7yENMzSOf/rmHaEtfl0h7GjMq1V9skBS2ahX5XHTBvyR6pDTxgi99vz469tHilORTFj1h
nDhYhKY/PX+Q2uSZWRCx2ShdVdMRYIfERE3DK/OGoX4NRcgbGaiDuRu+NJAyGJ66vAmQQVqRNsTM
zN56kcO550o8BPo3T3l++Q5DS7du9vsTX/0SaEJ7sICpAoRpmoFP4JapG2tH7s2jrOg7SYSDXKOm
/AwQnFDY2Nk51Yeh3/OK2EM0IHPaomWv5hkpPliZMJZBN4irCkxCmEFmWOAebabORv1rgazOgYi2
D+9ZX9V0sQp9QHefhHH7Q/Crt27szWZe8KS4b7RT+RhdUOVu5DhFk+jR7p2opVCELfnNZ0e6YOAm
R51imNZNYi3UiZYPr7emRioAG6ODr8eX+BPTG5D39J4KtHzAA1YaNi5ZWrJ4n49+ug+lUJs2w57X
C2HcvFMbN3SThqeuGra9dVWtn7/doFUOmRBRnIFkvs/hyxMaFC5C3bTBn9TDNvbt+6amAToLhsPF
S1jYfY2XOqUtWH/682H8iO4LpOq1Zw6vjJpioZEXPt3MwCS2IqDa3yQqrGMztSbIeUgBCnxL0ttn
JeUULu8sgP9sesTJ5pyr0Bp+CPN9XD2KD88hup60sf9PQyCK7TlCIqZg7W2S0PrtVR6dMv4OADDH
/8KOWdEBBtbQzCRHwYHdjdfYJ6it6MdjOP0X0xj54I0uZJ6yeEvXS3g04f7zcpWobKxOFqKBvL8f
WxzGZe+GyuDeZNE5El6lF+mGzivMcm0tDxw0NU9ERfyd1z4dtmtLU4fr2dvfe27sEPY7VU9QYgkP
4P4iIY/UJFuR4Y60oVo2t/9mHZkU24LvqbIUkhGK3rGh1LJIkLb3mPFX560In0l+gFlYpmV0/F9k
UxLarUvFsMj39hHaWcojagwwhE/mktrFLWyw9ZgZhu2ESclI04xYoqPbqaceU4tY7hKvnXLa+KWG
uEBdDWDxX3aVhoARswGqJCj/FRdY5wzhs9JpLXdGygrawySNKBYxBcXmHVzntKUp+UVrX2Z5omrz
l5rdWCShcWx39CY2KGb356wxkcyngVAglwHABrw5z5q1Ci+TBAcRQK4hptnGu0am5IOrl9NkhRNw
zMZ3WnnccaKnw7Jlhyb4zR+l52CkT7NvgjUSnK0yt16ObQxYPaCX8F/uU5JwhhkGWF/PiLL2QS/c
VxPKXxy2f8Qh/9cLeCYwDMrwwaiYkYa+/giv4mLz2nSCxSCydaVAQbAcWOMC+KNSPg2R3y8l+AmC
YG+XkgHrBC7t98OiNNaR9rJtSdSikQKSDdsLcmW/1P8FGpiw5IrOJZ2f1SGZoMiAkb+6u0DcnvKM
LexGiRV4D8MlcSiJ6sy+XRhMKR/u1rpgAXtCYNsX6dYbC5l7JsUiwC2LmHD8NBAeXqEVwI8JRWXe
vr9s9H1H0UTeBZuH/CB8nf1H1uZQR5CJuwu5V0rQxRRpxDMs2CT8EKBysLw7l5y5CQqrUOwQZ0uR
BiprrPUycmhjzNkh+WDNTxZwFtvoaW9UbEOJSmDSwBgwqURY1pfcEhPNSoFk1PIwT1CjfZZL6yd7
oulGVSIxCsOdp2TP94x9rO7tUJIP1earWo9zHoJDEt8hYP1Cn9MZXXtW6E6NVasj08op6ZfPiW9e
m6+S/YTlFq8DzUmpQvShlI70DcjPYGCpPHaBlQbJw0RWqYF7fEsLxRIw2azgAxMUXFqTJchF0R5g
5uXy0EIcDkJfsHsE1WUFX+JoCXHMaaKkReVFxJlb54N2I/vNGnr/qH88ya6gvjE/imhBMvVSe4XB
XaKNstvQN1B51AOHXD6B03j7UU/uX1+M/MgItmddYUGfaBZ9mG6xXOjv2f95zPqsYboTsGz9fzv1
MgRlPNqHeFf9nJzjD7XAD8DRalPfYVxt9zJ4KwJhE05scARUEfAs/yMM3jOauEXMrJ9fXOEyukP2
tCNMM5r9HUjiIhquBQR0Bk6AzfFT/1uyw77iYlYY6rhbmjCKXqWagPtYb1er5VthFw+eRGJSidSQ
01XMWqK4ug2dhZ+YYsR8DFxnBgUvcVBnO1I6xVdDh1GU+CRR/HEKVcbnTmbZdRa/XP7jC8fFSk93
rHhP41YIHfZqVxrSQdQlMnd3XzG/nfMJ77xWla68uLqszQh6t8flb9R0F73UzDg2iUBX07JDL89A
R20ElMBnbDLmBf0hriytnS/M/Q9mCEMNVF+u/scC1tP74VkH5Ixwm3zstCeRJ0IS0ruJz4yltRl5
mxYHBQR5IvtsWB91NVct21NQEb+3hF6OQ1TXU9wJYRZmFPiEAwfocKkjZOtjMKbOv3dKc8NUJA2m
EWZjSfwLR1OBsoehHAoGdUdgoeRpWqnerb8LL+p4ZjwgGaGw0IlUmUS8lo66+oMPb6AZSBZy80cf
JSXjsNV7OAiaOBkssPLmVN3SCR8j2siUg10uWXjREqTFW9FryDpwcbXiNmYPiFgPILpl6czSWEce
lKUOUqi4wqJzZkCiLBdg1Mq14unflZm+mcoMXscHKnEUvdHHEmr3L4uOaECm9EN4GPNcHCRFQKkS
HWLnj2enqLAp8r7fbhyRwRGuSx8E9aOumYafcOW+R8kiYc4kdmsRgPEMEP4fhESAqMJPdzQ0NWDI
bY1BnpbL0rTa3aXDSqKvAOCviteFaCO6nI2dhkidy7Ntr9A0sNiljcjaJZNU60gFoafhHd14HY+f
cT7SQ1JT/wbBCTp9Ady/9/pBbAbngbpJBO32fXw4H3tVl2xrjC1HHM80p6f+WXyV+1aYFc51UXjU
FMjW86ipibqJBjEsB+rFiEPtEEh55TSY+d2fdsIj5cWcB0VYipjwRNcZu2VO+VZkO1dVWE1skKoI
qj0D/iF67wpIDfqMYcfmfzfDdKsszGhFtyV5hDjdRy/+4Wm/bSzp4frCy6ipm00vRt7EC89HRwF3
zCiqsWL/1dJ2nXLRszfSDYZellhRfVr7soIWcMBhOWKL/A0QkV0AvJdjiH0qr9FEnP9fztppyHRq
0f+4AmlxooZWmkOLwSJF2ge7SaXRe61JqJOqllmNpbmylP7pz0O5o6eYE5HzzMnWPWCOGD3OgbeX
v9cEkE4oNhmvZKNK1XylCdyQPzue6qRHWz2csS7BY+vSB5GtnpY3hon5CvlK04SH09TmpDyyifcN
Zis/mNg4dpjD9+12zh+z6M8TuhpOrUWDcp3EX9gUFlfRVTS4/1a3iBq5D3SXJ3je91ISPcDXkScd
/3WIwhWL1I2oeARWIA3lJ1wAavS76uGEAWoU6but/UdTLHx4V3XVRI3C0Z8XzilJDaWPeWGzt4tI
Lzj9cLBC1amMyB9Rhj8LanaR+Ql1yF49XvxBkZfIGUZVd1yMZXFMu71zyPuSAIZLqyfmQxwVQrZA
3WgkDpCjnYa0TOdjL/FMSbTlTQkBJxGPUxWTuXQxXyuk+dfRWZzCj0tgP2Wqp9ZRpuUo2WgBdIEw
aZhRECuvUVi7pzrVJxy/hoj/z34KSy74cIsS+pMyKjZAjiB7sSv2yEAaWI1DlNlv64load45WG6a
TfpQwgkdTKkj0y7HZfIWHioOsJIzSS5h5ki/HUoJ5xUw+CDx/+I5ZC45j7vugKzm2uqo5lRNHgnR
kvYg8qOnpdJ2/n0oTRTBTTT3zkNGsZlbvo7/1K/UAyorDXdi0gnlID/PbtwDtN29IUXP2BEQy+C6
0rnjXCrjbqVpymtkZCRlV6YH067rDaqmo/PKjGnDFeZTGN7bHr6eHcSyfF4BiFoaPJo0hELCoWBU
m8yhWaJ0sbqcXnKK/f1m6Qdlk7n/E0DHlPJ3CDYGZH7pUB30z5KjsLw32MJHuZivq6BP/vbQAg0M
XkpBkhNXEVnWGQ1hU5/IGNrulmCYhx9hEBOOMzWeWj62yaXJikJscdlxWAr9HifncEH4zD2SQWEI
knJzgcAdbhD3fx8YgF89sw9KJ+X4g7Ba2yxv4/uB4H4W+xesFrk4s18pXExFz2mUvvCNu9htZ5mm
hxJv5AzuWnz0D6q6mLomnf5eiFUE25ocnx9pIJBrKi7AEw/r0uLKOxMfwl3rKk02Z4tk8rcVE4Sn
hmkOI69btj5RB61o3lf8zW8zKAQKBhDFIPtk/tivFZeRUzTrmEZ5DuHc1AwVl8jWTcAq9iD7QN+g
3KDXK8WNqteB+4UNQmCFneGUjK5S6EBV7Mp9K5EsIDa0EX1bb0hGJp5wBwb+xcWx513oz4dLtiR1
OsvxaepAws8tuQxUNPnxOI/zwv0Q4q19dvBY/s8C3dKY2xrhlO7QWQajWMRuq0JdrQgAezavgbvJ
YIdAXPgtu05zQXuNrI21RcINv7iA+W8fCXSmBHX1AjFmzuQ2p3Z+fHZ4PrA4uBSh4lpKwsJkBJR9
SUe5UXup5Sg8F3r8hYyaWRoglOC66dSrEbMGyqE49IRScOYpZi8nedn9ep5FglX62l0qFMH/H09H
To3VCIvRn6zy6bCuifopBwa/iPsQj1RGvfe+qik2J1H8mCycscaNJt8Dsf9U0vHfmtyJsU6v6yxv
7924NGNXynem2KFZN/pda79xgvCixH3qLoR21/diLUZrWChqCNKYot6ANtmny7NIi3ucRUJHNkkW
bAmNFyp0f+DnMv/nz5eVUT0n4XUwIkOL5dvw+mN56pcL2L1XVPCPAQhr/ztlEAJtSn5I+y4oSHC2
0WAAE8dV7u+1Jh4Ohw4LyB0A6zcvtpdCo+l+/BlZ2Xi90muh7PzlhsQL3DQI15T1DOQQdty8Jz1a
OLf39JCkFm3wjuJHE3kT1sqU4dtWFmBe96TrPr4RY2fybiRgXcWWf7maZyS0KsWU5nnXXVWq+OoD
BJXuiFuE3Z0jLUOpEi9fWcPdRKbMLamPUmoQ+U4w/rZXvi/9mSaifW0O2IIXc0fYm25h58dE2EyD
pJTtqrJtCOXQUNFNtOZ/iLHW93nGU1N5jlzt2cttiZ8vlNlhgup10oTC//CaVOKRYDY9Vapw1G9m
sN/g1DaWVBoDbFFfaNRLGLDKggtKIaLKdGcfzFzPSGpQmpgo3ZIusmMXQUHhFWl7A7F1vDqM0qDg
F60cPZ8Ij5S62B6+a338XlRLcfPWCjLCRd+Rt9H07ekOkXCksb2If4L9eJkNx2kTOYUi6r4/WTyE
qxZZb/v8RGrtF5V9pHpeLs0J9Gu2JtB46iETuxii//Ztf97kx3Suk3v+IeYp23rFfZg1sieEKQ13
erX2Me07MsqIaiKojH+VhJ+gUa3C8ieOxhe8qgoSuFQx3qsULn8xx5FEVnem49lRhGd/yBU7aYRS
vDC0fHEpXbaxle6ml5JPJs532Gv4X9mHCTenCvMQpRI2zd7vQxIHmrD9huiz3yyAwxVArH5d/v2d
JXg3IOruflgSclkoTnkdy1YBEoBpy+Er53erGX8PwpsKRdRDh8SAIS5u1pFtmEcTj3N32NiIOEi0
qGVaZX0rkv6YuPwejT4FzECs+XSYWVFCIocbm1pu+8YAQ8rl7rZVfSFX0mpRUTIyehkvlkj3KzGA
wfXA54K3wurACAVjnIni1srsbTtPaL473zjGoToNHQK7eZvE5Oe/pxATybMZ0IYjRZdLwX++mSlV
VUtAc+gwBUShUEzEsv0MTfshHhcPPnlRDg6gN42/1QIqdDWWKYSRh0NUTytdkxToo0ZCzV9WjsfR
CPcmI+BIqkaNLZu/FQSWD3D29ol5abaeGC39nuW0sYAbC24284Bg7i+SN+gIhDyWV3tT6tfGxHDF
v/yvlMF/UIf4Qtg1EmTQbH0E41ikBjm+0gfqBCmY++jDcXSnTOXxuzxMOF18rHtCnQ367I3ghmTB
ryN8uvjseKCwIFsiwksNOPLqiWkMHU50tBm3u7M8T8j255tiTmfIDoIXOg+/vYVG8rJwm1twJZaj
npD7L/lGf4oFxPFf2Ifn/Md2hLw1KbLWr7r81ZGC2g9p6Pr++tBnwcnY3Lq1hmMdORCUjCyeFo61
I++WmV7AhSgUnexm/z8db2453B56wbrcQcl0l7GXDKZpF/eRVi/6gbnhQn5sT8s0v1Pd0QhY5c6p
D+sc032POdSArFuIHxzLAtVgC7VBe83fFAIol0qObhJbxtGJzb6GZbsv68xOHRCDGffaZFW4ufz7
axq2UtGmY08p2Zpjs3UBR4zAKX2dV4Dg4Xm2023wTq6AtKSJ05JjxWg8oxKLGVQBtz4sPZQXquFQ
vOBuVV3q6S8H+5myWj7lZW8KysDmOOMippOJkT6KiUMSpM1tENi9opxtA68UvMKfBo2h3fxqG6Ac
nAcDdYeWXEsAC8IVMcJkIRTs/eeGML1VOwjniwkaEp6AZxv3THia71sxE/Cyr5AG6xTKUGaQgAex
vJejrZsc1wRpgg9SUa9gY1Nz3oDK9sI0QP8avjcdjSA/9/8Zh/xcjw/zLZVVE3/H5TFMW/oDAK7c
Fedgv1Ni41Ndz16OYeYMIn4jrToWvYzNs8VprY3rDmAcMqQ9U/dlk5G3fkPoywk9Rtp/QdSf6Z2W
lXm6fFcPK8/bk4Xg8VWyjNBj9K3GtKPommCz9o8nZ8mvXTlDqigsWGVlRDEY/Sg7BKXrEI4Md2QM
WyF2e6QmYj/Bq0E2nVVl/+i5Ar9Tm53jWPgpVLRXOTWbJ9gncs5rjmCViRx1YDO6SP0hta6yKd1Q
TOTigaN1vDgLBMlJmyezGVUSSkYsd2r7/wasFG0X9ZN2cy9ZiDQv2IoGCjh8MVB/S+q3qgJj/H03
i4y+FNIBcE7oqkMjzYWlZdvoWXb/CwFDpCz+8vWAT/hEKjJJsCPwzqREW7TMHRTtLMeM5et+xNwK
fVvkjD2g5c3HOr32j9m1s1B4PwH53fJtqAX1RGN1ZcnY90OtxJ5nAUjmCsNSqljJchqCYJD9CvHg
ogEJ0xz7SsEvHbEQfePTF+aO8i/h9A7YMJSZ8Nz2zDqSaBdw45IL25UzLPXMRClEYTWnzTuC/b37
3Mu6mGC0fCaXTFE07KYD+7Qu5bn2LhgsaxNT+lRyVr0k83gZSV/fOJdVLOvjgoTfCfkWwxn008nE
4TjFoqXQeLFdkVOJZj9hLlIM4ssuH/fX3L4kdh1DV2BjDa6gSiQWlOI7V7k1fvrUNMCIV8CRQMPi
hDNbF98+n+kXKC+lyuv1nmCTuZz6h5NQ1FUNkjRjUEmlqeG8g9XmVJtJWiCBuquzjo/PpQUWb+v+
cIn1twYAsD2mm7aoqu9ZO1S3kH6sjrzu+OXC/zM6msYeIpRfJNuzUo1ccrae8UpPUt/0aa2WkyuI
UMnnMCa0nIMnF8nvKFFWKG1QjXpNZdbS20UkU6Jog9m1a0+h+f8kV/1MYASNuhnWc+3AqnJRl0L8
1HhUufgcgE07IIaH52r/r0CkRas6LheUlSeAd0/c8iQXPbIUSnPJTZJn7GqMrR+MffnKwT2TjnjW
vxV+kkZZIRZgcmb0vybxQlJtOtfrg4HQQ7tak9+2cnTQymhuJkxn/KsubUdOx13BE9WcyLpNg3aG
TOAxPuBp96AdQmwtXWzkuCqmv6qTTu44981RiO1pPK4ELJw/tCUBpYFuQImt7R2Hc2j8whlBx4gu
2gZsUt8sOSd0rLTI2jr3APRh63/BsUoZj9KhqC9wGZ6nKYjMSNbQJ6hXxvnDMk4+RAeg8CZuXhEh
ducNjKYo3Z11+y0UxkZdFpwi3n96WvlzKGwBth8+79NwvcU41Mi29oZb4E3v9yMISsn75gml0VjI
yTcPHpsGn1KMnnr2VpXudmfMKGbHnt8LgkDJ9T4n5znBo6pwbLPDgrHv29msfmdrMF+8l8LGQPD0
wJks2m8ppUjSlhPUsEkbEwon5/gf8+CQ13h3jiZTCt4qNBRQ67muoU+QhUCbCns07rygYZMPW8jE
4aCYEQ9X07NHo6iK7/QlSX8T1WXbzvHBWqvlP99GH69gNSquJC8OzNN48rhhJznVjDRkwHPlLuxk
OBZ6mWEzZdh+CG4J4WGXyazveAzFhpmISxeqPewP9Rp1thWPgYuBFCYGQ5kgCebAj5h9mgv02cvC
GT3U+kjVd7Np8LLB9oLRZBxqcYNOjQNXelhE1Vznh0bFHuJgJ2QOGoehphMaKoMoLDj1MJJNtTlh
VDF28+5T2brl4sog02tDmjb3n9xZciDRvMgwOekhfLBMUVHl73YiEKkWovo1Us3YY+WkWBvjFwTI
IG5XCR89DKqjpnJxvZOVSuq6WDnS/CFRGIBAn+FJe7wyfzxApz1O6qFpcSI8X2udftH9DnjaV3ch
pVIRJEjhVBr7mwyqCqabPAWA+eimCIEysEBJkrTCbsJ6uYgNoPWZGVQHX46YtGRSd3VzzBOPisBV
i00DP+btFebkgDluz9446tCNy73yOhD21wgvAiDK5DZJN5ZpIsKSFgD2AzMGzCuhiHsebUHK+eBA
hF9bPSz/FQTL2Gg96APeZkTAj3cKpdJ3Y6vcYKmNyWGwVApB+QTkxjlQTWHiStL62jLMjPSPi/Rf
olc+5wWaqOKol30MhRR30wRQYyqDva8KWeDPrH/5QJDlpUxzkzt1MBLEcvqlTBnySs21k2SilB9u
2AVa0qG5NMlICnjx6MLkfQZKKP9epNabTdhUG7HHIj2/3LslWyAAHLTAUjmCRqTs9KkbB0ksdPyF
twPDFJ68ATjvJKisHNX0LO5sUWhW5Q/vlqTVmaQPnkoJsLBBVnmd0OCXlYf4Rj+zDWlhvMmP9bta
6boHLtM4vI8MUqmMcYBKqLRKlIbdVgbdjUOjsLIvt4vM9zG/FXx5gyXXfhvB/XPN2TgK/0HVo3W4
jJ4Ysd92T01Gp3BGWErgFzUGQ+HznSjgGm94BV1xTR1InzxHQ2l8qJ6C9ZxM0P9355zt4xQrfK7V
04aTFq83ukCmDUh1TZK69YWjnK7DdWfv7FVX8K4U2SR8NQxn6jgQDvriyjCEakNxijvHP60pOJn1
FsWvPItKBxiuciiMN2KKr5yJdovEVToIoqPCLm5+Koky+JD6ONE+3If+UTioWz0PjQ8IpWS6tNoR
V7AOMwY8XEPGGliM3epAax6cIBIbdmwCuugfehOHZ6eo6PGrkQm4y/HJS7mXSFGDVtNuQv4TidVF
l9gNY7rhm3pvn+BX/URVXltA4MdHw3U5swfxUkpl1uanRqa4V2jVjGhnbMgtdw9eI92KUPyuO2Zf
q9BKT7h3n27yiTOzrr868BUdi1LarpoBx45zXhUkV1CraNTxqM3TQYiol9LYXQOGka5b6UbbFLoW
Il2YoyGYtOAHVtOhnOaPpgRsqAzkVMy8/r/Bvu5BindYEb8exKXQU4FLmqLIDo0vgAjmwIzZtR4h
TTxAI6YrCWadgXA70XRpIKJhAxU0Fdx8sBt9tWTWMwcLBlkGQgr2rHwE+qPTQo2zHURFYGsA1zZZ
3aDt9roLBctgK/DTzBGpH05e8uXu/x6ioIKL8Ek3G1R+QTyMx4K7Iz3jSMJmLCr13GVMoBQvwvq2
vbV+HP+Jn0Dxye6vx3JvgmhnDnSnwrjZE9M2ysAGrC6dC3j5dg0+KRLTtIkkSnGqkpwG7X4VvNsZ
kNXiXzfQ7F5Tle2hG/v2/Sr5fgam2rqQUYF03FP5TDsLkcYpiEcnki/wyaIc3aX3QpNtUG1Ja/3u
mNL68UMILXqse6w6/BEFS3UWWXOyvHvjN4wMX1Zi53uDHVXWPHDK2CAy1H3deqNWO1QOngjMz763
sFENnygzFVOrAezTd16rudH2hQu+w1ISpfzIDHWmn35Gabatjf2CsxFCz/pYzPZwFpHeESm1Neu4
06jNJ5vahlPJge1dk9IPqTlYgu3XrCzxbhY25Q2B0supf31b9LhnbQmrF3Ryv/qW0K3IbDUXclvr
RIQNAdeZsvhHgeTTquVuGZ0lLTNO3dfz4V/b/v6iD6Wi6R8e+UzcZtU8bduyHpRZQ1htYeD6iKBA
4b965eVNoRBmU1aMlaIHf8eMOTvgtyWfrg+0ryqojmnPdGgr6xM/1av49H9P/QStS/8BQYKRSe3Q
6RB+M8XAHE1xkS95Y8/XHjv7hzJzMYnOCIgW0DJybTosq4VXeQ6WicgqIw2gEG4YT3X+Yk3dibDk
COfwL/4axq6vGQwJn2Bik245U6LGcf4URndCPg5t/sFurfAYiyDJLtKZwe+7nh08HNZOScqbuqE1
cpxM2+qFhJ+d0/c5pjliudL2hToSzJmm4uWJ0trdky9AOWKmiD4zjm7IBbCVyXfYPCDeVMh6AyqS
J/CB8lOXIpThmT5cbn6UEZRbGbtmrQq5FH9H/QDxB6E6/mcTPoLuQPbdqHwYR49qwa1+x1H9UZgM
/sGlnYjQr0VFfUbgtIU3cJ+etpHIChmyiOVOWQdX2Gq41yfV+IIEIzE22bV/3osCK0a+OimcaqZi
wILpuV2e0A6BlYqf/Fsr/t7IpoYcBMpQV3lxxy+Rsse9sQ49RqIqG0eGZMuZyOYuVIGk0HFyBxs7
manvTlP4yj5yauhCWwga88g8jY5Su0cn+Wqdmpeli3sLGdrgaJAdclKXbvXNK4Xn8uP2UYj382Y4
Vv/g7C+y85KCZ3gALVZ+gMIGIPkLTUdFp/yNJtOn89dfl8KmrnL4rppcbke9si2EfZksKez5FWTC
Kg5TdZvPBnUwiN2WnDgJoGn4MKLYnKsihs2fVqy/IR9nkHe5uJW0qSoSj9wf9o4ysImvaGtWckQh
my2uW43Kt1cjDBhyzZPA+pzovkc2STWeNSeI1USG0UKoQWOJBv1I1kom0EjDISZaDKgOz87JGyst
UMlGmd9Lx2vPALsDAu14XJPl8rAsoRqxzN5TyEXCjrL7+hCiPMmmpEirmmI3mt2viSsp3pMKmTKm
gfO91+ZlJht9ApsWAZz/syVxkDV38FUuPTKEnGIHcoOfFIyGFAV2sKbSWTpD0SaYpg2EfdbrYb2A
XLhW+2yU1y9YFhz+EAs5SxaM3Y4qlMzZHVGusNwfRZSqf97lBx8x7K7Pu9eMmJUnVSurHbsEUrj7
2VyK+xiAUqIpDCL4RsupDQ1hw5MDVCHjTukj+p2wutzL1lnGkoC5WZW7bi2rP9Iy1UUCtPXiV3Xn
fHeJjwcNvnQ0gtkP7bMjHJXrMoPl1n/1/RGGO8OwjHbdFl7aN3a2t1bnIPeg7jF2cc+sex1MqFs6
8gEXDeoprBlrIUpjGUiQO5HNVNEcPpGToaWfM5t9lXLng+3Mq3ViAmwm+Hsc9A/nLVRfwMfnM9xa
zPluWA93JrVqt7g4uDDe8T5ZMA/2ZwQ93iHwZdLdLO7u9s8KGQvReazht8g4qpzBqr0bKNgFcxVH
g8t2tD/87hMZK6KCSGAeoNJ15FpsaJZ4K4aPhRkZ0lhBaE0jlaDaH3vyqfCurvP8YuMMRzCUC+P/
+ahG3bG3OqcEg0wnD1pq+nU8slVyzds6Nhgym/Z+gW4SlbwaYjODm3PFYEvn+MTR9wsZMrmK1Xdd
v+3LRKdJyxyx6N56Iqm2gdJRPXqD3GZ6IeF1FT/IIE6CKN02YD19Fhk0SkAVsXEFp520XYRcKEbF
6aT0q13BEYk+359HeBFm+Vmt384f3SlJ0f4aQNvLNorBuzIgdUjwV3cuKqQzGHw4Sikix6ff/0Gq
wHjqsrIK7kR9b7Ab7ndbb1GV6JXtQqAq6NKy0S267oEtYglX5O8oMkWhp7q/6Lj9JSChjc5g2H4P
KNeqj/6HaqpgKJpvgUH5PMq2CLYsMes4v1n+I0guBl92j2YnWODIPLjrsK4t40GDWfmYnqXag5ox
OZxPkvwZnC7jEACDpBDzvSbUXJjc1yfgnHIS1bjRvcsCf2seFmnLq1FXLJjladlPLZciJULq+T3Y
hsHhHVsVU1IZbPAkD7DZY956Q9WRAp6a++ShTWIThwOzWYtclS4P5uBBIrqWRQsBggAWI1lSVF/7
dLtPIXr6j7v+aKx5pSvFgsvq8+lA4EMPFDQ1RVMYcGYxDgoOPmPCN6sP0o8WwhKGgs9ab8kT0plg
GhKzlUGzRvtCbhyYX+lM/vANNuGSJMm5DxS5JfZLBPFNoBBkxb7zZp2LwS8C8awBwA6M6LpurmsW
mE14fVBPlOoOZ3MucA5mgLOAHY/pPwzO2IkcpLu1RKs5ceLTe5tRGwPoLrg6i6WJPNSxHKFsF//9
YG9cc+6RgSpyCcniAmRRdnGQbtf8mBD8/3wDxHtB/Df2MgrG/zETvaCQ8kU1cfbKXeEJ0na5Zyuy
fIAdaGom33aQVFu2DPB0Tp171QKqi9+TknzvroCpCoLtuvd1qZWUsfKlIwy6WShxPajgtdivu2me
spy9eeWVj33r4p5Mn06xzx5/u+FmRIB2bx85ONl+cF22bi8Jdrm3pBM4vGZIgNaMDDehYQl98SR/
+txETd7HDuPwouGgyC91rQBc328IThTBUYtN0i2Z8M6n7N2CMXBKYGoafQ/q3Fch1HllEy1iT8AC
a2b4WzS3kUEnXlw+FZNRqNkJD68/h8/Tc1BCxnidpvqYmFsZ2uUG6bntXEPoBhwMY0uF1A6lB69d
mZOOfrjYoG37Y+PscF+WBBuM/avBC14dU/NatQXHXfoxdV24MGV1Bfha0NYg4BbRQukkD3pwTTAH
Du5nDG1No7uKED2QRmRZUP5ddtjB27v9OW2J00iZZhBxVsvUf/L7xLnPF5lAHQokFpcNAllObouJ
XU844rAWLsS5QdRdkmf4Z55zYqCgA/lg/HUaTztTnLRmQhWmj+g9rk9+xw+XRr0QBZPkUp5TF4BJ
URsL8n2TywpbETB121Frh2Pk3iRAMLAdl+m+5BRXtw4EGmUDRqspNW45/yfHLEJ++YSe67WXuPai
/q2Nu0bVidiH/N/NgvCMRoSwVIdCFI1QL+WSSEOhowqLNXY+kWkzrUGXLAgeoAHrIxvUzjU7fwMD
ZM6IWqdDsVmJf3XN6nND7edvemG6NnSLeJLPu5t3t6NnQREqZK5L5cuX+13s3KZysQSmAJ2/lzyd
LWl/ynD9l9pM52u6XD276tvHybNc4wAv9eoc2FWE+mLHxYKPXy7d8uzumB5w0nCWrn0kP4iLUDDl
mPinopC9ElH7z89UB8QUAhXZOGZ63TKH3UwnsXnaorKx/Ik/Ako7QqodQWq+179GFZNOvYRtbtBs
lsPbistgvIMdC2KqpNSkU0Qgb5YCgfNMkeIrgSheaGu8pvray9CRRPteVCVPR8GtoeDOADWZrtle
G2ZJ4RCVcNHluDKCcpXdJ+wldKF76lbovwIY7n0outst8qXQDodnlgG5a6CG3EdoJaN0slppRwQ6
1McI4pHIL0neyyte1dB9b6eHhGiOlDzFc1aMK7LxKEtPPHlNSWmA/kbChY0oN9oqvw0sLVbyQTTK
EJDdJ42czndiEPCSlNSIEqAG+saX9jAgzJWPSm46SWLxFkVgcg2r22FfEnhSFc7TmEXCoThilwj7
rMn7cSyPZcOBsesNB+pRpxiMDnKOoovXyfKRN+rs/CvXhYaSRWDD5a3Y2dv5tT778FH8W9Ol+6Xp
nyM3GxQDp/5h3JNBnOXhQZgPFEt/tTAy24KtYtfe0qYJMRkVK59WXf7w6VFdiYtcUOuvjukLGCw/
rG1YujXiKgtlUewLf/LbV0VIILVGjeenRmyPti92VZF5Oz8NO+5UhdYja9Kfap2m745pTBpqjCJI
L4IcJ729qbPeTOlAUhAw+w/CTh5qihaHxgmmub764xV9GUZndjNl12AjHACmo4A0YbknA6pUQTyX
xIIh7Y0lkTJ4gYdInkheKjmOVq2nmNZRAObJjX2bf2hwaxRnCqsRMvGdFCpZTFQPIp4mje4o0/5p
qvFNMvwF1iLTUmeim5x833wU894VK662MJFybyOdX7eI90kA0oZj9O8v945mgaHmAG+Zom2inLSR
5fL4CH/GdkcTd19IDdoXXBjApqOyDBCMjevcx+3ZiwcKRWgzhCu/higO5/ufQRZ3goOKvbXPY+zZ
oVKujQp3Oxvv9MMnqb0Qx6ybvmMcOt7DunbXE8AM9XBpYGkZ2rrLwgDvbjlsebyhvC4saeB2RFne
iYJEmzKiJprgHBYf+DHGA+nZm+57oRw+ZHRsAWWJWKfn4P7K2v2yslGs63TrvLIkCl17aoQvhv/L
gzb13ggopxp4mZ8eVGi3jK1PgmrSFctc6uuwj2KQAqugvcI7LX+g4NQcXjOVhyRcudeizhpJer9C
RdcP0ZIFNgWSXY4f9NadtqwJ3/T7n8a+V2gOq/gTzG0FSgLCRPpgNSewhY0mr7xv+LZtek/ofEEm
CXVd2lMrTo1rF0qnaKJJLAxUX85Hy1x93f/XEmeYjSP/XPxmG0cEibrz+PT+tjV/cBimtaO6E/JX
Mki5toeFUh6OBb79sqTh33ZQ2pBHguCDAqmmzLROaVFvjaNVA3oMCfnxXsOachaMfZCfBa54roQE
TO73iubNsnoicoR1MjgVtCItv/y575wrlRrZTDcCqQBdgzxWOpvutFe2fcqqUOKu35IzxmC5xKxz
q73VEI/m0CLRGFjCOnORmcnL/x7JyRJbmMpRUV+YeImc/G8mpVnBjPfTrJQj9k58DXl/eg5tJBhS
yOUFMZKZ0FnW5PqFOnRdRExQH1UezFnh3SXUZIbYKaHoDFyOjkxL5gYpiRqM1mAUo9fz3M45fbDX
PbAwi7dKCwu5ewQRYvvci2yHMyWK0m7uMqSLkFRBAr4fSp4M2fj8qSUujzAtElZY9q+Zoos2RT41
JuR1s/S0UeD8e/Yw/VfpH5N9c5OTBcMD3JTb589kTY/X7EuxSzeKXliLFlFoydGUz7nAMN1b5v+k
cNOUqEYsRcg3BVZlukmoKSge8I+tKvhNv3sYj+5hXJhErmUt3CSfog0E350h8EkRcWtICNh/9NlS
QfuufgVIbf6MI53+l8EQ4JHB7K04rKdUjPBqEcsUupeHvVCx6TxPXknXnt8UQFCARXaIilMF5e+5
cvIfXdZgCWoWuKCKn6ZSdZPXbAxyT09Z/j5kRIABl011nxF14uV4zt9M4UbDl1metmk75re5udno
iCVOydxRmoCmQrnyR915RC3rfYAs0g5mT/iZ25kD0JVGV83qAEVmCSCHmIgVgcAdomnmLWNyCnLL
6PDm53gNi9oqwyoBCVUFIwG7iMz+DYwU6WbHprbZpGra3XbDnt+Ii6mHL9Z5gZY66+Dtm85yqUNx
hjn+6X3KXHIa7M4QTqOFPJe6ZEe+KYMguTw7DEhqle14EcK+B/1OL6BA4HloJLuBXQGMtipLAqb4
PHroPccurRPDmFMPZcQFy1puFQRgFRtigVBIrGCe6egW83nQGX5BQwedYxtSHQN2kYfEwmkH5ZUV
F06xpju88Mvq2XpeBB487aSd2y0p0X+qJFg9QRdMo1PlOi24Erp5gtS2FzSN9ioPtz0Y7lAAVnNn
D3tvXbxhYeq8P+xuomO9yBoDEDDdzT46XTWlsAGnzhpvgsl7n7dCx0oQVaw2rHpACRzPU2hRRhtd
P/tvAfR/UdF1ge6fkSK/zDGL3LoZcqysUDVaxqaqewJhBHuQcZAe5A1iw0rzIApn9LKpGQUpkDJp
jLtC0Am/7LvIfZsVP9Dd/+f+eMxMvgrUw2/DYx9i7WY/GOVMfDsk0nXU/dibB3CA3MQQ8QdlKbNN
pS4EfkIDwAG6WOAmzA1h1dvz7E4Rdj+qETVdBtQJznE93Nvq7L+UmKCAtgBH187lWqxYEkwjQO5q
hINC9EBkZiOIkGX6x+Tk/r+YrwdZureH9RZvvmgIxVmwcYd0Pe+MjmiKQVMGL7AHt5UReT1i/+Vf
fGyy37G059W9zooKhuLc3lgbhR6odjrXhmRKjD9twow/+GRKtF3yeWKtNZWb3nhtU+vkSo6BwqU6
09tjWq2cviQ7bWrlqyqT5jZP7P4Nna55CAOXTe3y2qFmFZxNlfkJYASN12xPK2++b6MQEziIbS5J
R14F/VuQf51nRcrG5YVTz05ORUmnTteQNcgRkVSEqfLRful0TgfpTsj8qvHs4tfdb6DdXmD5m2HH
eoO+kuHNeqAMOPR6TBZFirY6FyUQ7DcPFk0YS/+w19m9P/IbZd3i8NZ+/jEbc/RdJTtZH2ZXaeIh
1cQFWYXfDwuvtc/P+Y073VJuBUpMFCiLRZUBPbZk+7ZTXduJA/+rByCl/V2r2BViCPbEarhyFEL5
1o5WTMh209lV5q0y1gr7JDnHFCN7tRwMKCmw2kzw+y7JYHd4SAZ5V2O5mDmlMzvDsrReZvmJl37g
tnARh8eZAJ5x4a9gn9kfalDRtgQe6Hgt8JG5NmFw2wwePtS7g/ZvEYRivyxA68So0FUcYjzmkNxT
LHtPFYm42QQrAYRQ04lR8tnQp6szN1rCeEgDY3NX2VDHUNA5v5y9zkggK2+yF2YSCrKj09HU854F
NAyZvLmIIux1cUwBPgF5I8wdtt/cc8Lhh5bZZ7+9EPnzsLMgNqmjI/B4+M92G6eFg1H0psReEA7u
iagiObUlNYijWDBQt/BIzrGx2X8C0TUyPQkGR24hHjg65AEGLiUnxz2B3mDHkCnSEbScUw2Uxjdl
GEDUaPNBFyLEkyMCWEkLzWB9xznw8UH5ys0af2jBLcml1J9qVx6Ma81a/q5uAl0tVTTqI3VUni66
mkskEhllQraKgvYH4qofTEOBL3xgAy96m0hsEfliV9NgKxpRkDa2D209bx7l3fLuu2icsGGOdrz7
l4JIVqnXiQK9cQA78YyU6TgE931Eqk1l52KkbM7MT5kAI0/YpFCpbCamnajYd5ZIZFBlw0EFeKfN
KYomxG4avkv2Kudt8N2U1TEbi+4lU3I+06RC+QSYs181YKA/u8y0MbQGMnlEH6ZrqdGTdpq8gndZ
Q+bno+7nZWdp7f8CJJg2KDwUoZ++/uISyI3ctIqF1S3izRfs6Ho2hMb7ZXCYtR4NYguqpLEHpFeF
yduqyDU39czS1slol+r+rzq0LyOMPjQ5XIBz0cHlHhwEk5+PJp4l8b/zScPwBCcFA4GDU9y8Hwsj
hIltsS7S1uJQzCmbHi8hSsD7ytzPoFPcVqLUPMbgtN27HuB8nA5V0LEbtp0kjI+/GiNt9pc1NUzb
bwpOoC7Zx4ilqrnJftrAvbip2mSnum6YocbJWlGwVHwNHj2yU65oR/+YUNC2fa6Q+sSfisFehimI
99zv1WCG0YITz9ZeDTuBdWRBE5d317UBnpC2at6/Cx9z/BTltLwgcIrRNaR76akmS9uTXsBiiISY
swONeJxVPCzElbJTuwhE1HNeUdhCJa0MZfl7cfeMRN+V1jMnym0n6ssX+GRL6rUu02ASKfOAB+FL
xTmEaaDadjM2POo45osdVnc6oJtL0WzzD1ZL1bFOtcTG27pRpegtefvcm+4n2JsBiAt/Amp+Wnq9
duQZNAfKRW1QyY6zVdpxcknWm6VngP9IUF9pw7Tz6BrTx2ez7qgCYXJoAsbnSASIn35FJeDLccEL
W5xE7DaFcTUBChiCcy4ZXeArB+pfObZn1pKnlA2/1C1QhoXfwaTTnHR4qcY5cLsuzS5P5uH0c4rf
wa1jEP29/YYVxq8qrgKMjW1T7ByDL8KkZt/x6rNcuYfULHge8NR8wkGFJibDTXFGB8/MgK8a3t+0
Tk9N515INsyOhvr3LXjPBJGwvqbIk4Oc85xJVGkfMIeA76EEXA7DunasiEsPTjelLmp9eEVG5uwD
3bSK59MZHQrpSUSrMU57c23h2xEB6qTysbyVgciWCEES/R5Ns/nrgbeoDTO6duAr6UytsgaYzWSR
V5EwKhUlo673vHH2XDkSa2tUVScRyqK6YSc9nlWPx3FELledkwrAYIjChzRC+DMH30JLW6nbyZHT
5APBLRNDUk7BLzUQ6Z2HresV95d4w/E4QNuUWBmEG+0FxiE077jdccp6H/yoDW7gQHjl0IFj1x0B
r6ody+XGMJg4rSSOUt8JswV60HYFCGOzsqAobRuOicVrE34xZ9jG83iWsACrvHleoqvCaRb4+3vU
dklHiBfB6HZgHHO7c71hSbp8HyyfQdotWoPQ4j7MGp++ytVN0FFjYp70LA3zUbFI6H8eJAeVfyvS
a3YzZjlSJSgPe3tw1yR7o3slYDfkpfuHiD5gZZvXJRXYbY8GKY3SICvcIt5sDsFtU3BiZ0LNIJX4
mgI2ko3mNtdj0K8XinGkLCndAxkp/9v8jTgo8e10kXGgrjQoEXx/KeHYy7U4yLeuztSJ/F9jKEtB
m9UsxGbuwcwkd5ouPGSGjjirRMp6LBzh+8uf5eib8AUuxHYkU9/AFeJWdG7rq09N6ZnFIY5gZLmw
bFX7XUTIPZqX1T3Yik6z8KoVXIR2kB9bN53ei3yXt9WyH3PVAP1VleccDw97TdoZmNNCMA3jRKsU
Ja+dny5AkXTa1HdzgWoY2UHDGaJg3a5mCaH8SYjz6ZM5/dhSlHtaEPHZcedV7X9bk8FMvH4kHI3E
r0t5sPERpbO7pRjLWX1wwgwfD02+iafgeyAUjw3pEIZY0zT4MULdLHcn7EZywOENoVvF7GwK88wX
k8Tk2BIS+Nl24OxyMDMegoxv0auiEzaehk9kW1zbRv9FqEZVHc170qYON34ETfoPx5/JRRV4IBZ/
LCDwLA7xq83ziYCCQ3LWfwRBqksTB6Cuv2asvRX56t4hP2O+6KaQyJUAP59e117NMrjmBDM6pEpc
mT9MsYMTiwTKQVdU+gMiRy909EQrg4J6hSILBy2g563y2qPyZlOKYNbBYJ682q6SBIKqNw+s8bb3
J6gc/velMqwXFJ0+b8IiJs+zTUE/iFsOvftj7KIeh2CK7V1YjCwSMfq4AhLMELBvDKn1xxfoCymp
Eo84/PG1uGMsBkgqiIC0+JGWsmp+gi/MjCOyaTAGqRk6ggvc8k6coWMzKWpQrotp4xX91qWzhdO/
2sVdeHOvwi0ibfJ79EJenz3vIrelOCBiGGM12mCqLA0gvRJvoJEJTNYjF1yJWVXIVPjKgKJ7WmjT
ReAwUJ7vEHrNyiW880WVZoAkSlYcAM78cx5tUjc9v5hyR/qoVoK7syQuT3xCcaV9GCl0Th/ZFPM2
b3HY9xvAetcYEN8M+IFBNf1pk8BMgY6YujWOnvaWJgHbkOMGuGJXZJJVEWm7s5HgTMY1zWj9yer9
UgM9RN4FVL/rz1+DZum8qSQM0W+JGa6Duwrpl6qfG0dSoAeSq8+I6TT1iFdp5ys/6v+F1/5Lk4vW
CKN0LVLNRkO7zG4DlTeBXFw/tBJDQVJ4t2V87r35fQ7t37zgK0wWxGPuwZ22hfmWbmjWVZCyG9MW
N96SatuOohDWyClFGKhBe3G9MRV7l8ovTGrP2Z7UEPgRDsgI/ELs1niFYBeEhuvokZM6ZzEDBrBD
DCtjpQd1/Hc5PfR+eW8Or8AKbCMRLqSn6onY07CeylkKsnTWk7VE+uv2rXx501thCcpOd5LP8a+9
DbdFos4L2GVU6Jl7eOcveDocQP0opfeUBjjCn3wpRq+YCiSlGAvD3FAzAsJVJYJkzWwBJz9wDVYM
SBqddvgpDQzbwzWuXaG9X/U+C5TmBOW6uU3ExvYcfHOigaHzRNcwg9r51DrFJmSfjEcc2eMp3WpD
YZVsrTQhmrXV6MojAkYzS5uIEHPP1Xd/lwJ5usUInQvprkoipDlzsSQyaYChfLr6BSunFt48vnFc
VsmgYgyH1lq1xR8tvdV9GS1bl26hB62tHmh9smVyuMNs3wRnjXi7KqSTZ61tECpFw3fIV4M9RY3F
Xa6cAeeY8z1aUGIy6Y+TSjvbmpDIeR7ceoYxGOHL2zzdLjGMTClf0rukLMf++LhMwUbLiaxS7Y4/
Q6AecO6NlGumyX8dAlnfiZmQe7mSfuxGKr5xR7I9LGWy9z2NcJ3FpQO58FAY03frx/n1dGQbE19Q
PiZAFELcfAyKArFSoxDJPohwt6Lh0PEhxGwrBbIaPqLg9VWgQYstOfvZzC0L3Wkl0Vb47tOTiQOI
qwpENDTz+KnMAqW4BI2/heQUWm4/lj0XUnhqVeGiqsiyRsqGTHO959E7S6gVYtv0B6qQyjJ+VFAG
hxpXbmIsicCWnw+dZ8wy6/NFniR0LRCUVHthPYBRUJ8w69y2oBLw44AFkosS2/y5qu05cDFJ4sKS
RYHKSbytOLdiM6PuUGNUhJ8+UwsHDuLWoitS2C3cq7kcokGmZ+EFXGJ0M6uQ4KpdU3KJWif+GiTB
Kv2eXVpLIHuJFUi4FXGS4YzRmPVHnjv0eO2iUGY3BBJu9yzvSbcbns78JvFHe/IHbLobKEWnqP10
IWFHp8zvrWxmgFBAI1foPPKSH1y4NnlWCww4nQICYH+nelsUba8tnTIsVj7cLR3axoFk9vQ24hMF
bDOL4hdwrs/l5NXMgRTeqq3LnIeI9zcH2o/vvEZKjG+GszXxvqIeEdZCMD0/UI5AtF84cD/9oig0
3oAeWwqZuzVDIc3Fmqw0T1+8ycrxNBUqfWmwkQyOK3FWTDfvmaU0U6uDcHZ54HK/qcYIo2zR45NY
QYEgItwz/Gg3M5C4bvOD9FblWvJd735UyIW5Uied9fDxp3iWueV8cwYWPr6TVk3UTShzmTT6V7iX
vNgqE/v9ZtP+iZjwBij/2ATVdwvVdzKZa66noT25esXF3J/pbVYRqnwBfjycrzHO8CCUss/MrRnD
nGDbNHebjEyjCklkpJGpnsaCUguvEvbPWcze/PgxZcg4oZ26+8bRtFH711BhjkyMbxEg7gvvva15
ppZhSscQIpUeiBg25jok6hWUR9OXhXCFe+BPKKAvqEOKTovQY4BQYAjq8kEV7/AOdJ4kQqoZRad+
ZgQP5LTNqMNLbDu+72AqeiUUEL7hK84pO6xJo8qUO9Fd8vpklH9ah435mSHnb+fjy7++B6aP8t6z
fN2/iEo1vUerGKQ/O/oxqOTZQyYNn9xOniuh/TJQsKgpkOpLx77BT9hux54zizSgSDT3w0FreZPJ
EeIXX9tSIIKsXyVSF6Y4mjAdUgwaig0vhdV/lb4NW6LzSfkGE2T0eaXCJwgFcJefzlTSLePC69iQ
i8CxMWoTlVBKALhD4XUktxJ3v6eg7Oi2XEfal7W4Lht1tkwrt6Oi7x8WU1fvWlyyr48m+NsCgVpX
OVWSpHXKlfu8RV6wDImD1ERIar0P1JsWNWBkW9E3bH13CIpRLLuHLb91EnoUhbA5L//u4YKCWXgw
MP0eUxpNgHVe2BasGSWqL740KTQ+bEPiAJuNczDfPH/ocCAIhakP6h7eJAkukrcdfqJTgPqBUnA2
2UHimUI+iSjUi64BjvU/zkM8LkomroDVISw2EEwUV4x7SxHID9RCzChCODWlq1gPr6v6QlwM+f9I
0RxiNvUJ5R1Dl6ncibwn5L8ZBRTQoU4uFQ5UOEECleXZtNHgN5DMH8M4F5c4LULu9cSFv8YwB/9H
bJ9JQeGrqDo0yPNuT1RNkxd39eDCiuX2mYvDqsEqQFP6HJDfxVgTbkFAmSPGoStqxpG6kFox6/Di
bkHWD0LA++Mjr6EKYVpM70q1hx9KqVZanc5O3VLHuaPp0HyfJk2eWBj5keks63E741xkufW9EEBb
yeBzyZ6SmFAjYvTPOr5misQmCvKlvu6hrDmPbbtfHgEuHs6DRzJ9Ho0Zgr+fHgbfo0heJAwir2oZ
5cXso3bE0mH7RNTmgi/xjKOTLUNBUDN7I7TbKbYiExRYVOVbhOWzSvMSRZyYlAp1Jv6lGZdZuM0q
6cSQ/+AXRgpZ9vAcqcLsP7FTpRZEY2ETCbdlLeifHrpG9YJwaLLeg2U+YNWfW6SXRBxYFS2eYtGJ
bQMFJLXeT1WgqKbPmyDmflFmg+XPGopbUaEw+kQNFBGYikH5V/U1SslVX/MzDx66S26i2G8jmT6I
PxC5EPklDVrdxiIXqZGTYfPUWVAEocii2Z1WZKnik57ipuWUZW5g9EA7x1GNn2A557pDfSsC8+E6
vSU+d4abRXSXjWMcTjtlnzQ03TOjsvhyQEQ0UH60g6ExElv5kvN9St7zUmDa9iylJo6WHdrexxwE
vUPluvmsfK9FMMTYgi/jF2P4ulKCAkxFFznw/wu/9NEWgvrbVCpiord0giWDkDINGVOKds6VICnA
2Fq2prWdFKk0Gbx/FhByL0BNsWPDUs5YM14496rk3VNZ+ea8N2SU4hU1gKuiUqiwKaSqPGwnI2z8
fryz5PO3yAmf9Ln0XNKV1MHzMJa570QdmBXZM33zclC0j7smC4lWZIKIVlVjPn0jjZvzEbZv+IUP
O8djqo1wfQukDElHwMxa1bVH55gispej9gkYO/s/h7xteMtNYIhMNXsDmYVU4NZ2S521tAQFa18o
/HN2s9OSqv6sY7zn0O0o0hUjTojTyHY7JYRr6KCvwF3lj8u/AUY/NDnVX+bdsWAog8yDNvd18rVe
GS/3CIOwiEqlEduxBN+XmmOu73DcV0bKl03v6W+TgHWIh/JUge4iDHdgJp/pwV7kOR60AtynnRWz
pdkGwnjfhc3jLbPQln5Dlg+wvNdqltE1FN17FF5+bCB/ZjmQCtwhSUK63ed2/BqRbPuql0cyoy3e
op/ApKZ1msigU9kprnsj2NOw9B8XZoCFsy0NuzOsFWz4ZlvYY359wWtOhfH7+aHduczyqljH8LnG
skESG63iXyg133CTuo6ZOHberi0Uhq7q+mt47hNWK6uklRHHkuekCac4v+2ZoAppeJesNfJTVPLI
zO4FPuPHGuyITG57ILrif9DHeLcjx6jjGvT4OXzG9huCfMuV2RvWkVDxdmda0LMZJ1enYfbRjKtD
CRNjFcGUnIX8kuYRIhev+usa1Gm2Al6GXEj++IHMbBKDuxFKcKKaVk74G732Hwb34+GJmU3Oe7D7
Gt+6tFSyQ7Ir/rhr38kcn/0H7vibfYHhj9Rvzmqx192upaRL4WrrGs3TCHPsAyolpSHjjB34aUmd
mrzPsjTD8TMq9pRX/08g9fW20A5h1p/6VidmuyzHopOHxfL+tGdU12a08Pk+IahG4PwS8ZGt4fEq
DjvtMtaWTpvpA9gucBsgGwv01wvKMoWkRBjDpWbVfvoNjTrYOtC9GmxAe1rxPWY/ElH7aiIorwrh
4xRBk7FInTeksep2BoJCk6wwAMwy6TAXT9jsII12EL3mivsSAb5YjEX1Qfe0yBwvnausw4DmkdSM
mDqS0Qx+U1Auk/G7x6bsLlwV+UG53DJEz8Oeofbu31UiZSpx6tFTjTDxcAR0ZvyRT867L/ofwfFg
pLNnjaQUjxqrE0eJ+rGRonNJ0jtd+26rNdLKdgyIrCsZ0Ovi4l55b377SLEx9iytA1uoJy6OeG1I
D9XSP8AyA6zYFTYyjC38OyUVbEh9ox+Tp+DZNeDjSpcq9KeeAwYlwz4r1L5fpFyDgpGAGVh0WiUf
Jz/hJ35+68vtTFkD3xlSq+1/dPQtR55ZjIVnv5o0VOVNsl/6C0nNo1Rxd9+GZELdDx78zWAVy3KT
9lfFmfJog6DfQKwEh1UPPM/MLs03VXyHkxvR87EJ41nAl4gF3drP5IBxEjbgLXucs2ay2c6LAHBG
sm2dO6UmpFWdwfRYz0T8vTIt10w3XDx15HE7zr/GSugPZNfQj3q4NO7pYTy/YmkYePWK3giX+NMa
zNWrQanR8/PgXBgWFd+giSY0eadXSU1WJtNccPpnvIHz5nhKQojHCnyXGdoQ9h4ZozsbUM1grOiC
0mjNQBaqYZDaR0qbKUg00X2inOBrP90QyhDvBP+699UelkPjEueOR2UtyXy0oHlFQurYQQX2q9cT
908nIjx8J2q33Bf1YsNYh2Hc/nwGNZnvT/OSFoCKG+c41qutXsoRB4GHwjEhvQ1+MgLyZoSlEy01
edE+sUDOXRqroaeokZBBKqhPcqJb/ooGVizXES7WMpG1lgGq1Y4e9DFRxJBouhNQmY0cK4mYyzzI
2NP3CvsmR4nsi66kporjYl/bF2uHEgwWsOHTHFU432vL7Obxtgm693m1mmP6LZfAJfqpIfUWXkSP
5gB7f6YpvMZtMomufx4+hkTYPGiRXeWLYzlIea4UNKL9gh9ok9W5VGKmu9qVyU0WqSbn+HujSjTF
FLasWwRZo4iAh/EeSQ0USylXx9NuUzoh8u5GYm/3apf9FsvRrpP0IxrphTyMs4/sg0GlBEgFAzcz
Qd3A98T48sLu4py1ajsxZNa5Tj8p0BsY6UsMJduG7B/WFlcYvtLpo4PeW6XEEuVzuNPzcCRyDOyX
8/E7rtsxT5PlGEjcaMGCkyMLZjG1RWTNLN2KiM01Vw4AB00Faba0JPpkeDi83Aw8k5Bl/BZIRBvd
GjP0d2jvHIcxk5e7Kr4BaZ+c8qn4lokFyxgDtdrYQ585gP0Zne7QgSqnyUI22Hwr2Gs1C3HhzC2B
7nsdlBDlnM9pPYgkCN77iw4GCLbM+funcBIBzUCx84u05CUiA/cZx/C5eHio6Kj5fJksJ7VUOEsv
LO1++ytmnm2AuJCDVp5S1UulLUzGUMCN2kD/3TpFWIkX/XsgmMj0uLhmBSF5eGeEK2sCmcb54AB1
YBgOX4HUa1hBHLMclRXUNg4+zF5vpa4nrklR11qQLEDbGYRRhNIcMUampeHp0FP7o6G3L5eXRAyE
r9xZE6Pf91AKTt/duZAhMdd3TfPkde0q7I6mNQI9aAQ2jl+9GzW2S29jVsItifbFKXM4A/bPKAk6
wKnOLxiSsADTgikOVAPayEp9TG8azd4T3lpXZnY/07fNOA/ix/YTMrN6BRQZGHFD58oUfH+hLP7B
VGAh34DrrPtrRRd2ChvxbSNGGFYRKLQKV1X0fF2PXPSRs0mYELRkbFS8ipbcoyjAnUvvvSqrMe0z
8aJc99IofQ+dqITIL6puACvqRiqs9lr/w3amGXMYcyFZh6xNchID/GHdeIYn0rssUgK1wWAmg5GI
VkwXi3dLp5Lzyga/Et/8ETimbf3jTTiCFV6tcoHwf+64L4M6TTJeA5rcuDl/Q/SWAboORrATMDV8
0Mwjnrmxm6ftFM64E2p8ljOtlkbNserJhgz/RYwdGkQt460n6WE7mmb0IeDx6UZsW20c+pBp+Q7B
8gxSTCG6OPEsul7cP7gZTmiJ5vIG/bC6vGurUekdxi9gbWOrMA72KcwmkitI5RkWwR1SjjlsNWi3
jDg9c338Cm2dZNTewMJWNE3EbTrdENiVePaoGm2DQH7oRiZKObuKv4+FyGdfN8jU3XEK/7HbIoSw
n8YV/hqkjmPI3Nm7sjVMOdkvy10tJfbOXkmIsHuua96xjR9NRatMBk2JkE74dY4T9jAm6Txbbius
orRj1JVubS8ipsRYHiF8du3RT1SZnZB1jLUuCC1hSaoUhB4yP7LAvR9zPDZ3wFC7ONMIycKcXBew
ed7JvWD4sVFdCkgcHCn58ss4B+o79Ldjd7LR2jcuuehVmtfc75mlfRp/JQKUPMRV5t+Quk73xKZo
CT7gL9obpzHA+Iun6RRD80OJnPHTlHqGTkVtiemaTmzO287FLG13/cN9ZmdD4fintgQ9jagLuw6L
ZcarOkvOlrQaDooU8mJTc7vWhkp1d5oUtOWbk14PeCRtj9tw/XQTeacYWmSsJ7kfP4X5hXymOX+Q
1JHgEBBWaB+EyVz70Qsal/3luKXgl0f/Xh8Bxx9/twN8CUKQIc/rLwf8cSTRkVWmFghnrqwF5Lec
BOKccL+J4t2TmxDVlL4EyLqFIj92BGUwXN34fbpClLUm5dKAEZN86V8IU+pHuH+r/XbPXP+6jBD4
0+59UJp6c2s30+fQYlTHdBgfFDrJBtziQtJ1sAR84ti4GWIf6laaMwTvCVpUB3hmtAeAik4v66uv
IvHB3USBKjFGWqNDpXROWu+mRk/kQRzUgVh3tyaB8Eo1edRx5HeWzEGt/qL4THm0tQuSuHQHn+/T
vrf44hYTjcCUSmrO4c6tUY48X2WT9BpJ5bYpR+ezqvpUjawvMzhJhVoNtGTlN0RqSPD4LwyA05Nw
SX94kJQPj7sa7HMLC8Qiw/4NzGv3zSGa2wmh8qEGp2BizWYnkr6H/1XGR9FEBcze+CFQwJR/2vS0
QWZpWGHAaLP0/O1MkhUw3XxmEeGNiPuEgWgKFwO0lKImkNm04CLPGkXZGXaajxSvQXz9TSI5xLlH
WuLMyGpLPx7vVFXFEyz2HNkUTNdIujvJyLlCAVCEh7R0MvAk1rlZmoY9ArKXQ5z6nSnjoj6Sa4m8
DCGGRM0p6O54cLV5xk7sypdJkyiJdV5PVQcN/VZuURmtGMqVd6Ec9sHc8pbycZSLURpJ1s8A4iUI
R5dGLv1MxB3RYsXpElSWXFI518pKebYsQo1ft9Eg1arPanFJvxUWIb0woyuHKTfVM5RJ/3afLCf8
8djG+soBG3f/ENhnwCK8rXtKX63B5Z4BKRYrU/4WzSXnn4fENlmFwaKwlXn2Z4otM+WgaF0RcjXy
kc0TFjpIQXEFIWH1hlgMgMaCuYZo87CXvIObiOSFFWvJ3jtrTjeZPd3Sg0RJSPJwIhQA9IGVgN+A
J0FcVfJUCRMg+u+BmjKpovuDO4jRF0k11Ko/T3xg68nrFplcInHy1911DYIH67juFlB9b+nPtSBD
SLtlIKTTWCMYRB4VyXeLhL9qzR1Muopw8sNcuC+R/izs2rLRbwttOD2fgB6dzsmcHIg3K8+E70qV
AhIph8Vbe7/VWibYOyqUu1wK52frBzV6kYcAXhHCeJxkt8+BTVYjR6SYLa0VQD15ubVQ9Y5HIR/2
ymJSoZ+n9EnqwBKKsMuPxiN6iqyzDaoAlYfgC9pLH6AhoV/C0ReSv2VluCJBxAJtnd6rSROYB7rP
667WxcBNFYV8dDF4ZF+C+J4TD9CL/PGqQZCXvUGBCOciSEnsmJyOiH9fGAg1CFCCHWf+psYP7U6V
cC6uULxvsgm60crrWyuJrSnLOflXa+lJzQGK50vnte9kSgVpk/MBfl7y5yfkJeF90vWqnFlbBD/d
KwRqvhed5fZOwtPTYqcsI4nPtBhJowLQT315tes6vNh//MUkxXdPYQU2W1V02EW6Inpuwh57v3ER
NRz2LtJ3UccbwLzisGiI+Y83/JcOhObgNQjhHd2VlaZ/cr8KoDr9aS/MzsHLyVEmvpunw1qmTyas
b7x7KM9bbIyE38Tct7EPmbbuvL/hwDvZt5Lkgz/UjEg1plc19coSUb1yW6ED0YClKOhiDP+TRFle
1zxIQn8ajVPgHWLxKKxSS+7JsMxKADTgADX8zIL+Jw1A3DBJWQprsWMH9h/0p5vP19LlI99G+WUw
eqowwtkcaTS5fMbxdYemMcaRkMHDMo1y782LODoS0ho5G9C9j4p1jTmGS+cs0xgbcOdg/HxncPWd
ms69eWANdd4BsZxMtbBTiUpprQ5dXHuGNbJDopkLpsoy5f6ByrJ3xtLSe2eDAMtc+TBjyn2j77uk
MgFWU5x40a+nKklzzvErg74EQW5TvucyyAilz40IK8G/MzDYmWInzfuM61rO1aoVUcD9faRj7YDj
d/Krs+qh3yC8562TcrkE0mie01cdJdB+7k35T3/BFoNAWZXfAUWaVSa+qUfw5yZNnientA1R+NSd
N4ZAJ5flZevNiMY0GE8BQv3N5RsvWcjj6IUAKNL6IHIkhJNkPjmToIgOAj9adZgLasw0ssDH+k1k
bUF4SqB2v/oh+HEmkn9gQeEqTr7k2i2kqjJCX/Rp+fyZbhRwU61zVIW+z5rbYsTYZTnoZAzG23ku
oJarXJdkibk5oMwe0kb9SJTuk1U+ksUNbonJnzwkUecFrhJRZLii/8rVc5feZ6E2JnLG5hgCCLzl
34iysOSCIdDh0JNxbEM8w2BkGPHESHb4lxkwEY9zJOIG2xTzEUIDYo5Ke0cE1HwALqTVoDQPlKdx
jHgL42T3cSLGPo/9OEzb6ejh8lOs+te2WlZO/uJKXv7NhhWstZxvDZSLsRLOEjDQuTGbh7ix/4s3
BmAkPrBYcLY1JSho+qWqjzMZZYK/fMVeVSItxUCXbJtAYd2NmpNw15czzgyOMdkh7RS19lTZxfzi
WARo9hKHZ9vzA5n9Fk/aoJFoMV8muv2gvkhRQ39HjhzaMIiCYVY8wRqx+p1NrjIyepmtAGa/24OE
q/n0M/+S1li7k5WQ5CWgOZxTh58WOUXKoKnVOIli+a2UjIPam0yoKx79UPfleP3l/w6OJGXagXvT
DjUjaHjzmkD+c7RxlQ1YRiDWbDt1L/QH8CH0GE9V49J0HlBoO8jak3x13cKjk39jhDX9m0y2vnnj
Crdy6bWWukDUVr5bxGyNZCkdlAisjZ61fEcFA7zNIGcD6hxCs9TXirpq9nB5kqZKBRMjmd66MJKs
pUGdyyij2MD3b/7jV+uAg/GCt6eHIpKjU+kq1cG+QS4C9EUUPGOoMdjV/P30J6fcs/gW+59LGOKK
eyUnGySLt8FLP36vJXFPL2N6gIC++Nn+FT4hZ/jVsbqpj8w0HaYeyj1mQfrwCYboQbxHUg92IE+I
JSzIUmzsN/69pnWJRTf5ucObO/iS6gvsvai62V8DmPuLHnF/UHxc2bLOLHIyNLbeeuR5Ac61Eg0x
YdfuiK2ov3poVK4sokwRXsmGA3Xrirz/oylARoe0a2HTew9fKcpRBFfVBEovnj3+rSZJ+s5t1aIq
9JYInNcplcUjgt7d2eYqfo/U/2r80gy20W+rdZ5etPcjOGwYjnqH3q7os5WDCLQfHzXnt8YEIZRK
Fzju+9YozawpxSK46PLuNzdgyW4qgN/HUiOyZsSG9xJ0Gkgc7Tihossk8u0pMQ7M+ZM7ANnBzIZE
jZ8Y56bo6jG6IumwRqHmb7xhupwO6RGBH5Vf5DUiyo74Po5cV3teNr302LtwXibPmVgA3Ji7KLlj
VM7ICL8cdJtYS3DNu8BKx+D6ByvgurXYu2QV7RP8gZoyOCiVWM0B8UyejPX3Rn9JYiJnpXf9RUuh
Ubn74bGctI7NY29S+mMKneIxR8goy+8CmuqLxNfjk9W0G8E9X+H8YOZj2AbNHwnZkfGn2VqRiAQ8
1P31jwgDYQ2O2m46k+vTxM/dxLFvX5rmoKLUAeXhJM9FIAeEZMiktWAyL6ni6IHG1wFXgknuV0Sf
L+FMe8+75Zuhcml9ny/pn+Cl33PEQL+5KXzbwrZZpKZqThYnxHrAyM7aCcAJ0cxR/662yOzvDwMx
RP/XluxAqHJIbyGU3agnDtI66xmT3w1VHvI+FJv40mIpBgVp9vtcACfKQ+j1TvGNTPmykkvBQjMA
Sw9UHL4GIVnvETD5z2s/GkqSazAy16BeWJps2BOdT9wT8jZBi/AmJGNc+df328t5MtPjL4HdkbW9
GzTKge79ZboOPZi4BTrKKsdXOK5XXz7xsZNaB/RT/aK4IhO589j8j59WtRfc7VivuTEQhOYewN2E
c10rLdd3EzqR1HseI6hco32/algRRtGS/Pxoh5XGNlTZXed7TAqJC4DzsVr+hcW6PJpWJDa/5Mcl
iyriUXoLwRmns7dA5SBPQPw4vcxz+2kx7nvSuEb513HmHk9r/TOigjL7hgJVsK+a2LWQdPC2ulJV
+4EyMsXHcZZK7XYOOUi6M8P4nanPENevcLK2HHRHYOhuS6MIAy4dNK36qJuuz4G2/VyfuJCBJLGQ
HLLYspMT42JU0qZf0djOnSMQDddSqobULHJjHkRS5rfXaoopKt7mH7d9EZBkDcFBBc1wFz67VDn7
7tWtnzHKXU4c4fnrMz/cBbxuUgx7EB+t80GaYAWdTPUo6yppec0nlg/En9WEAuvgASSqJLoUd3rV
78/gFygubwwO8NnxbGQ7JguQqB7NQgKQPeIJ7laz+IWeEUq1J8ULSoK6YGUc10l+0XnagcqLOvSX
r/2gXd1Th/whuSHVCBGiOavjBR35LSm/hV2/ZQkgAVrx38/hG+MFWn7TvYHjL4Az8fyYEgwQ+ldr
zgsCKIzr9s1iigM+8rRy5bVyaTv6V3CAQwKrJsdOtQdqF1QglLWK8FPXK+P/Ncu9r37+5h6Ihwvq
fl+p1krx8ZtezPk885UnKp634uSC82ZeoF3asfg9Z5Pd/eS1Sum+NnHo/xZxUK6QDHDfAMNns9qD
qa/J7mTJtNvwKLBJ63bPsB4jWJlp8vg9gFF0Pduf5chKklKqZcqMnnO1dxPJtpChO5lxsWoJcdfo
+ONoc0MIOaCZMue0oeyOzy5sXj93jrlZ5hyeJ39c6MZt3KR1LUeDA6/a2OeXa34HTpzF9DX9hY7i
RuYy1XdSMwHebw+r7/DKodYckvyS1zbXH4Yxl1Ay/692NftT96e7zped5dPwkgikdsOZfxcyKZcw
ceT3wxVZ270FszERGjwmv5sY32aLw/hVQhdbvIC410yFkUD0yKfCBQg9OvbZvKnQo47cUnBty1vW
HE2fnqqI7pYPCwemjagHKCMR/K9xjgnEIuiZmiKAUN8iMMFugZ1/rIhrbL9Hez0nrMG14SCG6NBB
yAaoPQUH0nwdhENCZzTVaG7SgfOvgrTFuWH0nhput5Yvv8X8RZi25SXJwsIDYEktDOYPWXkBkYAn
lhpBKfPiwPdvfUEj5m+woLm+UkXbrZzStrK7IA8Gp/dcScGM1Lj5HZh91wEzjSYITAkk/qmPDpyV
WJAsxKiblWg2J5Lvl2t7xNw8ri3cPKabBmqtPxALIJYkM6P1LeD2YzVvN/mLMQxonUJf4iU+58MH
fWVHWEHq6nbj2ulZFb6z59ZyOeYkW3c2z6Wd3wvaen3o1EO1sZYPTInwPfJh3mgC6yuSaOoT4MQR
FJc+q+GCIK6X/nNPS3p0rtSMmL2ovzu3/IDIi7lFH+63+bsFnRpFVn4/Bu6kCLyEb4TOHlEReBYo
gOgLoj3StZ/+bVymMLckeN1WiwDm0iJ7Eb/YDfgbb0PyHTU4UH+ClsPffLptW3bAfro8sO58T+o1
hWtEwE42eMGrwNyfooRTUpBqgIGlU75xpUJ5PXjBBm0wtsmu2kpCRWuY2KgKp3Bv2Xb3dIQ4sSbV
szeLtK5EI58j+m92yEkCKZNsQkukvphjlUxV1VB6Ub1zv31GTcDMYK9qlsN2hKS2ms6rPkwr42B4
4GIYhT1n+cppBSOOemfuLPLdNJR+n27Yj3qhpMKIGQIJ801RHgU453WsTi7pemPXlaw5+w76VHsk
FdcuPs7ZkSsMnH/OIWetEOPSd0aJFzxXq5wL2JBTZVLv4DHrubBlRznx6nxHvWRcALIKmjwv8j8N
3GKA3pbNusb7tMbY4MbJBGRfRLq9CtN6f93QtrGR/uLwpqmBphxJe6N7xyVfh+fY8I5AaMcqAS2w
AW0HA0LWXVamQC/o41n7lCfgau5B+gWL7fbUI94zMqfrQ1ryz7ea292En7mHa2/h/SPiXS9miEyE
JWr7wv9MYUpiXAFbWDkw5Txn3Ml3zBAYWfaUkeq6y1IUMett3hwvQFdu5v/wzE0exBQciv68wmOc
WwNwpKeZ79a02VBg5q+8WDBXFZBgcw7+SmHQ2LZ78UDTuGYE1n/yVoi+8OcBA7et+jdnASWHcbYc
WHxg/+42NWrGh1vdIVx6++Rscs1ZasidrgNLs1leIy30kPbmXBY4D9za9qc5hswb2IpNtER4B7EH
8Rk59Ws3VoeiJAhB8thYdDnmafCfRbysqHCzeF07gZLFn+1M4raka2D2peg8TAAJqi2rgSg/7Wvx
4w0HGS5MPK+muQiUk4CY2i24S8dp8TF7oL6d0Zt6hBKl8SPH+MVU8ygiyyjnFRzcjEEOaTwdqnT6
rZ6in1+Qf9p3WUW8UHuhPaxrGgcpD1Iruuz1/3RGxu2ru691S1naCbxrfSMdLt8jdhiEL6ncrFSy
p4l8nAn2yXhQi1MxzKt9homLfUrxmzdcZcQ747vuRTkl1kGec+SZA4Lexfi3v/jgWySHdyK2Hr9o
bgu2dPEEnjEBsQFcQTGfJxvwxQIHGWATwhUUZrNGbG4YJYYIKkPV457eRdWMBAkQLSQ7h2smjDGh
yXpm9tYdjpqchw0REs6oXmXJNu6RB72YW3dz0kQ2C5E3wyyiAB9E5SmHOpIJ2VzUc2hOQQsZnc0u
PLZ8uE0Ql0aenDC0EuM9wYrPeJNRyxrVcSFal9UkNxk/XeYF2XTIj7psZ/5u/sXbG6+2GtLGGS/G
yysFzqpAmwqi/oh6juWyKPyeQGBWT7O9/0znyIeP7/RNffdt8NXX8/IElnvAVY6dNxdyZWQv1kmB
2OvcCBTiuL12CmJjHjDWuyPBZ3/CtuhDei8hb4PpKkOle4K/RZrSAHA1K3glmS3GX4Arf2cpnadN
w5unTcieVF37E6/p+JANR47gu9OeYnRV+QzoXC74CgqKF7KTN8m6c5102L89saf3GoT29m7uSW23
4z3M6sVXPfXVqdBrqsuQV7+659XiXv/S0ghyv+PuZSzeZQWRAOPU/qsBr+I1IjmWAU1oUqk8Csa6
MPRPsWLLXmVFO8STRh+w3yKW5weyRZ3gRt3Ky3eyK2MCsu2fSH5BZAyvmEU5O7bsLOh/uiuWCkab
34F+oZHiT5WH73nNKghJtJ/uRQ4PKAp++G0HiHN5m2FnrVLFy1t0BPkcrZjfo2RkXkiFJOmtZWSq
oXK+8v9YbxLJ02b4Swd6YAueprfbgXGzJEkaMV57OF/8ManVC+phmkE0GvylDGqVWf2nKKQ+dbeE
IUXtRW1OZBfeTHC43jCNFpummOAOdx9XYrtCOmE1o4Hlkuh1TOUAPcak30Guhc9ZONXGoCvo4zuL
vJq2NubLpLJMrCqvvjqi0woVGXBqwAT+Mr4dqUx5VisM95JoB2SSMYTzCKCbbUnxqINmx2F9CjDt
3yxgOa70CPK/uSQAItmnuF2A7dlY+BRlW0vFaU4rHV6iMd4epQz5BxCQ4hripfzJsTddw9TWu0nH
WA2KckaNRs6boAXfoob5J4K8DCtM5wFRu+I/NJ6j7Fqv2BGevyrQ+hAvur0jY7JsH06t55tS8V4Q
r4S22+12a/aNkN6S+YXRLNfsbo4dy0THpNo4qvBKB25awoNUVm+RczO5kz1CtSrkFYSa1MeOIlh0
RC3GfZrY+GPRTQ4R7zlOjz2QM+XlGRDCr9eVDccPv5JfivRZq0jhEIkpfhcdFX2+0tq2FU+n44Ns
EJ1mJrkiuSF27Y8yAflnwmfyXP0nZpQMs0zgLBMHUmk3mhU/3jXWAmgPgfI9o8Les6qjKHXGlzN+
BMBedqMdkAv2RMqlYTHKDDB77KKtO5pXjxLLIOjXQoUX7/xc5D08wwctMPwwZZrX89+Ya5JKl/8U
/ghMgwkM7FgcgL7smC3ILIXeeXwsC9Rh/3EF59wLOQQQN9XUZ5SbrSjdoL49+xrqbcTFpqMfT2Rj
3VgrHeEKVqRJorkiPS/0zzkuzXIFI58bDdPT7ETPS3oiqgNctgio5RZpGqwYCWVPZxg2+a27c5f5
IGROVtG3aSTQZHM0koP1dTltXRcUEi40fctJlBg2yuSHzzIiML/bl9PktnJ7EVmqDUulivo4jEYh
liT6Dk/6LKkFRdwvdwy6jiwdpzvYBnKGwoIP8SAb6fDHMCaQm3ygHqbuJsua2ztyV9SOjPQL0tA9
c4UUENhDIRg+GPdGFKw00CFEVLUqpSiCIiZHa+fO3WypNMBtOdXztiYYz9CEPHUdmjQmwOq5yZ86
rDynh0FdISagl4ORHmsAwxV3cPCSovDGZd5NDk/GH0KqZwe3H3HRhhdNeVTbq3FmJib/IZKsgQRg
vlu9knK1rKli3T9X+OZNrRUOZnjpa38LzmDJQooANPMwH2nWYwm17aBSsPln/Dz+zxLXaJwErYb3
Ct9JG+13a4t1+8VMkqEcYIg8J1KqmUDGAwWazWGYJ0hWabnc//H2Ikw4jqDWn7T6MW1pZmhDb62V
KPgxfAiZPT/Y+k7xEngg/EZNGvhK6lkK3wV8+CldvTTDskxPRT15bZqiNhN0kS2uzNwfKplX0K05
Jzu8Wvb1kOFRjhV5tSAZQYUl1txEBjrRth7nbCG+LmzMLlEtCdstB13o9iIi2F7cFAT0fG8jv6ri
ToBzbBKfsQh11TVtYGUsinbsB8qQlQujiB+LLR6T1axcikC3DwJFV7/A7dKBtKlYZ9kepPVWFnkv
jtXYFSmro2q0uWSQavSKN/F3gMYppQcHYY+bRPhEQqmc0Llz1HZ9uEg3FuTygandZzRwGxfuHkcF
Vrk6I1rDXSzp8AaX2PEmvZ/4/a1pPTT4Yqf4evx05KIm/pup4HQmrodrruYL8DHQoknddBJgcHwq
aaD38xvYoIfA1tB0/SnVf4/fxmx492Cz9P7WYLUvHd1OErhgfZ9tfT13su5dUfVQ9+7j5xGWdVcB
KcJqiy9YBJt9rh91nVC8WqAfz6nOz2egtJ8FUFUKL0G3m5HFsdhLwbfivRmlLVccrckeihdjmn0i
Qm+x67VRVUq9TOfUiHKnNfpq1UvZlgw/pia1MxZAfTxJv2s62jTzmo0Dj+6NhDKPDL5fu+rQb3uy
zSM/baXVr8fhaiDdFO61etSr0qxi1l6zDNqUUlQhRapDRZWw/rxUpv5nGh0uBb4NJq4NbV4vRUea
bwi2umiYuq058+eM67ad2TRCGpSDEVrwqSBdODBQyL3MKD+5AvjLvLjIOkJokMdhUhkAVPpOxNuQ
+35XVdiHQMFXyOHZ+zsTgWh5xzadPIsbmXFliOIGSKY/IT4lB9L08XvyhcPNiqXiyOaz/gg/aCey
ssSD+vg8E1i4ydSR9oX6kCevDRB8xXyS8F2bWkyKcuUfrrAZH+J4dnZYQaGDj2qOC9vcgQSfjLnY
g/AT7TehlR0HF2PA53wgsChYF5/x1+ERScZRbYuItePL+zjLEecgV99G0puJTM40yZdbZ/Q5ighF
fuNjau9b6UnvHV6WNdibFruf2MBba3DrTJAh9IR1xQJqVsAdGsZNg18GT/1wznfQUiQkV4cMTnZj
xUMuzS0860O5Y6jG4Zci83K4SpnnZQuFKSSL6i9riszHDVVJKddrVuyQE2KuqrYrVm9b/iwPF2Ux
XRX3ldFnU03d2yA949+a8IfnToyARAXMp5TsDLtkT8aSLzL/H/PXNjAKXYLSt9WKx+IhPzhp2pyN
f7FiwSYu17QTH7qSIBKfGS5gAxoGaMdXW1SiCNfbE1QH5BEtFLhsVs1gye8lIM4ebSkFzqFrCS34
gOoiqti4Mn9v5Xvl7liqaHTBsx9I+nnQq974uHL0XimhXvC3wWVWFlLKgdUTVTtsJZDlWK/jFFjN
hXRcpKUUJXDd+DIHoyvnIBcTANP2kybcW8litx4DYhT/9TX2/GXCwBWOJtK5wbQsmCTO11b6XCIx
rXcOepzka0cKJDU9RkcBQZc3BtRnlysJmqRDpF+QMK5kykdPrWhAdgLJ7rkvYpfu5djbMVKxrVic
zkq3WwwSeFKMzv9u6dmWz7s314sNT/gRXPWENt4V+H+AWo2YGrBUu7hOprVDgfyPbQShKa0ZSnl2
XQOM5VSyRTfEf699atqEWokaHaP1BPM6nR9YTAHgyLQQ6CJ4Ks76L0Il630RikpTHdnG5y3rG0uH
gTkx/Islto+u1nbLO34aNEf6pMc9tbqZgD5+XAqsWK50YiAj+PMvTd6+cd3+ZvHrTgpODoXYQpCf
zV+RScACVK7eSjBIC25CfeFW+oIrzcHB71Z+0EPDE5Tta3An8CQNmyWL0PErfzUPONafmQdBfWDi
YJ0g0/Q2oUEn8g7pI89QbHlWs+riL/NIeXbaNBqsUCpjHBlrkJkt3aUFT9YNXYG9aiVwkXeclMwz
gJxXd9re8MiaQgTVAMfseneyTW+dOzzKHA88s8wLooeU2KbI+mld6FW2C0FdIIYMYWO9Q8JByvbC
iIrBVjyszibLLmMuzTQPAG4wK61ICH/UmVW6YMdkMW4XR9srKtp/Qe3RIEIySKIgRWGC4cOv0/W+
fCVSi+2VwzuyR0XS3AgLNAt/V//XeOlZEcVEX6gzlmLBYmG4RUb3pzOOMCaocxwDpXDCq9xC6KT6
0Tlraqk6bfcpNHYcqtuqfvg/4rP2mFeEPivf4AHLtYxLDV5EtUNmTrlx4ml3nbcXWVskJaNwIBhT
dFvJfU4faXKDWbkwNLp7DuVoiGNcRDJ4+Kxfa8fZcQVWRBhcx0sONZ85Sa+TKJzYuCGuleOYqINc
n4SenR+AK9FKTVxP/KjU5wT1ZFHPVMM6il3oKVG01kl54gcb94+uExrnlu2m65BpoVMJzq4W6m9U
Y+te6UgSLUttlAJ9ToDjnu3gi4gB/Mps0GYHKHl3C7I9oWke+0WpexMRGwOug38yb7iyXcHN+eM8
e2LAJu6xR2CbexIMQa7O+m5C7N41AkIZz/uOlCVzZladQ8hYXj2bqXCkCxFzgV4sBLqWkrvNjdqK
uA4yzb2yMhyQQauQo+Ed5p0g8cDhGdK9jFlSVGRGO0bNFCM3FaPTBBkOGPikvFniOKpn7JVHvV50
wsS0QH8IZ1/v9lb9Fni0Au1bQpRoIhn2pW1HOJbk4RydCbCh3w3H8Pw3YKKkIpAf6eq02SxDSKP8
AJP9DiJOH6ros1qeUU/dxoAhYXrLWFhmDzJ+h3nVmLuavy5gP2ShUPWqmp1ZRU+8rm2ELL63vF18
Hx4VCiDzVJ6m1WcigxzRGGD7kk9PKMrHJLlJDypJ2IblS3ekbXm+h8a+3sbfvhZioZyY+Eyjwn1X
bxw6LPbMnlYyNycEbn0s+ctqP3CB4+e8FGnW18qBnCUegFsqIlx1oEyAX/ZHxnPj2nChDYMEH33b
5dZXfTzBg7OSMFO8/M5ELiTnXwTZErfPAORyfNoQiFvnHyEXFajOiLDRENeZkRwnCFYWdz8P6gao
L0QNpoXdNKtuDXRY+za3EWDwMV2Aiwf6YZ50eKRjrJOnqTCJ3hZbEU0e9oOR/ldvu9TnypXHnYLy
27fSxcgquII0K2JFWJWh9yHAXIUXfr2Dftzeh6xeD9Q41JvT2521bEsT4BwXz/3aLXpb3zpc7eWY
5AFihkZSL9s+mrLGRa5dRpL6RjQ9Ig5WpCfeoMS6iTTVg8n+Lxw9HOB9At50i1u/rI15aX45phES
IvTpsZE5Z4qppf5Vlu+6ImMCMZyI/liUpH7ONxhnVdj6jWQX+E7vgaGudSmzl07peyAUYBbbxA0m
oPWmDVWFQcUfcNly/hdlSjYFTMEcv4J3qiNb6u9W/JAqfRgBFID/dOkFnS5dDPYGcbV3ryEyhacD
Xjgl+No30ZYLuMFJFXBb9lpMoMwtCrkZIX3dxC0KNCuKEoln6QI2Bxlr4Ka5UNda3+xoSoXW2t5q
V655fU0QoTUPAbwuu4IdQ4b4Te6Yfu+cWOOA3a5v3K98aypi81rf181DathXkZzwdM7tPk/yHu0p
nT0iv9qKQa18lGPfhrPXywdNagLn2R3mT/LgHWicMbQQNzRbZuMtAuamVgSKMJuaON/sMlU2cd8k
6YvwhbAAJE/xBwbMjZuMsStgWSjaLvuMC9YDiJlQxAjWNTL+GE5lmu0mGa9CWFWlVH92b2hc9y4l
v8DdW4cJjusJOVTFf6HA9cC/0mbTEev1OAbY6fQZktUoZyu6SbFZS+F6KVxKFOCOJTc4ixP8lfAP
87V6pE3A+nCL5ZKc2+l94LLZ3q4+VWI7+L1Rls/LFKwLCYWR0eXpAU4sy5ctGwviAn0+2FWHG5tf
AUnkOcwGKKhj/WEQs2VCMp3C2kJzjSfkULy+JolK4zGgY0HhK/JnZjsT3URpGa7rc3Pa4nfkQpyP
v/2zjbOJ+I4pnocKlbLKsDpCuMmzcBvYZmgl/uY28F734wHK2Hk4btpX9OWkCqGLJRSRHRY/1SNl
SazoE+oxET272/9cNznNjy1UYWdGsIY/z2XT7/Jri3lzLXYgSU+UoyCH/CTVfOF4RiHA55XIWCMB
oaKQMyxp5SgZEkS6U3xUfBHaSjRYrDxa7hijP2H4kQ94/NMLZJ/UdzoVOLNH2RcQZE7hSAkEuzR0
XOIHDSyuKiH8YEicMcJsXSGkxAwNDk6vCGXHNnRjAWem8M0xyqoNhdMiglg9KhK5J/s2DFepIxrA
KA9kZLu8fKeOG6GcuqbCeWyIuAyukS6KMxbpt706GcPbgDd7UrPDolU46ay45nj/QthWYxLJW61C
falOHYg0NcPIx4y5qzXGuqFZOjJktL3bi+wKFBEQkP74mzTyj0wTbnIIOKHPulUK5HsxuzVDRIo6
/SR1tVjPfxlv0ezO41Of91IpVT2vQwz9n9Vi6ExTUmTSGpy2vgF7hRszMjF8xZ6oaJC8Jsu+UENp
xsYBlH5V9T20H2sz0k5zS7PO+LvB4yOik+/EfYwEdUVqANi88tygMFTQtKSJyA7CIMkIl42wGtjl
Ob8ckHMiU23BfUohrkuK+Yn76MG7ncu7ZSwNONf90uUeoisNeWeW+VKxWB6ec8fFzeCzZ2dOJpcr
Kd+YSWJrf+XwnHurfmt/rP1r59GdtrU/dqiwD+ZLBHrkA6ruSubMDRcyeE6l9uB9WqdUpFKFZ+N4
R9G0QThKQ3jUlB3dulJDzi5zoMjMUqXQ4nk45yazmyH5XdKQb0JaaGgfOnF/Ewt43nrEp4kxKVmB
rVgJpvncn1v1aq8ArAtyLRisLqFxxsjGoSTvIoChrHTaoOspyI4ykphh008P0/cYwb3I38HBEaOF
wM5rFz140+9WDJxve/CesOSs7zZakOFWdx8J8/TPyaymjhiagqXG6OdOiD4yRhT0cVIPYtrO5eOo
Na+vIQYedkk1VuCDiB5q1IQX5kD0x/BPncOubbDRxs7VA6G9dkJ7VYjTe70Tw8zK65kiJiGnUraW
Cm8btm/Jx6LHFAJqxqV0w7pmy/CAqD7gAvKlWb9q9DwpoDIGWUqA59hETLBn205tnU8WqetHsyXU
jwcWMtni6WLnVPwq35508dd1agrf6t2H5IKgUndpY2ywEVwWeisl9ybQ0g7ZZpIFGXX4KPoI2IFr
nr7x1JbZ3LFBowTPBvabLyxQrWAUSJCT6+Y18bMMagu/Gcln0yRIywlL499xRzsudNUbHoYF71R1
udYJho94oH3MLLV1y2NQ2FoF069twQaGQzn4DvTUui59aqVuuL0XVZCMVcgxArRYUfOtt59fDicK
FdDb3Q4JhqE+CkONwWqV/fLznUDv0K9fRCTUNg5M0WnjfTmXdHP/wCM/f2dcHkJKWR5gZiMCWNn1
7wS/wd9AzvKB6Xa67Rjr4aYZc05puyZlymD/TbAwlrt7MSlWb1jKVAIXlhn4JOcuBvDKiKSLWzek
Xo8HjAtBPLPonv37/RDzfWPdxGsSEfWuCsySKhj37GY0MTmIG5MLkslp6xxlqyoTWG/aL3YKPCCG
wwdpnnl9hvpAbNxGQDGNgQAI13RXX4C5NMWYAwZwiq3rOF5/KX2Ek8rIOpg0dYh8bsx9xzy1t1wA
mFY4j0EO2dic5Na7IcDOmSSDqdbVX7bg2i2IrERixlMRmfuIvRyiNd1dCPPqQnmTF6plsOSG89ug
Y+GrBjz+aJfTemCb6m71D6ykMOnx+wm397c4+5rFAXRP42c3NCSGxV9PbFTq9y1cvZsGN2h8X2Th
e5mKvexBx4Md1DPJvtUrgQbuN5vXoGoc41JmUGUN4K4BttQnGSypp3+o7j68u/7LflprQ6NKjuH0
6rfe3C/JG0q2ysWf7cHnZxDPvA6WkNSuwVzgYaPLBbEcIkDZddI3pX88pYPhQLXYirHprcNhHTMX
YcZEtbcQlxwuNV4sb+nrrO1xhE3/TFV0nyrNBiI4zRxsdlOkQjX4uyONz0+zyjlCE3kzOP/tbwlg
Hhrtujma9j770tu4bjUOUyrTOQ69vgUVqO/izIs81R3LrDkO7+9PanQT/JjsIlN8m8Ns3jLCNPPI
MQr5VFJHz2TOBc/u32bR2IwSxe+e3rpsWoePt1slED3fNFFZJ7kaNchv0RvuMyfWvfOKRzoOAv+y
PGZjP/Y765Oho1d6wwT3GARHvgApTdkF9xNLWFf8htkOtX8yrWT/NMJP1IQUPtzGKe4GWGqtiFNL
w4NnTYlTh6lBt+z5mV8vd68C93+FxgSPuQ++trB300QeKyzqpMaZsTijMbQzHKOcOVRteM5A1mYE
U/wD9HwBm8JYES/E+ZHuq9u6Y3aGICLj0i7TEIAP+ChsKbp6rIyxKmo/U7TPfdz28C60a2FBuw2D
CXqU5jrOvBdRJmCIfu0UcYLaDbQ3y81Qcn+6joUtqCSjILqaGtxKkG+tTYMsKefHvXOfLx7tY4eX
ccqNRxfetabhqXckoolaKPun1/Wl/9vYwKaFntFvXJCXXYAV8gmk3lBC6VlQkrJWvQ0VwV+xWy14
9NAUz49CjoGYohIXq28FM6vwrp2HM0Dp3Shcn2iVtu6yAhm83ddpqSz8jsOhvqe+ot4gOtEXNx9C
27vATFTLV1+JFbOD3D2ctcZHWjzB7Sql4ZdB41vlyRQKvSPQHxFS0uBfPvsahBGaXwIDgshPsklk
TPhgU0eQjqAA4cb8txVutJYC1iNHIA9CUP8dl2Ye2rxQSf1UH6bjESO1qNBOXF59p1dPLQHN08Wk
AvDWG/yOF5WcQXVK2DLW+kJCqivBKYLTkdXxQFglaKEVlOR2K88Gq+QVZcthu+saLz6bhaJ9BTVl
11QjApYPk8hhnRCpbc/8hlBvnxcDJRvlnFwXxV9ZQSEcMTxYkn9sGyALy+ShTZHzA1e7XwBnpPU2
m6CNTlWETcDDZ/Vr2mIQyQDu7Lbsqsm6yxGW4sgdRw/EnaIZj7UxHDtHxU3k3K3e2IzAbfIATCmS
qqA3vKHyUBdc9xyAttC/R8lzvAbJrXel89iyQAxZslnGtUYxaM3QgJkQPsOJjzaFWDf8a8v1Qmk4
6JhdFLd2uQTwbhsjA7ZXRt45s1wdzrN6dSB4PKPGZLegwlJaMhZd0rT0U1eF2WnuQqk8Wi3Ffe+O
g+mfRzpyvg+U4tBBuXtWBVwCZ3qheQSpI7jUCbQBCdFtucMh7QgSKS8UX++STKhpD5JlTSTDemiz
Euxu722rD3+4v411HCeXj3HfUnp9jHC6lcBDNk0ud8DuYcp63JPAyf96/H/i7KL+bx8OfKLUO/xZ
z4SN8J8U9qFaue8vi/CeSaoARvzClPaOm8+4tBU/SKySGZBsb00ZBL+c7/mCusuKW+SGV0dmMaO0
KfCCWXCK1dBPMfwKRUXV26Hv65J0+aQVs5qoxdb3Zq6zZNc1V+VTfjkGyqQ4SQYi1ZZF0IIbDwAn
traDqVik3Z0a5NVT58/YTY1ghyjOYYls0oBqADRQo+i3UZtOD0EA2blbKFmt578hEecc2MdUvhE7
IdVSEJbMzQCYGZFOF2skQ+SMeK/X+YsDE17fMQrnpmwNlZr3+HPImHHlNohhdBJJsdzh6I9SY0/O
u+ui5ae9y9sXDoO8e3rXWtiGHUqqHTsG/AV2JG5B7thBoQqzOuu2t1TK3Anqk9ijWiVRN2M0GJSX
9t0zudzEwdhsrl+N9cNy+7eNragzHTIqYmVkl99vOgHzO9hKJtORPq6ObwmDQ5/gTnml7r0Iu/kk
6/kEkOsVfCP02gXsnHr+dNbnUnmoU+RamOpDKhUbhZR8+i3HsCIG/ktyGm27KrOip9vR5vzrJLzt
LRp/Wgcr03ahUsTc+srukf2qn2qN6H+tvDeScTjGpbchHIuQJKBaRvnpaWvcY1rbnGwwi6Dj0pY1
SjcRLwhooBYeRu8pycM4diDt+/w74SynLmoBCTmhdIF61XiCamluwJ7OwhJCI+xuGPvfDmpBRm0q
M5Vrx+hfb6MHicIaTdlMbXbINrxrmBgZxm0KWLWavT2j7yfawm5eM0nAKWqxZfQsQ1F2OYYjczJT
faQgpwMSat3m4lMPBVzuzlJFO7V1R1qegbCfKRgDeo0Y7j+xQDHSWLPC2cE0lsbnPEbjuPkWVFOj
dtc61RTbUXzKfEcE/4EAjUbHmeUstC5GZolPf00/odPwyx64//COB9cYzybbIAfbMh3AUkmc3OYD
YyHOHYkbbBUgmKjRy6zP6/TJgYNIOHQuyLxThnU4Q0zdwPsZPSHFy1dx4LW4PUTazYVk40lgnaRR
7+Md+Fftfxiyyan4FyKCJ8z+dj5bUJgZHLFBdYcsWjmRnKczMw50qzYkyi7mwVaTty8oSUc2Rawq
axTtIRKcHODXEnJeJcPn4QIpdxz9XwPLTT/mbPxfNEYwjAI2vUw98WBmLKXWnbufANChBtIuD04D
2KRWj+nQvSIPFUlQXsMMJyFAGLdfmLTHFNsB/8JfFNS+8fz/MtnjqNowiLGhetNH7V9HDoE3geSE
YSQfK+/ZOy8fayY1zuXV5Rg7Bww3HKPr6H1mA+cRgIa6KVqKorGZxn2n/xRpiq454gAlW59tu6Zi
9nUlOP/JowYs7JkF0T19cw/qNORr7prYPdFSh5KcUO/G3zEcT9Z9Z9V5eDPDqXBlh2ZNzHPRjZtn
Dy9VkoXPl7P1/EFobhE2JngIWSKITWtjVqf/8bjWQkaLwx1Zn5B3rTbAwg3nF/YukpUps/+BLLAl
/iLaB4dUZ3SFmrVDa+HmIWNpreyMYFYRB5PuVgWkoIrcdcKXk6FnSIomiCvqncMRFRuNMWYLXf9v
Hi07GtGQbVl+47FcwWlnWV+qg8/gglKm+2hYCMBp2bhP+YorWeQdDy7rLerEs4L8NMkHRnqr3SQh
RcAXCOmAjSHIZA7VwUHMRNLQ+gIS4d1MD5RQ+Z0U60hgKLry+/QkYziBAnllBAX7Y5MVY3kPZOyJ
/Uz8CVDrYJGSBkNqs+L3xTXLv8iFpRtU8BKZGTIynqoTGS9+5THBdCszSSwPYKqAAN0r1aSVS5vI
EX0QIy1qYel7VUf4MVRgbExRbF/HE5nIR9q0WPsEKGZgJmeyrAouOsznhhMBx64V/LWAVBZur4rx
/XvqG7g4VwbR8jtTNTqagx34ztxx3Tcg7jvIiwadyvHENZjrThn1tCWfycvVR0dPaCkAhUJKwjoO
UfV7aASQ+AGXBJ2u1Id441E4av3eb1TBswVOHVqoHCSDbQ2T/BLp1BTAUGhPifPoeg9AL8bMTuPq
ajwIm4KhgfzD/Kou8DUUH/7i6ZZc8ZnYa41Dnx+8Y0GG+nlEvYO/FObRWSiZW4lVQ1ijUgI6oahG
2hMWTF/L0aebKiU17Hm/fYaLTffxAv19HXHw4FjXgSXZbecZ01oeYIjFHEkItBMlF7BDxkY+cYF/
6i5WKDJ/Eoa4rVulsgmscPzk2/QDRu3S5PbIZanZSuQS/s0mCn+vwpPXGvnrqTrn2mSSudwkDYG/
M5KBQULAv3h3kuFLt6QL72zujlux0jgszzI9yDPmVIqamCU2qadRR2hM8AX76vcff3m9AE4IKCqI
MlPOMacFqobiRk96MNAXXgXkciVvmNLmvJfeAeTmmNVRDrtyPpABLGHvtonm38wO31EE2sI6qBtI
4jeIytKb3paZ447ZJ50y/9aSYJPOO6Nv+MQdP3Kb/w3bFcBMRtHPsjsYWLenj+ztqBEMrAusMKl6
2sM629E3Jz4cUvjXtYxPve6O4M057MdydbbaCbMrfMfK1MHOXLtQc7p7Q51tQf3AErGtduSh8r18
fpNCb1X6VtyVOhI2Hw79RECSy8u9aEpAK8lR1rLpUjfOFrI5A5Oa8TAvLQ9O2EvI0KW/P2I0AWir
Dpt3ffaY1fbP7ddrwseMDr7IgVivLnvXq7FkiRjAIhNjb3EcMMkZQ1swLJrc0LtL6NDlsAerCqut
eeVDvHq/5yqA6mIupc02NlI2m+t0gkvkGTH+uX4wuQWqantIcQ+xHI9skPr1gRTiWx6/l/PVc9h7
N5vj/3Gl3RH+3l3lPw6BSnE3IbrCLItlIy1q4gaUeTe5Claqdddw1odT9PHRoukm5s45jL8BDXrc
l2A1EhRTLdQ2IuDuwCbVcY9XW2ki7ryifCPJEZNSlLuTGyumGC0y7nVOICYAFrJrhp8R8qob+GxG
sqER2TCrUHU2flhokz5vw+Vv9ihWI1LH5GmiHtFIjpp+d9Za4+eAWyUV7NUy4RNEMVSavz2RLMfg
OPevuJB3kimP7G/vBJsu/rJe2aNb9UedbfsPLaPBbe3GgxKwAE5Pr4crT2bXsQd5MfvRBpC/+lsX
9RPfxhdndY41SNAmC4C4hkojri+nO+pB0UvwZqYM1tlkuOlxEwVaSY5ftpz4V44/YQCY4CIl7XRL
okBPZZvDH4BgTdTtk+m+yTk2X/5coqATLJB9IjBTVhlvENSiHyJR9EiceYi5mH+0ZeKBVNZFt+JO
ApNDolf7gntwmbUuOs5+exW3Qt8/8C6TMjabugRcBUX3q+0+MZRK7+74KirA7vFWTtiJVFDFlQ7X
F1lLkwP2x/5MLPzXw2l3gaIe1NeIQha9oIUm8Y+PNk/4cQgNR9CFQxf3hsV5XKYvLTa/0oKULc8q
dz3SFOgwNPO/Ob00Gf4XstgX7P8j4qCZ7hk2sRIYZo0y8wgpu/9WKq4PPgXacs5aJ8SW2315sgax
KOI4jpNzPJ9M4/rCVL0WOLDIOor7OVwSpTcKJpKwSeEsvWrw3qj1pO0XJhn96Z17CqJkqqBdNAJW
ExgXlQYmBm5AVtau1GmR1pGlPOZf8VnjbPhXKRygY/CEeoafQfuq3qaCYtwUp3WaupasCMCDH1SL
LTO66l0eVIMkTzg/oGsaGli45O5EM4goZVsSwWqCsoQrOAJ3oyZoaLHEXSojOAqNkXCHzP5FNNkm
yUVSQTBb/7x3SOt8AW/FQ/0r35Vx8kSY7lfQFoe+DCZ9Lcyed2Li2ZzJOb2e2w6ZFRt0OQeFqrS5
H7EMQBjc/wRojNqmL94zWX5Z1xslWdecSOGvUN+1KJRKNShwaIzsw35xHpxMmf/Wf4kczt4J00e9
QLjl6Dg0XyJqXTO2qSg6L+lXNSHRmuRNiLujc1EPTPHoTB68wEZ0+8I6mt9CXlMI7H5dWU6Roeno
s7HMpYO5bZnhWyG3JCqE/jbRgBP1Z0/lb2uBjyJSk1zzC+0hEhPlmAc47x8cx7BTe+nafhvm9PMm
PzDTGQVjOxLsDK/9nbY99+lVjyP7mzCt63YI0aRBYeoP67wfcD0ls5Jor59g42qdrrUIayB+LPwV
dUnQKX8HxgsFI/srrY5MpeR4Dil2ZxF4rnlztutkdSHX55ah0M+F/YM+nC1tPAsLBrX5zBDsWK1G
UMfoRQBWYyh1ejWXVWuMoycnq80/4LVHI9nIIFsDj6NcXsFzckxZ7zTN8parsJS3cnna8E17OTpN
/G8jUjwcOxQMBVuJqmeeIkPYHVJFHv3Ev0jZ5OA/bIgacBk4d5BUXdzp+UcAilpqw4eLSXo53/bm
xSuRr8vE3ve0bZYFZrGA2blXU5wdXHXatolLQsz9D6lw3I2akxfYZRyJ4X9Wdvq32U88nUVx6MON
Yf+syS+UX/it4Rj8qPaZeD2rhi4yPeHxO0cN6ms20qY1fGE+xQF5Wux1LNXBCkhYGPDTZWKpfzhl
jVvqdhqHIpgTvieNVD+eA9GbgaA0xsvHWZTsf300P6lWkKPNdJPxPDSDFzSuBnkyv1lbdpbo3iG+
QiBoEXtWJdprrAGJ3Qx0CcIeE8zWFl1UVF7rbsNCvbW6ByFXKQcF1APVrMdkGCDaoQHTbCcQW7is
PUd8ufRg6uLziI4E61B98A5p+At0WNB6CFpOh9yYYsm2fDalX7gRZnRrYFhZTvpNsZJR3Xubq1wF
uJoOOEifJ2XIQLcodXkZwWl/D9+hteSTlhqJxV/lplIrT8QycDpIJ4iITfXV9oU5METoZcZdaHeX
2fwgSg0jh0y+CJGcRjcVx0oMVG7TWXOPLm17w5PSgmpc/AH/3L2kOaVv72C1Th7armC4Y937EGvr
LeRrwzCkYUyppMlLwoRea35oaT6qHf6OKRSB3y18Zquiec51mQqFcIeRQCAnDjLAtjfbwSqPBfaf
WGlT2SmvMlQ/tklPX1ZK6vHhQsoo9c5r39i3IAQ1gx9UO3ucBt+R1XrMKVtUfPz0XBNX4h5ZSgw9
mEoNLSIIYtCTu0JvKI+cRKufSLek5RlzBRgC3pnwhcimwogwccI49vlJYq3vfjzh0fJXcYR9IgFd
e+OYyjw3/aZ5bBpBTm3Lvh9e5r9sk934H2p4XpBQuGTm7cOKUuj0bfP8J9hkhNIS/EPw3YyRU9XE
VDwaU2ZBoR/VwZ3oq07afGU44RWjAFbM4mkjBR5Eir04+Kf5eSQM4/2P92pWvX6IQJNwMC+z6VF/
6pNeVDnSsuMfC1Gs9m2FJpDZlk9FsBgDoBj8L17IwR15RiTvZd/+fOjFgLwzTs27iXqV0ExjF1A7
R8ehnUoZFybfgJGykhj3+e5tH6MbEiGOHHmGovUTx7kvvWq+xImVtyVrp8hfzsoqM7IE3Be/xyW+
ljlZne4rdfccAbNMRV3JjdDMGwHP9CKvg7XQcxaSEvNJg4GlrX4rZZSg7eHTukkYcMxlTOvt29vZ
Emn36uWFPo7LN0vxuj0P51HAQdzYTBB3ZAhEmhihhM3KvSlNUivZyX/lNJDB+uQq3RDNJmdltO/I
BKFnwOYOA6H4hfitOid7T2CyhUE+Q1e863rBUDtVF/u0OGlwC0NGkDiW2dPX+pwMFJB/VX6wf1Rh
WKxTVL7fLD67H+jM+5y38rGbPaq1wOjOIDcN+ZgJV4cTNnyH0T1hdJpWWr2vCS3Dv5ktEate8lyX
FteUYf0qdeS4szwF06XbuwgwzU/GuggDGFfdsW9Ck7xg88DSv0rEdnZeUka5DWL/ti9W5Qw4CkH1
ERDruUTPNtoFZDO78dU4cz/aZxNNlBD/zB4FMYMRPh/Hcag+0EZJ7O6dWbi6cNE0wIDRpUzT+B+0
aN33Kd3XFs8sM5GKQM91apNtYnp5moZBB4h8St5PYz2nUvwsQRvPHBYMwEvoO5tzs85Lp4TqjAP/
S+W5MmV1420gBCovvroXgwONIjKqgCrAcf+OarBwxJG1oGkZzkrr1KFWjPOJYOvC08k4DDZuv6BK
O3O+xw/8kMurkxgRc93TgxRvl+3zosI4U0etAvZbudiwaV4wr/VWgJCxmIJgBxHsxfGeo8e9khnw
HLYbJvGRWsDkFXqf+00tR3E8GT1X/m3oCncEgzbHenp6jo8LTWseB5OPa8c1Ct1yLgwGigpDnnOr
gtI/VVAB9tlNeW568Ilz8Ppvqt/DDfS/XOSppfE8x1RfhLQKq3slcqY1IEd8Y/TnZmraTUh7IfXN
4LNl8JmTWWpx+YNSxB2De4GInfTkPyVkNdmPlIYCqbWiSbXBuaL+iB6lLk6xKcHBzdU9fAvTdW32
+ZYdStnvtLkRDua3iibosw/57rlSbEnAkZZF3yuj3Qjt3UnrLc/0KADDsl9i0tsK3WI8egZvTAKK
eRz4dmpcZNlxZM0uwRaPURy6195r/dFcziuuVI3+zBpHw7e9C2hN3of6LqEmxXge3Xg/VR04ujtZ
QSLM3WD+OmTkh2xRL2opU+0CeWbDKztE88rybDGvM0OZXvK9E5iyir0EeLpQoCFkTq0JZfXDYeYS
3NhhmrcsmrDXWUTiO+BLDqb3rqfZz9DNascboIE3x/58WyLLusgegGQnxHrZzCqNBlh1fMBEmyaM
FFraklACmfPFFVkFvCZk89lXSvzomiyHWr5tTIz1nuoQDuyeYE35MJyAo8X0/d+62rU0l4BpTK/M
0TuqCpq0dqpexOS+Y/dlULyyhJC8SseWFnon5iqN7p9YF5+nxtXIJs9jn4cABn3UwVtlupJfLAYa
bo3bivy5oN8CGGrp9fg46dDbH8yRcoAd/Iz7duJlshUf9F28SVwByK6Ke8AMTDEe5ZrKPYjYei3J
QrrTdAOD9XbuzYw/ux8GH/M0DQE6UqonS7q284yDgERSbPTyd2pAxE1iOgdNryEFnynJTCqgj+wn
viME90jtDswGpm5Ou1yAp7nguUmbXthZUCiDocDZvjthpF9bRys55tEAnq+ergQb2HbA+egZhd0u
2yLAIFx4Kxs2nzPME9qm5WdzVV6A0zs8eFipbQW/OPpv6Gkk+PQ/+htwcPhIWWUFoktpwnoF7cUe
za5Gkgaka3aPVsSinjoGOfGcrHG8k5zlrV+0aVgD1U+ponTAdySnG0nCS3+kC40UmxdMbetZtQx/
kUU9DpuggYfxqEghFC18KInDHn2a3aHmR//7nOhcFQgHY/S1NS9IBct6F5PSmDValr4NQ1ffbmM3
1MZ+qsAjDSE0QQpeRrJQRu3mKDzh7reLOswsCdFcZ4rkXSGfcHIGXkaYbGtv+qafNWlyrUbV+cUv
vLIdHl3IgloRLRWzrvA0cENUsHlwNqP9ZLwh1NeJzv3BF/4EMEL04NrPD5FtDQfCcC1JEAihzsse
98UPq07Oj4EMIMENPZd0n9sdU5yitNU4GGR3KghA9xP5PPii3b2qLf7P5s9DOYnPNeWcJ2TB5sxF
Ahf60jEg2TqB6Y6Am92Pw5NLscDirrlWPWbq8U+kA9Au0I0xSmPtBNxsv6Y2HYu/RZbfJkws1PaT
fF++ywMSe0jTJVgSIs05OCbMo5uUjmyOFmJ6/2BGvFjZ+uL+n+r7Kngp3yh4yBGcP6oTJ1s99m9A
V8VYBzYJSt1lgTURvvTZF4zupFZdprbPaxWuw0jqf8frMfqZ4QTtotCNQRLQmXaN2UoZ03TMv/Aj
CbbzosXSI7DsHrhpYGoI1xQv5sDHBt/4DQZzDoBcsrNciTi0vf6nnMMNGXzgoJNMBvRpdveCLqa9
H9BIcYOSiHJCtB982PhOc5q3udxYLuB7QFhhV8h+fFMaXCcWYL4hnasoHBoo1sz2bmGTXstZdqjP
bMMXlRyMJw9cMouXUDB+8e63GacjZTyryVwbjtSAzKfwl2LEF8y7yxUivwatxZNUYcinOAcmMAaO
MKH7dVVzMo6D9wTC3Sj5rIN1Ccn+pOkBORvldD6OZD8LVQ6TwVbQZzgqI1oZwNZPfIl3H6tEL7z7
sSiqhFRNkWHzgo2uOMh8QYJVxU1a8N3oYv28E2ueNFH3taU2m9/uhV8rFMEEJp7M+sum6Jn4bd8V
CO8LvHR5lTYIG4WsczZZ07sq90gIcZf+I5j0YscuWxtV1YKbw7e63fBG/8bd5gYuUwRnFszHjkhj
+gX43GYuX1zSlhaBQBG7ZjekcHOvCzV1YwV+tAoJX3c+tIhPj5bA91KZVJPXQXgc2Ml83QZutvo6
Af8cXoI3N0v+QjqV8pI2nWApSrW/O7TFoMGkBbekZb3Z+XQyOffu+mrth6W89ZXGuP3Orff6mdwM
L76RJqdBOXvPQ/wsiUqdXVilr5doIZq1jH6756THj3tFjHfMiM4Qnao+OSbriSTPvcSM+S7zOGJw
Tz+qt9xadlpZcXyn/uj2g8lmF8NBftFTpHneqBV7/UP4GhneY2iODdR49TEEWR76sX/+QPOVXInX
RV526T3YsXUgGjyDrhwDbS8rdieI7PS9D52OvyD4iXlrqMK82B4ibSuA6QmnN5+naHWW6yktLO7n
a8Iv9kLtdFmQDNSYu0tRs1yhSIv95M2YzCt+0a4QL0l8B9wT43QBdlfH/NwXg9+nz1lHFhiNa+U/
+TlZ+fGs9uhx7GJL0GIVRaeiNq4+wwTJcLCX/L1bwLnsAL3o/uJJ4dGZdo3g+PThIqL4kS973BRS
A0bmryNjNBgX7TDm53nTzfjj7n0u+23uLG5pjvz+MkRT3NyMyqxOaHu9L42sgn9YNEQ17Jujj3HF
e/PmZD462XEmpFWE0zHW8ZqLWUHVaJUg7aQTdaioRyxvJxHbAB5ww0OF5P2/LtsW8A8MQCN+vxoS
xIBOf79aLowE+gll7fULjDnwUYQ1j7sww5f5m+k+qThNXn9wt7ya73QvQGlAacKciQkpEfbgkuAt
J1sBeFWRMG20TdyW/JJ1anoUu8XivlkExM7+5rAiyiDEAbG4WCSlxcglWxgLYlEHAInStFJ/2Wul
vyd8QXN7A9OLVmomeM8xBMyNLVXgB4eDFBq7q5v/+BWWRXaTJhvqfI4IcZusIZFCzecZpRy4AkoA
ayI4NoG12IeFY6MNQYPw5MN/hFFQ9tlo+FB6H21FL0MkqHfciITSLdHhbsSSHRvNYuTANquhzRI7
cjc47bgByOjEwtGw//pn8pKLmnLIZda3LdPKvxF4m77nEY1liNoAEvH99gyWvauIDd2pOd3xj2Us
MwppcVVdy4tDl6/18/hWCsX0oRTVnOomd1SkxJrTIctWqR8iatlMYzt8Nbi3TE0pt0AoPnLaNpZ5
tn6tEF1gfJcvRQYXQ0vMSkemg/y+Of2x6lpl4ZbfawYI4AEeN3XJIBfdPApAHBSBk6noQeoj9gJK
WBK4XMEt9Rp3zWt8u+nwn6CL2ekpp2WHsGrtlpej41GNaywvb60dkjXyET6ydINg1/3thXM0zOel
Gyjpo/UcBIWX3aEdnSWX0/ScjXAfxjhTlaYTHx++ehWlGz/yQRQDUHGb13lFU54KeiN9UjKDsFyW
OqW1xyFv9AYdZd/japnES0ZSlbegnnA8PTiVNWA7f8PFG4++RHJ1Pxt1w16Gq91q/OsE1FO0/gRB
om6OIITDhfaCCZUzVhlx91AioUu5uk0vvd5e8rmbSOqj7aiV0JN53p4Hd5gNTJTWN1rW/GMnlNWi
LvTq2MDoNn4kE54oChbzYbeTOXZ1MC9Ma5OhK0FvaMsB6W637pZUCWNRthYJgoGFI7/o/iW6qMWG
hjMSt1yBRxP+Iv7j8Zdoe3EIBTqrsmzeP+LLDtlRkwVji+9ou8FUSLy6lNjw/q/J4pspIdofC8e3
NGuISJ3p4NKiCsnjaa9aKLxUGZMvmGvYjQ7CJu5gubuC3lD8x+29ZW78guLdGtxUBYQdKta/IFwd
vCeFgR9HZQAjMOVMVXM4ZRFIB0YqfIDGCTouphvwbnMhB5lGL7GeM5L7qJ/6HTmI05JGZoZwVnyq
Xsst33kRTnXKZnqGz59VqFU4IRY471L2W8pxj1Vc6CLV+J98egBiHPAauds9Yj7FwRdcx4L8l1SR
Ii8KSatkMjxLQBV5x7plve/+vn9p0mTGyqazi4ZuIan8/CErAl3DhLq5U/FolXgOYYIXJr8iXtkU
M2x0ZnepvM88VDS9YKBzgDwMwGKSzSfnUUnLo1DJojQjd6KQX3r68G2O0yOTalIh+hBwt90mETvP
OGJhV7NIWgjKAlytr+vLizRFG/jDEoqoe8GCPVVb/2z02MD2rBIHX/jgH5RmQfFcKrzIbC07cw2b
HbnqnDIoMe0bLsvOeNHRxZ/yIIApQiAzQjTxc5ZpXcm8cKS2vzPLpruuOS10LJvr8z9juYQYm+YZ
w9w62ObLtAo/a0jv83FLd2PD1BkuHAoq9HUudRnmlcrLe0YMHEoIV4sQ6fQ8wDQsWZUee3RHQn3c
VTyFu18XuAGC4nGzd0msNYGmlmTar1/FQDl70OHsbL7ohwMIBMY6h/XOSuHbqigXZeMi7B3WvtcX
rzMgnHseG38chm87ew1zX80E+cuAYXmXakjAp904pN7LOt56FXtF5OGsmj5StBAlwAsQR+dhibWq
cr2VRSNlLZauYPsZWDR2oTSKl4t1iX2UgoiE4P/bty6PiX5GFqeMlCNR1CJY+GiQGqsXM4pmlowU
0Qz4FCHsho851O6NIu/wAJz3lA+un919XgKz4rREXvkAnnbxMqSdOnLbMjpey1t3MEmu8f242+TO
xG7pNDs30iOj8hcM6lWK+gA3YxT/Dc7QKf8540GznjT9AC+9cD7vAmjsQOva4ccVHG737lEySIec
utsfmnzD7vTfXNp6SiZjD9BoyEh7AGIzsS8xuLg/l5+VuecWJctEjHv46P24LdjAVDYTMLE1SwmH
gCE1bj+QLrm9aKQnVkb1iukgnmLAYDlRnpRloPOTK4kvwYMdInKSs/mjDZF46tnmS4Ak5PgqgAKd
okKeR6WvCINyNKqjHiUGeVdGJfWsMQOeRo5VynhqiLBj1tqrNiK9i0fuI4Kd7DquW/xv2vca1+cf
GNQstw2zRHA6UkC4TG5oX9iKdYIJiXj6moGcFUlvetcz4vDkyslNV5NwHU7N3RGeevaXqriohBD1
CeQtAH0uwXKYHxCIvQs/Ry5ZL/YQ7ZqAwEIqd7SWjaXg+b6AjYoh8w0PTeXMiaB+o9IuIL4PQkN6
AJgzxyjh+l9fzoceNkFHlYM9MeVPTvp4Vyen73p30Js5ssDQLFcqTfTRIQ29m9ZzLgEqPMkk081A
1shAnAezhxkJh41jwOV21+IPLHD+aHMUQRt8hm3wQXhE43tfpEkEWyMadaHmZDA0ZDPoEJI/EOHE
TkOwzqD5tpVEvg/8Anhzr79ztbwiwz4tnn2OVTy0p5NlAHKkGx+3oBhyg5KBQ/hmcnBp9TBtBpND
elEHuXK4lBaFCcUqx77Sk3ToQ/z0I/OyLpO5zGWJykJqIPc/t2BijrKCtIPw/En0z7ylrzhfLCxT
P/JYWrswNY9bKx/a29jLrhHoxhrES2LxNXIxgLUlxgOWP97Cp+ECLhVSb1k0ek+lDctj2gLObFrc
KMz9QVVQpl0AFeMIPUEs9HKeIuD4llfa9Dc1z/uUQZK83a579Y4yXXhIodXpkKdI5C32HEK5zvLK
vpSOryDkutnIU+ULqG29DdzAncBSixQvAafD1K9daUpPCZoacHCo4OGSCTQnUsWiWjt4YvIzWXCf
z7eB+fhv/XiBtSgUTr05C3Hkpk+xhVJoebnOq+LxGdBXWFswIJPuCBIaVnuNcZiQCwKrNQsWdbdO
l+lA0qItXvgMtxoa986rbcZ4CD37LUTUZpg07Mk6+SSG+UmdGys1KLPBFNYxgaw1I2Xb9kyHv52Q
hPEMBGAPrXkw67SI5Hgrnrv65rJ1ZMAgIDTXlyraGhpPGXLvYm0mLPq2R7UElnlLuPcFxGclx3Ed
Ko+2ip+82iHymaAfq0HoCjoy6CtlIfyfgji2prn4SS7IH9+dmdsFRWGVp+JCNuT7Ugs4s4SQ0SwJ
k33UzSMDzLF2sj+tcGRquHlCPw00+5itQWJAoMBEBsyHqdc2Lr5KtYYg/GLuCj3xGkX48009M0DX
/RvPeO0CMvVzef+o2C311sEFqqCTen1m5IeAMFAxZXKpD881WhIJo+tEhB5FT/EB1Z2o1eTvFUkp
95kEZgVku39KFYuM4FhYA5FCF+V1aZ2xpsbQLpu/CPm9NpUdeYZG7CyiXAWzVhnwN2z7fN8dJnds
3eyXYnBJbO7QkRDOp1BTID3FDAKofzTxTKzmsZHFzJadKFN849Xogi9UuETvQXRxysRrYBsXGgOy
45zJsoxsUHR5v5v0Rqu7FlCUfr0bv5IkmbQFuQ58enTvWVhsRb2hlRkga48iXU3NAzD/j/7m6N75
9DxNf9g/gLMlDnWqw7PC76YQamcjrhqgTJmY3+tnEXqB44cWBb7fazEvjiFJ3EeP8y6CAvRva6IE
XcjWuiBJWqhOjSVUTR39J4YWFD7SBtlqO95bDiBodLvmSGftAiuhqDzVGursxKtpXp+yFMXixCzH
WByBLxaN1yljSmcp1PzMMbWfiyFaX3ku4rvzfWN//zCwC2TxC13uU4OvM1bCHMluZaNlqvQ+ffTA
LpYlVXs8naIsptzwh0E3Y86VqBtcBJumPEmi0qS5d0ZSxxfJcEzZDu8TUzQN4arL/Xhs/4P2RVhB
CPgXq7hbFfFwynchJaNKCaW7onshV1gcP9Iqaowc0LgZ1T8usF+Qh+v55xag18gj6om/+fQTUPu3
LNRiFFkDDTrSsjaHCmTYstfrnbantuATJwSGBr/JeiUnXjMP6150yJI1/SxlnD10oWvQ+LQ14+/H
JHil1Dw+JfLeIz2k5vHf8UTArxHG+PnYGAgwzhisss/S5TsEXTf6Dmo308Prt5lKS9Mgp6q70RaK
M9Byx0h2gFv1R2jAjqrz6iw8DQXWyK/+NuRd9T8Z5Fb+WxpTn1QWHzD+XB+uniAVzbrNM7GSyrz7
xTrkkz52IRewIM0OXAOuMzjcwQi3kGDggHO/MPyKWlXgWFro+iCpd/6rIfxTn0s+S/Rs6IQgIJNn
855UT78Q5LRwjRxhS6EnblDkr7YCcN8764+pAHogIrZ8HMKBVmnYPfbVfpgnzqGTjnp+zXdicKFZ
/2/VwWkSd7jCYu8Ca3ljyKZJ0huGtWq7YNQQ+pNCc1uhcnEXLZ0CQyfVindmlwoOmulpx5eAyw8P
entfhh1aXq4pf3buPF4za4gWSw9fXUihTA7MfJdplVi6pbBRlLPM0yMtnAYlLSI/j3gf+f/kXo6a
hUfNA/HfAz9lAUgII8ahWedy2eLyk5wcHcVxhLr5zwhZpzhfhrc0L0A2KUIKoT9BNrJQZ3UZ1BDP
OjNS6oshSIjWqsjcLf7cSlj2RVAJPapegVGtfVXz+Noj6FgSMj5CZzeyiKMa83ynoqMkK5k8Qpq0
/EBqr3mVMyPIPt3VpdgWTb3zMTjNfxI88/8ix691jazC9iUlIEUv/CKU4nKxc0KDcDcJSSMizjLt
63CxwSgj4ymmtWyR2g52TdzPccEjPK7o+QmfA6g5mzKabl/7KOPR9/qzFQL8aytWXCBiUY+nOxDR
zgWlrYwbdX3hUZ6l7sD5scLqIbgBmJ1L5oK3/CHv2WJvNn+62sJJuaZ7cvQLa1f6fvb9oTW5to7I
X4ZZx5HVqzrK0WMYtNEY2j1f+pePhgnfvE/QLmwDIfvAnLSqn30ppMAZP+7d5v4GloacLJxXhPHX
qRHsab60kphBGTdGJL3QMeuFSOSDnGKVhKPhsWUs37X/YFJ8tL5xmXKr+wXQ3wK8q3D4Yu8OAy6w
07E8AN82QUpdRluu0quPayH6GBLve+Fzqk3tzIa96G5YtpRWnwIg7NPnrGilaoz4Fwa2EgWvrm3d
pAYjXNQbBmQeKH+NTIf9dncLHoMrzA753mS/jvgV0ExFjBpvEg3lx3ruepk4wLx4WldS4mQkjECK
Z9evzLnQvLlhwOegvOsMXaTg3tjWk6ac86R4ReH9hYtOEHfWJuQujHvqROKzk0M3Ce/wyciXJhY2
B/PK/CYQKxEcMiNQ5G22Y7T7VzR2On8zb2j9188NO3ndeTwqXzahZ3fFVUBHvBQfdp9TKz8yyoum
CUXO4ludapowzRpxvxTRCON7VsjZRUIPU2dHv3wjuLTU7TgA6obFJjWL6vmMdKa8UeFxbbK9irkS
09IA9wc8u4CWIs01FL/bUCtTsh+OIkf/+C2FNnVnpeOusS+vLkW2JAivu+W6irmggM4cAM1iaLJt
p9ECRgN+1wUly7aTvmzGbp3b4VOggcyJfsDa1OwJfcPDPHrOLf0pryCvrPFBeVxEh768Mywl5SqY
/X98qfIRu/3EZIwHO8I5bgmRa81KBpW9QOs2tvSY+d+bwDedYMvoqfPcU0FWE0MIu/Hr8ds7dcuC
9xRCoMuiV2nCMialMHDL1xXVaSijrllhrXIxRwsP4Gv2Bb2L7L9YipdYp39KO0yzWpiY8It9tGvp
8UOf+R57BlDIVVtJZLG2XEI7a3Nt9BKffZNUXtNgvHN/TGRVBZRCGdhnV+rLS7rwOZVk3lh3Hx8N
GTrguvS/VesMxyv0ZHA4Sdj5V4Uwe8C5UGk4F5WGcvAzRRExmHsni+bSHivrX1u7PdSUCwf6okUt
VLn5JZmNzKvRzzYI8/YKAT0GyTy0wNCkW3SZvkgOJ6RvaQRILg1fPGU+1m6C6OPY7TlXNgirIBtG
WjcZ86QvTm9zZ97eKUikX8a8xwdgYn8uYTFmTy/RgUjrPkCCHApDJwbPkPoUReXRku6kXgRMXXS8
FCg0GZ+kTEy9APoDAkYvd+a189VQ072gvJ2c9irajMQSO1S/d7ghF/2Iy/2s0tSrYn/vCniqbDSI
fKLgFQaDXeZ3sZ4j3Z4kbhlL0ge3EepDrk7jPoVWFL9LQ830V4Gttv68QZv5JoEbJh3nkM6R1G0a
8y+8BKNEPIxy8XV6vnphjuAR7o88OidxYdw0KDylefu74cfbbEg7h2ggzhOyXk7bAfL9f76Hh9iY
dB/5dv0l0SAmGa7LXIFBccfJ43PeImp+R7mE1KHAIBmhDcJTjvNYY/CIXfy5ZgV/wZuLomp7ljzF
+yf4wPxyWCDQRm0/yZl9rUV28k/6/tBEJxuMAS+qIJgQjg/ki8ZMNRo2rCeK6EGkOmgpphlt+ouY
+NZopvKBycb7sGJFeFSZKsYRGxsQttBke01xncIXGXzWyCqy2uDHrTqWmUbX7rSf86WJhOcrrlQa
gFk5bFEbpfTh4HtuvXkml6enMfuLVvPUi9I/9MOYDII2fcIpJTUlgdg7errxR4gq/43I15nsfqhg
WElt+5clSroz2fc/MVSam58+cKTnYs4dNhFyWyTIapKdLhl6SkFz1GeRoMIsQ/vJH4UGiND4TI7n
SVbxTwrkVrQSdcouQe21cop7/RH+4UJ/+27wsB8MVdQI4UFYUm/rC71ABnGZoBFcn5c2aW8sy8Qg
32P2KwH6fubldODefYQ6CikvFmBMHnHPL4BnmhgC36x3HYiL3IgbawXoXXnKKSgksBOAZzwgS6lo
qurn2S25k6ZpH03g9evkIaStBVe7GlqBmyRem8yoTxLzevtwFLnlhTSJlvF5Un1pEE5CfB0xnpA9
KkAJSnJjo5v3cCtEZUIoSLMPeI4O2nMFehHB+jRZ0yX5tTAK+KSrL28PHZ1kH6Wbcv4OJexvcQaX
JsCM08NvItm3X9jxjSPI1K4i8LVgt5hy/drYKGFrFr0DLz/5i+h5rF6rV315lEQ/sfJtgXO9Zcoz
WbKut87TVJEnBl/yMX8qBN/4WDr2d1S1rmrwOaSfjlXY6/VnaeoVnsdLJQysmYdf+zAZFEDC36nY
bhlqfNuK7mA4gNNY2Cy58q/A7LByjwH5BUWwwu9yEM/QEsRAjl6Uu/gQySFMftmhWSzqTX/79i6M
rYc9xPPb9PCWQrbzLEMHmjaNcwGijFl/wH3Ir/GahzIrMhDF4YWCmTdMB/UXs9DNiHbLB6zwwbb6
QbrCzWzw4gKGQdi2ub4cOesHoogwWLKSa0D2y5UyVA9Qu96CctluqMX4HE40jpqPrhIUvINtKj9S
1W9CTCz/hO2teF9/u6eYWvrWKYznNn3JcEYMBwNU/cFm5IsvG8+/QL6NcLHyd6gFfEDLQbUi9o66
2ot0xgKKxurSgQLsCJjttfjOa5A7OMVZamEF2cN/QfZ3uhVIFU/q2MXrD9uk6Ne3i85tqTBT6/lN
+scCICt7MGTJNTdCmiBZ4aq/RgIVVx+q7MHAekAb8QVx4u0RiTbmBOIKwqpsB1zU15ATk49OG14a
/qfmSGdx7CVKFfD3xrp20tLMGVHviXKzTs2pqLAFA+NfcTOAgxQgxpoRMju9OmR+8gRB1mSPSF+3
2HHJ+z8Cd8ybKyWe4MyrTOOGYObi8HYs9Ja7xd5nDeWgq6H+RiYIgf60pYhLorbncyAydtO6Rssk
Kf6fPP6eeVODLwYOuS3LUiiKEMcrXqZMbscUve0jxsMpHW5Nq4TTllMPHkPtQfz4kinyF9lVjPPo
EkKmHZ8/8LFRMZ0kshCjyY9Pl9mEV/tvv+AxZtLPZ1igrETfn1UBUBWLF9p7PquZzRT8ALn9thyl
pEi5fkEvBodauNpzdM02YEAzIIkf++gTzxU80iZba3L9gZdsD/5aC1y/QxkLj8A+I45kRUeEoGBI
iIhGm7daKG3y++VAjta3ydqcPBnawxLLlJjW+j1ZshycnDuVkwVbQctUmvvNfknlcwt8F7zC7WvH
tGqpjQCbTubuhAikjIZSvq/vMhgYPj4ftoiQ0/sw89xVDPWQaS+t5D00BRxIgCOj1MXzfhJdVBeR
jAFH24vs5B22p9AtPOOkCEOgU2eklxAfh1GyFDLaI4CRDnQ17NXUJmtaBNZpLBhzMAWNLJBEcf8D
olCNlm1Ecj21cNH/AO7jKZpHwLhrOVt4f8EQP3SGLPyAigjMc0Ayjef98tR8cKaCSRJ0rFjTKrCi
xh7MejqmKs7R3bM9U+RoRqTmoZ+wVVp0fA9EzXCVI4e292IxyyuJFUVbu26OjzThDV76/Skf/OL4
bI05cz0iAHYvdB36cs1nL8Sdq/delLz0eyrrgxecuItIFR7Zk3fngPQ72U4MAd5lvqbOEd/xorUK
/ZcE8uRd1lxkJhTbmsjt+KZ6Dg4n5LWdhPDf6urFilvVO5m4RpVWs/yJnWCfHKStyiug7WUSkXm9
5+HmvvXTM3QeXITzdgAlZVIKlYz34axfXPZj6IgiwfDAnHLg2Uj9QZs6iFKLSLPA3rn/boAF9tLS
SwQc81IzS3oIRwVtUfdkricYaiCao4UGCBMliFh9bUB9FtGNEGHCL9u9jTCXkv7IwVdPH87xAOOX
vfqwEbFQ0ewyXasmLKenlpcVWy69l587NhCBJMsdU4EeOlFv1vBB4m8bLFQKbz5lQ0VUd77b0olY
QNvK/indi+z4R+nih4Vl0BKmMR2A3ecZjmbzMWmki4naNpvb9spI2Mglo2N3J/UPw3x2xxK7eJ6I
cIpYsoUus60MZxP8YGtw18jYtAxqjBqeaG9ILHQfKZOmgrtizTYReXkZj+hWu4q9waeOrPD2bgfD
2lkSyf/dFvKow0svIiwJCPBMQpPtwDoNUojoyzPhMS7ViaLJEckrllFuRpH43hTNRXwPxp+4UcVK
yAgYbsY+IcsyF1/aitY8iiex19ld4xxpoRYEpD3MGdtkylk4ai4br13DHjwPn3q2endKaSVy9UoH
bJpySvqE5fXa1ETYRFtsdZ3PtNVT3ZxSQyc0FKUxHPjNNFwjBN9WIBvbpRJACZpt01OCPE1bsiu4
gnkur5x5o8AKS2BZM9NTfvfHa+43VRQ63Wz91gnBbSJRTusmw1CIgNTEAaQOWePb482JdUJD++rW
ORoh5Mw+8vriuTtrfp/FxoEZKQmuq8moH+4XxGwOB8ZBBWu6+r5VCeVXa2xuHOVg0POtQnPkLL+v
UC//SrQiqknmrE77mbm8MRyeinzS62bKOhFpZ/Tko0KE5IJ+b2iUXuSH8Ob7at3eOwUECrDrrmaD
0odiUl+xeU2iCendoRStQ2qM03P7Xm1WoQtMRWl7mRLd7xPlOqVi3JOpmvXOJI62svAAWjt3H+RY
MohhfUjmdh1DTyrEwrwJ8WbAyykJEU77QjH5kUhnjw47K8gl/Nl8vmnNm6O7h8f7ENGkjRvmOGe4
OYBuAfoiWXFbORWpsbE0jME273jC/2Ae2lGKl/PkLEdSOSxY3uuno/jOFC9FLS5ag/3F8miEado3
fkhE1A6CmGh51M+fmKOtlTtESpYhpP/Q+wEgcvKXtXs/+h7PD7iN9i/SVQkn+M1xxjnQ5etsbqpS
QtsdHP7SXHUE/+7rIFElE4+YIkG0ojJAcBREWhjxpDLSDBg6r61t1MIQVOVccGtRqS3zjYgsHTof
NZQiRMOUqpdGuHNC4pLQAcRrWquI/TJ5gZdTQkZa6OZDmpDlUxVFr5hheBm0LBuu1XOsBJxQODfx
g2T7Gr+H1WuFkNQl56w2T+/Qm+CS5yPLsAhkhUI/m4O7651k22N95tfRACH5xu8AADWneLQzkqcd
cxHTDuKYagfh+wDzCed5RT2unIGS3D6TVI2BsRYsUOpYzOSNIZHCOqyEpbLwqAK/1RveR/DjQodb
dkjSpKeqhMTnmG+FlqojlBX09i1mWAhixLf+T8cnqlOPvD2TKUG+jk9L5ApR8nvY9IB7rx5HEqoS
57sDMc2JDceCFaDhhw/l/QLKL8Yjt87VAVWDR1VSGWLCRecMKu8WzsrrrMSjOvEK/EP0zadxWEGj
boJJiRWjnqZGFfdFpYUHKpS62PGakOmRrfzMsHfEQAoR36F2910XZn5t/vzMW/VLNJwm+g8L1W/H
P+0BVCvD26aJ4QqM/dk370gi19c4/4e35Y9S6+orepqIAHIprqpBcrhbbO3mEQXyyb+4YTQyq4RI
A1+qkyNS/UWLAHK814PWr5I+v9XMD40WtMKkEtTO37G++PWPCqzRzqWGCxlTROrvSCcpQqmJnKqJ
5b3W3PijHYEdvx8uF8WVgpJtLscCQGw9QuIW001ZcM4BPbIguTr7V10Z2ONECkr/M7mRt3ui9wDO
9VesVb7Shvmp34e6PLdv1uYfPasfJnn21hdOQRh/6tlad+Ud7L6xje2uay0JM+005Z8xgDng/nQ2
N4P66++EeS/89Ytr3GM1rAX2AGsVnfFTbyrC94MZIRbLBJHH+lPOiQcK0dXh63amixUinQXvhmaQ
qsxakBIwYaQoDbyGZw7a1nf3T5nM1wU8/E18QMNweYKToYTkJtZyt6VpR5Ya3D3fVjGL2G5qKkMw
7czXUqDSMjjG+ioJQ8+aC+2bZcJYVMNxOH00NHooYRG3dji+gmRM5FhmPVONQNgB0bda1bm91IMU
CDiWpWl595s1BlqYTZALRsGqTOUYfV82BcXgG3uRX08VOUDI4DRrgELIWpaRz8CvjcKu6usIE/0Y
qAKfbeTI5XZqpGMkHyRNXy8dwcuIYPolEYGfeH3CWmTOyouJmPXblXGrcKxr9PBCJ0K+af+pHnhp
b2fK6fWkTYdxCX4j0BDzmPOWvvRaQV4rWbNtzjl7PKzvLUfA+Uh/tO5Lr06rA6N6vuMBpQEvBEO3
829UGuzVHyWHH/XR6LUbqGjyN4RtRFRqWE1imGXS31H5p/c7BNo6bStpoIaotS5RBIh8RvuHI0QE
b8JuCPfAE/QzPSVdQDXQM2R7he1Pxjj068L4QI564kN0e9yqBONbHx59UEBtDgFy3lLr8slvqBOG
7/aoAFnJ2T/O0567QBtgVlCrLTu+WunaMCys2WglhkD5NtriS46IBjfVs1RUSavYRCMjG2bodKV6
89Ki8uDlYSMrSj7gGfIJEjFFQeFTu6X0dVlO7jzJJdN9O2uNVR8F3UTYbRJ3yTY+eZaXhAYe3lyP
Z0PxsAE52VIiAaHPQz2lq+EAUqi6aUZ/b711V15U4rA6AK+xtPi44rt6UM94B0wBDSf1DLWlpvPt
zP7s6e19S+z3lCF4aZZEohBMUtb9NOnc95RMHq/9qy3uulp0HlVGRZxfvsnoF4j9lVJI0c05YryQ
wIa5MF3uI6YK7WDpFQK8e2HbeySXcKhI2g3KFFyz1t7w4r4P/WpayU33F/k8jeOGPwF462jUxEE6
X9I2T2QPlUJhqwxImOD5A7z8E9aPGKqhn5yAUbPxLeWCJUj8DYZA11h3FGeLB5nYgS6nw+Ug5Tfx
MAUj8BbuWeKpPJZi1jTZrpxoGbtre+UserNQG5exNrNUPRATzzP67drfe7HvmaL1CtdPqnpt7Q17
CjFdKeA/iM6lRWpFORqUFCx6L1dimZq3kzn5Hf78SYAIgtT8rbQDZLgWxCi51XyKlIuTb9ucqPc7
57xd4T4Yj5paiFJ04umYHEsHTkUUAMAPdvpiYWL9dVNlOeu0lusjP/Vsqf0TOBw547M6+9BiussY
7fB2zDuIFKADTjDVD/+o65jx03lQfUQFqhtHkSpNHKXNxn5C/k7aRZKEU374loBPXOBFNKH5RrEW
zmNmOF7paA3H2EKGNtZ8JizgVP8TpKZtfyNA6ikOyDKZtxq+9W17g0UJUjvDxTQRe4NX/4TJmo/0
G9g0hC/3EjNO1b15Iw1NY+8QNScjHalucGEo70QGQS0aOG4o3rSMKg+6gZc2pWCRmwtw5Tq31/+w
nM0VTHnoCATH3VKcLslKXf2JCs8YkrQGfCjj3VAayYR9DzjV8d2ZxrOYbQYpeG9XlJTtvYSVnJq/
H5B5M2gabYUpnL8ag2HkqhZSTQ6c1G5omc8+wQULtDWIerWrTLW9I5zOB/p9Z7cNsZfm/slPtQWs
oGMD2H+aYbcy6FY5sXc9ekVOKcRHtvW1R8pWz1Pqc7HbcEZipcW2QFb2trLByRFo2AzgtINbyYou
E8Pz0j29ciywEFI90mbqnNbfmCjrJGhVKrZXUboBIKUr7b/2set2XgCoVEWjQ1GGJgu5d0aMV5om
fzZsThKRYmhdoQlUcW5JNbvDBXBYVFxCroYTM4x/SckHpxB9nFiZpGQN9ewOyn8aTlYgtQOqEVqr
6rWONrba2yUAGef+oYJpG13Z8kTnY5VhKNODkTWVoViYvDYEXYhU5PxPB/W6/D8vyW4bKU5thqGy
AHSbekIPqaIGSVynmbgje1TzNMxevmu+cVaxtDQmDyDKoUEuZpJ5pj9g4uo78nd8MZQzGQDM+tOo
aURBhrmXY5cs/970rAGOO8i5h27rXZFJHuLXUd+x7QDQM2CzAFTEviQcr0YHvm8ol/IRKj9dA9TF
o62ECVdro6L6QnsCsiS3q3je4GxQtspazJ2XsQdJgJ2MRmjQWPduubzKMoY1rbX+m8SJlu15pGSp
tiTFEwdgcb3gocqaQANqJM+y2WFMY7XO09/ZptpQr8hALUL2sMxHFKPVMBrUExavk4Qsm/HETvUW
SAwayOr60vgJaSSLK83s3kfmgGwmnPnVGMt4zHDaBC7RLBlWHPsNIci7BQQtybqapZ2qV8Qm5Mup
Cuqr4EjAALHRGawCgnQuEyjt7Mlb+mne3eN1KcVlD+ihdnSWq8n20V7syPH/tG4dIOMcZrLyeGJx
hw+0gyA6ebHFynJ/gFy1iSlORNWK/4XF6MEJkVFy/yRFM6GJvqFBBRFrImAwP/7QegMEwD98pctJ
l3Mw+aNXFzaxGdwD2U7tAoqonyNBnH6lFm3DkvwPBsEuwhHkIZIxmebvWGMnvgCA37UNhsXd3Vyo
FRBOtJujCEhGiCg4VVKNegi6F/IGMP973mFKitTDTNlzPma2U7aveS3bPxEDL9zbds1Nz7SAlwKb
YikD1pY1C8yV35AN1DT44b2ueLFMLO5BSf+hbIn1QHvaSM2ahA0/IWfbAm0TVUmINvx6h7SGSd85
JNS5Qb7TOxGUc9XEElOtrX4LBcVu+FwkNyDF/wm19JnY2FkK4FWefIAO2jRN/cLGrvZ0Ezsc4wi3
fK2/W7d1Jfycv2WTbW9MoqMYrssgw8Jc4TBKkg8mpmw1eOh9ziKvDhm/nBVG0kFYowweTx4/S40g
mZHNG62vXbwTBgCse/mQwCXSttrtOLW4HbxOwqAFKNB1zCOjGSwmqhImoMOXYjR3RqBBVaN47WRu
2fVJ6gJ6bdgxHSghb27sVZJDyrTZoz/4BBU3Q1tlNO0l3brzdXwsZHLYcWnCUhsMRZCh5/wjJZM2
G892NDHRlfsFLhVMvtF72fJjpP06pHe1rKQQwbmoqn3YWrNCGb0qy/tAFPC7VxuQhgwWlXjT12ZU
5/TIg/6EYkQN1fuqQIOTa5bKMkdq+jPwVe12sco1jjJtlPc87fuAaObdWwoaPEcQZkf34Vw9j5Cu
w5nkvN4pq7RrmSl2NLvvWO7hQxhQz51WhbAMG26X6HitjQ5RE146Zc3o7GBi0ZIjjrK9SyJ7anCT
2O9OGo6FTpbu88QhV8SXwOWYVbATUXecWW/tPqF4fG0byuDRmlE/WFhPn54WGcnEtD6UKELD6xkE
9/62ZXSd+PjPB4VZGhft3vP/we5iDy72tDVD/coWRLJR6CcVZZLSdoiqd2CjqpivPrDzhED7t5HY
KT/skRJGwcPeWmJa9/SQViUMeZUWxpqcixxuwHWgcTmjwuo0phbeeSS5dnib0ez9VML7y9OW247O
WVLjRjjSMRApf3U5x6N4JNfW6sgJW7VIGklVpv2kphsPtmgR9NZA39o1bmb/X+0D3yB9FUcEzRIV
hZ3E40jH2OkMd5cfKTGvF7SGxYqi9S6Bw456imov07BZUGkwCMsKewklL4G6vx1xWW3g0ABokUTD
2SeHIy82q+LHH2CMOOkdddLxUiX4oXQVs34sfdIDeGKea7+7aNwJNskSWOflTxB2Rr+SVxZru3lc
H3jgZCcy1iFOfSsrazgTvDGBxkOt/vhq8FDBt2A9U/0/28MD3/Sah/8RQfpjeP17uJxB1ob894Vm
JVpFyfm6a6Oy7BQlAKZvXv6wHAbA5vUiw4V+G2xr+Ae42916JkZ0wQXtbtmb5bpudhvATswRQFD9
/lr7ZG+Ebqb/JjAaLUuVpAFKP0u6UxBDPJqcyvrQH9ohC6C3xF5y+ZwfTL7DDglc2ray+YW5egLd
zdWble468FOamfRXhT2QGE1i0tyLR+jhOTjKON3WD0hqiFidvUbIfGqe4VvDLX5Eo4j3x51YL8F8
pHHZrJl6teOMR3E4+xDNQIiZNFxhVzNImKmVKSYup3LhCvz2ICQlATQzrnIb6mFFj50GInFYZPzF
KXDNsB46IiP/hE8lTRK9N/z3YfKjjTkDrDDHxdYPZy+5mkE/cZorZJRbLPJvZNHCzPjF6v6fvvdC
0KDQg9ck4RXYpeF8BKl5Z0675G8PzylGMlvA2zTJMRaKrQaV8d8VYxmYOAVYQeJ0i5PuSoWJXvgs
n5U16Q2zo/xGwbwl7LiMDKTcy4VC+100gkMbggSYjDRQrVLHvoEj4SCytVrcDRMsZ1P/LLRzpX3O
GHLkfDtCho+AECV5F2RPw4wt1huW/dwkttSbzeYPQ+XxMhtcxy7lOSYrCCv1YSotGwYrXEFn/EwW
L8uxeNReJomuKPhrzo2OqrsF8YX4PLdrfb1zVrkECW54gwaMft7yyRtBo/Y2gRarzKixi/kB1Loz
hMYh4WqKk5A/++Mh0pO1IhR9DkaSfZ+OGWyUeMNP9ybVdMd/+Nv06dXDUyKmBNWAAy5I/HkyFIxG
o7HlsW09UTNvLgIXggnZgMujazrDd7qaRZrnXJwbUH+wa8T7ugIa5kG8wcv22bfgXK6LwK0eQ93g
gMWvfFaaHT9CvmrF7GpCVOinHqN/3FbakDMInuM/CQBhQhrRodzp2GwM2shS+/sycj5QcMwt4uL+
8tmnRgqE+lHz6VWkf5337yi/u9hmGJ9t+SHf4dLvNbrcvrNzusqDBhDJiaq8pykdpW6Pu5JDQ1My
a3ybs/69MpcfcJG1h0B86X9Rv+u/HNJyy8te+zzuN5VWPnyoBZoCdMQR9j0AN3FQd9w0CWn+/FmM
RKULea95+Blju0hp4yUZK4p8IA6C6WKKAaKvLobV/Isa7whaDj8PqmdXORT2HhBk1bFtxLGE0ITF
Dvr/9FQMXFTSD28qAPGh3Bi21jn8tE3Quy3p9OPXNpaYK6U/PELYzxPS8pO9yFN1pWRGywK6mWlY
PtXxLJti5W/WpWNJBcsnX0qqXUH7igtA6utg0HasFSinj7eCDJvCoDL9WjiwKlMrakAJ3Tzq9AYa
A2MZPvGMb5i2QPk4FpElSUGXVZGH0uDmV6UKv6YWRYvNv9MR4/ciNWmcewxUouJ4ipmJDgOAPBqw
vgbBukRvEihfhOS6lFvdBCdzxlnOw1XBIjuXXWlASQlUKpomstzR2Gkp6hqCLvIM0ntVegkQJkpN
csqvzq/eb94Uw+m2pMKy8IGrFm3gujJoYTR3KKRn+uBkrwupqi1JcjL54ecOZb+MfQItqPkecWZV
FQxtAC+kutchdvl2qHWpJ7Yon6BuWJfeQOgo4JT3DFtcZ+Rj3vC/OEdJpvyC30mutf96siZu4que
Kx5Ij27uerRDNAdmxGvvOOrsHh65AkjFfV7BwfyZIIwmX+cSITabiH7BL+JbZ0GtEbX6UWHaa0VO
cdYyio1dwdnY406MNFq2qE5Y2MfgdcRmKoSdgodfvLZncX8iWBbmYQjRYlNhnDeM83cg192shM70
BWoUz7+UKR6joV+pjV11vxXdlHKczm/gdPr85XEgrcjJMiqtUJGYHfQzG+9Dq/AxqdCGA6I9Lv5P
Z6facNjsYbhq6kIEZUe+kOJBIVLqg51H3bKI1im3kTKxWHdHlP9gHAJ0JzLgMfMZSp+k30p4zqSz
SYZ006PtWfv8dF/gdvwMD8aeWXZpbOW7btfFP97yyRLDEoDlRKDl6IEA77flsRCyL8WK1wsBax9w
HvpmrvZf1ymTXzgQRRFeSptnnBLupA490hBplAhCIAGpcku+I6DMB3v29mwtmJ0p0NsuIrgwpdfM
UhTLXKamck9pU3CWkOzLCIfXATfQfHgPhbf79h07WlLcCiu/Juf3Dt/ePMZkYTTCyOmh7POMrfb4
orxwXntkWsZ+sCrVbS6Rz6t1vzt/7a216whJ7j70y4e2ng+Sqmxpu0p+Y1IG+EPo6E4bQon/LQXd
cM1pfsE7pD8ai0zs1enfcbYbAp/SROqmMOIOsIXvD7x87XeU6nZmkIKwMqr07xqtwiI0a23gbhYk
innElxnShpxwX5wSONHqX/0FjsW2N5qUHAmSxBEQ8VWtZqJ/MQ5mj/+dh0PJ4cBz06izPjZifrIT
fOmYgrOjYs/oi0P5t20Oc+D3pA0Ry1OamXGdBDs0tfy+muZ9yD3IAVFDneBbJAgVAOZHGnxLdhtu
66xQSwGpv075edMQycLG03vbO+m9YhXgsF1EU2PeHMm7jQXO8i7bcbVtXau4+5jMqU1Sfa5xLD9+
Q9dfowdNe/gU7RtVlur/WrcYICOi3LI+x0eiw5ydUKVX5htpQ8kbB5IRoOweJnKLnUw+95JTLbTK
fHsfUYOGycqXS0wc9e+/JF0Cjso9/n0zaGU5/gP2g5Yuv7yMS5zjEvuvrrA9IL4RfIo5QvX2/Uwv
ESmYMe1jv71PGhrXlrvdu8PXk6I/oPr2c/5oxPfWFMtVy3CXYfDhukhr3VtUoWWz6KTEQbtkgQHQ
n/2KwkU81PtPM75nX7khbPd17SfSXmQJRUzoJKN22D9hhG+/ncl23U092Q5aWlPxj7oxp+zznRNY
+ZJ/0mLq5SemVy/vnMGSlqs/DjAmhba8c6qPZicgvZcOQQq8tnsPL4iuHLJaXk0hAKQO1zyKhGEv
rZ9BbX+5KL8k8WHktCZyqe/WcdSHv2sV32H3Xb30ePDaTxKwLg8zGEOKigjDZgmxymcgWTbj4gpg
DvTdrQTjFYEDJu0n4b0acQyjvB+LcHRXQX7X3+CjIlZOgIMqMdFAnw7GJqjIH7JS4SXMZSOcs9Dd
WkmM5J/7B6c9VAm0HCQ9RcNXINBunKT0LYy1PBgHCFWn4jeIxcIkv5S3B85tnpXfP8gZYkXP3qnL
fchpo78SLb1KV0/08yjZWZIsEhuE2h+zpyH4uuaHq/Osnzl54to5MWDphKh8NoXlD752wOER5hR8
SVfvwjolXQDOtBnGbIRGvlpcLTrrjyoDthYoGT2P2gWMHBXGEdJv6ymCtVqMbIDOIODUTdoh9FMT
nAufrhxkEAhM8N3AR5TDjGT8Siahbanp2UifWFhaCRAgKKnDe4zCppSD2DdWGQh3u0mjFrZ3LKy9
RidAP9HaP3SgenpAGr+MrcEj5UHaNXHsEZJIRrcytFRsosNsb+5OlDPUemvKBebxoTZm1tLlkyGH
jDH7YJVeYqAcmXTKjSoJD/KhHuYvhC6bFK/eOd6WodTEdwCY8rk+qBOQbo2pCApK7RLzdB3Ab6pG
KljmOGrGzGRfvt1LdlB/Re1jzPoM007ALXG3/rU04W09XmA1g2ptdGHTw7o5WiZBWTmu/K0ILgVg
19PaikY/VzL378kPVmULumsEDBX0k/+vzXRua74Uiq4QaOeadRLcaRnzzLhXiALuzk2Z1xzdbaJL
qA+wFA3X7AJ/ZCDAE2biIJMVUIGi3YWm9jpoNyF0KFzVOwCEXwsNJIHTiJC6cebGF3iGeWXikfqE
pPT6b/ptAATkAdwHfPvytLnn7VYcgd+Ok06XASFng5kCdBjJQb7CHIclmoeaTL272y9mJgwxkAQS
OKxMnSZKW0IquWiBmKwELIVOUnlVrU9DRoa3tknOdtF/MG7/k84p/asjFVU0koLrRzb6Ab5yQ5NY
B9lhCadqknhG1ULmfYbzLOJRz+HMm7i4+r1tAid6/zZelGL/tz7ldG4g+Wv0EGvuOqFHwApAXwbB
V813rlq5Z6p7sB4rZb6x3EPN+0ZiyICYbC3O/GDUvegCUZPpR6uidi64uBPeLyZFGSKv/LZjq2Ed
zjGltGwcBihh2uTnzys62r8Z6aBTfrFZuBZEiAmJ1MSS9b2C3iz9mODL9UKhcHxBveAJA0KQIi9h
De0JKAg59d6VY4kEeg9dw1HUaPIfZQHNAwctNTt4O6WY99gvrCYsf3R156JW1bdMA3BlRG3aC8s8
mhxK+yUQXuYn445bQXB5P0CNip0urvYEh8LrCSfe0FHRlaQBqQyPq9e8DCzcUy7X6BRUvUwHBKyq
9ZCo+z8yh2Z222YtC3agk06sKgrjkbm3RuXbzGca9FdyNFuvAZ66tYW66aLY5cuNhyHwOWnSjSBe
MqlZCen/5AJB90Y4E8A6pw+XHcmzSThHkqjQqgd7DsUOKuAMfXAkkYpA5LidNXyfMrW2YC0wYsoD
WBr6bJh5kNqOf/E/sSKdaOnKoqWJlTs0yitkYcbCQio2U3/Jt/InsCQZcYSaczt6oMDq77yZ0k4+
rc4H7S4dlkI6Lx7SmBndOwcXbsCIDILew9b27GmqoFG1y8RndNMkpKPLT23SpnZMaE0iepXVjirf
Sl89yDRzlkptbSF6J8hJRTONB+PkBl1TO2+7N3G42FMYFk4cAgnyPqJITmQHcQ634gzhV7akVHLT
RLb1aL52TQYK6viCU5Zgd5pgcrDg1bRzQIeWndE3tz5zZAuo5wbGwOc3RvlMzq25kVwtWY9iBtkP
bSamJxL+c+lvUi709S4zmWHv2VASeExmLBMiBnWTME0DlTMNLKSkwZmgaW5iQ+CoKf4T878QhKLB
Tqr8Oy5R7g4KycWzJgdBmYbD9xlO7LU05c3B4qG/ZI0f4rDUHFXVI9x3+BLRL5NAWDymWHfIw2Tq
//x+M7TI0G+jeYloOEd13QBwDzRb/oT0PlAuqB9NJqIJRE36TAAn5aM1dy19BIRZq8S3DdWiNoSu
2fL4/ygvNHVyinJ4cp5v31Eyg8FbHHdQ12jkQn20892Epq/cVVG3I9+VPmoRBDSON8IxB0Z+1Bdk
i4TMO1qABTEVC4t/VcYAZ1K3ehDSEaI5Y9ILjwKUAKxZfZsU0qT1ovCkazfVFSqkZpuNNs09Wgcd
MsXV4tvY1xqYPSFUwpwyfWctC8rzup9pjJpVbZwMszButMH8amDv4wAVbRc8b6C0Q2eJlxrekAHH
w6XzAwneE+R1KNbjGOfJmPc9Z6L/3aH66Z4hK6e2LG4i32kS3va/LNVZotUXU6OuLpFYwHLWF4wJ
eCSAqxV0rFeibN3E3C2Ug5/P92B/o914xjJaWqS8Y/OjHSMwXBwzTFmM7XnDn+pZwV266LklB2dQ
1NPQ8DP0yCDRa39p5hNGLUrWe1jKydBEV7bPL7FYEqu55FDXR+n66nmDOkF6AB336IoSbVtrkVRE
vSjcH9CmUObnJxCznLq5iR0LjoL/htVx/nBqvWI1c2QKyigezhUXIs8qOtJ8TWS/334+fu896A69
VynymX0Vt1YEavnl2CS/wl3DVRO8I0PKArufKdCjvwE7V+IDtOrzio90aIpnSoKsRcQrt5DyjGEL
lpbNgfJZmnXmIXTC7G/2/ueF7qQupb6DNJy7QZDUE5LlGYG5AP7I4TMdPeYkOMgq0zEn6PE9Auhv
wVQGMmcnUnCisR8jgsUxcZjokvvVYyIXCE0Ps+tdgWxsz04zlkZ3yj15hktwV6Rnhychi1Di5irc
8tajCvQS9vBYFqS6VmlwwpG0VpY7Q5TyfcwgKOhK8PadS/F17svwl4UnMNxilyvd9H/hZzAdC8B2
O33Ls5w4xSPmGViGpB4tqKfpH1RLYmwnyjaoPysQuh27PX/B/eURG/29pZ7uWdltpXwz7QHwh5GY
lxfIBsam9FeEXXhJBcAhkSn0IsVH468VZxZWO+pzfXNlJ2/mWqs1qFxTwthgpH/vZ8vAl6f3h4v5
vCBINChDtgam2D07YzPkxdFNk1at52LpWB69gW5X6t0OZvK3DJ4KujVV0HUMXsCDkFzmqnvp8PIg
epXXONVDfMVZDne3UK6ZQDVKOGe3E20W3ynOGg9Y/0uX5c+cRpuZUj+1DThj8VRZsGiQ6Khbo5E+
3+VpK0ALGOs1SCKb6SdTjGh0qbLmZHcX1uRDZgn1Qxo3l8Lo0ucCPZw29SdbD7mefTExK5IxgQK8
+7BTmi0EyiskcxbNZ1ykRJe1AczjfTowXZhzOGrhMPj804gqvefTvgO7QvGh5JhNzy9omD6Mo+N0
SwjOBTIzIR6tHHWlXRQ66mepiENG4f8500npFDG+erXrqO9UAZwjrNMV1V1Wyw23sIuXx9AIvr0C
3YCVOKUIJnWG+o86v2zA2qYjnuHq8kXHbCrmzXBbvxX01Bugy6s2piOTt3P+FbZ3rqA00TU6TyGr
aTZUtDhS5bsv5VTb38ubxUKpMnqL53g22FK+rtGC72clpuW5EwsVYIlvxTpiKGhlNbTPpl/tFhVs
sZb0x2biENH3V+x5ghFIwto+QgzT92yqY1jbsR2Z/ILYEc7dVbbrzEdMBCauMl2+oNPzLNelrxnc
wYxxem4JB2a5Y3P0NxpMH0Vvz1YlFTYpNDIp0vk13eLPQTZ+U9VO/DC8q4GTfCXlP8UVbW0NGAjI
szvQs5o/YfxKy7muVHE/IE9Aman69Ufj+7d/mDmgWPxscTVxSfxjEHXR7zkiVgvCgVARmTGDXa8/
tEuMvSKXK5PgLlg+il2fRz5zVq50127peGs/kk0K4mlMRWaGyD8Q/R3abYbxPvxe2+Rb/QWYWDor
2R5HjjFcZOMGxKoiurRc8WSX2ihskSBC3QOZ124SjYusHKiCFnrA/4daJB+5qurGcVcOr0CIPP63
tim5yT4ZD4kjS+A9wIGl+oSgWrSKo2jGf5ZA61y6ta+rb4MDxoxRFUHy8hl2i2cVir3wXanGackl
8HKC+zHZVyny+r4Q0151zyt3jrgJQqV5Qg8Lp9AwvPxMjx+DAAeLMu4sfmtUqEzrF9N6ZTEMLsP9
RCV7X8LgKeuMwoa5YZ7QsbcIDkLPs7KmVe3y9SI/4O2Catzph/KaCbEqhaS74+6AvovVe+Zn3iVH
3E29Ae5sW/qGmvjJDOHUZ1WwYXOp2KCLBkZZHuzf0zJr5GDsztyZwHkuUFpqccWKMzl6H9QY/+8c
IOZotBfZ9caYSGFs1YyoSmCqpARdEDRK86akDVOHmfYhKzfxaOyg1D6H3sbun9MuQf2bb1shJgGZ
uhtOqC/DTcAfzPfgaDA6KJ5oDIND02XutKlSX0lgmNKlYbMopcyB7Q1agGcu1n6Br4w7pXJFqqpP
IttPFebufSyyilT7X42Qp44HJHBiCBS6wz75pQEQplLBXCNwvyuhLxZhbKs31vlUK/0vPLk3jcU/
T7DskOaISwfJWpx8BwPPHe1mijFQrEPQhYcVFh7DCIWK7sMjNcxo7O5rshhC3y+QFQ46LCcXGUad
uIYExATEssdPjwpCiG0ydIn8CL9YehkTTSBbq9pnA3PwIG27MtY6k9a/m276NUqDqtlHp3aSqR18
u1juN3i14q4vFsS/u9f4rqkQVcq/8DR66mIzgIG+XPN7c2WUHNjGtY7ctgHnrUyS7FgngbHzaF2w
CRXM852qToK9aUD0Mr7eKVLWkWYhS7ZiLhISUXyuwABrXjA726Us5lbZs9k4Kk+vpzdH7ShSWEjB
GXFHWkMNDWoxK7mtukLnEGaRomReFIr1jRjBJiHtUz42XB6Uc5hWxoBcuZq2tPOL4MceeBBoab+D
ra/KFSpkwUlGUl5dmHL9xXkOzqTLb2G4+zFKM6P50T/N5be+8rnAZt2jDk+7r2HvA2e4jmEWaxba
m97uv87drgukbBYDDK7yRJZtKOONzL5yCFDaKPplB/JAKlduv4ciDvTYKDe24F6s8kcEe+gVSCOv
IbjHMn8dzO6w4BlUTogp59mLXFjr9vAMqWRkcY3CGm0mKUFoS0wOI6SVdD2GmlLA7gFy6UKD11eS
wRAegDrQv1E236rreYpFuEBHe7LX76sy/zR7nexEt2yo9rjflucBgI9N3gpTZ07En1tg/gFCaSUf
Ku550FZWGrjjlrDjxT0O9O1vHvELY3jT7tK5uEbEs2fG6XDHQvl3O1boQLggCAo2J+G2XewsYz2Z
wNbWT45sDSnZg4oNKZ324UUhXlJ+woXSXXwSlbqr2CzAUYmQJHRPEDYwO1BkgZDnPvN9FABOCkmc
HXpxbjBONCMq7Fb+n8DYyS1NgsZexQqDArGp1/W6wZ9lzumMvZkiDMKHBY9hrLCbmqpPJ0coJN0k
1+ev9ekzHJb2KAWsDRhE2DsnWQjn4ybN7XuJoXsmGxVl8AuyEIJBTpLVi4RIRY4VbdQRVUGQwnx6
qSEmGESQzjLLbnKHW6JsJfOSDec2mxJx7pZGWwxMrQNujOBBXGP7qOMYFhv1U+bxJ20cSSF/A9pQ
Ggs85W82UEv2MG5shRJF3cA1zAuFZ8SqRH7kn/JrfTDdcvJI7K460ScA1odAYaq0r1z0fhmO5AcL
pa4BzjAeDu8tM7ujZmxM1+n8bEk0pGE4yJ8Az9d38pGIMwIvO0gj9V8Po7lSu7tt2doeyQtdkls+
kLMCA9NS/6FMWQ+9PNeiyKnwwUaaCc8elp1kSxAaKFpSDD0PALF4hPhw7RLjQbyRak97xGWhUs9Z
6oIm3ucLlYZr1SFdKj7TgvssTey7WWv/zy5Zw/VC4Em19geZspAP06BXeT/dTmJrntE7sX0UPXGm
P0eN0xmaUBE6oJI+dosZ297ZL7ucJmVCLmGM1tWf1/mLEVDYslERltR7cNdapjX4DAux6dK0fWfc
2vv/hzJA3kU+b7Cu/WKW+CB/dGlIjQMsGxhpoHk15ah2hTW1O+WaXI6telKObga/xOKMVpJcQ83Y
uUhtylufEqjmlRjdVj7YsDIDgPcxRuRZbPPD5xl0Gqh2uPodQQGStOBTTDbpGXFI5MMpQx1D3zeo
ffobyR+j5QB0KyGpeTr2L16P1mG6O8XuJpRTYmYjmArrQGhV9obA7cVmKbGUBI84eC5EekgPagNg
PVad6ZiExbZTowSe0pUzAtHwM4k0RI58ZsMxj+ZSLPwGrr7FkuFdNJMjM4BzW44JfQ9fIgiebWmh
08mcWHAlQSpcbGGEmUUeSYNR3pH7l5M/E9lWnYPGzCHsID1tqdSz/tJXKq6XBMqMOukCANZJiN4k
BdgT84DeK1pTEH/xVgVJUwcr4EIlw6ji2w5ZqDA2cPTEobMLaU4W1pwMiP1XXqFyWuIcsFZ84aJs
C2FlYxEaXz1PKl3u4xGSnV5gSbHu2wNOL0Xkqy8wiB0GQ5GsvGQ8hxjkXHWLqUWTDJfyJlNG6uT6
cfUNFYPW9BYZaIJawzgyQ04ele8d7nPGXCKfcRmemCf3uuKwgqwR5mWGg1CTXQTZF8UFJI310Tu6
jd1d6KBhpnd/vWnlA/4fUILnQt6mCdWby08RnaxBp9C9WUjoDfpmTFDZBhSLJ+Rzra0znmp0PkCU
cY4nCI5ZIS/kKFHzQWS2tIWAdQEQk5zMSREeOF2DVnkZdRE570qPF+vSCcrbwhhngreleVhKyIEu
3VWsGD6eXP5QATV5+jXRLxJpJ+rbdWM3MlPFMrt7zi3ycIbE81aPflaxGYYNZ1kOYeP4zrN1edAV
eVgRbbLp0eyjBbeKPgg6KTyYYnCCPIUZ0mOY8lfjw1imWDQoFqEV0kKJ01Pf1w5MQ3lbXWgxmb5E
FRXWWzFAWX3H0+s86MY8/S4lYsUxHUTy1Ew+jWBZXUjqQQw0bSu+Z/ORhLdLnKlM2NyB1hz6qKRR
W7nN8LADoNOZY/QBW1QqxeGrnoW8hxz1nlzG6o67cHJs9kwKQkg7a8OBwZglaPOZq0J9YvirJtyz
izUaoNhEze9ntnLFDIUpkLLeWWv7CKoe67lTaTCtZoiUbUefVn67aXFsckJTVxFiAJKIlfTtDEc/
V6JrIzBK9Jp9Tu2iBfGvMM3Ehdu6+TLS/ylnmoEvcnfu5nd2Uw5i2KEU7q+Sei3ErKLpyWHclVDr
yUmG+fhUkVPVX3XQytz+BSi8BZwnAAbwnQwVeiY78rQkUReVvluhKqxTP785FxODFtybrfzTrhSZ
h6sGVRNKCquuC6XlfTDjBaqcJk2hnoUBasKZEPWAj9B5LrM33qHmVDMZZWByQG9q3kBwBfIMG1W6
+WO/JwnjEKU3fsWGf9G7Hv8ixsChwOGRrE/+MZyT3FS1n9A/6DBDZNxKkehACkslusa1ubBQnR0E
u0A4hMz7b1Bd5hhVIKqT3I9EFEWPA2pUUvZV6sydugEBNQyUz0+vIRRbjj6QlB8R6tjhQ7BlQDqB
G1JTw+H+wrO+PovVC/oR86a809M//YEl83QHA6crJVCl6qFZ9YqcVP1LU91ERF4B2Ji0ysD41TJ0
BEGa02b43Yvg+IGhIFENqGM4NNLjRpBcpALpuohrA42zGs4EKrvAfrqq/EMmGz1Da1/HnBJDWIKS
vZd4HHc1O14MEMitDGraGRA2ornQhkq7epVuo5Kw6w/COsCfzn+2mLHW22Y5wDWGSt59vE05WrAk
vEi7PzTy72tYcSLLCFSIUXfEF9BjAcHwB0500JDuyWpIqQbrZzindeazKG5RiLmkdbQXCxm/q3TX
wrjCC5VwPKkX3dLHy4T0mz7AZMxG0a8FXu9dDjZzbCEn0PBBx0ZnWuZJfO0J6MI4t1QVT4Rzaj9V
iNRzv0tnRvPNIEFREcKx6oUY2+59ksQtf/soeEzqteEKeWJiTBQP6TAqrfyR10uLW+Qwl9gVtXJf
wwesCsmBU67IfbxceoK5/w2RPf3dvZjCqt19ubc9vYnSQhcQg/T56P2ozmmESOvnLPA1xUHRtgu7
WPRnGWgvBZi2BL/hH6goS/9SrGWY6OPuLAok7alRJkjP8kT4qsXvXd01RFDU34bfTAk1KDJt4D7z
yAYfXER/Lyd9UtgUVauH6ksRGgelapP32jkJ8aFd9jkAsDi4GfPFcvs8khunHLSWRjYZ3CR0UQuK
V1l8CejZk62z8BkuKG54iju+2tOijS70+sXgBcBZJiFLSGKxs7DShA+dLR9mT+gJplhwVkkurib/
Qw37zjw89DChoiL+50Ybo8yapVwK3+QeCOCUxy/CLFIBmTVU/4aWTvKUDz7uv8lNTvDy+S5BRPh2
EZzCP56PjOkKbOLyevEMnSx4kaEH0jsoQeYjA8vuMVj4DIaX+2dkhwaCXQfXpI3AXkyQQFHcC/y5
95xoQsr9li66r6JtZeQNdiU2fN+6+hnvVNVJnIUJkYcZRmYwv0GZONo872gf6ka3XdQguPM+JxKM
YDVSaW7Cp2G+GRdAqt5FCyso8Wwj3rVz7RnUdh0sG9sWN7YsDX+XgtfTCQdSDRL+XJT4ggO1kIg9
7SLL/YlkXGh6mEdcoR8e5W7Qi8PQVYhoSFNUYOamG6HTeqz4YBs8EEQhtRv3LtCVi5YBYXUdNPmj
9t6M7BUodolC1NExRV8JAtzo++2coA+bx3t3H2a6f9mwyskPPuW7V5h+p7UTfhA7gebqWdWyyTzL
IJQHWwUns02gUXB7+x24ubhKQkQNtmpoqBxz2ecWhJNN70rB5nzWT5UXmCX16pQrDKeq2hY7Jeuk
QAknq3AoUBdxIUhsaa8d+RK8w2cJzRHhwAD8FZoUurW5hzU6oKCMhPjP6lOMonnCRePLvpcq8OdA
/kl4ALhWIU6TFzSid5Q0hza8duYOd7mzj3U9/Ht9odrQYFq3XtaGuCOZKkeYLVnqdQxl3dsEYOex
LKqwl2HvgGY9r245jWguP3HFaEj4+eWV8tuLVS19cBs+YkpfsrqEveXjYaGZTGdcGJTUe4WFNBc+
VujlJMXmJFEGMDEdd5jtZh0M9PBJTkKR48uFBdVqpzJ7PiVszG4QzsRWJ9CYshpjjujHYlEMSVv1
vNfh90r26yIKL5D6+Ldj2NeM6T0hFwyBD4YMAI4AZ6hCgBG0ULLCQNJqGG9oL7WpbdRsz4FAJ7rE
M7lgrqMxErSTx3Jb46sf9Fv5TvAbNlpWCCkQ39m4qNYUduWyVafQmlXdgFykL7Zkl9GoDaZo3AdW
n4hxk+6GuwmRIPkRYoH5XCqCGIgRNiR4JIevGTKRK8z2D5xUwwocJKCiMXDVqc/C8oIdciVkUk/N
4W8QPx7wK5TfFxwwbF7N+Ma9IpnVX6+pT9v5mUNEVvyIbIf01+U5wHLDi6tLcI+36QDyAKgRu3ka
GrbnvomOsG33BO8adidH4/d8UYmyhxnrGCs/gTu6DFf0u89MILhk0GN96oP3KLkA9rQUy4ZlPj/N
q+w9Zw6ZxyPWeuAOhUTZO5CWoPwR/MdbDTnvnTuZD32lBXl7cCubZ+FSG3F7Zxea6lmbgwvcHCXk
w7ZflyzAU3eP3hWeIlploYZZS07OgCW4HWIUIQ94zsnkeq71dfyl3gIggERhx6ue4kueFQk23mIC
EyUOY+RbdrvWqjDRFxbMMEUUtNUK5FQwEq9gOoa/OvMP01wuL6pcLSLWcCC1iqGVeNqusKjwpzFx
Jqn29HGhgvstXmO1TOcozipDCSpCQrigqA+gLxlRCVwuzhocwxdnHc4PAAy4TjYEo8VDHP28P0Zc
acLdLQqnvG83c84LJncwBn/lFYvpXR4eLMj6AF9AebLasFgyRmh8G3VbveEY/05bL1khIIR91Xt2
vm29n4sXk7mY7eFEiqX5ILpSpQ0y2dg4+89nMOXUxvGeBrpxBvbNtJadSdiP6oSzTTKTBA3WMdeZ
aVoLEX+myx7FHbQigk6C6pbgW+jgX1qTailwEdp9aNgYQC8n9ewitceVDX7UFqCzC/jBe0l6g2gg
lQtcU6i653fzA+X+xGQxwpGW1UFyQRRZpNpowf0L948kOGdlb3CYxzJyPr+dCvYcmwFl+3kyOUP4
tQsLBgciTX7wXRFgE5rHz1s1sxcFhSXA9da9vBzT5Hb0ES0s8IuMiJjn7+MrMBbP8VFkukMLjazF
2QjOSumiCq+VJ98tXaVRpHSPHqCsw0Fcjbc1MlK/FVCsgXUuQylmZqJ+aoxjEhmrmeey8+F9RTog
w82jMLLhMvGaAxTxInqUJil6Fe7IW6bmwhf3wjmzcCmIMb4NbfGKCldT15wPT4Bj9gg8ogzIV89v
2W6NpUeLIh9vKA8UAFWKHZtfFLeHIZFMANLijNCTufqqh3T/wmeZl59gPkJEzAyUBBD6Rbi/70ho
yndO3wlxV/A7Z3QPD72rHKtCYWpDP65EQXd8WJ6HYK29VSJEGE8W+WDTC+K3vYneawd7PBIjzaP2
DiN62EdygICHwIwi4vztxVmR3k1MqwW0YA88hhkyd0QrksstT9NXg2p6sj3CjxpwdK8hhgzXZ9CT
BGLOTFvEhtjzcMU+G6kAdeHg9ZLRRbx8sfHHFeqVxdpfn/1WfrrZySwxD3H1aDX5jWxCj0WDbPdC
ddKvhahNvhsvnCYJfmaMryO3VufgvxNdmDfSsu7wrNQB5CBmWy+DA/YLYow0G7CvlJare6qNsg4B
DUa/jJWXfx4tpXTVzkQQMIJ9Rfr4O0xUQvpyz/PBLhnomt2s/n0tDo9dIE7q6ghlwKzvVsGwAVRY
KCrW4BVu9mPdO6Zmvd0gE0UBLz7ZIBALdJAILXtqk2l3jMOs1PYAxFnSedVbhsId/ACPLOqvaU2K
FbepwEeCZxVOojoEIQJhsDq4mzXMuKn8KMu+97QcBVf61pxDsDjOlI+QtM8Zv5LR4egYvREGCOSj
NuBmALt6y+uRGROhR7WtI/YU8BVFFtc7rWm57akReYjDKxQ26yBRokqyoJr6WQ3sOBzo2k1kGtVK
PV26qiQcontqJfnbQ9xfBOLmWzfaETkF15U6EfbRG4dvZ5+Vs0sSiw2sFAfKxmqFUZCJIesBvyuG
9KH1/zomOutmwGP5f0U1kMCk064mQsb6ZvV0BGEw+zavYPAoiSHUJ5HT5+/MJjJQsfgJzjG85KRf
F7i0IkXclJb6jHFBBbu9owgV0iEoDMizItRRpnZWv+jOiaRaO/W69M+PQ3X4yGesuINsyqTrHCqB
A17sPxbg2MrCkWqURlK6Dwqs2eZA488F0PyXwQKzi3T2vmeoQFTgapainoPE4/aBwAS1K6eIlp4/
Fhbry7eXsudP1lpTe0LIid7nPsHH+Ndjuq2liy8qGhRAp3gxv2WrPzrA306iy4Z+Fg/F5UnHtVx2
pUEgYh0Nm2wIKRTRf9G0ss7xqhKyNPEVW/EFDUzsuIxBgSYNCz4NynpvPocR8AzcxYUUMzgmzgZa
nP47JHyBPEwWEB39Z7ur3SpPlzm6avBMAiy5iG5JzhGy7+MB+0jno6Ux4p8bIqw2q/G6sg5NcWLB
0wBFH3TbT0zvFm5pF8RvQLo+okrn4QEnIC/9/sG/EVMit1s8LckyIIILmo/Xebv7rrifk3D1aCU2
xcFurTIvQjiKdVcj7DyVtabUtAv6TsxIsI0Ptrs8aaETOnBSIKW3KXoZUqDLa+y34y0K05IHLN2w
Ww0FeXcUgXTYiJp4rvD+nnEjieS2ZphOzgZ4bA1inRI0n71jm5K5tKbLShXc9DVZ6skZM7+xOsr/
FpZaBR0WKwRizTjZd8CvfuQR+821P8AjyKtyzwfnb5jNzFTOJLEVKQFdp30NkQPzKOTi9mGfiCuO
jPsqLGq9wiClZDR3LuQE7v3rG494AOyd22taeAEWQYw/cyG8CcrmplWvatzKFP1htr4hNPuFn29t
Srl7j6yx67u+A5OfVn34HhwR+J81TtLPDloZbkMQDNMVrh2JjhZj+87okr6d0sqUJtZEgLZiiIv4
X2HY3XcaKQm9eMt0MQ11m2yWW0tg1uG3jOI3SMA1T0bdQcNg3x1QNe9xgTvWl+XqwAmmIttwmukL
XN+a2Am9QTZo0rej0GC10XMK2d5FBNsAT8bryH7Y0TE+eMNENTbJY5EY9SGAvvVJOayyhqpSlS1X
Ifd30Nvl4EZOmT1fsNr4jx/y0TXtCE21H6/Ab0DSFrj4Kr0zA0QnZH4HB573zymf8WYtSSrJnpGL
CMfQDBS01qzyj2NsdHBOKpTiv4h8ofBwLZ9kOL1grGe34QN3OQyhqkdf/rWMn+FwQNlIkjr/INA0
Yv9hEDS4/7apwdnp8uXEckkgxM2FMwEijTmx14btchvKqIsoT482fSzZmpmkO9P0DXmgmuXuAcW3
VwvmtGQpp4k4W+FIgE3Dj076xR+60nou1z74lfhoe0+ns0FYKUh+SFYIanmArGtRa/5Y3jpLZ/d/
AWuf3tRWNgopCknGiRqQzM3FpGzx4gZG90MvSnlO79ONw2IPG25gEdHKYLdXpBdlVJufJZK09X79
HXkaJGNTh+KMQs0tjdOYipyCyE4f4we2rArxc71K1dk0xZMMF6mnRMFmhAg7PuLxqBIcNh0hn9Sg
E6bK5n9Wjz77tft9WPLVkrNu2+8Ip+VnfKqRpa/zqO+3N/75fT+i7xdp2W6hBi7B37K1QhrRnBsq
KdVN/krF5qOzpTvW7R+KHX6PgNSFeUvWLvyIWuYBv/1LrANyz7wGxR3BGlasxIZ03l9edz18cDZz
2Om9ybKW5nQrvyv0kt/DxCVdEd/o5QAxFsCI06Gj7EdZR43zEUaEhrGewUQX5FqtTeO+PlkwxHAP
h+EBaEEbRFGLREMWyR7e6LjPvfn8rRCuodJQ7lrkjOUlDrKzZkWkL7bjFTOsEWcVaoyBdVdqRZ04
ROIWJtqh6SNfcg3N27B2JsjVZMUVBBKznYgugBXH9fp/LTHxRnnAWWJSMcba2Qm7W0JpfGEwCzwV
uVKJTIKksm3hRFS7CiUyO39BxS6lM2ThfQDc4DwUmJrfNOG3zReBa9K+F8A5aqjFy6JpaUmjamDJ
4Cc+3KF72yZPsvnAGRqvvjV0NePQsGKlHFH93DI+77vl9stvwUogZLTyWQ5xGZcawuXUKOdmpI6B
h3ct/SwhkHsl1+JsZTJLTEzNyRfvzZYGdFr1wuY9JKQe9Vbom+x4209yu8ZYC0NN+2ER7unpR7LT
LBMisvYfCwAwi39K08KJlBuwCPPpRD+W0N61yk81+aFoZthAxtxOSHe8gXmQLGbxJv1HKQpt5eMt
moWhSMz03GdnhaK+MGtY3fcR1kXI6ex8OPSiq0XWuapOemkOOTZMm9HeUCghQ5rgYq8kBBhRUaCA
uI+E54wTiauplAO1WNIrjO9fSLwe3fybbmmi5oxBY5sFGo1aa7yQFSExdidQHS25az9yj2db4682
oQsqf6etV1EoGslFvE1nAVpfGEZ7FDDu4uX+QmJcmvqfVKowOhdrHvJT/ymn4YWSJ9q63saav1zK
SWYs7XvsBSi/3gaxPM27IAZtNfonHKvQ1fcnKXXC2z2u7WitafKp+n9e2RcPJYyxpdFbxaMUhC23
Nh885+b0/x/SedtDNp9mrn37FToGwuAOBbnmYP5049TarsNhnhEDk8wmrBhxgBgdK1R+qAEQZmzQ
rf2aK9JnhBGqGmabo58kIJrwqPeKPwlEsklXcqkmR1VrREs3X8UQV5ZcYLa3WINp/YGWzn+lYcrB
G9qD4YxmERA71VGdHgNmE2PBEwyqJSD5V8Dg1nhFVtKdT/qJyPfU7QfQWTXA2gysp8sRSsXkmFum
WavzGF/PbZfG6Kso8hPzltNUOOpyik1GWN5fErAk9UNEPwjxb0CAHcqQxVZKNxEGL3sVcGR+By4H
wGdck1VtxXhMdjA+rtFT/YBP31h+YEkjkDMIQrengdGHxQq4ZPE1sDAXg6+Dc8P+jMuiw2qaV8VO
KC5qi4o4rwu2/I1OtNJC9aSVCMKx4zzcwGREl0UNwcuI5V55/BNjkGb8uQuZL4YFNqzD66UOHkle
PZ9iFBD1PkF2/doeikx/GzmWM7sMCicuJ/XX2q9eCNdebxeA8zjn5XqIxXS3ea7eyNVOV2f+b9KX
HXZS6kHE6Nh7IPt1PKD30N9KRthT8CmRfu/oZfHjN68frgAl2GprzGcJTdvXyCyKhsw21LbxcYrb
qGrx/3RyrbafunUAGPM0T6CxF5/F8LlzLNvq832eShER82PwEOMUzC0BuSEo17SC5QdlMCbKAiRo
puEjSP9iMSkNXNJCzHMROzr+EnLKHoUgV6DeccXlsVqeK1cnglPquAxmlNshs/MMQHHfCc3R+4Iv
96esi/LESho9F9TKSUf5aE/8pKPTUSh0qBoLFadicmF6FISy2TqU871lAaX6tPw60dVGUXl6GqK/
sNnxmEkbpX06zE04PyTSsBNiUuDDeo8nHkccaxXzAhgg1lU31v1tx372TQYX1Gq8vyTvXmVRfaJW
w+Z75Hv2GCwyusquzF2qfykCESO5JHBw6rrWZmKsEsJfoDyGpFEZ7XxETMRyLHG9+cFw6fOt8vho
bwo4HELqKv/zzj8ltta2IWYIongWwdu4AGIIWeRnlFT/zQPeM4PbBKy/xTglZP8tZyUuHsKhlKY7
oFSHTWOnZTxNkKfekzB+tIKvxVcQ32WDn3XlfnjZMVlk1d7RMFYVw3g2By5ZWNbZF7AeK7UutGIW
jANFAkDDtK8pzHeUeSSroMgxDA+R09GMYw72IUmzHU+Rn/Wdsk0Ac1IetEhXNURGDIoHRcqaUklA
R6uivtW2alEbjXidnTMlEqBtBKV2oWwmK1tOq3f3sDsVuacxayXtsHnE919J8BpUeVYH322i0XK7
KPzgMaVK3LEr9USDmV0GyzHFVXZWATPsPjfDoq4/vhYIWJKgnwBPyPFtSx1IVjYBoneXyPo4pKBW
dvDM0GKe1Vezv6tkumEXFhuTKtyr3Nwvz7FWr0npJin6roaoOpyf4GMVQ4vw0ytwQ7BAItiaiH9U
L92VMpU6sUSbIxnIGMvYzp+3W6ecqlgxLrlFzrHLIr7gkMHlOqGUe3j73X/qjRARDJE9y4Xljl6W
4nI3m8x6rFhW5ABKjxXP5D3+7f60TTBy3bS5qEV3YlPJmJ1u5IBCbkYT3xo+38LM17YMgcOVAgOb
D9gMwHwMnQoxPsXYQFbmy85ZR46/8ODx9IO2ZXaXYDdQqHmwt4WWOmOlegjfqIOVYb//lYFA+7gQ
9ao6E8C8YPIWX3RSSYYpi7eSuhcH9wk0SB2PaGJUtdpRgay9OUqOVzRDnTLjGR0t34G2yL4qWL7E
yzIP8iqraUVS23Q/2XAwRIcncDtJWycdyuaw4d2tN7EMIeYgLe2aEJ2FKyPuF7dqpoT/rhvTjlvf
qPym6XHNdeU9SVgPhFcISd2Ryl4lz8ctU0JVyNV/y2gSXSLx9ZjhlqnreA3LrCjUegkJIGqynmWs
goeaYKw34w1PJJvCvn85l+2KPFwpXFP5iETqDAWNwxJ8UCGccUDjLnvn0k9USgyDD64qZv5x+90C
OagPaeVNatuauq5qP889CDkBM4FoYOfcT9HEEBoaqAG7JjpSJ5ME05peqrGvAqkTXmsWROYxWo30
9T7075wNSsixGiv3K+YO4EVH9LKo1cjjh/uTzPywlH8sEvEEEG5M+uVmccSU90oDYwaq11S0qqFR
NjMjsAtW7MYL2e7nxceHtY6RmHypTxw6eVevvobYxlnWX++nhAqv/En541vGcwCvu/t6qDP+2Fbo
DvSIN6PhVSfyWKQf/an2KQb6jXGOm6z1Sy5A0DFCAKGbwZwFl+aFD1C9IJId/mDTXmpGYyquBH+y
ovKP5TPafSFKIR4oYulq4MiNtZ+1WjlVRWkfw/os0kXia+zMgISkLBXj82bhlgAJxye8Lz9JGtKT
CVZeVLBNvdn4dwedjN5WUVNg3qbbgTGw9OLEkAPUHH+NZYlV2T3tzrGQRB1o/on1utB0TgW8192j
Ifc3RcaCmCLUMImJDZgsPNTUPZyNdTtIgq12wQlecQmaqe/EI+VAjpqoTMhSsXBBB2Qx42iW46Jn
4t0H2b7AZNRS7QqxzW4Em7LIeQ4ML/vczA2T/KRDMcnJbmukkH8E/zJP89BqwcFw8YLTI+wJeYDt
4OMLzuvpBBJJihTAbCpI+HWTd7enVANrfnyzZJLqwMmM0uEvWaQBuL7O81uNnJg+SPAgP5AvGls0
tTvYq7osW+gj90tjXjJ3p977oxKRgnl5ARnjGczoFaPaDvHropylIY3PcUWa9CMNIo7rh2QDWybq
N45awNBXLgSUZO4hodk0PXRO8MlQbbjGoerY9kiJgAfpoTk+SRzqR08ILHqPvUQfLC/ran3isl0c
JZNJswDYJw8WAm1GGsbBA+fTazQvgK1Vj4bEQnmoHjSUX3c242ERmLiRyXtTyM0HUS+0x1Xw9tpg
zhqZVVUbKlew+A5j6fd4WN/pc2AggkUfYAVYnsFGylucyUO6DSZblbHNDtBTQfC40GUSzpgjx6UY
GEEnPcH0v/ZoOolnRmla5FPZltCmiEDk9pK5BEpS7MEraM7+x5yyCD9IkeTYiKvwVKydr+ppMhyE
wAKfSNuZlu2g4oxNMfXKv9tsnjP/TOaCyx9p5xoXj4mtI5j1yXvlyE5ByqiSqiM+2py2CI/pJIqn
8XGyJNt1lGkZOdhyAiyFpH6GCmbSuKeX/3uk3vrCvwG7aLNVmIkRTrnHXpT0c2+1TFDBsZ/gsxsV
+lh/xNC1d0JtovQMWc9YeGAwSDAW23Fp1T0ifd93dfxmlUL/upRex2dVzf7gYudfowBhJCpBKPmf
swVESyGcnHDXLZqJQujAyzo9W9LxYRdLpP/Vkh++AfVynaEU7PGJ+J1xSX9z6cj0g7DRTTHAfe5M
9B63qutcSwnBGWl9vIxHoGxxsrD7sig5Z6luGiPdyv/fqcLRg72F1uYtLjCQ5GgtrKanDfrG7dfz
1QNqM8AQbu1Okgx/X0cAUXFvFTckHjcalrDzXCLMMrblnLIbcW/RS5YdICgTS/+aiu2oOUJougAK
YO6rLJrQbcYQHjRaGX5H/1zGkT65NsSs9TqCz4DKy7YJ4uqaORwNxl8JrMHkCvN30JhQm9243kUh
fFQ2pOE0BGLxtVgTFDK+a7Kn76FdtPnb2raZeHXKtj2oXPbo9+rCs8pEfabEYRaC/69drwbPKnsx
sX0jnCZHAMKyuLwnooIxiYDWRqcc1yyCy13jxkXHeEsIsSThO18q+dJHze0BefOI+k7IJ+cd1lm/
p0SQnw1b8fJocWDOM6qF01lqRTCohJtaeST3l+k/zJvsvlX6XhQpsw7zqGvwwp3qMn4HQlspTE4N
IrHDgZRgNsHFAlKEj5t4I5yq/KymepAQjek8NLG6oQnv/LmxlTSkGpsPenlg6zWJdlkeaYACYxX1
eOxW1ehSllIl+Bh++rQcjLTwQdVVCkzOslc4oL71K8fiF06AiQD4W9R05fKifkpCClYkxQ1UIlCX
3K7cEubFbubGSBCS6LsKquy10GpM17xwiMz+xNdzTG3GqGUfSc8ZkOI/uM4fuT8B9xMAi656xYAW
EUY99jVR3eSwFFEimJo7CptFjS6Hi2gRFLBCKo31gM+kvEAjZACtMLa9rxagWO0IW9sYPizlrt1a
sLgYGit4krYHXTnbuEdWys6addf9nHz7M98tj1UtE+lIvCOaX6cWSXSjUHCOwhlzn2xJr50On7ER
q5133AA80M3Ckro4mhql803a30/9K49Gd0DdTvMbxZsT8yQm9OmaGG7a4c1Fxyy2zYPUJaBBkzl2
ziRSylym256r9Hc3SkoY6v44iz+D151vyMl11CGkxGDbEWgjqa48cNpIt/XfeckRjHWV6O7eeNVB
SPkD1A261qTdlDm/4TqVumtJari2olJX9u2oJWHsBN3mm+iIeQjfNZ7MYpbKAZwv2FaloGUiA26C
utn4eBGVllfWZsgehUDKveYK2Elr+5rKmDhAaoilFCTB6Sb63gZ+9E1kwyNpU1H3evqgkT85lYeQ
2XtqFOGlMXj/M1XxqhQwwq+J/+gKOWr5MNC888pNxQDk7+9dgbqunvMiHWrCZygG9OgVYosVDnVf
8I99RGowXeYJ0j4l+Tu3CXhWF3cDctm541zkJlrIKz/ZHwDbD1EdXz6cpTaC6TTXIc1zDoXI4OyU
Ri09mNvZWZzy+8/IIuB83tt8bFXPg90lwJ0QalN3wdfYNcGBJFtl8T/QxXSvxtavncUFnftbz6+M
ZxnPrHN+5OrbuIczUEpyUKbK/WtUtVKKyQj51M/PXBIP0bYlIDDJvv20cQkJK3qaKlGRm6p4v+Bx
ehN+K4+z3OplkdPDsq//TiWSkv+YXercEh36qev8dKu93cgveU9RAXT7Fhbw/07gyVS2WX/kD5wW
Tf7J09G9BmOydlF1aXWxt+Ch2gZ+Dj/lSaApPaDUi0DU+7rl7nrjm5j7fX9n932FPlRhLaHRy4Cj
3NzLZIrmhwYHK/5ld3sAncvSFMY2fQMSMDPScMMTEEut1AsDDjFi7fYYJtD2viylmoijHsCvCuLK
8iSr4MxC7FuQctLIRBUenpfuSpDv3bAr8dbxwPmq0k/so4z+7eGNMDjJMyoBPYQ9qvgxPi7V3Bv0
B/oFiRoD5QsnrVdMYn/ShajsBioAm2IPkzY+KHvLCToZAJEjTnybHegtvqyxrmTO9u7A+0tdztxq
VYQYp/9MSIlc7g4wN/lLAfJxHnUm1JN1t4LtRDqktS9ekOeKvAEuYAb9YnlBKNO0YErTfTwU9A7+
9eJnjYcNUv6b8/j+A5lyKlCwLUON3nbJzFaw9WB9S+jQTovVuuT0zuVvlN/LK4cTr8tilgT/pVYe
1qj0QAAGeNtNHZO3i0HA3YDtCxdyxKK8fngkpjEDC0dGkdh/flLi4lA4u6K+KpQ2sO/PqW19FTT4
YJlNFv/rq/pgxyvyq6RIfnZZoFFG6oblHl1T1bsUxVC37Zf43DjC02kVW9N482eDLeALk7/QePz3
m6wLMAGS1PGGjk4doev+EJ/8ZhBesA1mpmo5rZWWnv+g5Apa/+pzDzzZ4qykKwhs3tVJvvL31VXh
Lq29DD9G1hcNBraS1YrbF80e/UztxTqrBq9ld9qy8Rx8r++pjmrn+lIQIeZ6UEhHRPEDbMmxFsot
u9DZ/UVmOtZTWu1Sd0FIJRIhSu3EkcBUrDZHf+W7p9UACPicS86rVgOHT6Mm4JtRHkB4YNi4MKQe
T7EiZySVgedPDFvp+LCbbxcuOHoIXk0YTaUwNU4I9eiMRFEYlboVbz8PXMvbmgdSUBb6nxaSkIyY
g0Yc3dClp8/qFVCEgQAzXHtJB9SjKSDMMgOKmaaRojgC8agt9t5WqstdME+pDnSA1BSfMrD9R6UO
Pzg4SM1JXWPWfmmD3PclsAReoD8i3KHEf5AmhCSGyLDhzxp6RIvvPqnhF8bsxnwNttxSAb4kdijw
xEcZHhl3iHj/GwUIWSQmAD6XZEafMEniuf73OS9P2++ZbiFH8+sPVrP5o+c84TDkdJDVSf6JSHAA
7bpZ00XdlMwsCBj4W7VDIUWzuX1+gWjFg4mcm5nPQ6OhrCQObWzTeQCCKV8eIxZzxXwRPhc0oDK8
GFbMPFcCVVkPnk7fsdohp1UlTV6huQLTVTXwdEVDM43bpnm+aGHXDlDyxB0UcjQkTw6lqBiuruSy
Z2viUtC6UBhqDvW5fznPS4/MqQMZai+jQkL7ImcijFH4ochXF4KDm/07E4HqA1Dkfws2GgbzXQKO
UnSyox6pJm6FSby1s/AHWmCdLdWatOI3vYiq0ENTjz8FQ8kcKS6WtPfnzqos7EiV40PlTXEVH2ue
6JWFhU6fRAfrBdbCL8T4YtmtS3nJTsmaezH9QRfs6mguarnru5C5k5PfmCsVSxPbKStQc0hJGoYs
VGbca7pt7fBvZzolQ2B2gyGAPbqA16m8w2Xaz1vW4Gkxgzw9vXBR2uSRZs06oBhCJRXVheWyGhzC
TYskUjhVMM8XpunxWD82r2mC/KZGhRo8B7NLpz6AnD00NhQdQKH2Krbcao6ycKnCgsPc100x2YgY
P/++NeqYR7DvfiPQtmn+5ixhqIqBGJYCC2AivvJg4lbQnLesBcz8EOAPq9x29XURVZEiQWeulgVW
FLVgz4ZztGTqxnlNmHLhTdkZDC6NwiJ51emgT5fqx/MuBxLRRee1DK37c1kq1gkkiK6275Dx0sCF
1dwzYktCR7doUjlSYktpPDidAacjibnthvlxBPqdNLGuSsSHenw6EgcIqDOOODB/OoLk5t+nHrwl
si5gtAA2DlvqNGGH39pps+dQHpi/fCbLL7n73O50p6n3YmLkfKSZviRnDk6+TgIY4+DlT25L0Tih
McNMCu6Ic0YzbaSStCi1DGfkcISFRI5zxT7j4UqWS2ZJYFud34pLyiLxpA0y73hAjarC4AGO4lZy
Ea0w+MboUSzIsblUU8H3EXK0/+jWZ+5eoioPpR9D6sxSCrcGQ0cUoP8t50AdLPhgj4K+w4seVapC
fzROckdpBlhmKqxoHDVVhw5LyRcGZ9wYLevuui+wT6W7dEM+4uOJshcRC43+oN2ZKRegZK6PedEg
YrVUs/Ktqv0zcHjaUv8bVwp63+wOEm5dae0xOlSKLBMLQYU/vXpS5uYMJhMxnrbyWnzTip/6j8MD
O1Vzmc7Z8B5A5S+HXMNqutKeBvQS7QHz6+nS5TzR+/ZUAmNfXeWyDwIVBxhGLApfXABJHR3uH0Xm
HpEDH+DIjAvT4R9nP9Y9tLKNkU1XSW6yBJ0MqlSjcu7s1z+CXdwNGUm2oykmRaBlhhSQd2fi+fL3
HKnqELH3xLT/gOGO73raWTSJkCymY/GOnFVMVWqwp1tr2ZOZ4DGymxkNKfoWZ2MRVhQHFEeweeau
rZI3ZhQSogz9gj7ctYiR9H/QVj2BqmuoAWP9bRa+afB+0L4SkNJynXGZs+UmZWykmcPxgCsoJZU0
kCGfwE5+TJRT8HHGtWPPrYtTCpqCPLOP8xaFhNf/m2RPxZSpu6oFW1A9skuXoIL3Ylp5kZOQCpkn
uQX9c2aOugt2OlLliOgGp4W20vk9Ecas0DaWhTIfjDpZxG9T6K4TQdhRUsXUleuwtpfq4mQdN498
jH7+pjEsR3ty2crOsdWxh6FsWMxKzki36nX57C2wLsG0OX25nuO3XS6XnhkK1c7m6DbbU91IrCLt
sxKg8pBkL2dws/ZbmPhCrvI5IlhZeqFPDIsFHDzkm97dlNBXiqi0LHct0Oi3dch2gR5nP/3itOTh
jcCcJ/fteX+IBVNWp3tU+JW1ttZgSU9A17FeW78gKz8NNJ67mjweddhjX2nB30q+pzhb4HU1m7jD
p3H50QOq1JSw39lgSJxrsOMXQrzkBPzes87MBAMOabavAfxbAovW/iOyPJoMVEsvJdizowNG1J94
wiKZK8gfqVpThQgfYEczhD0GZaHA8F4v79ebTNQYJZFAmjt2uBIFSU//NZM2yGUOMNm+Nl9/aDMh
2f0qsp3gwSvfYM+J8ejcGf2Rg9Q1nyANTq7qvjL6nK1UoPsSD1jxSBnieKcXY9PpQe3OUSdIVJR2
oqFEtvmNVmWAKkBlnmVtBROOPS2Ibsbzb8vmOfPdW9j2WIYUpDhXX5DK8+blPV8pDmIhkL0uMZO0
/0WMDe58wTRX2MSirYsWC/kKqYDg+1lPNiHt2AiG+e8eUJsCudyPY8zz3ctZ/8h76fXdEk8dUFNl
am/ovdOPlWX0atFicxCkSMVB0hb4+fvmg35XeMxdiTdOPkweGhdZL7UueGSaxmxwsGCjaTwG5N11
mRXaQcPVEl1YJ+45IXPYoyPX3AS0AR1momSwU8T4CsRZfnuZjwzyjF4BKa0ipbCOXQhQM9hACZv7
VPK3S49bDkYJgF8ydKYm0HWohcy8QB35Y1aeVDqAzpT1o3W1gAtI0kTUw2JlImgW81Qfifxtt//P
Lg6ruePmnd3htmz7VUGCLxDtbnVxqoR755oxQcqp3JYswpNQPxUf9z2lAOXbxB7BXg85Yf85qsKl
isA4C8lC45aczDnnXmy3o6zJU55UMVWcQHVZUAiBRVYlAEYvli7aB2261UEIeVIn3R8swoAXasKA
bztRIGDop/1FSAWDZODfblq7L5Z13paswX6AgbMrgFbQhembjMdYvwD6+urV3Nnmq7yVDsKt4Bch
DXBKT73qSzKnvBN+/40ruBBxbfzHVOKKWeGvF8gBLnv1MBpRXoB0oTvQ2rNKfs2Tdkoy2y80rx+1
zy3+MOAz8u+7oubIphVbIF0wDVTGZwabbjeF4ZjTDheXqlsM+aFYbB8GS/VNF8pe8UnwuwlnpzWq
IZOFLG/P235gg4RmmxUTjO6Ds4uSO7necdDC1SVIRjgjjjZC3xxMMm4RKIf2dZVa6CWol6QWTS2c
V5AhP8nR3AlmI/5eo6qrcQ5djwQZ1DdoOYl2HleqaoOY87kQVk9Hk2+DhSYT6W7USB1V1jCqLZax
G/7JZuI4i2uhQLXpAnLDX5cNovg8p/zOLk95BfpYFHGoeQoojoniMf4JiDePb+d5Olk3P27VXdK+
MrWeTQUuFwlNhii+ob9WaOYT5Q4j1jet1KsGEJJkBjzT+WEqfusLZBaId/Dy2pu9bIG6g1c+FeLR
Kbpb4faJmadWVn/3VEZ45IvMCFOh15iaX99ehX/LB+xlMA8fHWptiQtjt5meC07y8CILHpuEat/L
4UjmcleE1ivBxjpKk2AGrdS/mS3dBDqRQiatc8UJG/W4ZvG04op3GpdF+6A3uCw62vIiSwImLGcX
Cyd0fZkjqy6JGUxLKkiGt5ivVRcqtVf14B9TM2hGcEMCtXoJ1Ys8cnutzo2UkkS8lEkGc1nQKaP8
9izuQYFz4vN/I+2wcwzkm+/5sD3nyg9hNXUYBJT3LzIEKFRgsqd5jQWx9ixVjwlUIerh4uydz+xi
ylM6RQIoZFGe8zIBQqN4/u1N6xTlHp1IAijypjGpMjfzKYX16ubgg7yUEJ7+ilo6l+dBuQQVQ0C6
KlLhFcOEo581iovvLEGD5Tut/Dba0RQ290Or5UP2tnxg2S606ygP1iVOOIxlF5uICzj3wzoRXvwF
RayJq3OVmq695VvfRBgHpL+rzd7zN9QmJbTnUIfaZrwUEyCQdLcVDg6hTC0c0gyzIsSaac+DfPgt
s7DltsKFokP/+AlR4+xbc5057CIZ6UjXIC7ygZLq24d+m6gnft7jzzrEzQaIBlzU8KcgLQHX0XnA
j+YYnNhwPzYgTdElVW57rlcAqpQjrh+MNgLU4ss3uPxY5MPHNtilEw8L+0ZXo/pggSatFnS8w9sI
pV+lZ+k9Bpr8c0jmDHIrs1Ur/s1q8PRz98m47+7Tw8DW8s7T7bzJVqoQdQ7EcONtul+0cTNK8soQ
9hRGuwC983v/PYVAX25yu6XhkG47T9V7fR8Oel4gNsMmOgj0097hqPmQ+flc9NSqkHIyF+9ldTCV
7UYIK7c+/rMzcmbRaKZiOGNoNhZ/kFzJ1XZeBQmXntiTXdymQbCmBs7csaAm+KBeh3tehQB6rWBC
c/mXVeIK494ri4qX1jlWcP1EKzngJoFLl/WHucSNeIJG0nj0Ht8dA3UUrL52gWmvl9FtX0C2OL5B
8GLgQqktANyo1FKBnZ2p6Q615Ew5KeMpa/ClK89O/zTC/WSuCfcwCTXDNxOMXrsnw6W12+Q/Q7nW
a9aEzbH9h/YYn6gon42aKCLHXYgmhQPeKHG460ZN2xyfpA3Oi+q1OXkj0PyDqeCOUFC0aZ/l/mQ1
AB8NMk7qi1sR9+z4R008mgXu0qWDsQ4GQ4jB0i2XomjPYi+tYcPJoyMelPA+DafsdHnqOcfweEuG
0eCeQYwQfaBsxnyUZQ4jaD/wUr/ZNavLqgF2jIDJUbWcTxxC203ciqe3cdEklsjUohgbW5r9zhD2
+zaFffHdc89+iUsF0/uuWaAw8sCB78OZMtNysvnGGTmk/nx6WM6VUlFb51jv/pNl68rUcfn+j1pv
IXCw/9vzG0YO2kKnsotqvL9BhoSwjyfC4rLwSdebeb+aduW/4+IN11NHH1YbIRJlhcxzJZq1wV2O
2DoR7x1f7NJAJia9CR4/XvK6ITqgMlNonr3rYEidWspaeL3wa9ymb2zVgWqedkEiWSu+75hQt3/B
Pm8DF15U3wb4+Fva99tByhqgZth8r1z8Wc9T4LUgnTKCGs78UNB/Q2xkI+IDYa1oqdqK08ozptkz
DhP1TCiVUjfVwbB3boZcO6/jnBhRHKISLySPrKgcx9wiS12vfh+GLA0b9erNnLzUXt3DiUzBz+4Y
fJbD474h+ZD1n/KhKgYs8wmsW5XDEGhhTOYHJs318Tffg5SbTiLoVuRs+4PcDfZK/6FSG0siNNvL
RiyeWVXpNPTqZ3iAxErbngdTzbbBXl0VbSo9KPuF4XSgF1T1OV5L37NzUJT8f7J3F5zx2VKODUT7
HFtT9xEYutUnWvOzZoByVpY8MJ+GFdYWKug1N36jenk2ZcIMxIA3uYA0ob7SHsnbAIEiif9AAHrl
xaqof3yzUdwTx/fnkdATGlj3RuG7Z7gNuDQ1Ek0e+VxskwHDaWH5lZ3jUFE2Hs2e03pvjtTSdZ04
dIv8tDVqz6wA7aYpwM9OF1cqLBHEbCXPjq2Et0Vn5MSRvtt4lXWQPbRKNHGi2baxdAwIYzBn0l83
+hKKl01RYpA4jxKCKHe/s6PKHT6LoCKPwxvEkNiCgx3YTlyKUKEnsrrQf3wlxUIr+PEfdaLlPzq3
BFXsIdv3tJm0jkBHkoRCud88FUrWLB0kZEF1pBgeOlaxgXRc6RwStJCfLO6QUjItFUD2QKdr7MJO
0MUE+FCvfZy28d0g03/UjmYO4ISI1oM75O3uGhCj33CE1Xu/Qmlr/uCnhhBtOd9kBXmATIXWfK9c
oZa4VadHW+yjHs/pWEmK9uXVoFNdzl1FkCDstVuubunnsB0n/h8Am0LTLe4jFWKFmqG4YHlMXr+b
KGQzDrDw4+s3Pt5i77YwGk6Kzkrkxr32j+ALVE7OCw5xfQO4+FJL5HLj4y2mOED1W5bEIsOad25n
5fF6O1JeR08M2tSIukov3IVxtWuKnCx46c3fMhiXEHeS6H3Hz/uX8E97m1FckumKDHebVyBocKkS
BjwgLBqVQGno9ZptMNoHTKMbyNwCjKcYgNDfp9YioSOl+jiBiC/G4gGWPlBkHMkjyGwQGbrRoLTd
+xELUgv2FL4Z5pFE/62++YKC3ipMp1wTMODDGq6qllKjOOhvwl4TG/obPz/KtMSi9tfGAXO/v1Im
/Sa1sEAVzKa1S5yKE4TUmN2ZMVPIG6XBSj3RsCK4ZR9PNgNKJ+VuPI4J5uJlNNQ6q/3vRfgpJVfy
UDI1wr6J0fsLUnhmuuTmKAMQWQdjQ/88bRyVgarL29+YIC2x4Faa2/hEyBhYYZkCTJlgYJWfaIy+
wTPsmtQJHishfjTn1tMyHJ/1rt1NJN/ixNCk71z8QIzpZkRaNScwVRVVIm+K+cdMFOB26gIjUM7w
kaGspiFfhcfeYJWOSxpdrLcrxSQLXPFaOpY5298v+W/VkSDLgrtjRsmlaspQut2210CnCYKi+G8s
HYZgU7VmTyRn2h4KU2ZsxKjlyKG0tNjxetr5hAqiLDAYfxFU7SrrWj3HhExeB+76wHG5AQ9MjVhz
nBg4DIlBFv8ohxJAY4pS/qq0kgZCvz1laRT53+YAmORHJCP+MvZsvynbkHhSOgfljgUtOdfNPMMC
L1X9IjjC8Y7a3BkD3QVFp7N58eGBym+xuHpVdO1dpoIxP/ndMnKkejqjKMSk3Ejf5E3q/WbDyVBj
0kLA/qG7tyN8nIwfX3sjjp1GZkCXnj2Pn55oVSflxrnoId9NoO5Gy/boMBGmWmxELzYAv1+rgPo+
N7MD2pQ3WNhgoiSvHbum0rzP5B13kmdQp4Kv8MG1pDMyHNgITF02vz83X6nwb3GMvNmkXjG7xzvH
QKagdHlELA9Z1qheQ9wFB7IuuvEdRp+hdjNeI4DEGT2e8nyno2CAnelAddFbGIsQACT63n/yhUIH
2a3MHTyVBY82bZJZm2+pM+Q2SQ1E2qXLC1kqtZ7qjWz5FnP4uNIGae2tJ0/2wYCzQwjv+3xP7KCJ
NI8pnS+j+s2jIm8wQFmPoQSFWdromIbKfUVyk6bFW7hPrpR5n0ZER87DiCQEd2VROtxEDqH3JIP+
m5VkXXvK7E58OP0h8kqvKzrM6urZV24rTzAyyM4/ZkmQvx6IbxanHM4m7JBu2UjEIJ1dElbg76n3
iRm/fPWQBXh958IkUOiERmHbwT+qRjD9hUEovrYGsMO+6y5Rhldkys215zbQWml5klGVHdxT34pT
exaw0MOMFHmWQkp9oiYjvttdv7hZvLF5wayLVBDNJ+qj8cMAu3BOfQCydi/tXXiMU58xf5udjzLG
Xerk7DkgUcVjLc1RJ4ic22uJVyCOVJsyS4tkx0gFPsVC3t17u7Xiwvaoowows/aRJy2rR3gJQGhR
x5fgOZoqEr1eGq9lIcrQzuZcxgf/vkG971eR3t4TY1/b5L+Y5pUX1jVwtFVB9l/wZVUBfdWboo1Q
7ATMzrUL75bIBFMY1j/UITPHL5WCTDdDtj/sJ7ddQXxJIiVhua8B4fVHqvb1ELAcHQFEs3ijIV77
UYWMQjcgfZA5cP2DIkSkgExt/eV4qh9LSUW1q0rIf7v78cs0uwdpLeQIZmHeQ0VZyeGvLj2akNNZ
S8KyfzGSM6TLWK6gI6LsgvYmLoD0x5T+Ots8ognzCgLD6/A0Guhvu+VHGgKTvk9rWNNMRAwV/XTl
U442w84Qkr7SH8c5P52OC2kDrv6ljvuCt6FL2J6XNHOB8e5o+b4tINrkYc0G0MsIs/oiQQqGJC5q
tn7D+rPw3dfmjxtMllu3CduRhgMueFwCdM/7YH822pt27gnF0haMO0BFplxDwNHLG1rEcaVwBuhK
bAsQMiJFXtVcvm7w2OVTeqY1YVmJSaWjhthkOV2lxDca+75pUVemR/J+Z61Lxl4ldv2ZsGuLWdIY
f5bLdswT8o1bOILyb4BuOIGcp2eq3c8z7VceRcG/+TvqJ1Ww1adthykbiI62j2kJGiiQJTU5AOqs
KeO5wX2DDczR6lPD8EYJxO9oYAB2+Uj4R4V/6NEuUc3rkzLGYrpcWXOdYJoMFM8zQhrvTD67p4j9
SsW+E/4LTzwJYgVKJbtCZBm0JXFhaPh+aI3dV6aZuZhZDIOV0V34VgMZRrDrOvMxcssec0evqjlW
H9pwI7voCTLkpqS7Kf45n7YlN4tOkUtG+EFnidPgnl5moJAkchkbzqErUcEn5XvKmi2tc/BKKLDe
acuskBDFX4eMVQydny66mpwFOdj6kn80cwYnP2XnphWplgNJ8k+g5DkS0ST9RGy5z6q2nKlLPtoa
Ny1fg4Nml5n8F8NjG+GmWaDr0/H07C3AFbwQKeQr5CHY/XB6qbV9lRXsHyrky/+2I/PVtEQP443n
2HaD8HFPCRKQ2jm03sbLJ8vZJCnYBoLFuPklMMUiRW/z7EkzK3VUeALhGHDm8ObjLAP+i7s8x1Il
n7aljBCS0/TNqJWTXc9ExXm93nsR+6x9RDcLUAudniT6pXDKqBUnA+0qbF3FqHNWUgO0li+uF30d
MXNhJWYYMchw2u500qYhvZPj7/vIjLUGent86FFTrcwwF05QXosxQoOgKffAjzK4x1pNYDp8uSeb
MIBVvLy34Bsr5WnNYVAFqaEpkFhtATyJ/KEXl27Lr92s2AIwFJxwFEsHwgIAaZlA2THY6t0xvpxX
LIx0P2ap0GPeORrU8ILYZa0HSh6tUXsGjAkXn92waAohlHoQPpvXocXMfon6PtVnvZM1i38a38VF
gwDTGtAFfwRofKm+A12ldyagnEofm+hFBfSIShSnJzLhGNx/r9qyfCPfpYOmfCuG2OxDNSC60iy0
RQRbHhnXqo1gv6D7bLN31Y/YP4ohM1fBxGzrloCPHnrr7V4oE3xFu7iMREfHKgNdjejmGjtp3QnW
TwKwqLvJTvZifSmjoL/YnYVOZH84yeF+cOeoCBVtFAbdsPuKtkUo4G8xAtWWKdBaEo/I7KfYGwWo
4vnaqH+z/d5RGhP42YBBH7dNfbSCOV88EDoMdAynDw8C7xVzWPxmHxVT6O5c9ygT0+I3z/GMHpTA
wahZTUVYKzZ2dD/Qun5X3EqtQCRm6jQuU5BFDDmGeJlnaX31R11+WbeMJzjgmxoCwJKiRMU8fQ3v
1lWDsjOYhG1fo6qZrJIyu58OmMPTruX9GcPImqseNPuVF8sLGOylB/uwpi6vq/rtMrzVwl3oLTfC
LWbnOyC0uAIu/2cdh1UQVEevOTA7yvJ3mK9OTO5oq+NrUXuCPRjhXNdV5XqBvR/Yg/A9tXT6FGLO
V3Uox7V5buXcq2hHYAmdM732KiZF0dx6jO0iJ1FGOfw7exCW3zNEzO2XfICgMmLu5az89euRH3Wq
DfpcsLP5L7yyZknqFDcyufGvpNOqcZfSMS7P+tGYanmiwPJPhFhAhN0OnCAjitHPM/PIWmblBg5u
/HyXfQstL+IPlF3sc/+s3DfEHmQ1ahqIIgMV5AHyRZiSuuZGVAJBfpIa2vltlmRIuUNtlCJ2uAna
+R+L/4mO7/Gw0bZV3M3Ditb+Pb/GajmWq+3fqbGoP7pFBcNlYH3xWz99ZqKUCg4+DTas4SdKHHvI
GiYVhpt46yTj1ZFxJrjrfngXMQE1Z8xZN1hs5zPB7dvCyXOeKDLz5JDADZp3ZyRXqHgYwHaVPmfj
z3PUCF02WBeXhIztIAgGU552qrHfkSkEsW0OHGgyC0PCrB2DgDMFzuJaIWFIzIb8lvZqrD2SyB/V
EIw3J+M10RU1eAob4HdBz71tPPYH4AAHpRg4Y7/Ug/A6FqAhmGvz59345ZurJKf/yfipoBPt+ZFI
TwVXKIJE2eeeiqI7nVhfCjUYq1WzzOeYQKZ5rJoU8d2GbQjUd0G1JmMtlvMVdc9reGryikAw9Tdp
4Lxj+Ru5qCsENS++A5l1A2r+UhSKc3DM9d6TRFTzpTrWFFgshf3J8kMAP5ljtgJ7dR2xXjIzoCAa
Wadgb3ftXaTL+6Cx53bMuceQTGlr3bhywAbRZxmNSSiAPxn5ar7whH7jJLnVhW8O/I2eNettJoOy
DfI2eUNgxgKe6RO3L5mPHXFhlakYK6dp6GXQ7kn+6J0rJ/IlQKneffzq8Q4VVRXI/lXQ8HTfniTD
JYV8C+HFBEAHVto9IkwlD1tqN/qwuAOVBCuRlZUs84YxNW56wErHF6AhubdRlZjFMO5BMX0e9YYt
8y2dFhF4wK9Z1/r9nqDqnm4/kcqNU1JzqV5j8KV0FXakj6Blh37Ux5C0IDizGIvugTV+AU0ncofJ
9NZo241WYLlgyRNyjEbDPIba8Zv8Rde3K9CcUM2Q+ML18IYH2heZlshxTHclklXANimcWvdt+Z/z
vpxsimlUcpJIoUx+oHZmdHdAo/+8n6FX2gq9KDx/GZEWdyQr5MuUxkOPHWHhd6WkZfvkm58X9P77
QJlrjna6C6aDdkEArZ6AmyEFUZu9qzxabIGfl0CdhRBmzvTfUdNJw+qvYsc8dcU8HgM3WodFQeWf
QO6JJDxM+dsAzKIipGY+6aueqZZE8xjsXT7xyis/651YwecQJP3Y1fA6W1X/hojrtud1f2kvQR9e
SPN4Vh8thBaJqsLaPYYQW8tnLjUHWiHrhNVmdUMmKX3yyA5L6WcLYAlbh05It4N7miRRn4DYpLW+
XX8YLdPkj9+KuC+xuY353927HCj3avnjdm7i7NSNUbBnWejUl2tErzxTkn2t71d8xw56PUUGZtJi
KoL8+cays7tqCsbQB/0J5jGgwiQltF+sn3EPWtaOzTvqoT2FMJxTDlqJ3Hc99YCKpMsSSFIJLiH3
4q6utLiOVV0qKIQXr09nE3dtAtQO2qvmsm6L2W16lCMBQ3MfcT7mqjFe/9lABIIIO7sC8vhXbTsu
rKK3MLaarJYybGeJ+JaZL93fAgwAggiygtY4X5v2RnGMIvLdt7ZVx/zn6J3AafhETzsyoId0sVml
xX0oeIKfSZI0guTY2CaivIVxk1BQWKhZgtPQHgTuAvEf8d/fN69w0HJJdArSIhVmIAv1chACCCYU
alyeP7f/wiV2qMwPY+aIWuaCbWmg0m32b7anTXJuIRhPmwj8uEBsZKMZhvONnzwU3bRb7DBw2yX9
BUm64jNBsdx/DqWGoX3f4X0XfuGOBuNfHQtSjKCO0XYdSKoyL9uROCtP4sg52hw2zkC4URdnrnbS
i6sZsmRw4cCQWrsD+/ve+kocAQ1bW40rutjwBj5btCXJyyTf+CCLQ5wO9XG4DiXvDQ0M/7HccsqH
tPyt5xYU7a2TZnl01a18OrH0wUVRpMdivKQ/YAHRnqwKVz8DsJQHZf9JFc5a8CqgDhljtSLzBqlr
01NPpjXJ9BEcvxEx9Q5IQ04LxsK/V42IlKtp4N7KvfJlCqHXcnlJ5m7dK+cgmxQ5Blcc0vZ75/OH
gq6sqiHK5TkWOc/mlQzqqzR0zGZ9d+/blfpjsjY+PWHuUHcDu08N4z1aFABn64W0inNt7HyVp66h
mxectcUNqfnPuVNj3PwlUZ3/mP5lJ/0HxlIp9z0F+T0CMqE8rHxNsivEO+uDfd0Y8h3aZJEtM9Yv
OXFFwGSy1roKocyxRnqOa/PYbsPji0Gc2vCWo4N50FnKEu+PebWY01qiC67e0hHsDZsXlFAAOLOo
o5kGrOPvote86JKmeL/uMH7+iRTUT86VBPVrjCQB1MfqW4AwdTCf69ensAw7wOjvXs6yu+wMA7gc
Hvazw7SSIdCQt/G4YC5VNFvEUrEHK1cHoy+sRg+E31A64Ttzya0ovLnw8GoZUoUfHa/+acgdoCFD
lB8dNPR9ITTjP2vO8sUbFCdAk/Dvr65ziUc3CVFElLXROQXdjUywpP/PHTtmPDpbS/n19K2rIvNQ
z7Bg6e9/+CLSKvkVdd7Gg3NfKjD5Ji0tlfNkX2T3KZmZA2coD/JGLi0Sol8Jbek1VgATmermf90B
yfqUbE11kpl8Y1hF3TJXZMjSEPIr3G27gmn1vtk0pfmBxKe3MkXuOMWSStPGt5xiWVUuTgZBBZsp
x3V6HqZR8mGls1MIooCu+7WuX90gacWeSvw8JVNAYpIxg8ml8xC4UOe45O0lcxO4gvmJbwqorkff
TKCZTcW+BUHLlTWXNIudbagbwdcfMCNvQuMkWXh+Djb88Ra7Bngvk/R0Q6mk65L3xrCe+oIGXCyQ
GmRtSwNuu1n35LKbXEtwlp1k8FLth0GyIyCGdPDban1OCFH/MQib2lk7qEI64s/dt0EqtDJdU1Pc
nse/o/fKthbnCK1R0POMG/5AR1kmRPG2UedXdlhpyi/HJkMDfM19UTGnrejneztlNCdI1yJLKWnH
VYe/zA/7woqo4Jx5G+k92QCamFGmvMDbkNhkvuPckqSCglyQ6PR/zff923+mykOApp8poryz9+i8
HG317tomOoSe7tlbL4jnvZJqcSd+U/8+PWa/i8aOMkR6DJBLbClyPkbsbtfS5p1u3EHtLAJZ1R9x
QYxtY0JTVmzGBibUHDQh8+qaYRmZUvJZDPRCXDKmUK5Qw18YepsGxflj5x3FAusz09jIsRqKrSvA
EJ/lwwWwgkfp6nXglFxDESlS15DA6PB+xXBkI6IU1rF6VthPyU/+w7/5kDoHR9t7RH8HzsDTsabG
lCfTXK3zv8vX2xmlYZZbmtALxDTZIDKGeDlUVXmeF0YBcfVnE5yc/f9uTrcz40b7ndRzB4CyIuPA
OkBvj98VYyzswa6/cgrQjPzP/qKexeN1bXAMmW8g1cNzVnUlsTJF1deFQaGnzhuORF0DBlBw7AY9
QysAbY+o7EkyCVM/V0YBpW4Idx2oIR2+S1yQ9IVws+a0WvzQZHNtDF9VhfC/sSxw1/xc7qbVZXNd
QEEptkMjG9Y/SNOOe8VHNeMgVJ1Ci5JWBT2/Uz47SFedYOprwiHRE4GySu3w0HSDC2xrtrIpqNS5
3XJDZVb1KapV3OWPCOLXphs3t2cQWcoVj4S6NjmnkhcSjPes0of9E+CrvJUOikux1n5LBXQBJsIB
s1LGbeaFbJvGrk+s1fjezesfWocVMHLPVZ6ElkRVjDoS6hGqbAWohgxD8NS4weDD00VUDiYEXCpd
aKBsAxnXPdVFHKk0ZNEY5qMSkPQxIpzCg7OIXxI5YvQ+Z7Xeq+mAyqpVREb03lKAsHHjopJwfzfh
hMo+CpkcBCw1jFGUhv3hDKcT6ubl9Sc0TodinvtAuCHkowIK6L79aeNaQEjyToTP26DFc8bpMEut
Qka5P+wO7fD3Yl2hqUwH3rGTtOPif+WTGdZ5bfp5BsDn98RhnhJ3keji5vALPpfHVqje4wSIexML
tuiOmAdpZOFfxhVKSqw3cqS/4D22Dao+JR6GdfmdXFl5r8gLv7Jj3wHM5qsLSPd804owFQnwMmPZ
DOsI/YxVNOxDuvH9026VfQi6Ru4sGHKklkjxdnfU6lDSzsY2jkTKNeXuJeBSlz4qO9UFT3f4m9YJ
mPw1HtMaj3CE3EOe5JATeoiP/ttj1QHp8v5MOI16A/LHP3RLiA+lDM+hWI0VtqTgmxNgM2vi99Gj
VO9xGFoNFXPjKhL0yNqI0C/xAIcZQduynnHpvmkPfHG7I0OL1hjbFXGlFJD5VMtFdw1SK4XWoT/G
wfGkCkPy8d5gQZsmgtbB+GTI26/Zo/GTKzKqp+mwhLl2vFL2q3iC3xgw3tyzEu/OjwAZzuoVvil/
HFmey8LDhU4w0CRiQvXWgtywRhkCMU7IcFxZNkYCN9csmMhkBsnLwTDzs2teTpLGWavS2nkL1vox
VZKWtN66SdafHEh8cBgHfNrYDgbRyiy/E3nmuFLLnttZ/Hq83zuMuqM0CemrerBgWUyqXJemdPgH
NfV+VdQXpFvL6xG2MJaaNBPILiKuJmS+zvSUBJgnghHyFGGi3/r1dZTo/mWlEApZK9k9PdSxhHyz
xxgueMySx8od5BTYcBLsjN9kBUmLty3DKXPwasN3wpYX4xOikDT5ScjGQ+kYmYaV+yYsRTCciz6J
rPXDRq4pVNwtKqf97OJikvCWhaMgYzpTVwCDHchkDfaaURr2DhL3CFPbv4JS6v10lS/I9ixpZFX3
G91fN7mZlKSIN3dFENqbZcjJz6FIQO7XhgffvNf7eE6PxiQV/A0h2E+p5V4uuGe7yw7JnRUnnnV1
pKjxhvoJymDA3zHYX8egxwF7kYZx1ImITzgALM6dvXHGPO4GfQB1eZnEdGP/8/2aLJLtkUKjioPq
jBsCIiuRANjAe8tM1CBo//pK6QZEccxsPF66J6swa+sjT3Cdnl6UPdUnurgEyU2vmm2rCcbTe+Gt
tFD8ewL5m2JfQUCHdHPZ5R3M8gRof6fMMEXFl4qrwQim1zoAfQTaewgKbtrXpvvSFzoPTXx7ubI5
dONvXn2NKjWCTwzwvNg5MFOaQXfpJUDJ8VdlvX1O1HQ/+r1YR1TWNfZdkhsieVQfJTIQrkQqqBYc
3WJQbiq9TQfMstz2hTv9DnIblCXsOaEjlZGpoTRDZOYLHpVFH2FksxXLghSnOLUSJ2NFxrBv5/D5
wo92ZWHXmhE3/jek70SARz5KvLAyBvGLMPcptfBxvNnU65u8v6rzWrjAzu8gLoO2gu268vnMe2hd
SYuJcAPMKKiM90DZpE97ZVUC9v1IppJ/f6hBJIq/vFRs044245NK2v1OxE9f5DchroXGgXvQDtOL
TNCSpvukBHntZG5j7DxJkllLKCgRcYZLXr5Xzmk0s6fz1g14sloRdc8PCoQM6po9JGa+1DGoGyLx
A8CVvrjRyUHiMWirRADRdD349AI7H9tCPz+wzUr+/pAgYXJ/FeevZ11diSvmi2HKVmVo4myfSjHb
uJgw8ooCPKfLlFMYNXgngYHazPhgiqMuyec33+CoA9Fd8Q6eLdqBkCRhBxkVTIu3FTzBW2LzZehW
kb6px2wplWXb6jVsdTUiSDY9OEdSOmyPTh6eAq1oT6C7j+iz0gtFJWGjz84BCluo3sJOkFq4VmrL
hyuSYjtRWRuQdvcQbDlFJ2T5k33tcAVzNMYfLo2n4/uJyVsqI63OCQ9fo/ils7kEvsfvRxyntCAj
ParwXREjd82X74Jfy6P1jlEKAstIRHd+hL/Macr6j6vfBa+pb/fBVMmImFMpNJ/4ECmS3tsPO/BB
ue7H6+ttvk7xEbfJ49gsWaMlPKo9HUD9Rt/+GAaL1ibih2LEYkGzCVJ1fiGDD4NYHRUrVJGpSXyj
t5gGpbytCn56+s386Oj+nzyp31VCNHel7//81lMyGdZbba73VPCSIoXnxM44Oi5yIrZgJq6SkpBF
12B/xOnw9vRJHa1j9Vqe2iIWbOpMetemO6wp3AhOs49dMD4SgFory9ywzlMS7PVaO78Ui58sc59F
iSu40ee9xX53f4wlH3BaFC97Xq/XUig7tNVxhbrE8IYihynw1+5YTRWADU/CzJR5H4nD1H35kNDS
acJ9kU/WZfCZFEXkVPEjVCEYTJAdSihmcdU00SIybFPX01wYPC6dQitmxmPgZg+lCCbhFGtqLCuT
cMmkabv6gOTAB9JqzarCWCeGtgFG+1UkzZN/SJKqsiy62ITtjdFaw0di55Goo7WJx8G37oiYvj90
pjThU8oD5zFpj9eqX/BYs5k+6TsQ7VK/eVhyxkrrLfM6t12jgNPjyFPAQ906GrYDR/yvXSZpJZtz
1ylbeatxDA7vU00CwUPLPiAXlKJoMUbK9XvjDRXjpZ/1dNpw6cjkZVOWS2zMcApX9k22Z1wTVF1/
QeRjuq7y2ZOfhPl7ihJi+ImfzHM3QBQ/9uLGtVZM84wUlxqVdt6m0bF8dXHykymt9tqIyo4p69a5
/vIIkTXUMy/CHsqs38F1u045tDf6YdV/+6tf+mYbwXdB5H3CDdIH5+dkQQ1GSw3qnhZ+Og8Zz4Yd
NK3QszhGVHH/9bhP4w2Zc3PQeygsioqT1o29UEXEUdsHXxMlohyyl7NG0+qAAvhXnp/vWXMXIRw3
IWRON4vhEcOb0uP05Bnl4bAUqKX7iF+Byo78+LWbUp0NyRYIrgY8shF3t3OJyQb0/wdbBN2gOj9S
+2/CduJEakTjXZ50TdlrN4boZoKjWMsO1FFANXZYuzWTlENSwoYY2tuy/mscg890Ym+BqW778ycT
87eInqFdpAZk15bliFH0AgXoVLQH/sCbYOoQr9tb40mvM0ayKoRAyMhoGW2ilyCQkdhd6i0z61w8
wEMsP9QAh/USwqxgbZ8jVK6J2h1k/d8U+5IJCqHK0umeAL6aSTitiepbqjhYqPZnc5KBc38SIUQZ
4SINz3+xyj08k58sCQJJ+s8n9TrOoPn8nXp+oPYLzQeJzrVYmmCtkImXLOOdpanMQhDz4AiteVhn
AG1snYH7EwEL7vTlMwjHL9+HkGptc3I0BXNEY8PvL3jvSnWE6fgT3yRXMrs3/NWcbIA8+7E02bhW
vDe4cKLn2l6jhtLJrGeb795CppgP7w1rMjQVTdKUea8CgoE2Ygg6aAEYDAiJ6RI+Jk70W0+7WCw1
Yg3FYqfxt1C06BnRXVCIynvOaJn3sMKt+Z/P7qQ8+ftYqzlHALbYp/ZLXe5iRJyItAVHs18+AYQy
qKexYlYDyYeHx24VQtetv5Lovr7A8DbybNXw5IKJp7yegdzi9T0u8JpCndNsOtVMypDCAIAcUzEF
f6zmG9oLt+GlLB/1qaWa6OzY21i21WH2hnKBfftDGrLuphP9DM5694YWY/a4B61sZ84Jx/p3KEtg
gTBpvjD3F3toUZQx1vb/9YjbZc6S1e69DBkaai0lSyVhlltHji7/y2yVe81+at2wXK7LsRZTeLUr
1zXeAycqpOZninyMppfeXODLqDQUSQQbEgHwPxMMDqWHBAltQXzGkTg+pEmBjz14AP3Vz/362/Kq
uyUi/zrTHbe2lCtIDF0ydQkp4mOi4AeqjwSHu113tDGI+mkosW1BY1e5lKW/QO0Fp8JOxGyJGmSw
frbuS+/SKh3XrYw7JJsApBvgogewHxBZep/2w/1mtZO8TBqmQLj1IfaAv8ZpYvQfpa8UK4YxbukT
nmfYjzSY1BmDabfYjaitEbuN9OPSRnG49gOpTcIkgPu85JrZPNGngvy3/gUOwUxY1obQ4kJXp5d5
LS6AfUtVVYmzmWhxj45kgrFCSnDI3KeTltzBM95fNMZNFpHdWfGZ1uW6DehkaThfMtOY98r8oetA
r4RWZvs3y+ul60KumIpyRybkju0GQ8zstSM8ols53RlaRuxzg01iVQHATozROI2JYsEEQf77gPzF
MC5b0FYxAvJUUTwBmeGArZt5o4WBA9vvS6ZKoKN7kTlmvFKunyUSs/y2AbHiEagYqQJX8pjOfG7U
DqhUumwU277WymLnVjZVlPe7JQNj9G7u5ZkQ426dM9QPWmmMKu+6zJJNuWdiVbNGIdkv0LXxMgF2
U4405rjBmFtIoqdZFw9/wZpGqrxggyevHYCeLpNvWVX6XDSCJIEUh/lUmuWOReSruN1DsLdId8II
ZutSpM1JSNDBCBZOyOfQrX97k6z/TiGS7U1zQN2Mzg2J2pi1iKAQaMtDSCa2kZFV5msl/HEQfXbE
iX95WIZ14jFM+7cQ4/n5T6qgIEl7zqaaMPybh0kqYQjv805oAsia2CILqJJZE/7G4kFauua3aFnI
7Rq12SomFEQlmgdWtGBWAzbRLFJ77SFfioe6oWAZxGPLKVdoyiDELjsS8uwn2H41urvky50Ce9Gl
QWa7z/piA9GZCHLg4c3EfAUkqqnFMHWlCWEt0lpGQk477bKPquxzrsVe8JTMCVTVEUEfLtRYgliv
kOYJW/OxO5UHvf2eg196CT4SG7RqSBEIXXrxERS3Rwz1QM2qlKcaFkzv6D4geuF6MV/PQzw/5Dq9
GXEjYF/0QsEnHTlezshOxAWiADTM8IEvGptiMqrFt6jicWMOKWv9cISDhOurJdGsoQ0G7cqWaZUp
mgwvznipOpDkwq0uRX1Wk2bOr93hdv8Ro3MDESwjJapnzYG8QhG9w0XxS+rszICbAz6qgY5oIGpK
f/bBvxsWREp/oKUqYdtmaKK9eIz6xzDXGAmuWDdHi0AYwmArwSWzofjugag09bDGelTfztNnktrT
UyxJMEyCubx2mPopMYRL/ckep3Ya37JFfgwabNi39f1gAl8UXJi66bD4tQdD2ToWdBZVtQcQzWj/
NEBS5egR6jCIJ/rSwRPCmx5B6Fgymw+4ig7fJQk2VkI0kFNWHuxQRISh3CMOMB8yj4mSuitOnqVP
yP7jPIWjCC/p5aAwRdgyHl6sRAAuoibgVbSFTVY/4GtfhrqajnhSLurDYPnzmTYqQ8k4DUlOCRCX
+oF2JMx5skP8Tg85n0VBP9z8z7YQyigowS+N+FaK5YR4qwUrJlO5XKoXlJPC+6gwaPh9Vke00EGB
hPwKGxcyqHL2+cGqedRr+iqX++bGmXsA8pPVusDJHwkNmxdFLOiJ43j7vkx5nY9jPcJK2a076g2c
qvAgZu9XoOMzDXF3b4TInS85dZ5444AIFTCJXOFyEm5Z7cFAPTGRaqhhiSRODqXc3yVJ7mOFSW+1
ubASGrJRlRyGGnjqoiJeWzJoUyVY/otyNnVM1kLVhyfHTci5o1sMfxOf8Paf5+56kFsNGQieNN25
yA0itQd21By6QXD37zWOY2ZhraF/l8GpJKibUlE1Q3BvVt54qzq1gAgyZIg1w9X4roMgkXSiQYQv
pJ2+YCpS5+eaubjZ5jfxET7FDAZxejX/cKnwWqVl9Fmfxw44vbU5wlA6zVPq6bGbV1YroW2xxnO2
5KGtZBhd1zO88iLAs0imW3uAYC+6EvH9t3SsyA2G73vfx2H7sA3aGuY3nEd1O/Qdytzq0SwHps9G
pTTk4LFbHG55ltLAppAlmq8iyRB3L2GW6YIzCFpJQDMwrN4+ws2GPq/aAHn7wy0QnzSX/j7jTw7f
NDJUazVnw62L3CK+pGgUqEkkxfAVoi03L2J8QJgrASzs+qearb7rAIPMmULy41mHOJnwhzTzJ38+
8Pc038bSPptX+mt5svk/7861Qle/BCd3QQYpqR+g1DNxbN6G1nTslkSUM919tTZZaRFj8XifQXj1
okZdJ6/d5y46c5NKOJzcSbEffqIy8TZMo4AZ6jYkqdDJPPAJMqJ8YiHJSY02z9ulBe/rrVpO+yMe
0QtCNepcNH7vgjdQGYjUVO7ThbRZwun+q63DpOS15OWeCluggwBJFlM5JQmXN2dyGDZqhSyXQqtU
6q0X30Yt6mvNf90QtxZkcKwjWKPXnVdVaaAkDYAxQVB7nnJNXuiwR93+6885px//3GiCJeqT0YB0
vMwF7z+VSyYvrkmSOlTgv4UFawSccO+G6XMJDN/ndoUULdHXK9ShbD+27YdhQjDWlZ5wu/d6yizP
nAWs6ozn44pYy3mcey1jbCis/lvFXST2t84uWUYPme6kWogEGThEy4ZJqQ6UDTwGljNqzImmfhkO
S4a8EiL/ZwGp4P+QxMle1fhkTE0AG2ih3iDASsQ3LNCL3sYh/tNeGISR2EK86SkaZIai681mKe4z
Z3ceXZ2OxkvSjFi5ApdMzIpPwKcXodnHCV6Ad/MloV9bDciEYVYK8fy4Y9SkDjbx8uXAsu1cLmD0
icI5F9TyoY/k8uz+oy1KIm9bqKUFTMGCqxtDaGN8P73UY2WLCR3ysgB6Ge/QVWcBx+ZxWugR+/r0
6DSVPKTUCZO3P8dtFTaBdUXqRA/sMaa5tJUcb+eyDBFKyBB/LtNugJE+F2/F/kusZB69uLbxIyA3
Ug76FKg7LYsMSicJMg+yetqEbk+g+zaZdZhY7/a1K+rRWUi0IEOuGdimPTG2qC9upp/i29q9YU5h
SXQcnl0jnWeYe/kFzGgKU+6RmEqVo0JeceE0wMU7VjGe7DzBuX1qMuOhSuxW8chnti6popgiqjHF
IGLqB/G6JGdbZPV5+7KmiCLR5euaAh9ilnNEfmUdP9fuFX0ZkTjGIMcSpML6ZUFx9GDiFzhJVbot
2QA71ydx6GtMEHqOQzFlD57flTAD6oVpxBVXW3LamQrpmhhxEvofAlm1IXvrRt9iPvWWx6W27xg2
72fQfORFvMNtnZpDmpxOnJ9ejmhpJAxaKSpAf97lMM4b+niFvDyo/MOz/Boy8Lx0ZLY9NWQgg5If
3kMGG2rpWJAkas2tNXpXp+UckWlvwlfTk9bNeDydyF3L5Nq9nAQrtXygwsu4+NyfrlnSvLaP6GDi
IrlsS8yHwSHWrQkcc4zpahgwakuxoohmo/S5OkNBxYSoADlYl2BTefvUNMFSXnbEBss6Lkqor+T1
mHvGI+ujBcXCof1NmnYE/cfobJoSXRgj5L9Bz9y2b2DEEsc8z1dYDzmZdgD9S9CjF7P79MnWH9Q7
BMiaztkAiFwUumEP2jnEvK2D2JHwG1duBApT41HAiaZtqGgXk29uJ+hPNqa1/YyUA7OjgDCNvWVA
2CAPkzDYzcstNgF/m3jUXsbM0HsriQn9H5k/4dj3hJEpqY03wv39WeDClyHP/GHmCUI8lCkJHPFz
qwjOSdKdeIhyI5RJj/hU/Pu/U9nstB+qpNIF0/iGfBpoUE1EJQNCb96dyvCr7ZGHJA+RJ9SVsX8s
44+G8Cu+dSK6ymodO3628Z0yTrmaL+VdBx8wYylUtfORA/1X0ZtGV9sexhV8H3N1WS0u4WJswb9Q
MgGI/YcnVRLDslQCgr8dzQk4KGSIpRnthApSsDbVDs9FcvhThguNrcrTbFWbBeNarKXPBUTPun/R
AIbken40VFmz/sR9ca5gTbv2KQipQoD09vXnk8DV/+4hU5e5m4co22XgVlxb6s3uL6g+S3fj9oVU
HvpDRX75vnAGfZAnTHapSZnBzOixR52QvC3+j3+LAGvpznOMXYKANncMNqV1qO0DeNxth2zL0qHt
aPwr/MR+oMy1roAzzHAEcU8WGoUimHf5TNkk3rXrt3o8jEmehZ8k0x1KA81fabTAIGEaV++Fd6oC
+qiFwjsL8pfrvZTt6vVQGHbdsemetQn19x9eJf2aVHaDnNh5A+0fAQO1gBJwnm0PRxq5Pm1ILCXQ
+NvEeTfx97RkhHbrLlfFeg+L3g9oe70a5pw/Qxdmi+DSkJJ5NRV7nyaweV5gERaepM5cfmqiILpX
bXT/uDdD0o9HP7inB/eJX79Vfbw0OOSs/rP1Slzz8zPmEqH1NKjXRQQ1cp9MZhHIksXd4+kTOpzw
VflQJyHaeS0g3995CpJL/LHbRwODR9TRTeQv4INckqHgRgBtIWV2SCZup5Zv1ojpREXA0/Q4So2j
V5QgVO/XNV/MjiIMO8rJ+0U+RHr/ji5FjdHTqkiXWNu2kQmbwsH0Qp+knh8ZGwVWfRnEAXjZToty
Yc8kxWcKT+F7cZVuNPFXs7Mkn6B+R32f1HJnGlIE4PHEOeDjeLozvZkA514PC8LIRlBPGFcfuNW0
Ki2s66w05xJND+frnQdyPE1aUGIKZUWYdnKm5sizR4162KX57vz/MtsiB3nc9BYkitQcEe2+sduq
zJTb2xLNX9HUMv3HTeFiB1citlaqAEzL9D+Lhf4o/o5c7S+rCDPq4egE2PYdzcIXUFm09dmwlU7Z
5UyWj/QpXtq/Z+qk14b6CLR9/k2XDQpswyLKnPCb2xK2DHxph1o35/cB9ggu/Ig4nrBFxXn38jKe
4zNFUstypd25T1O6IVaS4qIvngiXrPJzHGJXV8sLCFNnBwdcjTnEKShxZWC4OMvNKsnXNgRxj3Tt
FPH2P3VsQpJ1KlLG6e/VoBCtNRHThiBo8oAL4sVPeE90tR/13ErMuSDELpz3MAlVWxYWLLwFZ+ir
M1jLPdn1tyM/8yMKTwXXXooNPLlUzrpg0yG2s6ymmuXtBFwrsKFlSmhsH8nNK4QNwylkJ0V6ZhAC
OlN8H3nU54yGaRhZheWPhCpN/LH5VEL69DbA9+Y9Lqu/aV9jslCwLMBQ9i6rIFBCgbwIDnmjCRT2
gsA+vDEHBU6w4exM5Xj7D8ET9+ucxZhvAwngOmw52tkydhPl5AT4BvkrW0P+fC1UTTXwW/wEL5C9
UA8ZqZDrps66URhL0ItYUWuUsJsvt5/cmHma4OskpFryby2lN5XFgF3uACcpfzu+MZ4bT94lFdVm
YmkYqbrh6OjRyQTT3zsMIKr15iQmcrp6qL1vYJMaKSwOj7Uw1Vm3UradUxcJ/rIkt8rd51SDraqF
BJ5bqcB3wf6NOo4iAEUNiXeR2BSMCWvrDrDZTRxONgdA1Sr1Ddv+uurSdF2A/I9rBOtR5Bi97qea
yWPTDvzepbV5/aawz0xBYC/58/DZ+Q7dOaAiNWS6Ud5P/gXUlFPTbxNpif+gb/BUD1+71E37OYwG
NBTdQOkw7Is1KLEZ3KhXA+kgicYSsRl7VXo8EAaZaYlvGGZO+r1m4Dlcrr8iPtMhsIanWaIqpnYV
y9ECt+0G42sUDG0JJLxJtFU7SY7XBGnckcLR4xKiYrCrw6j2RpTFaNdbkgIBlTbfxLncSphWy7jG
y9BeMYUGANjj+4s6hCoix/MaUm0wqB7HERhwj6qc2ZSUdqzuDzNWAiUrca1qgejp2d/Ikd4h/5YL
uI8TPBK4NAN96N9Xl4at59GgS//+XBdUwAeQP/Hs8ZDmNrcz/O/kU00J18ymdaPXKpn+EO72iY1n
r4vtAhz/9B+PutZVmsIRXG03Zp/TsHxRQZZm7J2EaqZ5McIzkHs/hReoKBtKesR6UkJmdAI5hyBZ
PuMd9LDvwtfSQHESS1XX5/qvUrREJZy8zynouVsEtVU73OvWbuHgDhfmX3L3q8OpTUkqti2ZBGEo
XHuPjxs6j0XYa30cpWr6VS6Pe4JUVGEFsgfmsiw7d1nOlkwR5m/BeLNdpNd9X/+sFK6yrWJDunml
dcLry/y0gjOYBTAefhiPXd8erLSIeEDlVnYLSj3hsQEW4mHVTvWCiXPyCB/5NJD5akfEqj85xN+r
Oehwx7YlewK2NbmYTy+71Wpz1i/sIcf4icfLwp40tM8j1snVRPw96b3tqfqreWascTvQnltP07HI
ATAY9SbPRRyv0+bPU5322PnZyFWDw5eI19AE8wUQDERvv7kGGhTyw1a1WCRahajHPUHk4BGJAsVk
zdR+SGQnLAh6/M2+9Yp/a4yESGOJBRfKb96zpLTpHnt1Jrlk6+3P8nREAt6J0kPK8V57fBFH/Hci
dQVjpf/PjWN3Yk7fxdOOxv3ItiOQUkArdW+xl9NJiFjlRXLOaYEZCjO5kRLG04DVMBqXbuUy18Kr
oroWeUX9EDRo7pgA/SovWmc9SdsasDZ3xmavoqoippjBNuj6YAy2jFDtHMy9ZO3TXtfZ7i/1JU/6
V7sGyUMq9gPBKrGoDTPnuogwXzEb57TddkIXvxPsFeQ+4kHzvYpCnNdCc4csuz/Z1mW+rpGSpsj5
RO/496j5y5PLjhOh2+RfMrtK0UHTpmuQ6fyMpVyDn/51N5aEpA7B6npeL+y5QOuuvN/LpUp/G7/7
nQlPIyot+h9dfIG+ABV+JFyVqNCjyK6APfMdfaFMBMbGDseEc/87YqrH2/s20kb3JLM8FxqZncG2
yapvmRS5HlSVxyLo3CIaKOMYOm9U/hZUiSsqGIzybTosnLpqhWC7LoeoaWWmMZX1y26l+v+gU6JO
HeG/AQJH2+fIcAkCMPap026xRlBZMV1ferrytLIsKUDAp5RSKF+1U21toZKTjClcQvfS4N3gd3Bf
kR3HCvmlnb4hKpMI0xDCc1iNh9zZLV1gew8SX3FuvdjVN4B/JKPcBbqnd9itSJLCrvwTkQc9anpu
vjmVfuJUR5xb4wZry6U/a73WcZUoVYw3zqNyovrQRe1jZmS8d9bm9A98TjgCc/TkUEHyxVetvTO7
kV8gzr0/G801b+aNIX+GP+k17ZngpEnEnd3LBSklCANm2X1m6tjTk3x9YWC6CGkEfcNb5Vgx9YwR
Rfp19APSmWW805Ee+4u1cBOpiOPzPFvzpvc/OqEi5r44cweYp4WL4rvNnZaoPjTldAeRl2JkFxhM
bKnYVMGCCfWpLfc977//52TbyJ15UCZjyWrOLJuP4aPbt3+/5RzV49Mc+XmyiknBhfTm5/I2HxaN
rkcQUKOZ2FUcPh5Vpl6PRjprVYJG8MB537LncPokxfoceCHdOxzhmwyXAeJXVMmT4MT30Hr0vAQI
r5sk/6a8yyq3qRYUWhvqcubf8CaYbScPgAvpUy5a1kzXfba44IdRdi2dti7xkKQq+ReY0hU+LgBU
pWi+8LnT1isiQI5RBmdSvAP2TJzLkvsd99c0yvZlxR42faHEKFGHBzvzGJDFQvMUC6xABltwPxzX
D7bojchlhzFro2lrDaPSFaJlalLbzDfsspxR1xS4axLXBmd2qwCv1smiMA9ozSvwNZ4B4e4BsIil
r59QMOr3V6L5v/GSi7vMg0ZPpz6AUxQWEiOmcGJk+Z/+kBwneMGrFYEHPWe5YxNDVnI0ho2xAd8e
oTlaA5JZbphwy1kyX5Rm69gP3Tx6RznsFFuKkn91amy87CnSrs2DM0onnCenkA1BFZkeNu2ctT6O
lvUQlryB60xFga4J/cHsOtUMCn4JNxw/ASfALzQX2hsBxAxo6Qlfn+lv/31B1ryblrnYYNbDcQaK
rFnBG2WqdOqYS3V4v9X6vHS57k7+apOTa5HdqSoRpo9qjKITTqP1lHsD2tVMQEwJwfF61PTjlJIX
pVI2GRcG2MjDdjGRudcmmFka3wHfy3Of8XtaQ5/JvbOv0LQiuC2YxnliediIY8itQGdfTelH0r+F
DDlL8OShEDvFn/Li3ODmgZ70RlTnZWdFrneczQwpuu0Q1z6xvo5DwI6unLky4HBFLqujRUafOom0
DgJ9Kt7cPBsojf6yTTmRdOVUfjxWtWKgZOVYhzhtIIvLqSpkcBBc4r1nvzUbLMVpq+E1pBVAYowF
EofrlON0IJDTooTvKmr/hOmdHPsqUcuiN6JZitzg/GDV5kD6Oy6OUmIwQDZxC13glR3ryU8U4HIP
0iSgU4W3h0swX7F9+qmt8KMpktbm8O51d3+G8nNEDhyjWj2rpVa3BZYeC2JvWX4AUyZbRjXZQw/i
5I7HoSDpwxRrAf9dF2xeSDnhNLH3fKf/X1gm5nVx77z9ps3n0j43ki1V8JsUaKzgAk745mhRgcBJ
1Ff9ETLzY4WD45l7P0Xbl2Rn/bSSO3/cj1ESEu46zHl1jC+6C+2ccVZTkdoFv1j13Earbua9Elft
MG2AvUpZPdYuVEhM8tpxkeF+Uvxp6/SzundR4YShWKFDcns3J3n+XExyauVAp0zR/A2mEgVy5RFW
sCCg7Mq3aLJKDMz9nvCD5W5DQQoht4+pfwKbZY151bAV6esHab9nTArh9AiRb71PQoVOd2GjOdA3
S2WbYbMgAHJ8HjiDwSDUuEn2/Nwhyzyb7pBQ0kSxLwWZrLwRtBGdAEPwisX7CMaBQIlQ0SxzgmO6
PoX2EfL0k1hjd+59u9Pj6qNF/+H5EeSSzyFaydAQML34+qc1lT8NxYiPJR7OFaFi70uNRWo+N3ET
XOXFdbgq/0iq4yHTrbTkghu76W3ee2HI4yS+5cWDuFUrXQEK54QD30bZ8xoXKaBTwRjppg0BVllX
t24RmWy47QTgZ5Z8No9IfMj/fXM1tN8Uibz05ZvyEx3gXI5OaHc6fCSlLNTYF/WFqBmjjr7m3auh
OUu/F72s4/rd1P53erWvCCgBoxvaFbqJtOlIHdie4hEEzLyDxQ50IntLnNp9hiBzhAlUDhXN6F38
yYb8hO+ATTvYw0zM4XfK8BBs88SSUPYSXIt0bjto0cPOfuLb0IwKN54bIgNcpx0KHZKqV5TCTqjG
4RqbnhfCA5pk0tEXrCGQZp/ryj2coMUIWIh0bUJ5vtNHTCZV4AAzwZKrIMzOAIt+iSzN7UYOlUsY
GtYaiDIUy/gVR6jCI1cF/CsG4qj3xyjOsVb9dJGSPSDgAg18pL7S2Kls8RXFiC2f7KxKceX2KvZW
ormecSoW8u2M54I//gPCwlbyDXOQerbSXPSp+15pyEdr/aalt2udga/3iHtBcX+6MPwZRDYVmLOG
OGYC6758djN10YZfOocJlHWtKW2pN1jn2lhkF5YTyKI77iqJDlstlR7Haacd379ukP9zrP/YhfU2
0NPvZkkmcPjK7bVgici/pfJ5kv2k3V66CEPRSi0FYg7p92ohgqbjfoky1IJL2jLl3cZ+ZJgIJ7hU
7kAHWWZR6BEtNLvPgsXcQIvkH/1HJpVWYlpWmLLWqtwr3vu4jPQx9fwJKRnYXz2oTB5VUrB+9GsX
K8qPAccKcK1+6ocEzHW7qwd8wiuwE10XsbnANw99rhELmmDQJGJBHrKKvM8zOE9kIXXH58rOgMbx
Q4PAXrLOM76/Z7K4YYRw7nw7dG7SnMSyPMdJ5ArglmPtvCkdas6wr0PkhG/Nep6Jf4YIgMR5usGB
EYFcQAoVLaeV/lKUSK4XPUsGsEtaDMBCZxduzZBqXRPJq/6S/eVb+04e5YtzGxADTQn8+minL1Pg
XpPW9IeIBjHlhZ5tW/VviiCo8WkdaiYNmZXtvITaSU4dLfHdA9PjxjNBVPlPgSRMPaHvWXIl1nZi
dQ6Pgdp4tOEjidG9a3gh0rvyO6XOwR5xoTfAOCwG5mx2f/wYBK8y5PopmYur7O0dbTBRK3IEHkSt
TFs/oZWB4Zt+tejEtBtR5HqLiyiWKidfxP+0ZpfIc494OOvhOeClx6mOigE2P6sZZ4TIxhoGblpr
gpMg6bunL6TysZmizizoght7OIMV0523iqxyeU9sR4utiFLSlyngdwd1aXNto3GLm9+pQOrTrlBc
4AAWDYG79Rlx6LkPRbb7dYR5N6hLfLFR5goaznaf3YCW7F4POVJcg5JxCv89BhvkzeqIdH55WMEP
VIGPEDUaYWK2kAU8aZkPMA2Yfq9P9BKSicBmJLJvBuUh2AkfscGfYTpraTtcxK/ugPsJMjs06VTy
Z4bvQjSjTU39a0vFNDGXNg8yBt5r4Lu5MNUMzrqyYlpiSTcrjoep0nqbA/aURXoZx21iw/dN63Rh
YnhXBzBJMCUpAgwBRmeddLILvtw9zLeFcvtPO1hsNBg1FpoeIbTwLDe3coljuQtCOP2FEdEgsqdL
lY6VbZR1rNuDAEZjonzKJOqo20xyVuqkkpie0edjsk+l3hfJozap/CDGw4NyzLzzn38sfgX1EN87
+cAUszkRe2qaZGKuVjt72pYlR/FqbFlGljPbbTmWaQCUvYSioDxl5/iVKyPkGk6a0Y2ZY/jNpJui
AF787J0JhdMue3z1aJQfTIqkMA8r6l+/HX22+HHkeF86836a8RMI6I0seVCOumrLIfLoL4/SK7EV
ngikSZPbwSuuwzmgwbN1Q9NGG1QxWmsZYl4v/W16Lkl2NBF97VGxQf5Nkd//h2P32xyZp9fPiR2Y
MxrN6l6vzoCjzD7NAwocFf1iINekgN+Pxrqm7+XYYc07RHoQkM1SWLd+hVyTmyCjvHLQaYTgDpUm
HOzEc8r6oz1tmd0GR6pdoa2ZKJsa7RxOz1fTsWbD5X5UpLOafAgKfS9gAtWGOfeNxp8aRtgeEWhz
V8EKFRwTEajIlpWwgJ5gX9fOjKVlOrcVdYiMRBNNZALU7fl0402rtVjTPfw0P+HKeZsORtW3tpDn
Xzqp+4kjYbriBsS3zXMyK5iOfcWEfteRz1R6xhHLjkgi8nqDZjx+7hmQJNNtJMV7Zsgeo7UDYy7K
qRhOy5oqR36Tw7/XVkYo+ZB5E5hGAV8y4zi2oeHRBUX9bb5ZKRzg/Ltwr7Yuy1ObbMN02vEvU9On
HsNeRqzLo65BJTAmeubI6qfOp9wjnKc60FymSGUA9o6Jq59dCvHfpkOH+k8TDDAs02FoqjqugxXY
KLCsir4dTyDdzHhCAFSXF69TNe4WqphONYzGAd1yEuJslHhfTfjUt2AM/TZVyLc02Cq3HNqQ6MN9
uhVE0CtktlUGG3f2WiETIrSGnCdi4f8V4ZYnL3IsFJ2SCSVjXWYuMu0PTvv8TZLj7oKMInul6R+H
N5pBFHhTAnybU8Q0L537BsgzFe/5JSphLUtPjJn/aPpmf/PEWtn2sHAo8tM6aPimjHd84zkwvb43
23/f36xue3Ez++h7P7zC7HWgeFRV3fVXWrrhMWLgXvmXtZufIZW55bLY8NFlLzHvG6BOKkdKLuut
RJrmdrh0puZYhyMVEhgndj4Ac1ba6ILeS2KnWICX8oSLR3H9WFCepQrTbc1DyVjXutBtfAA8zilZ
XIGnIKEd5/v2ZvfFDLDqmqfDRJyLpszlTwdy9U1vV6XLW8Vw2ksoSplSpTXTWsKfSFGUDvgkfMgT
TpLEI+VvcpChuOrT/zFLLkSMp+cQTfPiEpq8AT9TaPiv6xw43DMO04FS1TEcLM+axdE/NCc7ekg+
3DV+uqcMPwEqw7ZcWMBsA3RON2T3s2aNB9lyv0zYs90s6ZRiWnulRY62RzDJOl3fIYcs/CsUqhQK
nmRhDZElEHGb77RH5drDGteNPsTQXTiqP1pE2kfixUS4LJBoK07QV9onpo/ydMYIJdNc8L4JoAx6
tQ+JShQ6222EI/Uw7gyhKeBuh+gfQhbNQZWqYXVXnidkgMfRVqpeATsjtB+LvlShCRA9cscF43U1
X4HiErL0MVZInBpkdd35ujhFC9+WO63LcKomuXBup9ETxot74/FF/BDOXql23K5Ck+UMz1rSVq70
LWZLbATTzRMRiX3dAQxUZvhm1PlT5RlBDhyrxDWYkNb/JbXR8aOGh/z1te4rNneG1XhMJYPlq+M4
UWjF+FyAhgEQxfmV2mK8ky2/MVZN1dnGoSxiF+XJpE/dr9i9udHgLyZDSTD0mNd/fGL8ABjSrg7R
MebeTZGEpLcLs64Avfl4vkVNxT/NVJL+cccDIAoXt78Lt7HTSok83Uz9wFr/HFNLUwtPLBjvpqOG
a0jGh1zn+Busnoqzi0MRJces3h+HxvvuQoAF1fzEs7qkKvM6gRz6c4DSpIkFCnYFWcvgndUxgP96
OJaeNBdQ+FKy9MJcRJ81z56Fx3wOACxNhOlWPIQesbYHj52C+1x4ecRvyQUaBmGauvgRX5qiR8kq
YGvFcQ7JdPAzy+Nnoe5H6YaVSAtKje/M7WQ3NC0Lf5r+zEalL9QQ7nV41rUkSXeO2TC/BdQTLpZE
7ozaXkWYeOdLgbMq1mFp8qs88khsewZ09LGC2hT2qGTgM/6/BqOOmEhqgmuLfKqaWAPOxkX/Kj3R
yjvn3uOUw+Z4Cx27o9t68M17ftmCbtBBro0r1qeqc9C+T1HMsfcTZm5dxV0jZaF/p/5bgaAC1agR
OPdyKy4dUkenMWErtGkKrN8takc/z17faQpO6wDLdxJS07pEF5oJiYVbiwUbKs4F++JqVyFMrSCD
bIbPdvMrErIfCP2d7w/dhd4Pb29eWjqtmWskUohc9Co7Xx+OFy2dvJNDvr8r8zUmS0vwSYxuhd4+
eyEdbJrd1xx4v3TBZSGWWGSTS0ZRE1i+tWrBEWJg/vAILS5XNCwQbKCdqYDBFbyrpX3fC/MmE3y0
pul6fFeOSLGm/UB3s2x2KiaFs3GCKwRqFbKMjAyF0Cq8DJoBjLBYQOCLtpTFkvpHhD6mREEM5H8Q
lPCJARM7Kgy80Jqv8c+NNCwTyd4SSweRxlwE4pGJ4ynlqaXPaJEsuTab1v1HcnNdu5RLaXcD/cnG
w8hRpq7VtdLNuX13qFSaaCacrHfJz+g+nCg6OJdPR50hByiiEujlneyocD8XuOSTcw1zfx8aUSIb
Gi8H1sf3+f1Xs4ALJWo0mR2Y5AGfPwnnbhLrAiu63fU6vKMB7lBpAK12V13r0N1L9KUWbUjfiM9n
z9kUixFddYiBfDWUbWOEjCu5tMDzmVCaW8FpLY2Dz15eUWb7D1RIdKuB749DOCqyWMV2thRuoKOj
r+sNgiY6PHFUmGnYmtRxrts2xjTvVg5qUTv/Wu/hn9q95YluB5ny9hw+gVuv4vCXEy69VydmDSt2
tPobiWWb7mPsZAs8PnUpNhOc4T7J2XuXOwSwiRB0zD1svY6Y2SAWIwSzP+q0HJjNYjXReqmIe8lI
0m4W1szBDI8iRCf8+4O5/nqAbqY0yeJha+jkyP4VAczhfgDbpKsfFnPUAMQQQM6e+F3MngTnJ44z
hiOCNG+HMYy0sHYmPrKAfI3Lu5iEaQAEyjJBLCYNKkMWz1yQjkJSxPsBmNlsuWJwcNCC0sYxKinf
7DzJcPlAWKAtNsIOchfOV1WG/DmSJGXDlbx7/rPurQxFisNCaWwGV/MrYZQijCAd5KS/0qhwjbIb
OoDvFN3aWCtdKmbEZDw20pZPAj6KxKqSv4GuHCOgy42/M1+LTlT/ZADZTDPEE1YgXsRcr0HPNSxT
QKHC7YnHv70Zly2ZR9E/jJdAXoCMZSUvMMZPbKFilqaldKaUnZguQfuOBzgGzI5A4LujUD2yHa83
6AXXL2QEVVG+MELm+emiD1DzLzsW47H+0reRlnvxBFOi9SywP1TaeFNlKtO8H4hYXrqdbU7Ajmz8
qKxPaXseCKtQG8R2R5GtC2bd+FfAE2X5Sx8c0suHdQsK8Lc4p6ayi806wSSAmbfGH0voL1tNn3xR
UPQnHbPBT31HEhL6aJeoq238wefLE5mCknp1iecnRQ7imZOn5t8viG60Bylbpjs263p/FgcR3Htr
PnR0rm1Wp1iTFqo3gSpjJ03LhSncer9Uhh3lDsnIsUi9fTS1DyxIRn2OmISNn9R7akJImhcJebpk
LOy51qHCPdmpiPZNkFZgfLgd69zTUgs8p2h8WTB+lYUl4h3Vbb+LBF5nHqkWROClSQJ/KkkW5173
VGkHWcv8GY/SV6Gbt+bCPjnUQC0GoELHy0+PUTRLzirkOiYx3I3QEjPM6DOgGiVKCrjYzc3jm9tp
8dyd1kbeNaVz+wSu0Fu/0sJn0IRAU+4M2Spk7vTOxNSam37rlOVlZbEm4nqrT3riDZczplZmnYMJ
x5UOX76sS/JGkWunMlpcGV7bFv+ejbomNAR/CTxkvJ50FO/aDOedGmJmRoQ1ClJm9y/1BX1p7sH7
D0RnJFEoSVplDZwZkXU9tPsgpFWHnuf1cEPMXOpj7dxDifAjaUiAusfjNmTRElziFpX7XBFZlCHa
XPXKV6ReKuBKZ0NXbZw2r1tpC/7T3WdtYqWhjBvewH89LDtuq4sSJRbr+Y6POHB8GDfmvKzfES55
emO8YrwHFVxqmiDQR8U/W/bPEDa7Xqrr+oAdt5pTwEuhUs//ri05PDeU/LL2lBgjfGMeRHn5d2gW
8KeL4RJIAjf1CsML67adwBw8Ti292ClhcHLgb1gKhMPYFSPcIkjfqTG0ahPlPGuNtnzJTjybjBRP
t1RBrKa0sX/bTKJFPnWbJKhPUpvHnxZS5H/po33tkRag/249wzYCaYzyHjZzvILJa28yiEfktqur
ylyG12/i1sihGodvVuAtVK457xMkMbOk7Pvcl7Y82H0+aWhJAHtjXPDF7EAFTDQSR+JTmqj+yWQw
HD+Va0xraAH2svCC4CAQ/afOafVC+VvM9P/QbZ4X7/PxVXCs/ou3xNjayXnQ1rVCgqTCt94pawCs
U8ZPlmOidWnKrz/soafehoQH3eDtXJ6YD6lbS083Cfx+HOXeTDd6vY5u6E6M7NrsFh2sLfgYnYGw
Km9Bb5TDH0DZq1kkyTx4RneJHjHSylTMLEBNPO7QiK7IcleHfcUWWbtqP2satN2hLdIQi5tvRwgr
yHc18Al1VXM/KACXvFTcS3uQf2XJskM3M7oKJc5rwnTPlt+7QgtU96ug3dOZemo2JFDJ7mPt03dP
WFBU/jySHsdzFcj86LZ/Ni7dZd5PJXR2wQZS62x7FMGvD0+hp9Fb6yaWX8aYxAQEWTPmdSt5HTZx
+C+csZ9CX1b2/DcdatNQUupiQtAXCQu4dtUP1/09WmmP4fMVDDVa97nr2TvIwSlTUysG6dATVgBX
wEW4yUgo61UOpz8MOgGxuAjJJP3MzmraK0hVgQFEPRdgSyKLtkZ3udU4zFMAUrqSP6K4gLW9kOVE
sUKsvIq0d90oqmou3K3Odiyaaz4I41htbZKXjTV8LUU0lYRR1ZGH4QVvOCy0kFidt42/7TaAr0Bi
yMEJl75FT3UoRKqXG+9POxvtgB8cOWUms0nBQgAvGyjFNBT6dkobPXb09LQTbLDQ6zYv/f9c9SNF
gBRKtQSeP5ugd7Xji4GWnPUFSS7RlBcuemblShfIwXjAftMNK/L3V2GdfT1bt5UXyVNWkXaI0Iqb
jAUHgzQfC23GgEffNU9EIxtugfwA11ym9gs4338zMJgF49NHPAeDTweWb19DzEMs3BvmO/1k7woW
pRJ2PnE9Ispsco5TiDfY+teeqJlHpjjUPL94ed7eMh7ZMDLD3LJIQfUhtbNdLZSyvB3lzafR4RTy
K4621DOK87VyF8MPL+PFRpqJqwEF7qCVB26kLtZ8BZ/adCsTjOXTOB5REyWJ8ZJ5rgV2vWg/Z0kU
HdpshFrX0vBrCIMd/ShmwtMmFmZA4r286XcTwmmv/tl/9S9KrbESjq822rSOKs4NXKHCCjyIw+Vu
e3YtBkuYWf/Hb2nVeEiSlNwy1eSG22EXbUfV491suCY+v0biopvGBTZIzDdR7Y55C2sGw4hBOY5a
n+0XXgt/Gc8c0aj0gTz+JN4w6Z8yWZTx1ATC9k0d5ERcfUXdsCn2w4B7RIllc6GWehyWZChIUjLY
Cfgo+KXB4m0916OUGCkgvZQRDQ7Gmpus7SnT7D7TALYTSA6xsEivfPgkaeneYP+gic8Jcd1BvivU
SCivD+pMIyrdxPvx8qLYDm0rmrdDd/RgAMZtpTQJA3VVqTUWV08z0njrPSJh1S6oNxlAFffbEALG
0EUg+3Hlg+DcZi4nqGD9KciFdR5KP0pcHbSn4oowFnsXRGu/sVIV0RWulktOlq1bklv62mcwcnHi
DlKycBpd1jPa2J9OgxLydfL+6j54GbyQANgYu/sMMkO8k40wthJ/eQ5qMYlb6WvyNRzehmKOlGzz
7QXxFheJEVgOa+BXkRzd5q3uyvG9+uSsQ8FZvpwtu/V1F4HSrbTD8aKP7bZ0bo+tFeAus7psPsAe
mIo0G+Nj6xrQBc4lkiki47XCV/dmS1TVIrNhi1XTyxQ1kNd41203S58IhvauOGEbjNlvyv2YB+oQ
xb3wfkED2hgmmkfsRvGFTxVqemqd4VG1Ko4ARGgGZ1E7qKenaw70aW/qG/ioaWbuhL4BKDbwdIdX
9OBX6wROJP7DZAsPjuiJIUyMAvYIbG/aYSn6a/JFI47+TsDSZt9dyRkz1OoobQwhMuQmmvdtZmJU
MJA6N5l5s5NX/AkWOX2sElvD2HCrah8op+F3RmElGF0BkYzcCKkaKYInjk2pCSJFQ3YwxqSlEGxZ
yE+VbnyW4yj73aurCsah0iTgz6rLs4KBr6D3vFwk/3Je4l/LfZxVTmVa9h7pat++Y23xoD+J1i5d
d60aVp92kgUrw4X7BnldZugceRNKZ6TqMMdWpklbigyggVjbdNk0Ix23mhBuMxOrE00hh1TB+Nkl
iiE4p5s1UzoJLU4F0+kSXu4IgNwchJ1m+DSO9pN604EDbEZ6BvmHoWh/invyA1Ng1ZygHZxYfL+J
CCLBQjbO7Tk5D1aluRgGQqvHvnTk3z6/2356nK2pJCsBZRC3NzXl048YpBgk2kEC4AVQnFA9u/GQ
Cuy8Pht3DPqBihdaiGI9KjprRQ2RPMOLbBpzOA96kTJhzuBKUVs5jXGV4pM9WYd3l89/cqL77hve
iFRhNWKOlp0DBFpA7GChBXDT4ywrz+GaDLzw0UQokY6dwu6a8/ZV2Skw6XJvCND3odVcxuChSgaL
KwhfgRUJHZ/iA6h+uySLrEtabIFzWeKAEi1kq/RWGL3Jd+mEkHYG26uI4cBI+eAM0LA5m7LEcPnF
5GPtNcwe7mVlqTe9XDyS9LwkNKWBHtqC1pimkbRAtZ7tmcle0/H/HFXAoxlxK5pt9/X4yfPjpdFK
h4mRdheS5Nl9F3IgjVEdXLNOowR4XComEz+36bH7BdTy/cyb0Vfti6dy4w1uckm2Mr9CR4oeQvTI
3M4tEaa1wGlw/7FSAoNPgTR9ZLxO6WB20cA3molCr8tj+FPdM/r9BuAkiexnQh8RSXNVFpJk0TWH
eTibYa6AoPdJE/+tYaGDuKPkNHusihiuGlB0c2jijutEjU8gATfKXGexFF69jHQigDiAKaCtdZy0
xxf6HblOF81l2V7vERlHWAegybuomZ68pOz+RxqoE8dbhtKDLw2EZ3q90AUhZ2qg1iCFyOg/Vdpj
uUaeYYZeNjWVBU7YT/y7xE80A3bgyD6uBAeICnEUtOgQsOu6hWVuL+Sxm9LdQq1gvxnN9w74X39B
x1pNERhepJKQGkxbBzKLBJ8xpgAPDBil9F4mLXbzqh+0QLnvBkD2Ez6u91zN6N6vWyZgo2NAAZNU
iIMsar3ZFuvJMjapYXOYzmzqu1ls2hmaS86VYQBbEuRfMU3WaHyOrd33wTjVqKpQrrGZSiXgR11y
tUPw9CkjBtolvsH2+SMVhPuyHaRFaGvaTuoT4L1D9wlZmKhc5IzAE/6LqcpF26Ldw4qCofnTc+jA
/HcdAATXCD97ycLngPtdSsmKzOoE6tPUqStbMNnuyotdqz7h1bt0dSvgRYU9EyFJIX/DMk8QG4Ex
Rwuw+3IVJ3qnPX1DAzQyrTMeDwHYf3OF0QmV0NGBtgvZ00P2m/iLB7j7GB/idLmdrGOLR1Y867Fg
bgODZRU+7irJN/y5Dh/tGRj8anAvz/9VgUMLg/aEnjcDoOFkrwdcyXc0B7PxkW3QS80+l7k+Eudu
5w8HKO0LKkikzf/aEfJEssjrj43ZPX+nu1vV6IobX/joAsH8Nq+F6ovMnm9UcTnWCO5GTinrTpim
WxaIsA5uQnAUVxVwKeEvFtRbn2v0D0Ckdfz/yNFGQY9x8Kru4wiu9+FSvXxKDgGecqTYjBOG59RF
/LqU2twTrfDSDLwUUsG1bpjfxcV/P/Hf1mo+iSG3q3ZCDFdyt8Acy6k4t5bkk/xiaDWkLpISNZRc
f3yDCpMUGmErzueQro5LVSRJ6r/EDIfOpnJ4wFEHaxvICuZW8VH7DzGf34XR/Wq6qJcTfpirXcwA
2fTHQkvpf+GvpV6l7OHf1G0FSEsyvfAdGJiTQpK8mnY3L6eUlZlGR7iTFw0iih0lgrAD1Ut6s3fS
pnmKkIZflj/Xk+mNleK5uSPc4TUqVfWRPq4QKBsAGLW5eUub1DW8Rjw4p5blw7BVKM/sK8qEhw+V
Ea/aUfXHFwNp4bUn/mVuwho6RhUOZOZldzcfpp7C2CaiPRRyUPI2gkqziBnEPzIxvApk+fSyJKR0
h8EqeFtEy7FDvgLvD6NC4MyaVXF0e+rpLqfNjlPX8Sug+yirrQsz7IQhh+2L4oAExo5hfHC23ys7
s/lZmYrzXCylyHazo56A8zj5qoN2zhO5wlcAyjugrrSZiPNyckMsXF0+y2O3qVa5HbnE9S5nrsUy
qNFiu8jRcuXpCa8QsL/WkZaW9kN7Pj/ZBmwFp2NGXc0dmDUZ3hM2bnar4wULzXbFrrKG3/2a6XNy
+InN8OvxsS/3dTBGsXkdziRWMJm63ZEnIYErMtTJnx7KzBqXD33thn0AtBtRCuDghb3EkaowrNKJ
aFl1FgJZ3xKoSUHzJdjT5SHl4Xde8BAx+zY9QXxf9oN88yvODGm8g/JxCYYEV65M49wiZpE6p83M
2upd+kW2mTIjTb0+mINDlHEr5uAD9sD0R31GYqTfvW689OcOHUtc+4/vRCip9YwO/jDGCab4sTJS
q2aS8wPP+DiT3QLTcXt4RTcI7BD+1VRS/T6oRwwtSf4u253PLN0RuJubX/el/Kvodc/tjDvZkty9
W2m2J9Sh5GOeVifp/++1UBmZi29nr7BOeqI7WODUvHPZ2MSPXHmzYj+IyAQKrTLCBwSuegkO2uSn
yW2/g5bzkpoKZsPS9efor5wAXNi7aqiTSZVv9h1OZ55yIsBZOURiptWZy8opEvM4X6MLoDblMcjt
aHr6obrK99CrBkNi891Ur60R13vYgfg9ay9YvFxREciAxC/rT9alupLXwmA33MNkCRZCjgmEfZ4C
mFia1XFSsJIhtarCXXiwHzlp5q8nm2BCCTJDBuTkfdyjFjtec4mj+xyCFzCmWZQK9PWsEhgMLcXF
xwxlj7hVD+R+PZ33e9Y3uxxe3CY1uENUtAqOO756PRz8oqCnzTcoo0oQQ/J1PYTPnhPLS7V0HJdp
9xv1K4e1J+bPpii7tGG18DSqg0UuAHiJRs2t0LAqGQ3vf78+ZV0EiLQ/1xtVop5Y69lHD3rJS9W+
+6FvF4HdEuL18LDdpSTkHcvBrvvoNLTLBXf923EiASLl+lXg7Jx8AKeJVHpyvATr6q3+ITKLkYGT
U7QgUQgu3h090GiDY/pLK9Sodk7Zow1BVcKCJN/m4actF8lJsof0BJfomzBIXp1BLTtniA34zMw0
/EdQmEUVE05nCcYbIrEoHJufAhZsUv6IUa/jWlBQqDL+dXnyIrGIDE1NzZAgPfWdS1f3Yv8Ve5de
E/Hp5cKVM7wiLjT0q/yp6PBY/arE1oO0+129YoCpzEB0vNuEV1cBmBewmPLetx6gzzo6M4TV3xHd
e7jR0GtPktwKs4xoytuPFzjQihMSZJkvXurB0+mU6ss8D5eUH9PMZP21NdXed7hFD/VsaoKPlEXA
ckrgVxXLw0x8fzOSZB6mjs6NUMv4vcpdX1mhlSKIoGlcQd7dx6FqfTGhcK4gThy47HEIsKr78uzR
yai+XBV8pCeF6DcJAzcJ+UEAb7An64DcRmM1VvI2snidOsmTWUFRnf/u3STGPOFRRuBrFncwCbOb
dLqBMSs3o5418mOMp1QbWlWXVcMmF1QNyApG0RmyieFb2PqCUtTTYeukGgTPb5sQRQA4IDG4NFHO
qANYHN3QfZGyR5YZvE0ve03NBCK02SBdr3KPwbjXizkoppCjZQcwrDRReVAufgq/93SHb6a7d4ma
cKFfmqs685Myuhs7yfo2s1XZRozlB9LMk63iGF7NCtMJ/NbKEMUOBIbYNVw/Ic9yg9x0HYynUf3+
sRApC+VN6CxffdMdXtHazTHRn5xIEYuSUixKrqbGvGv/X5+qKPOuFnkICMLInP00qVpQy0z1mQFW
ogc9GXVlNXW0k1gZhVuzyGW/ARQ+8QawGRFDn8IDenVnuLzGmqbMuhKvyP7/H1lV+iaj35KfCUgo
i7Ub3JerlvYVfO6b9C7wPjhbfE9KLytOXQ3RHLTG54I/s22iBHe3MTL/8REw3kESojouNt8Ko6J5
ZDu0HGBREfvx1AvK9XjC2QwlR9VIzA3WltrhInZQ6xFWMS01cSmhCniggF6j1oWKPA+zv7fGGLrl
kvek1cP3cmAwfgkgk7RE131Z9zvSaT64EINS4dD++P02+C5yUt3BEG4gvBt+9rOECPY2TVZdVrCR
BRDC+Mqqsu2PE2rXxG8cx7yfI2gL6QEBqDe31/9gpWb240CFxw6fcnshj2SLvHcd05b8KFqnyi6A
MUKxV5BQ2disr5kJbYoW1DzOGqEDVuFZe7ZI5jbf2hgSF1qXKDQ3Xojp1jsfiqbFLsYoGlPdjIXg
RxF+PNo8vxPqKBh1GQmTFnzxzAdr/14VJb9/YscFuu+9JLg50D18105SdsAQMtSFauq6SbLMe12D
BzkCtsoAlUQFQoupFQ0ETi3NkM4IcHjsMHyahyLlqdoD0HvHDYtwTOeSjl2gyJRbxqUm0I5sroSz
oa2Rr/KBer11BQR2TaVLWfT6aLHUKUUg7K25R6+ldVYXsufyU3Jowi84io0SRfBB5sUKy6LTXwfu
4ht9EB26oWuAgxbzAuRsgHr+78cE1JyQ14M/wrXb0zMPjSe7a2Mg/Xu7GZYq94NZk+0xwRm0fTiu
rBiUlsXaF2GIeheZ0GKnVJk9AihQ2suRYzT2/zBNQWmthvNe830/vL0m+vw4fGOxLNUHM1GBq2vL
URg4pHnnX/FbDKmCm5pQ2U8cE5Xjcx8zv7Z2FyR3Rx1hCpfUZN+td+aq91PIX1gBWb0XjZ3Y5Xlh
249uOgL/QGtQqidebUMrGEjhouxXS4/8tFsamLSzbQqSHPcK8bM1NbtyZclEGPVb4+s79xMmXJ1m
jLBjT+GM34k0dr2WYdKBezfCxngtfOuIk910bkoKo2LzbBbLDZe/PkgJm00Ndq398n5qGtPsY42k
hZvITTrO0Nc/6t8P+oS4qGg0ZXFa/EMqdKwckXC2Tcp5bwBSduVZ6eM3oeqllyksFAWORuPf/X/Y
GdT5jSE8F35ufCObzG32V9DVhXkSdwTb8UXxZ2OuPVEifQjLQRMMeXWeRWDGnswFH8RTadZ6tYuY
0J663gAwBKaiQNYvAIi1hjD4k9fd657Hja3tah4eDM+rM3fKKiR9VX0XQuiyPvyOSXn0uzwIUEgv
08VcQPo98cTgTOooF35yKhaIRrKTtCznhXiMJsud/sPpJsRIa0kU/A/jCiMxvqwi+zDePP2FUAaL
AcuArZSH6Tft6H9ZGDP2Uz11PHaZ+kOfuTV2pHDiwt1Rb14Ve6DKxHTNrs4R91x4Qx6NUNFegcBA
8MIX9gr56DeBE3pRBXhyv93J903ic7FFQOtgFcSQTU4A3Wkmt6aF1dYPG8/Q7avIoMfJHk9gPgpc
wnv+20btnkjt7Tr8wD1DS+NKMSmvaGjKQ+YQSEMQJTAi0Xtq7Qy1U2Ymn9D1G4MGrTqQE+3I6KTd
4JQetGgGPb1qLdC07IMGWupd68DFC5NgvvuveESvcE52RDtF5hZ9veZ39/5bH/a7DbRpo4pb9tIx
HGqSUFD0vVjLWLi/VQs2iA1jKXFUoWZAAIAri+RWJar5j3oQ5jLmIit8UWuc0IEXXkMfe4ADeNNu
ZeYcF8i5D6UtgYXtoFZPxbi50jvY1/ozIdvDLnJyCIxaRmcHlBgfapYDqQ2XMy5RVw5VtCM6sO6o
v3NkoLSlDAmLaO+qMWIvHYrjZNJLf9Li1nP23kMaEJg3fS3oP19WRXOidbgfxxsUyRFreRmY2N1g
79FFZ1SPDq0i29c95ivPh5pYdn0OCxpalHpPlu+idZ520maNL9/EDV3TEJfFc13HgaEGYWVzj9eC
5agIwvspEFsowailwDgVhQyb8w7oXJgg6i6ZxCrWW071OHnfWRgwiI+UZVmtHIXDRB7rgsrcya8N
EamAHlA/xMYt31Y4O87bY+mORkADXWNspk9yT6eQ53FzgNZZubPPLBXhCRXknQwoz8ifcRClXZQK
3CG+9lzmQShf5HIwr7Ht9RItNr6ZvXcd6neMsGgqCU84nl5IXvRIXmdgGQpGLGnbID4i+fbedSFb
AjNoPqIcqsY2cbq6wtqhP09dg67m01km3NA2WThl39zrIQub7bL87FyXzRFd6rLO/XKLkdgwotOE
SSJmArEe+MzGh4jCwdVzG9kYd0QsGfyoR62u9Ao+MXaL8bJXNtqbJ3Z6zS7Q7jR61ROUi7/OQs4h
En0XKVaZXWVc4BaXniS6B701KnOtnPjHtRHzpw6O0WRnLDN0vtBBFQqGst/YwXi0a4hemdh/USvo
CR99UiitDiYNyFMJsLatdedIgs8YFSoite/N00EHDX2j7k97EerjUBQ1AAG5WOo2+5ewE/SZi+S5
M/g465NfjYwOftZxxPconGkxuBnyVy0JETxRvUc7ONM+yUcAEqFanEg4772XUkOfvd37tIqq8lvc
dsUzGn4gD1dFnPSi5dYpMWxyLdr60dO704URLoTxBEtxucP06cniIK+X4nr7mILgDsnhcnd/iI6f
Ddn623RKDhNVQEDjsA2OxJtfDThnWcvfpJIE2XZQg6nmVD4/dAWj+r6AV2GrbjRlIRbvV8mFAEvy
mAu0tzSu0IOgB3u02fe2JWDaTwZIApUbTXxKjMLI2UBN4s9k9WgotHR+157RdHqKl3pIqIDHGpWc
acWlIauJzSbTIsgNYnXZLESJCsUQ3ff1L9B+dYIuX5wn1sboRYBB6zgvhI2+8MCjnOxGd4EteTce
FbKwjo5Yy9KPkLGyGURmeNlTCo+BP+rcp6Ut0kb/+8A0f7gjx72IXCyferpvRJdlkyj/1PmEerxX
/MrOrs6KP+0DzkFV4cT9mN00vAWBVN+JjKyDGygZe6WSAqFbep+BsiwE7YjU/m+5Pciq39l0mRcj
0lgIFjMkG3UX+u9PuSdVhvVUMVPED7bcoDv2GuUnzyxuQxtUjXlt8H+YHvGxMn/Zi3FaSaDixr4r
uZkro0OHN7bVVP4F/Fihq7fAD2xtQLwS+i0gGVaLUCN7O67hraPH3VGHyr5xp1cFQRwUnObAGmOZ
YektkaddedIrC87PU6jQIsM0hqr7dUcfA4xdLarvbf5sK8Q/EGlH+X/tQJvAvfN6bgwp0TkAIUSm
E/iG5BXPDKsYGb4hwhsnB8olK6X5gXyZ9kZ7aKmycD1ZtZDeSr98LdooF06Go/vBxG8/VJz76JmR
VoVBnSCuBfr6xWxeNTGAVyU8AWtnxxt4aMsQUf87E3a4+jC0QqjsEHb7c2Uk/wT2TIEyGDk4M22n
APm2HtOD8sNPFIJPzNnx41qs6YorR14zGfI4h/dD6IS+qjVBjVB5fFimBetf/JrzCsoywohsx31S
wJ9WgszLXZiqcUPQal60SPoZ/YhZ4hstq4tOtNnPknIlikP2THh4IhMnw9V0KPGn1N8jwAgQP+Pc
ecOI90zZsE8bIP9iuGs9kVNG/QllCNNJr0YYFuFV6fDWliD5lrWW2ln0qDGjJaOB2MR8TfQPkB9s
S1LQe0IiFv7/O/nNAklvJHMul017H0qn3GPhnCxUBMenss3vJkJHDBopsA9G7NSODxnElh//ewer
DLYBHAzivYephIGRBMoY9SrPsC2pEJ6Ks1DVL/r6SpefOlrYc/eG7g2cZ08OAihPZXcdqoaSOUuT
qVR1qs6cWZzaUZjRP3CpZy+QwhXPIQXIVqHjEBgSe9KW5FVuLlnHkeZkDg2GRiMdxcQ90xHkdF2O
0Q7bzKKEUllut5PhHrzdCVtG/cTGWWCO1wk0SFXd0ot/IpwVZmJfE67C2yVbI689Gi6g3c/47/PN
1F6Tt7SPuNqw5cosjInG2duYAZD4qahfHVEBhYWrrBPwG+QSe4Mcu8TJzhUlOlUVfjj9rz75QGAd
V2T0/jokazXsnZOAFK4IPtk1BnC0badcrWy0DoOJoRCIxlICNOHW3F3AzFoDGX4KFD2Kjxd3gE/s
/JeHWqi6b9y0Y0FD58503wMJmPLAFU5UzGf60sshf0YAKA675guldVH7OTrtwvRU47fctcSZzujz
WPF05SD1sDjaexxGe62M1C2VatMoc8LZsGTRWfLH063O+8pjbA5gI8xT8Vs/hF1XipjuH/E8vEyX
VJSIxqtGgtAxab1bS4w4Vq+7sdis6US62GfQzJRCM1eTvhIhfzgsBA19l6Vx78Fx7kDNJUVF+kUZ
its7WSXHNsij1JqsmrQJwtFUNrVJwZ92yk2cR5cgnpTs9dJ9GLuhA+gkSVTW2lW1LMgIOK1UxFBL
xjeI4cYR07UIdDmYYiU87TCkcqVP2qNbz9BCDxJL56wyLid9+Y7pw/Ywt7kBTx1DMDBY/xbdt6Qm
bo2cSYlAUsKPWOL+MA4OFgSL7J4wiIs14S5f4dlVDInMApEyI5lXIulSQbibKeTVSPA0vgYMS4uA
F+90+R9bHfbUmfffiG1wtw0TU5+I9vbjOvqAvlbKhL1/4RnJsuWPAIxM0Y4m/rNuUWo6wyPpNnWh
V25VanhBZDulfJ16s+uSYlZlI2gkSpWBBEgmnvIrEFb4+9Nhz11cJuYQAodE+Km0cvarIhteRyHL
Pxdl6KsGeIYhUW+o7s4pd+eU4RD+9I3K6TYHIXpXNAhtoDf8QZDQIeQrDLtcBjfs+pq1+eqmHlxf
d2fllknXpDTuqglPpv4xldibG0j1CmPH6kDWpeJK6Rjo8ONTf5L8KXaJIcCjt1uFxmksFiPNO7Gk
e9/eEPvWsxoDPQrVqze01zFEKd7WGSrNHcJ0bWJiOi4yPxYKtBZblXxY4oJBRyfv20jKqF4DHTIj
rYDKAXC49gS/gRwmfj1cPs9otuy8R6pHfVnLJx9Rkx+wT7EQaazTv9TLWLdaLMlVBrBWB+UWWohm
osPu/4qnp8S587dnJPb0aGke+0wk3WN37+kaqnOx/etDED1mpbm65VXNXYRuvZntb+K2OLfmABny
BqET7ZCt+gxEjksuEtV0+GqOv2DPohPgK/9RsPrx/ehvJB+ZQ33EZ8wLPHBf9+rwfARSBqOKH4wo
rcmzR1j5pKg35tn7GxBqzk9357Iorke33TyuEu6PFSmQezNOGF+6MJkP90JsJouIR+ae/jLA1xO6
k+xIY9ZHRmCQOqG9cku0yg4WO8YUUvPyxcTR0zpOajIbOMLtH64BDVQAi0wQjUbZ3TOcNQFSGK77
pl4kJRf0jmI7WZGU1PoNWLEolX9yZI0QK65ihWYQz6ejxAoOiFPTO02NTbwBvLRyRnEE8KEsde8e
EJuuz0bdCdRFyiBaX7gGW+B9ZXNNbeYQFONU3Wn5SM5LlpV/wObpTWbeMhguIKCGlxJbA30tXbj2
6gmkF9tRGtyyKGSdvWKW6ADAC/VhkH9YEULd9Ko1w6WRtbnbMjEINheE5kRE5GekKC3QeQigpmD0
byhRjL/MSI54frcVBADqccLYhmbMnTyBr1LsqZmZX5zPBP8MEex5YCeslfwF/yEsDxxSkRoQgPvi
blQ9EuA1RebVhYmz/NCIw6DvU5Y5NyLmd3yZV4wA7NRrRe5TuTENtl5gB2F6lTV6R2w+QaMUeTPn
j0ClUo1bkv7OehqHGxY0wnO1TYI0G2XynMk+5xjTCb4b0sD7DxyoqGiaquqAgi6Po6EmzSweCaiX
1rPWf0ZcDxTrJoi0j1hQ9kd8xIPU/LmO6nvxyHUsPnVNd8cBpwJSly0By/U6NiwrWz5i0omKRZu8
/CD6Hh1YE6GfqS7r7N1fIe8rTzO0CLLdFpBGhIYaV/4tmBqgiaGqQX5Fpc9pp6En0Xc+TZGcx5ST
+v0zJ8wPO803Gm0H6QTmCq2iCed+Mrj0/DnWqUcgt8R8t+9AHxN5i3SS7OUJz0lIKTZvz8y12SbS
Umyympv15RqPp1hLG3vyDNbZ2LrlDSIYFG0Sd+nBZ2FP3whQOCa5KbGOVRivAImI2zOFxKotq7Iz
OEN5WhiPM+16omGdDadB5Nl7A8+izcZaV3QEdTVHrTta1fEnYUhgcpDNeGqbxonfFJxWwuibhhUf
QjadzRSaI3DtKIu/EXWgtfjjFvmw8aANIdM2o17eLluOw0UYhw443fkZcDxjNXKqejUP5v5/w8Ug
8AFZ89ZVQxErREp90P9lheMKVt825L0UgDXvYDdYRLqBB3GM/iewE3zFe18OEYIav3quXgoxD9nf
QnF2ZJL/3VKVUDj8Kj8skDkPvzL+ahu0fjhV+V35ucqsoF5hCrV6ysIEvRE3vPYz7li89XHHjeZe
8z3IPlBycjZTY43l5wHuQE1GzJfgarEV+4DVlurBx/NJ/p0lIaVPpqkoQWkYmaCA+zluJ//zp56u
3/OcF0fbhj5KEGWA2jOgauSNvP/QW8x29VFXuqTglFt3crfD62dRcDtsb8goXhZGiX7zaBKCKF+V
7ykvdf/9gYYATsXHxeaCj6o2hLBjZFPw1NuwyUN/3KNu2P3v5E8JpRdMk48Hk7XJ81LFUow7jJTu
jB8yyJpcPGEPG88Dc2GnuipYQgw5VolzHQsJkp60nG4Erlz79cCzZ8Wvrzqx0h9HQEF6mbyppy28
PbKnL4HnXW9CH5OWrd1HKIKXMNuCNNWcgdyih0dmKYIcrpACHaiZFl3tHym19QDV155PB3Nza0kB
to8B/iA9tvCmdyPhYsMTbCcY+EksmhcExtW3DFtAa57smK5d78Gp8lBMgTjUVOHO9H2JUxhIx9E6
865Rso3EVM7g4xPaYdSQNfxZsRmja7gJo32IARx7WFZGr4sJYnclnJh1ut0iL5BX+90uyMQJ6NYr
qt+URMfWC6ESpuT99G+Ld1rv4tZCQnqid+DcbyJS5TZi5DOMRtZMqEor+HGmJSpDgGbSUgvJShNc
7PNR5TDKmrXtPgnUOX6+lSQbOCbxGgl8v2J1ASGK+gn1Kg3qUqBLrYKSo9toqAU3tGtlyLH4AYDq
4bwdr5CVtv6cqJKVFXYCKBFQXDt6SLXChWLoZpiH5n4OnJLEF+m2KcFKFay5l2LbMiTss8uzsXHD
Pjo8hQXgqEdNCPlT0Dolq9BtC41lPucEdFgp9VaklLnlfUQ22/bJIjBAhXlYbauo1M+s5XaySEs2
2QHtHWp6S5GRHOd/2Ay9gjyQ2wnQwh/WqxIIjirTluy5AoGbrdD5WgalWgpw986aTV/Mj5WWIxNW
tv2BT/KXpinJRlC6z9GUFGnAayZbf+ACjDFyOHP5ca75wvukW4vmV4E+CfbW8zGHMobcbEuQnuGl
YYnUiQO4sWx0WA3r/TP9qcrxRkEpNOiGetwRLNGVFy2kM4HYgRQSgVL88JSbh5KLrZ7WU5D4o2Zm
FKHgzv0sdw7AI+XVUkYp0BRP7UW9iKC8ulWyGeNHH3ZiUdZqvHE6j9nn5fOOQPU9azaEAXoySYfb
k5Kjrd3wI28eCcyJprhjTuHfhlkGO46ssuv+S/uCywXno/vXZI1f4LllUA/3De9jJCc2Fh1JHJUj
uVrS+qdGFt8a8noXNJhY7kgqeMFX3Mu4RmPJZSwqIufU/fcbRmeC3F6U5NK/dJ/0/DZG2lT51WAc
f0ZQ68m7Qdw93+lIjdSjuk49zOIGsbvCBlH3S0ZVQFwgeCiHAkFALshsP3i8RaZkJqjbqkgbcAPk
SCj6/qT/GtpSEWhijKtLA4PNuYh5vmcDFjLSMPoX3PmVa5keYlxrcHmv9WFtbLN7JL7SEs7wtAhz
k0yyU2hloHIWCmc8DVBtBTqk1af0JCIcnl9T099laFwiIuN/s48vpoaJ+nKbGIbY+CY1XQRg/MLl
sHgE/ezH72s7T7kJvKqeHCZF2NnYj9lGqGhc9AMVmuHKhqICoArE/iJHFmro9RbVXoH4oFbEsKFl
d8aCfd+LYZ2DuMhuQG/fyuqkDe3HFn2Z30DulhY6K0fxpmKR42mvN//doMMPe+so28tGRFKKee75
1kX2yFtFa1wOIA/QG+N6MUhNUYufMK3Hg01bFDUsiodGw2MvvGLPCi3v3Pzxx1+ASQL/fW5Hz070
nAUPUtINu6UNoCeZL1SEndeu2eLmQIHKHkQATbyen9WBDCJ9COmng4cxIT9WdaMyG4vddVPE4xRe
nAICyn2Yn/kO+Hb/ny9mR/9iVatHVCRP679RxRuDcqOnRBDkR+9Lcvs/vI83l/G3YDrrcLbeMbIv
XeD3G3IFf3Ru2zIp9yhGXOXan2/oeDLGD5LmpG5quf2ZzqLwToLaT5b2hSFnHTLkIQ81ZJy87Ny/
PuV5Gf520T3l+IcwDZ+hRxflyiRNPhFt/7NXK6ndLJMC+uFfZT7C3GmSA9AcH2iRFCM/dogOSNzH
N4rpJ55gOUlx0qbPpc/oM85+cXgsaJsmruA68/MfEz0b3FddV5bA8nZDR5I/chXI/GH2PgVeHvvV
umsxCDZklwwxocWqXIImKqIXcIEBdB/6uh7pv8XVyzP1IRcj6rEWQg/xCBfo6kTeghZizWX7osTR
8L7W6ewk8fs7i5i69tZ2loSb+lmqt/ma31ePxnlrduSrPQrfnSGPnXAxnguC7K0xxuzx87zgntcX
CfRR4myChRAO8DpU3PA10YD3r/0pco3MbFLHC/9I9szKqNmB4TlFbDRiYSiXLHoxKG8qcBEOS2zb
vA+kApriXDGBuyfAfz3HsG3yD9WP0HRVyzktAY95WL7z+AidAbBplCPrknUqfcMNsgv1twFX8MOo
vai/UywIHZe/A9+OBCq+0DPxgQz3Binf3tJDzyEa4Cs72ZvY3fgtBaTeiNNyUIQhMUYljP4kHNJM
y53dAzXBIQ7SYvHtzIzLz0ie/8VKq1y8nwzHNzyirQzEI8lJ7zAWqPp9fL6mYTkz+uAQ2MhMjfJy
jNId3DkH4mHCpxbg31c0fuMqEJUgZOQDK5V6LnOsUJs/iEZ2amwkg7otvPGy4PCBW4xk3YmgFHkR
AiqIDDAwea9FCohp1fJcrfWviVl/dSgxkDCPCVkLRWodYjRGWjn7Xen68ztokacNZmF22qZwnJSx
+3ZXQITB/vlxdNYiGYfk/l2n80aljfADJPHgI3jAc1qIC/KcCRlCELhYL14GUEE1L5A661/mWYY2
3FighMvT3lFxCDmquxC4cJlHlNcpFvD1Kw9+8rdrwVsBhUCejCKtAHHfb+JbgBjW0WImthh+6/UP
qg0MjXI3/a0w3Q812IkXx3hVs9/vW5NNAlA70iBgRQ6YZ+3C91f3SAeh7+KSFbAsIwsaQ0E0/Dzi
zG+c8q4agpWO0h6ENOLtYoHujTlC0WS6wgzOzffPMTBFccpoZpHsi3hgBzcF46t1uyEMoB4CYhHq
vndYhUoSogpKYv3FoSSHCvDQdEVbkDR3AM52VTFj/g8A5IrZ/U/yRUmeRXZgWT9z77yOTeI0uFDa
IHyg5ql9c+FPaYUn0zrNHjopCEUi3gUK/BBHDoWJvoXkq6aDsjwvlOuwosobbc4D+dPKDXnpSCjJ
VR3zfETLGIU//VhAnMHOEdlemOJE3q2DZkZaccL2LXNhyfj2BGOqMmrDWC6MqYBJqkEZTRB9cCc0
kZ5ph8Jn7OMKh0CIwmz62hjllgn1yHdWGehyAXI1dGpGxzmOg6VEeU5a7AcC70bRIIuuv7p9LGzS
Rlk5hB9L02fr0frRdFSdfHnKaJYOiN3g+zjcyuVoS7jZLt2QZ4L+eaElIEVLsgfF2u54MxWRZWC9
uLWIMBz2EWO1yq4IG8qTCr1ce3DFA+GbCNhX3TZcFFuO1QdEm+cd+emLHANPlGT38hkdFdDcgM39
juncGbD4U0mTq/ENf1RcgciyqE2pE7UMX0rUbjYxDsdHcf5IuZmKAvF/juRHe86Nz2+6xrjKGlPF
VIn6+QQBIFFtztK49PUDnUzd8D/X3dOH3qCfgmENiKSFHbFAUQE1NuGtBX7Z3shx4wEorUZ/0pB1
cOFxnNbkhK4m2Wu583l0HxVO6/QOFTnBjROgbmPc+MfMNy78q8qAf2iZC8kqLpF1lXaSdzuYyhob
qPNlHR8LSzAl6WP1+4M/QgbKIcpDow2MkyU3rOB9mFFhxgU5yTQ93BBuu7BHO3q6EBdw90TuNLhk
zF0tU+Z0dAVwtQKPgAqtAx8j2MC4FoNStPc7uipt8es2ILo+YxvNCVw4TTKCi9VwmsVu1WihGCHT
qd/Zx0ylalMnr92SEIKPt/Ro9+4KP5DePn7Rejj1tdjsq3vt+tP1swhvpuLY21mc2KuZXR990NOe
Ha1V1fhn0WHoYkixZXsX2Xb/tLOz2V/kgu8w0MMZ8cGYxxyapIIz2UrLIM43dkmAnBCUdzRLNA9Y
avWXp3ABoupO0fgubAlIYSLhRtfpsyzbbbRzfghtEAEP6pSecNYyOg0LXXyEVWchXrHRLfRy7UM4
eb53NvzuEZOFQ9r5WjOaf/S1XRWywSX6fYkXMqXbVZm1uSgt9FtGtPmpvoGakF8idGQoUutK2K3s
0iwsajCUa77w7smgXvF4P58hmci0C3bXfNlEd/MR9aQmuLIcKwSDZNjsMRIvGb/fq4+p69CV1/yu
Wf9ym8fTs7h9F2WocQ7NVPHecYppatUtPsvhflsWAeaTUYz0/X1azFuUdy60uLbggAeIi+CtzCLi
fGawN78/ETamn2Ei1AJGc+8Brq20tla0dA6qINf72e8WBQOhtX6A3I/ntPhCvx4xgsYCpVTCXOOK
vO+5CGPtvXv9xLYifgmE0bve/1jtSvlzCnbw+6svwQdrYCCGjmYdTlU1cqPcS8Sri8IrDiTXWFSZ
4qIMAmrW6XUKOaej+SZloMK5yUbWid+cNz+3UaRoZuey4njEwuf/jqOoTTKqlUZTa2hgJPKk86Ch
kgVMYbbhINt74wmCZ4keqmdtMCQDIyWujV/jxIOHN6w3ou8B/6vusvHYW1NepDntpB1/XbRpQXIc
VUVTj2LwzTUCHsOPbv+cssFqPcqN1va0fkrvaTEIi8xVtAvMTv55jz7KVcIl5atyA+CjnIhK3rXH
x6maixJ6tR4FCcb9aCD1qQZG+iS0EcpL+IpT6kd5v327AVROVDFE6ilePXcVddWnqxAujsqQe49n
P4r04nd2Cad9eTR0ixyMhNVo6HNm6cqkNiiMyFm+dOfkNTRWE+Srg1JeDWAmJ5NshH1lZrAbjCZw
CGq0HPfIjvWWx9TpyJYwIQEanOo/dRte6iMUmsi51Yg60+GM3NTGHeO57rcU1orzP9PH2n06y9F0
n+ntAsXv+P6oKLIaCYY0eD81ATQX1dbubfanXPxMzjv3gPWLxG1j1aQtO3QqFNUDExpqlRU+he5c
r9S2kDSnjAVForz/v1xepXLvdP0MDOauiQSYXvRz6wu5Uiw3+jZilDDVzyEsK/S9NB6V4RWbR0Xf
sooEUcuoaRkSBHsGRoI+/IO4DCGUX11dbK3O0QK3s698AG3upqVL2kIu5QVRy/MWZJ1KGUFEZ4kM
Jy2n9pAbk/Fg0wZF4ILUzPOmNSPsfJNgv/MekRKyBqRVsXVnbU+tyWvZg8fMjKmHzxB+VnC6I/xX
F1gVUARtC3JCC5/CJRgYADxQkNBlSbNHlgAlXv75aZ7c10nXhvUuIARTAYppm90UMaadPSnEiYdU
WCW4ebofgK1O47h03JoXdaGZoJ9zeiyPVuDoqZ4gddjXg5qlZSGFjnTSyKdKZiskmM2UDGOA+Wru
9lRRjydj5zR61lyExOiEFFIKdyQ6oQKBO4n9XV8tx6yYD/wbKE4taTszW6Ov9FCJnC1xk07v0SAe
6eeePixUoLvJjG4gFvfWC32wvPb03DcmnQAKjDf9hi6t8tXdOkQ7gMFHxO+nS0DFUz8xRspDzDhZ
Kw8z+oGglYrKjJ3yAGyOInBL7dzTsDR613WV+SWx+7hkIO8hvJTYPEkEskb3lbFyryi2qFWvQUir
QGMCPQ6BmCh0XzxR5z2WHTFQT8Ug7DE249eNm9kMMAHzbNXz2GALqgl0P8OxxmXnmcp1+aADHmKE
8vAdldJsaPjYW+1f61p62+z3dKJfjxtY3SjtJ3LtkaTSsIT1UZ/7MTp+lONY2RABQ9R3HTXSYI84
ewotmlI77XSWh5rzglJGrFFajbd+SZIm8y5dtHT3qakBr1tq7uab05zgndIlb/N6Tei++fGWip6H
oo+YKqidnRgQG62TAko3l0rfFvBt0EzLNG3Kq41nCYNzywI75XsXDFIaacKGS4GuWU7GsYhsJnak
+ddONGrHeuw62zWkDraQRU9aS/qvITdr5IFb3eUyG22djXnfq2xaMKn7dj6DuYC5mjhqzJAPkucY
4a8vQJMyTQl2OxKqMFPsjEYlNZOYW6777G4t0W0K6UcAnnKY2zliizySD9zD1oThIS9HSROLnOSW
BMgOvUPgeNFYWXj+hjDXEIwMxvvWYWQ55LG7AG7DgwVUwcqKhP0eP3276s8E6PkQPaFmRdS9lIQs
SKe6DXlPhZAHakfqJzO8WdiigRyUyFsddXGWc4eY1QRcBUQ/+vBzYIQa7zCj9O//RK7e8A5sUZ8B
XphwYTHQETCdGI4mNLoGPUaPi+G8AiwdHLgwmL9yrYaMvlTFEoo3r4VYZ5C5xDd/umF++A5puvOQ
rui0maEWYx/8R4wlGSfZNLl1b7cZyavPvjLf0KaOdtgritzMGsTCUyT1E26k9CV8sTlJjJF4gHU+
G2qK2V9NGYJJukIzHhSL7xwDlQsqOwcCO7VJkgdoit26zabtDkwNoDabSMcvB1IfQzqX4gSAAq1S
TFaCXEXUUL94zz34UPznvPX3Pvx6IOPLxwRLS78ZaeFC8uNWNLPYonqSFExLdbyJQs9WE0YmjqBD
OePJikYyfNDpBY7Y+lAcUq3mquai9pKYI4xALTOaiY/TfGSPuhD66YXskY6BIYx+O0tvAjdh9IqK
HJw1sp0OUazrF0NFolieblbwXm7XNuCxhlXMfAiASiXplA/epcaMIOQOjI4hSeWeJvyIvehzS/FJ
KaikAvYog2gtCTHL+AD+Plv7+o2ZfNMhve4amwUYx5WdPIs2Sx5VS6nnDwp57T7KwycTXbqDjdVi
UCx0KF5qWpUTHO8HSxEjIZvaVELWTE44QeedNEX0RtjeewdaT/eRWThmHYtRwlOJ01mwxw5xLQFO
BRnQgM8mZCOw7v2xpzucHTKLEQfl5F66bKZmR6hboqJLNxOKjztLOASpWBQaSyj0k2g9u9uZsNx6
c212rbwOIw4ElX7qgSrV5IZqKHbgyAsUnkrXK7J5DPqx4R3EXbksAWQzvirVjbp7TMa4hr5giLYy
1wUGnKnhDMK5Dz/IyzAGpe4PVWA/SC2h9RvF6HG5MKmpG8FpNX8jH9ymP2LqqZe8iIVmvkTR6wUe
Rd6FvoOsHtlTP2oU6Hs9vJ1VwoagcEQLVk8hvPBB6EouttwZ/61w4PaZIUkdr0U+xBiBWN+lk3GT
Oz46CvAD0E1xHMajhs5Igug3Vv0Q/VM0HIcO0g95gVpHsQavdEy5aj1kI+tyBDqTt9vwjLIbD5qZ
QEYjoID+JL1sZujNP0wRVmh1zkR0/Wi4YPiT+IkQzLwuYDdlrRAdpyaPOb3etE0kKK+bCjdNeVtE
7zIZsJZzRCOBfcALHHWkWCcNtS1a3QjR18DsiX3W/LAIFTkXtUuR6E+7ESnjqI+inOpXzdKjViLu
lER1CqSEtUjMpKqOICgm564DqlX2fJCfdOfii/180HUEVaf6smmLkUsjNhWp8uM10hTCAsUo3/1x
BJDc+Vdw3d8FHaudn8qFprGBfc4HK416Et7ThdTlaCjx4TDzN3BTAflAA7X/+IZ4Gr63AXtbLBC5
nFXcAXE5YzxTonW3K64vblkbX8g2yLhjU07DP4wPmXg2IsX52JopXqzavl40hyeAtR/GKFG9SgSN
EKnzHBeyCwhceH7IDfQtbmP2lsPhDVxkuS6EdrqCJ7CZhnKaLwEa3YYoMzBYJzy/K+iwgwMzX5oi
8+bSUB9qvy5sRlIRj7EvM84sR68vRAchAIbm5ARhgfhsygfbyQWQnGK/3BR05oqG97TXuW4TLqld
hpGbZPlLIJa78oH6QTGUlJbvN+kigU11r8nX1GpWMSZOcjZXZAlBAh3f/oR4VKGrE6JiDNvyce9p
v1qiunSJuKm69ngonkdZMbNIa/xUj4629i0IPBwxEC4DeF4YDvuns3l975iS4yolDTqrn9y8EOuA
Arj1RFQDiTROVAFKRwEDSEqnY7rI45G0FNt85klwFNOv460wzdty0uz/V2XSnAfFgNoEdt569BLv
KNxnLe/rfEeg3uBmi1Got1yiCy7slupyh3EpvdE+P6SAY4+HzqnztbNH0dAAsVvp6w6K5FNc9uhF
8bcXdDvBU9pKbnvMN3DOYkBkHst0xRyzmYCQnEW+VzNny1bzIglS8kQEDCSykZ0mzzHwTua+QzDT
gYcVY0U5JKGGFpoctsvLimPIdCIgUBUh+j/L36lDcOYsdzjQ0YEd7XTXeZpH8ctKy/CdPWp/lVEN
+LEJgFfSBcLG3kdr4cyQJTk0rzB/EZm/yDsPzsFulj18VzuZrTtKPix+AVZyOGqfxF9X1xWnO8A/
ewdS6Pf5o4smSA639Kn3hbHDFKs5u0u3FMtCDk86clETsaUAPxTwXuKvvAqxpMXv0YG8R4znnEpg
MZfG17rbOhNUW/KA/aWgdoKwbdZXU9otMgbjwx1jN9roIJrCIlWNA48Wdd3JhzFqUGsr3xzE5e+8
3Bgs4H2In6wBM8ueICmMTVedOyXl3pfOm/5guyiFhSDqBXIj8KAK8YPb5I1crghoXVmdWxlLlh2W
nxCfNleCJDx7x8fSRxXsJEkH9i2Zs4BVJ2heB0WTc0+zcsT4Hky6z4M8IGF39FTUpRjRUhEpmGzJ
6j+uN/2uEnz9lOZDz+8QSjVDTah9h6kgitFhhME03yMUh86wptxVHmOHFsLYPQ6JMQ2bb9kz5USd
hkEuhAV+DJh3aRc7UjyBZOkHAOjX3HdyadwV4GQQHPoemYm6ya9sezTqnLoqnfe2bkPvxx/MOMG5
QvyNveuFWWP+Sq+BlkZ1S4Rlq0pagSp9/BdxY5/r0OrIvQY4W58BW0i5lmitQct5FMZmBNyXPFKS
lPKpgV3NtxicV51SU3c6Fqope5+Jl4K6odinisXb/ysuPuZUBE4xJ7GcFdSencMMUGAxeBXQbeiI
xdgTGb2eUZdiccAWnLAoL9i6vkILE6bHKY7gJb6OMhVFfo1Aw7hk6SiROzMN6XyCNUU5xVRZz2OV
BOBvEDP3s0jM9vVM2T6zGQUqYa6iVvaSvqMD4kVPkS/BTir4k+KX/v/RXmXj1dt8bf6Mh9pPY9tA
9wPy5PDYiJFyKrCd3pQp/fNfHhlgBg6HscWf+gjE0pQU+rKkEnCVOEPEyN4JF7cE/3oeAPgokrRl
mxeqJokDLB1LkeAlueC3Gou5ikfGWyxioOeIO7CqLFn7YebAHjxzMGzt5tR9WPcVnI31ZrM1+POS
SmHcVCwRI7uUQq+GjytUyFy3uy65B+7Ib3zC1zh+p9dtfgF24mpHcQi1huNnCuiWBvU/v8KWrYvm
D824VTZhWFGiyC0kefXXKC5mUppdRKsYRcdJbIVo/Tdfj/n8gHugIlCmC0gAfJiG7aslspBCpwbE
SQOaTkX/u4YrJ7noep191pqZ8ul6SQFiORsknOpUIwWKf2AQd2X/evT4MRbbOdxxfF9b6HqhraE3
50imEmo/0O/5aboKDF2KWZ18WZcnJwmd8aHL2hVbpjVK2hjoU4+UDRuWqlpg6R5mIuDcdvQHo4jG
P9ppSD9mrwCbR50FzDY8fFt0RPqd8WX22dHDTXNqolJ3cYdul7UBi06npRW8oJppzTXfeCXindOc
2q1mNfaguaWJeR60N/rB5yfm1FF6v9R94p2iIjMwoK8pea/ORaQ+jjWrUZ8unEeFOZ4pHtIkdZ1x
rwNKr8cb1pIjhJHVyR1k7reP9JWP/ahzzp+Bk2pLzimpD2rReEpL8UIOmZqMwzWufG3GU5H73aTF
eixP1Fxfh5o0b8ErZndU1U/ADBxrWHhTV65PAeURdRk0uhWQvsMwHiw47OVSVxqQJw4hyYjV6hNi
hDF2NSje0SHA+V0WUlAPhTvj1fy9Jy/cG2nT4s0CKq+zdLB6eGK058vIIhhD5r7XjnGzesJUAhSF
cogHhR24wMNqJiJanFLvGObicwupHbwwgVi8nuiRmVTv9e75iljdNIS31G/A14ED6qpG9lAlo+sy
xwDBaHgMFQchy6CAGfHVyM3rkof9TJw/hYowANNbpMknR4i6i3LvKKKEcURlN+oONnUinWNN2l9b
R/nF1Ht2VgYdfF4omDZc2b0UCAGbHsW+NKNcoeWXA+9YDKSNcONJ6xcvvbnaCyIM+jNLqg1NBCIe
u4HcFGFKBT8aHA1lU8urYtiFtrBts8CxsH7aIRNIkwUwn5uV1R693FU26vcRnshyDYwdPZQqgroa
zpYOHq3UlH8k1z5McgC8oabeswcFS4xYLei5mf+9qUsgzLLc0sVD1q6t22i0oK9or+6SekhQ247b
rEE76VqgF8jzNq8ZU99uDdofL3V8O0z1v/7TUZ+L0BqGhQa/ElOixOMXAjCSPyac5IUg8gMnq45K
xxdN/rd3HBBy8WcN9zblcPwedPJ0hMbhe/FPAIOgp4MqvwIQL8gQsLoNidVrm8M+FQ7coTw3Q7AX
3PhYI4A+e/aae+ODcNZ+Fi7IGlOZ5RtPtr1Byd8WgfOa+ZK6sTU2+imHYQrKP/4+LlaFyumc0ChY
3GnKUTAnc1btp5VNCB5CZUxXNoyr5w1aAJ1fYyQ7cFWmW3HvnHF6jD1LxWviweV/C7QzEq/hure7
MYGyDpO7Bh/ZpXx9OpUckoY1ilhQI0XxsY4RfQa/EjU1WLwwpRnmY+snyznqDOgnlLRuq3CVLjrI
yy58H6AoqIGcDimkPg5QI2Mj8YUW+PdIh6e06bZeTwea8Z0oXX3PmXiDYu4PMp8L63vDCNBtAueq
Sxk3zU5IDsGzDQQd040uishZuwPSsQ45T+JTzLfDFuD3SrE0h0SYTwrUzwQf97MDmKtTi2S3ygrw
zz6UPPdGebl2R65IafSUnwQMTCZe01hH3zr54UofXIIBiBU3dyD5ze5rhQMQOU96+iX8rZpMg39N
QeFQks6kIU70ThlFU5h5Ta+vyo7Bt9vrK7uYuDWN+6FLf2nDojB8yUnbO1Yet1wiH71WbNWkWKt+
CdcIHU0a+x+ue7sXNJeoKOWI6zAa7V4CDRsdfvhnAp/IYjE8Dq7Q5txd7EQeAQA+/uJ+Hb/Mko7d
B+peuoQTwOWFiR7LWEoogczoeRcGnhyJm7SfMBjDyd6tJR9xyDRTmWMOThQM37kY1Niv+EESNl+U
bhKUtUKE4vW/pW85Tuxl2wqTT5ax9/ACXJ6Sc0iUbl2G76GnKLrYrpnCOGJJM98eQCkPFZBuFVYA
9nDLz0RZZD8nqPJn6UflcCISwug79A/mryIu/jdJnX/YbGBZStQVh9vuO0vitZNg6/bPc4JVpvh/
GJPrnDl4P8lINV/cPne7wC1Hmn/rvlGurxZ953ktHKPdV6aEi98mynEmeLIsZ9lihyuEbV8vxy56
TgzbplHwLRcYOKBxfRZAjBHH6KrwtfT2HcmVBZyPgYyuMYFBPFME9CEdtLLL2Bk8tDddoQDz9J48
18HqUjifbSS/pIX9N3vUNWqErkriTPEEtM6NJdMGFS7h2ZSx39JtrU6zpwneVkddqWtFm9J8sWnu
ywNYTEfn8S27a6tdFCF0i6VKknJtiasEq3oRgVTGoeODGv8AsEsOnm0+1q8jdUnbYyw55TEOB7M8
bNXM2OwmUx/xs/Z5cZZuIEhF0lYcuwn87faHTz6NhLyW3fL+sCLjIwuj9zX3SIPq1f9fmXeG6t7s
BU9HuGZd/qgi0t2ZT+9dUk2UWr+1aXiIN1hdBIC/jku68YeZnMbBlYukwXpoGxHQSum9UhMTG87N
lrUW+7HIAdQx0AqpnVmM7AdVZLeymZr5RL25WnPfxsIelJ4+x20+gH6v/zb0WaJFlKLG7t0lnufH
N1AtSsqgLxxuNJVTY5Sb8+9u3mup1kHdKgRKLF1vDXCzCy6q4eMIiknmO65UPUCAVQuiH/SC/znK
MZi2pKHwK2nRAn/IfSO2sLgp/lWSo6xDgnhzWxK2xNPx0uz6HxETCvxE7GzqbRSwoTzxsgWyb5c/
djI7Xjs3S4BFNk5TG0Y2klY6hQL/nTuygKdqSg0n1kAq7LPufoNzDFmdX18GkdI4Mpr0njNOCcyC
Jwd744qUyAy8v7ERHuXZhXRmHZ+8SYbih7QqmD6TgicZkWGZUsKmCN9TE/BUwkxrMf54NERIyKqA
hY5ZMAI1ZXjQZWzf6bpiU335IJmrxwtOQCoMjAAxlQGAQHYrGro0RjiEjz2uN6gkG1wLn6rJNlDy
PPoYWtuEpyvN29v3HpSfzxyh6PvipOWtV4U4xNUINIJkt25W7WgeqSzZpeCcS6UUDFcE0vFNcQ0G
g2/l6NCE+wJ3HJZnljtwucusXNZcp319T83PUaqPUHjq3m9oNE6jQky2N/Ab6UfMONnR8Eu1bqLJ
s+w/PufePWKy8jYm5Q13h0pbkdbhKmND9wQP6hjxkzH291C/sMjKWf4zxqrzzkX2tM4NxcEQYv0a
XdFnGgyxs5BD7yBPxxnqp9E6Ti/zKrNcPJQ33inAtgh74JhRoPyTql6f6jNvVBIlXYcoafR5gV1/
yARu89yvTQSy/+e1bxbyZiX69tZTfBlLDu79PWirrwppmq17MtFyGBlytJ6IPbscx+/3OK5yPgiW
2G6tiBqikrDFR9dniktid49TeSDqgzHuInsb2J2C7WyvR9iKf8yQhY5n+l54PF2sLKsWidbpjepm
CsrcdbROj2GbgEy1P19NYO0upmOXUW3ZPWbSM31cFAxrvhfFeaSR+Vzw5HTNYZu2YoDFwKXrh1Xs
hJPvBJJS9SkvxE/mIjJTB6l6CRZQmoZz5xa0l5SeR9hvtpowLG/du21z7QYfCLO5tx6YmzRn2xs/
mO+QSFfU8GDH1pe+mBWK3LudtneHDgQJ3smw7TyAP+3b8YDsOvU7kMLRYjD1txSYC8t9Ub3n/cUQ
XskBhGEiItYL4D4Brkiqma9ssu9jJd534JKiZRH7xvQgLxKjpoYQJ1c0zcCjFMGjw1cSuCFJcSn4
VG/sD7RZtP+0j+Kku5vF7jAYdRhZbaCR8/wsswp9BDS1Ju++/GBrtmB7neZIUua3i5fLQDDoSlo0
Us+DAnXivSVtXG6g/q9Fu1iYgUK0fo3Nn7teXkC/+VNopUHLrl+YCFWu5fQNWOiswafIoQkIUY79
JU88fzICLDbvgbwCpvFGJKGURFvLi6bo/cNs5e0AHorW48buLHpNzvXK4/Qv0GCHWSeKmKoVwRuk
5Dgx1Noyr1ENVJMBp3miNeo1RqH44zMRoJgSpyK/oIOWgv+i6k+L5Qn5gdVJ6ECO1kJwV5po6g70
jwIvtjth7kcprcT1ZD8b9xl7R/ZBrKHAL3U1cWPaVMOfCgZK0Vjj0ZJzQqYoyRFOHNGoV626SKKV
Z8iKg0/gBbU7Tgk6V9mznP3TvgPmb7BDVUMRaPa04bYm+obml/wC4BjPMKyL4Y24cPdTkLNCYPC0
bkGEm14VkxlXFSf8Eez0xGAcJ+7TSwcqOvSyYxU4/DZ10piQvTQ44fYg0OLj1A5+tQ2t6JXp5Fyk
37llsAPwW29Hjvp7a7Q9kA4aU4RzLCWxgEaCu969FFY6TuwF+XmYXDEluEIIM6LS85G78U+NxDLx
x5zfMXAxrlzCgOeXoPBYNoAhvwifO3WQBQOidHVn8XzMBgxVbxVDNu0k5yi5CTKefyE6BbZJA7KV
gfrpkow9l/yX/2qngpw1mvSYrF6NCS1flqFhtdyN9zm5I9yHmW8HORm71FZ+gL5tIIlKqnXDsi7n
WfrtcHlhmd/IS/1pD3uE8W5P+w1zwYtkkCml1meJw1mpmFQsY6KEkL0wKLz3u+G+fSOuVlwWZnIT
mglSLYnfPcMPHrdT9M9xKtwNxJQ0v/oZpI0PXIyprFkD/ARym0AR/QeP01fp73b8atdcC1wPM1kw
YEvolRp1Uz7PjvvIKBFUlu1YNq6EZyJJ5hD3ZXTOtje6oKKz4iPKy4duaCHt8bl6hJizQWo9Py0u
hnxfY6O5DAtRksdRNLPmN80nAtH2IB87MQ8jZvqybiiANnsT/Q7u7XMxHpLVl4EgREIwrTW28I6W
C1VVcMXUA0re//L14Re5o/CfwOfC8mRDakmknp4mkgZeRVnjaxuFrGCUHNRRZXp+W9zIgUvKim/S
3GUhJRBKI3TU5mJAVTirv+fX5KIzQVk9F9Yhix3SPGwzqzEsrBOCkq8+eeKTMyXVfaB92htgh9k9
c2ec06j82BYjKQwceUg+UjIKtobpAHhd4KJVNoZpamDqMY0Wxqls4Wc7TzLSWkhnyMxPYZFjcM5o
UJm8cuc2T8Ba5UOF4LZemjJxzE20BMzUMkFl2KolbTs/RNhtJz/avN7WqXrRGenEO39+0dQqv8Xa
+iL2uPtsh5Qq/DJzT4qJdsZ0UIC9lsu47CKK1/mzdZ/g3NiA+lXqTNxbttQZ9CR891fMszJGC2Lu
qGJZOezTdB7Bd+msOqf/2Io4ZpYl2fiPWgYGwgr5TwHS57PzbnAYj1XC6PTdE68F9xbjddSzCIuD
dv6ZJorqGpN/HiRyxC2QgcmdoH4tRuCvyNTl5Y3igKUqa3SJ3wcgsSQou7h77fZORxkaSZm1fqW6
aMH1UNt/GdFuj1tfXNKVkxbbi3e2oIK0EUcsTd2at/KgNZugIJfpC2KjE0bHh39pD3HNoo8fFJpQ
MvnB9IK0GBjDswBvHd7tg7v9RPNV1ZiCGV3kisMDtf5Sk6Cw2o+cJYs1cCSuC7VtLfom8CH6b92T
bnATxuQvDJLNRFxgWrIpmY9HaWz4pYB1LImqtpZV2A3QCVRkLwTMkWEi5wSIfhoDm/+NYkQT/PIz
7iCOaJbnE65RwN2eKvzkB61TKnlQ87Tk+URYDUVMquS93guTOUrazEmFgyFxMG/43DtYOc5cn2n0
dlOH7oTlfn72/t0Sb9U2GdqTiDri5VKTvSSGARx3IOu7QQpt6VnPjTxgoIwQnSEiMAjxg0ViV3me
wtrJC9zCL/CCRe+NLQLnGFBmvOtxLYVjoiU0XIyDkwuzzYnI7Va90QlYfNcHRwj4+7A8SBtt/bzh
t2P+jlHczowU0zMq86sfjIxlq88/1voUCuR6ybKYfbQMxzx/NhWWmMutP4GvMmXdmu9jYtT97ORS
J+Y18UW/6btRqpv7ic7gaXtryuqxI1xXk+upEtJ8/1cXwFpe9DA+emwerLqqvzkLjCp2v5f6X6ny
yb9/+zqu3ZmdwqUsQLalzYCZtzhOCDcIdBTah0G9sMUZivfyKfyEpNQOvoWOMnD4nLPMRJMjM8xp
v8o7iU4Nkihy+kSYS171Xkm0xs0+nQ+ZKYHJaF9agkcD6BiSwyEiX2N/rlC2ZwgVuF8zhJDnCvdR
Z3+5RMen0y9h5bVl6YZVuh0C2P/V9+4KRnpuKdwSCQ04J0rZkkqfVKX6be512L2RdKWWJCihz//F
+KBwpx8APjLEgUryQkK+H3rEeZRnkLOKFfca3u2xQG4VFrI6yTl/ETMwPnhC9hsiyxlJ9hzl+rtx
uspMXdRJnpxowdROK+et1yho/mQrfAVcDh+Fu1bN/VAsjbvwTdTCTaYKS5hdAO0xvomJMi8KuYI5
ByR5WOg6ImjQWvnhpD7a7pkdHSPIADvlKLFz5MvEolNcudM2F5i4JXhXS3p3vfSXTaGnFjrtOPCa
dxl+BiAiY5DsFZ4dCiOu9yel7sKUb1eXPEqkfSWuGSWwuvm0fkrv8TMeHRzzjDRJGubPs6wSkMJV
j6GceXrjxwKUpdGeYC6HNopg4N5XbNz0WVTVNNx6oBt5coIZ1q0F3y9hx33RS1HKwc9hGdSeDGBP
lNvCqLfXuR6nrfKv2QonASh55bIfaf6iCn8J03mRh/DaezmtBV/oR7ZAESX3G/w34CkIzzvTFC2H
oYlnkhgb8nCXi3YMFnWI4UeyEqYqDk8Hm/4GkyWw7RZpPXNGRSN3nt81DX9tj5O531XGJvKFLzsx
BhKH9KEqOHxd1gIKVNDB0dWLnZoDqeYGKMNQS/OqXDuBtgIF2x/8dc5w8PP2cy5pY3UtXI3+VtmY
L2zjbXlktycTrPAKQfYNvbOdSSlo1HcgyZfpTEzyG6WJltyBXmILiemvqVmnSzl0Zqb1ngwEzi7K
oIk7o9c1ClxWz2FRBijnu7S8duGLV+dIAmrw7y1f8nIRqqL4cSugfzKn2ESOuD2IA5OXOQ0KAkSB
eFphAigx/surZHOfCHZO1xJmDidpPy/vEGjhwHRcOUAfnPAMp36cuXiRcZkOOKw35j/jTVboKOqj
glWwVGsVQSKxL7Aaz9jUi/BS9UUdrOfE5IxFnedAMDwYlQEIhKot4ODh44bEpHHHk5rRL16Scn6T
O59oO6tlKNvaVVAYMCdgicJM0+YpzUPaSii4JPTcI2peGRURkkMVUmRLlDKw9U7xeHBgmr/qrNNS
qCGE+oGcJe7UkJC1jWZAex/Qss3gU2D+TzV41pJKhmRru8Oo7y2KrC0CGfrcjRY16WDvxFONEeVN
Mqslx4/TgT0U1yOgov9O+NYRpDsY0z3jRW2y9xGz8O8vqXjuNOV7JAJvtZUnSXsmNUXGyuiSBqOO
YmAMQ0ZccR0WksLKgMp/0a6XrFulOhYrpJVqGn2YMGvsbL74fAPS2WSw2n4fU5WL68cwIHNSFUul
Tkz/hxUknHz7Cw3hHYIYtxooFyEGrd/7EjhYKa3X+48hA5n1TXwkk2bzz1VJbfkDQFbavzxWlaK0
s/D2kIhhTHU1UHT56XuWt4Da1nRf9porVuSWqpiaBHGVIADj58wykEPqpgfbv+jNjHJdQuHCkDZ7
0E48zFvOB+vP3V/G2SXS5ttYVqjGWbqQwtymHCO+ysojWNkKaW+sVwSgFIwYzKmP8lUkLMIroYoj
R/Yixygr7bAq/bB5Ps445/7v9401IiO6EUTsHnijs6VUXUsH66lZTrIs45o5ZgA6W/y7TEAbvg79
WdaMy73ZW1R/fmERPxRh1kst+yYVzC+7HZAf3ZtDL6MYXncnbuXy1AObupbQGOygmD9IAxjhXF6j
zt1hXjYRqq3vnfciYnQGAmChGdyqhr25vx0IIK0OGOako5k+iCBd8kg0aPfrGVdJGQ9ENSb3aqoH
38NvmclIHHZs6xMkbG9bEJiq7c6BmJsoGFTHqtSs3khJ9IHdo4LecqC6wjVsovwOcBqTx2DG9dcB
uWCyxNisz2klRIQ0XoW7eMjJV9XOJ20r9f99YncpzsP74FX8aRMbQugwDNoLbtGVfG/3JrsTVwLP
sNoSBzIvMPcuIzCAFCMoueqxkHa5+EaUVpMNdMdHzijPNNRnBe1xfyRH3KmrQI1J0JxZ/+qjdQZj
N64R5wF7fw8CxBLbIwSJg9W1XDeR4uwOfciQDSh4xeI2Htu/TshLijPHXE20BtC96wZk3w3fLThh
Yg2xUtRa1uvH2SuKDkLelTBhzRGutyQZkboZX6jZYdRxxWbbgoy6Fr8I2EsnWJoJ3k9/bmk0g6M7
PZpLKeEAxicGY/+bm9uxZUJCJdTU/cyPAaWRFR6zCTvoDbyFF8LDG750EaFAk2D2PKnFo5xUaQMJ
J9ChFOnzdH8tcwRJFUofbNbPzi4X1lprnAsmZUg+egaYiS+xyf/0OLnKedQfDatWu7MPxznc3Y/j
I+9u+gxlfDCpHtTvlEjjS/IFD2s0+DtsSs3VZ0n5IoMC3Zoh6m9sK2Lyn3uL+Qf3SL538dnkw0H6
DgKYwc6D7p4J7vC6AKONg9WyPL6ezQPOtmaB7RgSJQ/cNV6hkGnYAwHFuJ4lLvepz9Zg0de5bZiV
ZzirBqfnickqgIeXNLuAoA0rLxVSdvwUb9jX8wZtrXgTHBhgB3UhZSjo6jWIiqfF/BAdrgsi0aTB
RR9kKPrA7mdq4HFdRD3KT/g8ksZUUW7eWyXNWgBm9S6E3hMMRW6/W0FoC2XTtxYz966QPK84eIgf
5Fk35KECAbVDdE+7XDRwWxU7Wpih35Cp7+a9nv7e2HIkgtRCWRE+3w2+VWQTSTcIoSkmt2LDZVT2
m1o1+WKalNpnbQ1UlgjvVoIVSfC0KyxOJYsntbUZUDkokaCpCI+fc0QZvMYXT9O7aY6vRXriZJCw
WsyK33zbRHsirn7nIFno+MMS2DzveyyvIzdP71xJVLYfz8p9GGD503OeBjJGp5MGavSVjY3LIh80
unnMqO9naKVWiUc2np5mxJVo/B1SORykXIaIf3RRgTlD8FwddjZ0kuPP0N3gCU45/Zp5FXyFZJ02
+prMCBIOUMHc2VVmWQ3cJSC1VRPn4ToPu2CeOYEhnFxNUuwCazsFyU+Gt686G6N314d/FuKDh7EM
cnHZ6wkmXxFoRTHAXpQeb6ncw58FZeETb1t8Eu+H6KlXHtbTT/hNfdM1LJV1KYNbNb04SYF4E/ur
MVJ/7SDSa28zoegQ5wAhje7cbQv1FK3IA0wcB81o0lKMpBQla/Ey6gK1SDCn45KOr4rUP0sjj7Pv
HhHo1/6zG10c9nniRSEqqOhmMGSJzq6fsWPF3qXTHZ3eIascnbRJk5dT/gkVpPAR95god0R65xZR
iQWDGXDOec6NzkQpCyszWZu8WnGlHGcLNS5SMcGRMwHNm7SjdHOE4tau+Cf3uClM8PjjLRZ5mG4Q
vTu7A86Dr4oB8TzpIbhIQJ5NdycBebuMS6YhSF4E8n4GtnUj03HTqPrL/DSK0/cDreYeTxu8C0oO
cNPM1BJ1zo57zAhU1dJZI9ohNJQorp6jiYW4KnXiRN4PhTfUD224y7WCZGFuRMjM8BHEv+EPQO/y
Bd7zeWseDm4oMl3Tu+SciGPX1yud7dJSfKnSpK4fTr6sle+4dBgPrX8oqz0jifpEb1hmxH7xMxbJ
WgZWXophmVI7jPVeyhCvEf74BJUv+FJZ67niqtiWjdiAN6pmNRqUp8kppKbJvQXS+rJHjHuyfhSQ
3ofWP4FH16uddji0HUooLQZs6ZOyhRjqq0nI9TcviG28tGIHBvuzAIadDDTls/M9OUoabc1hMoRZ
Fl5QCeMkmHUmvLCz31Z7pmsg62JwwSv5i3YcQQ53Sqi54QCtcE5Q43m8B5EXO/kOGq2U2enpT5XH
Iz+Xz0NsDbe9EeMkLsUBMTkO2NxX7JhTXPchvh7DEOPKkA2SGVr/mPQ6Q1RSWSupb+DE8FdTyXh2
DxwreayU3eyDrPPPZeRgAeBJaLXdCm9QQDmxhRNJ9/bUAetTnuYtqXFE0fBI/X7e82mLTFI+ENrD
TbNhZJG/C9eWUj0gmwQbh71z1p4Ai9pjVAsPMGogYrKd3BFVDBp+dSpggl7pkMrj4GXiF8Fvvmep
l9a37RZt5X0xBjgpdDcqoAqw6hr9oFx9KDk44Wq8NRX/74uZiTzf8e4nEszkeKAYfzKCkEQYJiNp
pfEE1Jt1Jj5twExBToAcKr1e7k1cTK4vYXmUToX6ydcRu0VUlCp+WUvnzsBUu50gMuCfisSZ/wPG
KQx0aC+8p9+Bqo/upWueW5SwBMIC848f8S/YPpbYElygj+1U9hcIQTXH83ziE1he/PXXoxXix98f
G5pd1hMZxB/r6yRbKPZJ6KwPdX5bjF6vRnPnRni9GWbsWMc6iwTJsJwgxNS+rVmeQJIU90f61u6R
5qvDPq1sSXP5NsDxH+mYcf3eKX3BUhMwRf6ACkfTGjIDrMsEqozyCUPR38mBNviEHOwbv12m1s1u
a1ZksX0I5b/WwvWjirIQLrBnWioJTgNTAn1jFo0PYeItcvu3D2AeKbRP8B6H1rrtDEs7hDO2RwXI
ANjE9rNNZ3Brv9vf+0TnN10XyMB7oI/pQw+akB8xtmdvagBlJkAby7FLs0sRRQv++8+GYXlU2/Hu
daOnTSluEmeVlX1ssITALQQKnS9wOyLGeLN911Kr2Geoi1ZTLSsxjoZjgc8xeFCe/dspwZF1jvrP
2/1gmaH5MHGpivSlcmv/NXG542PxkDUfo+M6VKI4njuunc97iMzFhs+dL+b5bjou7HOKfR/dvpC2
kV4ung45G56A88crXeADOGeD7apH23+JYJ0FtUwZIRI+gHtGoNbQSeSQqPD1HISgk85cMTUtEq9v
KAJgSZM+soZhdfdnsJZOFdfy2gGe5nu9GYGlXmYGqzxbyO03GubKigEZjdumqGZFEwD9D3/+Z/e5
YeWSziR2VCHel7+B5Lpvt8cGKl01kgPuNQzzI823YRsim0ClmRWafFm9FtqedOFqKOgCSerBLlXM
CIuluqJ97i3yKwGFBKUjxiGqSCi2WwN/8aEpwn9xJ5dNKdlN+E+l+1Doklq5cGGzyJ0ED+kDJjmh
YhxS3R94MRTWSaR6N3LXoxVAOwwgsZK44NId5yfEOmb+1QufN05ZCPwxDJos8ZzoS3Ivhc4wHP53
f0zt75p3AHpLFqA39locFRMi5ZYvw2XcXsxxIkKWjHTWi+qrzvTGXI+wXBpqSZH/zAY14wQbhQ1X
+vaRyGKpSARLR6+crIXnwTOyv7xJLsFKfU/VP16Ub8O0MO+0e6E7zwsaDGk8nd4HEiWfEd2MSJ0q
sPkIxlYFN0t65B5uY9L/fY81O+d4BzUi/9x+aXdbbXDjUyfkuJCMWCv0WA6S3jVOimeZPIurH/Nw
v1WHkmkwPeXqoxPthDAvTwdb0LGCwwwlvEmmbIaj5heSHvHuqvT37u+kL6jaB0U6JOKSPT3xU/YI
aAb+qt4tJYsQtzSi+ioS/nfZPUmSjqA08mxXUDpojYRPuQh1dcYC9eZ5yETo7kQrGUDWkCdVA5s/
Zc+SVLfFEqpA1a7imAvPv1hB1XqiGsCFPbX4e8VMqzL+4nzQRHQD94Hm0gdzPrbysMlugrCf3Pw6
K6oltaB7iipJGZv14esrtAgWWAbjgIgjt/UBMzVDfkLY2hWwEsQJklfca42Ovg9N4nA01AarGiaQ
qqeu7luelslJET3Lna60tEPVH2TF4v1V4ATDZLg1XoomoRCjJCyxNQCUtF3qhZapWAutfhDq3s/E
Whz03Zmx+F4LU623KYu/yANLU9F83fRLtpfCY6ps5lC6HUCLGgsBMFYU1jUOHaPL/KT+oP+nJvK6
Lmgql4ZUuvcTEp5HHvmySxDXtvbIDwk2G8tcXgom7CGguggiBOqWMqCcYX7+7VeXvCOzx/RqpplK
Vys0JK3BlrjRnL/ca6SR7xxAz5DvXpASWo8v4nAcjCmpGv7i/OVHlgzYLwk/G0bAelueW10LuGjZ
HNPsKYJsip/o0Iifv9+MrilkZenmCrayrmEpLO2KZgcZ6Rkvn6dq2VYvOL3NBQdNzdHo0aChO9dV
pqk4eubxLch8ATF3FOfexmf6yo1enCBfeZ+dXqOfvHjyjj1GZnzp/otBbYZ2Sn23V5aWrvnnkTDL
4zsAXKsuLYKlNIIkh0EUsFH8Tfx3IuqX+aVhSUtQ0Wvvk0N1h2D9SGmXvZ+1iMLVmcXNBmUIYr3I
3i2VKiTLsg8O4442Vj19cuj3d/jEXPST2aHbv6l8DVaxhNRELdm6m0YoYXNXyMa+elF0mi0vTGor
wmPqr/ulOi9mFiy52sl2joLpGtdz8E0y5csMiOo4Z4La2DLgj23S0iD8wp2XhkGrYTepVX9ufn52
+LGM3QpKiOUYBnyU4fhY9LY61HYoI+eJaIHLOWTBs+cSOnZlXfyBvxA2onyR5GLXd3p+z8S1+eQJ
daGDHy46Ur+/30j90MRUBbbun5lRCYs8hpN8BcSMOgeWLv3KbushtnCeCytJIilDcJka5LDrpB/Y
tjtSff6ZlNFuS8MmvnMyVgAw66tHp190XbMB7ZXmvNA0mfBVsRJsuFnC8C+DSCXwKZmNlkTGBGKh
xTdB3gOBuvUUYmpQDd+8UsWZ8EHYJtbQitW0R59d24lADQoribpx7BcOovwHa4OIo1ihSUsIPMLw
iT8GMkepmYYtrWo88eslI8BCnHJfszdpa2I/MEGmYtszWNtg55pVRx0zifgEzl7sLdz+ff86O9fF
zcZ2qA1PbcjcT9nj3DTLwWDqbeXcxwhj3ka4R8lH07HKwXa0hSI7ZTvk0Sj8e36TjCyrJyU/0s2+
S+Qc57NcO17sEFvM1SnC+nvCqDEX4rxKWeIIUO9Z+NWAJvjnXJJww1TvhpevHXZtSpiqIkEiM2Us
dTdDU9z06tl7lvK79ErKGsfrnV1MIf47aiO0dv5+Hlwk4FdeFhUyDWNFd+bIzMtVUHqLjwIJJ2tg
NUUGuaCy2SbX7eSCEZ5mTGFfYLH1kv6OraY+ocgGFxkSaxi4Hr2LibvozpAavt/iH5nvdt5HUr18
PhHw+5aLVeJsZmGXgDQL8Pnu+2pKGAf2D922uskVrBQ/BNido3VeU0IG2uI4//JNKi+6XPvhw3iY
Xi0bqy3mzQcwo8ZUuEDQW/pyKw8Xd4DH9z07+skMCjRTYW+e8/4Dnd9NGrxWcOiQdLXfmf+rTCJC
Y4+Hb1cgviNXm0Ga/f/1DmStKkCxNSA/F4h95TsyL8qYOn63v8kkwkRrXyrHlHKS1Vkwm1HIoRe9
S8BN2ZByDB/SCbBUgS6r9I+Zx2RVLKwzVBRrXhHi5drmDlqFwQWtv350iksBZnnCDz7+jeukatJ2
nSjmCvyB81+RlBggIiAZisUIaxFZaN34+8Yx01CUbg2BpgIVHt6+bKXb8BpcApgEKRM2ihYunUT0
/x4hSSzFGMKF68uKM1enePogxaASvut5dWezYYCF6AAH5CcY4SolWkdzcVsjbUmYcDPnpZ/pTC/M
wzT3V+8+BND9jzraY2O94ItHDjJ1UI2FAgZgAiUvgI4ujA2Q2p3x387phkzsuwSmluvt4vG5c98L
WQk/8qu32cnXtusv3qqwtWsBpEgfFg9hDM4IB+1SuqMMRoK9OZkzmPDr5QkpZkSlQxOTG0Gls+iH
S+lQCZXvPeHzG/acznQUwoXVrqovP4q9hPkrDf6xZPL4nq0sDlPA2dZxnZiw/DQt2EdJ5xjdmZIO
sh3inQ9O8bpZPz8Iwkg835sFAoid2j8YdtNV+/WB+3lbgMZEXCkrOrIHCb9scuACQHGh+lzN+chk
Xtw/DndcefzT0GGA3BDklypb4BFHbI9xGVbRmuIFIHZiK/ZpqDrmBnc3ZT+CXtVT2faLhigwYLim
Uo9flfkavf0gM08gVawzbZy8Vcr5//oeALhcG1HRyt5KA0EGERHNqil8CDw4z+nokeeg+JhMgeQg
u+9yIsRGtNfpC2KajT5JI3oAOalCOVwxbtNNsi133/pZhLf74bhyWRraofZgOw1rXMim9ahYW2vI
X5yOmX2aPYYY7m/zz89wq+ZQDm78ZVIrwO0R5aRyrp+zgUwa9dipsUvniiQ68Q4ZR3iK51l3pxrh
jUOa8r23dw+T5eXTg3jUNtQFYiPxIG7t3f1PAqXJrEUbNLRG+5+5dIGX7ryhLHQG32NDr0aL9qfF
FMtPXjPL79KQDeQhYBDC3mqZ1HqrMm5Nnn6U5zGqxWw5l+SBODdDgVpzbr134N9suv2SOh0T6Lrs
vkDASscPXKh09O29zj3IggOT7hRdSE0HhBXGq3HXLg8tgyS+kxza2R+XUroPne+7VMoZCI8iY4xP
ulONTtq2x7RSxndvm4yR9/fVYPhe4GthpL5DEdgaDcrwQiCPQMmt54m5yOY0H6dKsBUdiyOrgEqQ
ZNEpPFl5KTTsHTAomNYBggMRugEz6tYpn/gkCEXVUIxFIh/isc0r5dJU1n9o2WYKi+bpvZwnM4hW
iFvdhihqLlckdha2Ilh6P21UC889BQWPt8A2FxFslY0p0iXHiF/jGryrqDUb71rv7GqhdlkJu4s+
FalAEpGK+7nMrREQqVktgeOBo0VVQhhpcQZB0K230YkCM2zkSIMwrYrWm4hbzkUDHdNShIFkG6bO
wk2+jcmRxrp2dTXlFWWGRp3f+XoYryhIsTGBmjyQpUsaB3bfmi8aKrFpUVg037gdLcXshrTt4a5H
StYwQ7KEM4vBly0NtMniKPYttEqBXtXpAjRJfVLB6fZZ41VloQry27XSfbawbjiUTCrEI7IJvgCm
XUiMe4wgCfDkoCmLmts7URtf8m6I0DmRUoTSsc/iw2hFIL+FeLrWwcgGuDG/3qywo7JYyfcOoVbX
/8rAJHVg9J9B5xdsSvochMEITdsvAoiG3gsmt9DBGvdX4vcnF1/xb7beNSwS9VPZmVRwWDD3N7E6
3jPDLFyqjtSOnKnKCEuRjPLQ302SNUPjmqMlfMqhGeiHFrPjVFy6hdsjAsoFU9SjOvnhBHDdWxLM
/coImMVJqOjIdUGJ9DAg1cDM0uy/+vLEkcMCt3iFE7cvFARtAofyLmgYC5rwoym/IreUGHj9XtAm
0xZdXyt0rmNW+FGagaKP/j9RHxlCcSCCAhKRdydEQazeF9hNx0kTw/2zBnAdPgWJh3KUvNBbn0k+
Kyuvo7ssrrGAUNrplAyyfc8itJ8I9hmWqAWZYm4U4EgIqQCrRlTnzxgvoYJkDyrYau16aEmCn0uC
zXnztfVQgDA89JABU5KNcfZEg5xZMBK/RAiKCn+xlkYOJ1KSZl06g/ofy6LxAU51pnf+Ua6fW99w
QWWUOdplNo4hO8AD8ZmskGTRdfkc3wZv+ISkBzAUM8QhcTmBCZzU/2Svc2IaP+NPxxgukyPyht0P
j0m6ULAqt7i2431Zr+tcx3GEmJogSkCCPKT7OOqG+Qi3i6DCXFvam+P70YTOxaG3CRQOascFQej1
T8L8o20rua/z2oWZcPalU0nGXg3fdkwW6Xiy58gFelCpn0HrpZ83VUMVQHSt8Z+VtQf09pBG3crJ
zLjxMXmhxnMHyX8Hqwft3yEAoms6hTeyhB/raLBLre25C9pcndYux1zma/TlPQinzOFci4+/wnuC
LauXe1PX4wFQ11e7vDBjC7K2xtmwhVreNfF51PHsn/o+gijfvyYq221i86OSmAvlld+qF2c9eoNQ
Rs4h8X2ppWka/EMM2LuYU4J6LmBODwK6b/AUguLjs9/FMbOGobmCwfcCJtyy5Ikf0vB4i2aor+xm
Ow3B7Mqize0m462x4Tuec5JYIOF2gpaFsjBNjqYsjjjsGeh+Jg8lQzUvJu9wTDJjY/0Ra853XFrs
VS2FkfJYV4HPCMsL72aoSiq7otCoRm2TbPzuCDsVawO8TQOZY54Za8ze4UrKbbFumUEW5ctCedkF
CDV/0MjLbJvFd6BVr8PUMc1CnTvqEo6Lt+aiUmW4tdsETW6ps+hcTGZAnc0pVrPF0rlCMZ8RR5oO
GOmb10yQHypBQdyW5AvCy+0WII4GspM+um50YdMZ0fONcMP+XZ6fwxiuSpq9/ogIxZRSxl54rUvk
//dHeMBiopk6WC4GU3e2ixzxD7Ffoq90GGtIIrbQ3NdAd1rAULWHIC3LUyNUWV8rmozT26L4wTP/
SchragbDrNKQTu9W6FObg0LU70Gegs4mPspxHjaR9FmS45s3AIaHxG/g8Z8iypiYzjLYP0z9koAL
BsnPFNpgW6eeKZbpgr/nZ39gPjll/zOvgxkCoKbLzgnJUkbc2akiP8hhBb2jVmolXgcSyDHnF+Hg
fQkgJWj6C1wWV0CHR73kpLl2TPyJaZFMpy+SNL74AiRdHhzMkMsHzK8tkJX9kaT9/pmFrL7jisn7
k2shxlc1jL6cJ1CJd+Vlw2/f4yA6/+KO6yRzrsVhMELhh1u5k7CBXpRAKsyNdK0Mbls7J1aRTyv/
Xzgnlt61GRZ8bFVRjfh/3vhqP+ahsG76q10ssqbslCG8Fr4i6uDuvsful5+cAqv22xhBuXuBdJLy
gR1PY1EIsBTK/y9+cDlmNiY+N/FrJKqNXmp/FuxfXfF5Tz33zGK3AJmT9Ps857d9HA9n07lj8agM
vAHq7zY9nzOMBFlYL7/WtF/PZzBQjHUO5NzOi50TFnCd4ZBTvVlMVtwJWALa1mAmnG+pvL/gHKBt
Pm+U9bNKCZWh0AcGMkb4XpU0mXsBpjMM/QvIXRLSmz5mEIggC/eEzly/gwc5CRZn86rsYnnjpJGI
kfNTBJZXuy3jdGsUOL0Tcn3QvFp2g/dtnmikbLGiespm7AvafWPbaPLw3PyHF9EKieloL+eWv5y1
0Dtdf/ri5Z/boNpPLEa/VHjnMW81d0q0w+It44J3jNnSkQ5bV7IRTbGF5IXNp9geW5jXOhLODTwl
9ZupL2oLhuUw8yAkFuRnuqLy9zI8M65LJr+8u/Kn+YXlUB4+Dgsm9gyRHHbSjPAqYr190VWXXsIG
BL+x4V+DZxWkYDxPQnmsozz96Ooc7kjQ/oH2UksDR9CC8G8VUc2VRsjT5G8a1pNLm37dkNr/FuYL
R2Q60SMdyIXAZr9YBSjhJsHY0wIaJHWRX/xgQXMP03ma7dAbzxbIeK2WOSSijOKci4NtoTChwOek
biHU3x7iNsie43goy3fFIqiBrXd2otSy80ce2A+CHaKJmKW8fyLD81yKxAx/pGbKFZUyXGgcKoOC
WCH7jGVYmpMA4nNkNF5UWd3HfE6UweSukGZF0ml+ZhQwFUfrYkd2lVVGTeKCyjV8s80uJBiV+nBZ
rO/SqICULvqv98Ysm5JYgv/66GtN/jZGMWB59uwp6v+BPsxtVtTBQEh7WhfX3ibPM63BoOr7AQ2H
X8R7crtf59i+2A9TdnOKWF12t82j1/J6i0/8hjPhqxO6XP6H2eEGqHsKstQ9/JNCd3VJFt13jKzs
7p9Je81zp+IA+Z6A7aJmjGUJ6sTglkApYGx7H69Hw/HXs/67H+Re8uGMu9rrUXmJFdvPQ112cVo8
Qh4JzfjuBBk8dbZm8nq/kF2KaoyhfYldnEyWB3qZXj9TfxZxPsZho2LeqdkCPLoFjaRRYGwDIWse
NZjkgR6MyZDh17nppTXSI0HIoT6RIHB7nSTh0OilAj13aYyHlAa9666tDwGdsrl8DB+pHI/PqB6W
3a3nrY1q+XBIa0KRYpmPYWdpC3xCKx1c5dddZ4IWvi5zr52v9VxGSZaJ4VLl/aNeEPydYEZAlANU
oJAxDBng4EMzpbGAIdNBlPUQrWW/4Om4o+2JZ0TeptKULFVMf9sRBajFJJAjUB+pqdjA3f4oLZxG
1GJxpwME2HHrHX/Wb8HCtf8QPBMSpSsMMO/4TMh4FKsc7dqEM0kK+TS+fD6XVfAowoWbURmse7nx
DSkzju59rc0Dj18cHz4GxEPBGsUdiJc/2O8lldXWCpYakKbx0qryz5yKZgbQcxB7dgk2KBlSPbd9
hkikxLxM7Oa0lmi45/eaHEPCOPazciSNXLk6uS7h37YP82AgZVqskAE2WK4gjvMJl/OYWHK/Hv1z
gYCsiMGgMUlREEy28MXBnJbGf04qu5xCnobH971I0iN3AXFkjVnrfIyUyyb3sstCh2orS36GjvXg
FwFRrBBhN0Ztbk/eiRL8qkmM2Ft1975QnXT3cdLFda0/fe4ZQ1DZvdbK9/zOvDaZ//5rEoJ4A56O
YNhUV99b9T0Vz5OAF2yJhVzmJs8peRpgeXTmQ7aHW1bzvqz3MYObATmhU3BGmgODtlBSxsgGEe2F
Mkwh9qUx6wY47iKi67L43m14rnwa3c+biHWqlCyDOBtYE3N741aGx74+vqTjeoq5guZQghz7SMKn
KKEvjMm+58XIPDczmQh9p4dFkZEpYAYknddbFv0wnLSPlYZQTBk/E1TEf11VBCjecIO51YPMR9zy
AdXI4wtibt/yzk0K3OkljQSeaqMCOeWY2ZJKPFBtlVBLALWUFWlvF++Nu4F4P/r891YB7QtPgITh
zp90DYRbaePZ3xxveaPH0Sl7CN8nsaAUoj9PgeYgbrrVmwfLVo0V06TLpWKfPcfJxrXPJPeUyJMZ
rJYVAzumWWkLX2IurTxwfkZ4u9VG5N/uOPgGn2/9xuMXzoQYeJuxwy6bdrObOlEq85/royOW0W2L
8kYTInfvKWcKTNeT4uaF9i91uGS++uEON1172lPMcBlbd8/u6itcBskx+rKMG7RXhcQktHpE+gpJ
kwREtqiuhCNnmStiNRaRrwNin6gYxg/Eo4/U+/nqecp3RI1ucZ0bdYKP4W10IXnrYLAhvKRDBqCv
eQB+yHkEKEv18aqWkhibi1MOheuYF6eqfPkU/yN3hKemCdm+IHUdztCnLn8Rh0txWyRzQOmg2iVZ
P7AfCGHlFexfiHjxNKSQ1V1Ra6HXThEnQF4GlODFfcphJdC9dyuoOK1qa9u3QBufYHAWoP6reUO6
G7XbL5FWJQJpleRdIorbpBKa0lqgEc20vRpZ447Y2V4+MAYaU9nYq8xFuTQ3yesVG3BjubjWCTce
hkrBd9d8CmwK0lCg4M0KsnYKzYyUVRdx/SGMpcJLhCkHHF3GeLtIBdZ5+zEWD/UK2bXr0NIx4z/O
4TYouFN4MDa35YyAebSs43boptmuNMWZ4kZlr0uIoGlBze2VgjXqVZmN1TxYtRCBzusSWZwpaX3m
z8NYZx9j3TO1XFGgouaNzJAbFRk70+x+W2A9g/kSGUs626/OJubQxErI+FKNN+cJ5ilLq2IEtAg5
5ci8UZ+z07gRnSYSpUQ1KwlJ5Bb9+OdF5He5aue67BJXwE0wGicA/s5MIxiSpRB8lDd/kf00P5yR
rZY+puoVFuo+uSx06riSfEyozU6XF84/dNwcupIuAQZr+eNKcEX34rlcGWwDA75sjTMi9ie+lmmH
bpeOdgFUrdOjK6+hqg3puznA6jJRl/Yf7mzwFnr/Zc+gSX/FMQIGexeY1R0/zsZKrsFaIagmTh/5
EgFDRYz962mlmGGdn+Yx4s8DdHYm26DVIP50Mve14AwoPB4kpYv2AxHNEI94PvXuEPBfGfZKnHGt
IjtR7GI5sGfFOvu3yq0gIfb4NtrV4AO+1FQAJJbvWkHKnyETVIV5ioKOBdmoZLsqj84GFdRf7ILs
oOvs9e62MaCJBQLvzmxcoG+NI3UsOZeSZG+Pt2ZvsDFL7lOVgaY2xElENJA1b0skw7JegsLhdxfR
pPdCyMSuWiHD9lw3eKNscc+AtVcdP3e2gNLzxMO9IGCWVh/UZX7zLFGL0+C/xhp6eZOIgl9wF4Ac
qeOwjry0MiyUCK7ufNkP3sA0g/tVoqdkc+GAY4L4t7EEX4GZNEaCSnqgi+aG2AOtg+DUg60fWdcV
8+ORGe8j5rcmLBvjhIBW54XuIQlGtDNvSC5gBD4oVwriLL8dQKB7rwaJ53F5C8LmvDLlklW+s9Ia
0UQ+n0zZeCFBL34Z6BEPi8O8BM5g02o4iA9qlJQcQgSTpc2K1Dn2BPoEU3kOyRABP9ve1hUA3RFG
8T214V8D1DfeT4fFvvqSq5r3BXjGrenD4b2UX1fhAMnFJXwLFUrZW/AwCKA42vQbDojcBmpsRQZH
gejjU2vcg5TuCc1d7q0BucxbJ0hoQ7SDL7pvv1FjVHP4UZwAsG6c0aZJeoMGodFTVNYiioIJMRHs
mS498LFwU8a++XKyYqW61xCBEAATPtUZ4GpPtwS+czcfN3XSE5osfdQpQnit0+V8PvzqB0La0X1H
beC8+7yEW4Y2M/XrqZm6463sWYUW11bv6ZlmqkjWqGpO2Ib8BYgBuTswQgkv8kTqrzxAdYbHEypN
EIkPi3/9QWBy3xv10imJXqjq0jj7OZQvyUegTJI0WDYmoYgfCYVI/+jKFTizgxJMw6/C5yn/X1so
9l0MEZiLopc48bIUScbAM3vrWX9bA0PyS0/zFkdBlR7DxaWRD7ka3zA4kxvSkv4487jbOosikVlC
sDF2fYQKlsWZifpu8p15c9Ma81qxwp6XDgDWM2yWw27WXRTNx7XrIFDNeYvjZwNzfnI5B9olVUXG
OezJzia9AxsbtYcYKRjdL+4janvmFKHgMIBSkEsjs7ICw2pHXM12AN3c39cXiEVQxM6zCPfkajl/
INaBbZ8M/Ci0+g01dmzUKMylGPrGIzzhfBlfpHj4jvTu4T5miO6LRnKxbntMUCsQCIxD8GlYhnZQ
GH8cEXxxJEs4yLO4WWlrSb01hTWh3ybi+/T43++FCfoB/SKXhe+b3Rjx0K0xYH0qqIk+8YZcpr15
4WyI645F1g7lWZjwXuB/9jUstcyAT/NqbHQ3ROLF+96SKtxKO75AEBCnEuKs6GYy+167BIS9aUIM
8kPAPnotN6GZjnNW9TGxYfhBF+gTUE2663PiGW++Se8042gQV21qFND/fkNAXb4kjyg9Z017crnI
7E04mV83E0CO0aYSf8Wrh+b7Ep2RkLCKEoHDmz2F8bzZcNQtIum6rcmng5Gipp5kL50/UI6Q3xTP
uVwYx/d6A2MUCKx8dx/9lZggkI6904b7EW0+5h/UzCfKfUCBxLOiWoPtwJdKCjb1pgTsqRqOVUxt
L4edcTBfrFbzMaYltvULyUj+VGOpefN9AQWWuVz37T5msMP6KAfzWMjqtsoDAeS6bJipQO/+TbjV
xbLX3lI0OAayMlSWNP7QNpu+HRsbs/ZtUH3ZhQlKQ6GrS40FtWdOVL5+NC0N6Qx2La3PUpiiEjxg
Z6B+w1kIm1wF1NNPpMJNapEDhZPyBm+o1lN8H6I/07QtY7kovoBadty7gQNEs1gCet3y/qSrRPeZ
IXaOboSCy8r+5cf7l+94T5vMPkbmFd1tQ3Ww4+RNrVC0CFnqZ4TNIgu5U/dSe2yy5qAaKYkNYWiT
WCDvEcvGf+qFCO+iOzAkyaTbr3l6Xl1xKGj9OVAWKCkNbCFxyTPnaZDvCORgsCZbfNHy/SAcKJUY
SMTgJXY7thRURkkKxIUIyYexNSEC/HX+TYXa0UGC8gOTKUpNFBz8bZzyOjsH1/AgD02Mv5D38uYW
yVoBqWG6me3aMgUHFNQXOETqwnqlyRevlBIcnxlAiLpRKvMVhoaZtr7euseM8qxSufOobysRkhCY
7XnQsQYWltb/wBomr3N1aISmcgBX7Tbutx+fsw4w9UZ+d373MXys7lKk2KKE/I94TGbQg0VnMl33
PYAoDLyblxp9IQ71QBd3yLRwoe7QJbgCn5FjyqYxs4dSmM4IkhgTBCSWXzY6KQsgw1C90wlRsHCE
XDI9roJFA8MExobBaD57pRljW0cl9GqWBOM3Etc6q7/FuDjolqeYFr0kF/05Cq3oHfVLDUSBQwfi
4DVnzKaZy6MpcOKnMuCxPGug4pZB7iN6K7HqPRite1OgRBSkERwZ9v20x/5myfH++LDx6er+2GN3
ftp3BRAXzubHt0XfTi5LChZNNlkFtGcpUuOhzX5VqfNfz6mfxDkORkvHom8O18XdaBVnJoa99Mw4
pxp+qN0kOIe3Gtyvtxtzs2losfe3CXR/Gp+tt72Jwh6HfgBAHzCKY+8V6lU/yKNJ2rgooVbn9Cyo
X1K4fL6+9b0MYdEGfjc8vgetwmejK9sa5JdZZ6bWM9LaMQ8T1lz1s7Fzq4sqr+HAadF5yuN/5+Oy
QYVKw7dL6ij55zcQq33fHgF412JjcBUZRbsIWKruNETo5Atsxvr+pDdPdN/A6fbHxNLZxcrYxfRn
KlQAq1Cw16Wogw/t6rW6z80bKtUGK3W0nhzg59KoyXK3jC+3brMr6IIC8iJSni7AP5lKrMtAMHij
2oW0a3knMPCGiNo3OfieayuYOOo+C/BARoXvTRQetD97KAIPKNuB4vqaX30QCa9DkfLDu6A+aeKQ
YZa8VEebBhdSb2gZPRicHLTJlzVCr7jVwhEMX5FWEoaaqa8a6tDK9ut7rTQBEYfax9H/7EcW+Ihu
nzl7dxX3X9YwRr8j1smoZ6awVnmHZlldP6YZ6H3sCi4ZVMIvl01v4+RntmxEzuE0rwwJ90+9jl9U
C5+8sjJXUwxSCVTzM6J+RHAWBOGD4oTxv2PB+BFFdVMteyg5Qgqs0sI90OnfDhLy2BZZgfbIOrlY
R2iKYqrFjTCUuK2VXGDudoKSyuMAZfSMqwglTOtBVNspD/i2wQoGltBOBvvgPbuzIqcM3cmCtu0q
0dALu/cx+CUeSaUwzgq5+aSRaHUV/hP4gOdiox6lkh/N5aA+eif7nwRFuaB4fZnZM15yISMQK4fD
8rs6jh3ArZ2/EKug7e76p8wQ7Ku3mMSZe0ZE0B+A8A8O8kRg0oym+bjMX9xHnaeEWyUQ4muvO3zk
XqJ74mcvVU7D+RH+rrZXwhVHj/sDFXPdc/Oq7X15qsypo+L5JjYvDInraZsJYePXPuT3lUrFFzdb
jhxUgHKU+Q7repWDDy/h7PIMO+vUmiQg5dchJVBWf7xWHl3lYsbX0h4Wxw394nXSG7uKYcv3wTsP
QdxmaTS7U3vDGNSVvO23obvlN2xU7j3yVUwq/7FhT91AeC/TxYmXJ5G0kJesUTnrUJOyIkxjPQhR
YlVmlUKKWWM9k6nJyVsI7PMOT5jUs6rIL0oqsZUt0YoOQOZIc2QnSsHmd3Ifin4YFDBacAZQTyQE
Ysc383sJdLZwdUx8iWp3P8BjAPl3rCQu9Aen6mbyVBykQhU5OxcaErHlzur5kOPb85N3bycDCpaM
oO/PQEDTD+iNrU/rG84pSDuGeriWXLRvn5HpNccWpUVap8Hfx7TkZ4PKul7Xkl+EYyr5J8/KNO4W
pa46roYyabkZSe3mt7bt305eiarqX7mPwAaW/G5Cx0T1aQ+W3kDVrcVcIrRJjdoMph4mPN+eTaIX
A4LW0ecvty/ju5mCiOruElY3WqstXvTAzSAfWnLpU3InEN96zLjvQppGjn9BxG1Dbunvml+orYNX
gekLWvqdDL4fCs2faYwV5V7Tz7b33jy20TuvMk/0uYd08yMd9P6WMn3P+t0NqFVdaEv74acKn3zk
v/tRQaIx9dIJy3yVx3GNOlkORVj7ieQGrokwugSdCx0EsNIpn8m7ZDsbDYoPq1PutJE8zUCfeHCs
fRiOT34Zzo5pFvmJiceY+RblZGv/3p/lC9htp9bSKj7/E7mcrLD7XawGbO37aAbYYh/SiODtlOrG
NyGXEHTh3P+hUWKGMMPqkBkR7ykWWBy8a0iKgwBKyfjB89PYBOVkAdRTPIDUPPUJIIsPsBLPOFOP
3l6X7VVOi+Yl9EMRqTFPN9lq7UdJRI1j4RU6ny7HNsDIKD2St4017hmmGVGMhdQzUujdSIE195Ka
41q6naLosTksWuCBeXpiESZiyE3Yyj/zSJ8k7sQnC/eRAoOKGKtdSm08JrYY/RA6cIxFXTxqUysx
j4185JwOV3Ywd4MjsA2dTPQNs96gVf0sK2Kutb7SvBtUkADrfRs8xCaKELc/Y8ApQ0jYoU9hDy/4
SPQEnMW5m0vhTFL6VEq7tOnigFWc/OrMSvfG6EeiQaC1G0U8bnP1heOahYoqJ3kSc6SjIenRk5M8
CD7xNzIAc4oxsIJqqxk/5Faas11Yw1HQvkR1M1TSl7Oy8Xc6SgA3qOze225FyP0F+gwDhwjEEp2l
WeuvJaihL+ity4XQH17+IgS74xcW7d9LurEc6mwwpgw6CEv7TF//Yuk+Os3+7kp+/4eKzTSZeTSm
sYN767FKqckZ6p7NV/ts/IFY03N1SwsOpXS/xakMq9uFC7uzvxZaBSadKwGgS6dVrTvEZDC5+fSG
sCPpZn52NmaPctgESNWMh0B96JvQ3fbLL8Q0pXpNinlITgn1diGewHWSrCz06CC35dbzvbvcExpI
2XMHYBD/XHsQJkwfRNhNI//OrawWrVdqz7Qc37kIReluIT00yyKIbxQcFKR0Xe262NS+A98rTVmC
gWOcGv5dxN9kfdtQMkeey77VJDfzgxKS9Epc/Nk1bOv8II//FwghajlS5oh+3iK29Aoa4FhBok4u
NyT8DIikFkFJ+f4sVtETEPaURwkiyaav7xWTiSdJqLmG36Q+cIBuK1dxrvli2Ic36wQH3MevzxaO
+DMIl5P/vUsdyy/aOieTkx7i4nh3rXGaUROvYg8FEMPrU+DXYntjK4QP0j76qFJXHKK25RfZ8bEr
8W8xp8R8mE6hcppr+jg6hLgkcxl7sXP/xGo+KenmtrRQ6aOGbIbTu8Hjwil0GdNkAIZwA6XR59XO
o3qwwHzhsvvg/x5/jJcrfj5S/OGiBItLDIhfkrr9PlLyGkflf0zQAzvkNnEt5TvKDqf1dqCdoUcA
YsZ2cEZfs2HvXAla3IuZFGyxesheySo36YyRREstR8YO7VHPqqgqpDXju9c+8Skct42I2Cx4Nz0u
zXE8h7fCjYDIGBMED/oU4ewbO7MjSYq/e91uGkv65bfbHvBoGAxv7kiAXGoXRqeP/EZhrW5j3xEX
q0St2EvEm2jXRnNF5EiadsB/Yl9aj4uI5nK/WZvXk6ypX8ikWpb7XcIlC645hXLzTuj6sxjDV1oC
XABfv68KPfIV9h5x2uBPhHUm02HpN4D6lhcVuSldmBXl0BAwaqdE7NHpE0L0EP11J4joPzldZnO1
9QyrtPIYhoymkKkP7S8M87fL4E0ZdJ9wL2X1HgqTlViOpcJGmvGRCOXkAY3w0E3Oe4ZTIse2D63s
FN5MPDiTy43uXuRItl2Mg6XNgIwcxvdVTDEgFMBaBZAFzDbAaKy3x28rdBEoHYcbuF7jNkxDDA9X
6Osd9zWcgbz8TCNbd+EKyLVPskZ/K9JNOfLHYSgledxOekLTTrOfsgtJBNOyE0Fs0KwM1nFO3U1o
++KuPNmYDtvJsBr8zg8xwdF0inwsQ2Dqwi0QILICQ3IuVpVo8vxWjYXfXnboU2LNj71VtOPGFw0U
wQy7bXuOit584Bd//3Dp+c3ZtdglgQvdMICfoDw5b4vArDSXbkmC1G9USLvy7PEtb95WTuMAd46c
aZ+XPIB439jXOC5yI7NdCoPi3ZHsHzeaQtVH18heDocwwGWnSzz57mexyIFbH/gL9YAno9LJBgwq
SstLJ6Ls/4kzx4D9RJbISy8Ke+q371j9XmaZO/lPgXC4mUXU6cmxFu/5IvJN207JAh1fIPUwKCu9
JfQZ28oJUaltH6EOhNtdoefsEi4O2r7EiPEpIySXT7XJAqEfhd1iGVukAAPy6LOpFjnwOn7A0kJW
zoUr5nbhlHkHSym8Gumh9JlZACJ5KDdTIQLgk/6cNFV7yv183BaREPNHq3rb4doBdnXldWamUm20
U4bHuwWNRBD1IrcfAb/hOkEE7F5gvtsrXtkjjCIYl6+rH2or26GlTfiAJmTpmCotDS0y0JpXN19K
Bq/7DAKEWht43PdLp3Q7zL+za07W9LrLJpveQu6wQjCxANXYyFdvfCMZlF/KlVqLlaKrAtCiNQxM
En1cUuvoHvoj0p1/4azl5x1ChKkH+PLCLqkRDHX0QUaKuRnaL2Er+J06hKkcE56v4hsndNmBYhpm
8npKp1j/ggP6li0hh13kSsYVd8zdXradxf68tkBUWWkAH3fftt5Ww9nvj0IIn7LfWg8ZQ/JLhrHk
AJ5GRHYoWqAWD5niOw8VCMdDlR0ZeyMaeZWZyj2i3q0UcwupfL+znCyEPa3T/ZdgyT+XILN5iNod
FwjbsiB4SdSqTJ4A2uaKI0J4RJ7HJ9mDzKiUbSVUpgGUw7+VdCVSeSj3+w1uiBi5ky189mH5cSB5
Xj4dSIyFYYAwcwC3BgFLVqPu8sZt8sEIp7my0Ctfp/T3wRSq+/iNcvj8bd+mTgiR1r8kmVbxeQxP
sk4t6HeWE51Zz3/XlJf4Z2jZCkWgGqMzDhbgNgLGuTtSFkNwHojrYO/k6Xmixq5GofXDVur1KJfI
QUTbg+DrDAJZVbm9gMQMBGv8EQ9jyf5emHEG5vUormQHbOZ23rb2rgqZlR0U+SaQ501v4vEuuLJc
DOVjrZOjWkdQH7Ep/TXYBeJHRN1P6KlxezzAfQ7gI5xamitnypwdZ80+PUomtKfHr4Y12p6VM1+f
Jrp63Tv+oIKEYSUUfwc1y1O+jrffQkXdiuph2MSF912ecVLXksqGvf5VFYZEysJi+I3IEEqyKt0R
auZu3ieRsLmqLGadABYD0a9eR/+gHNbPayrkrY9nY2tm3sgNXOHMnI0cJy/c9wUUrapbw0DAg5jA
KUKq8swbqNExR75vCYHVvcQRdZmIM3YinZYijcN1yM9ukPDWDThqykjKb+CcTvktK07X5jWk+Y6q
nJpSak5C5s0mkHoHJF3ndiD4ejgxEPYKWvOal6I0azgYO14pbxvXFvaDzjW4JR0LA2ukGwZpdiIF
SG2nOwpDKWglzUlwQ7Wufa8AFkp+ePecgyD5V+9asvheLKeHYs4yBQh5DkAYkRARsS2b75/0TmMY
optuSXRuObrqn2CNXXVXcD3exzoOD2Psf2tWij465TWjjaU3hgExgbyxQb0PvptIQANJPJqSs0lX
ZnM/hP2eFTMRsdyUM4CsI8GROKtgKKQOZrGpTI2787hcTxqu4OhoiKeyDVlVoxLOIhP2w9VabuOP
te47juH38FCwoJ/ceWjN0JScC3MsIpBzAFQzV988Dxmc2kbx624yNI9LEaVm/IJTD6NFC9C5fWm3
o4O4P29dUSpYuLx8kULQdOc+j7DsQ6fE1ykt50k9myw3FogJU6Yjqg92GEjjSiOZI9otSROnb+gd
tqLkjQmlso2FHbzS5XYSfUgqjDWQeOYtxNjywUWgIxlJ9eiuIvvMDPw8QhbQ+d6hWJjtI7LDBGaQ
mzrGWRWvfJU07hqduulWj/fx0lZbPydwyTWqbaX8wQ1Exy6ERWPZ0NQLtW6HFlOmoQjNghzSxsPs
9dewWGblHf5uO2/ms83t7POZfbNHU556tHFou0NmlvCdArNS9h/7BYY4WIZf893HrQ4KT8P1tblh
T4/JkburaAMXkM6wvUtnNpuz4x4CIkIRiXvTgSECice/KEEzeCK0+BaG3nzfkIP/jqzB8ji4/WdT
PPErUnvCqNQmItrIszqmixwslnwAA7p7atgh31baEoggEPuQq9bfopblc4Gg8uXXXEQntylzEnjJ
Ii3dDrcMrTasNzpc5nAmorhVLITwZcZLX0Tu8KddfkpzFkSjgck5AsF9CKEehTBHWVlZD0IbuPSF
dqIxy6k+CtZ2zdjZsjDt3ch6tYvuynEa5v05PlveKwSbJUQKOwCORZcMwj3iHbgNzD43PQS58d/d
b9cPssQQf7mGRKSDxnV1OBUrX4NPKORIn/Y+M/Zsw3XGORZt5OE/p+f0XMwLdYqObZ0dkEu6ojB1
WZRbcdpFdQ88qQM2LaRbkCy/jLm/MfUh5NFEEB7OT5MyiCQ/P07a47+2waUdKB9qFFGwoVPSgeTB
zsg2pel8cQfUvVeT6ou1tJzFbozqPN9ynQSJQ90AT6Q7TW34imyPo7IbOm4ar+8+K74n11wjxMcH
8avAaC1dXXK420zELwqdxi6P+7rQ8ouWIK8fYEIfID9ciY4OfzVMbrJ2btYHGK3eEKX2pCjPnHLS
Eo1+spGfgqnktCOnPyyY2y2yC9gVowjkcDaMUEi3HhlG1K/EwctB5VfRx1oIKeaY2I9jtTYz5J1T
lWZdSrJVVfclMugKrLyAVeNW3dZq/8PdHXwZqr/sF0Pl+sb8b1OyS/KKwzRaJUHQaG05SGsRrrkM
I5y1qbDabBWZTvtR3fZfYAHVuAQFB7/WsDjArwawkNdMVxILn/r29dX+E5thIfj2/dL0rCVmT74N
SfBttuXqFh2N8djc0rhsiZ2ow1XsH0WIq0g95okMue8HDFHEK4B97X4+VuXsyRYP6vXSB8mzXq8Q
17QBW5MEH8wIXP1BKo3AqZ4F3w7yaJ+yMFRHtLEAS4QojSEpKwc6v+B2siB//4edYvGLEANNKSow
P4FKsMaBikrNxCYPFBuFpcxHx0eFH7rSp18crmKDl/SMWHgaJO4rEJ3/thjYNAPguAJqW8mS7xq4
jIlsRrbmH+Mxv38zMUIFbby4s89tNt0SgBA4yW79vTh2Za5Uwpci8S7cpntkgwyquStL4eBQWgVc
XiFk1cawT3bXKp0FI06efdWhpzjQJ7IQW6iHeJGE3zgPTkgK3dbKj5xCxRw3DGqlbe6MArbOlxDY
zbvpdMTBgnirx1a/EaBDVAJuIcxVHwPVVSN+lb/WV4h5cvUlngPjVOfAPBHwXb+rafNTlbSPGMD4
Zq35F7zUt8KxeF16cEEeBFL0WABXIoapqofVXp+TJSpA7uUMIvjK+emwLCH6u/TASvTNod0WgJ1j
4sywkOzDjMPWlTB2bf5RZL8aY9Z5rBZXBEguwq16Z1dqw8Xii5Dstf4yZJh9qYUvhijrt+t64d2a
Su7oF7Pey4fRRhcT56/OfqFABcVMnAPddYVNwATRPzC3FFvs1oaGRIJ1CS2eJeBGMbMNcvA3yIm/
8rNI/oxNHQxvlHh8aE5vKyHbcg9lDdfslasuj0Vyaa1XoAYd0GSmpKwyLWkcihHDOzNnBUZ6KtzH
4vZKNYdSQWTy3MaC2CX/X84sUtUqFqkihGTN1v0E4L9fVz8I6KZ1ETrQI7ycT40evz5lu9Vtc1bM
fpAzBZ929ajE7D+pZ0hDbniA2QwLvV3xKszUzXdRieByXCrMte1suHPc/udlBu+w7wAhqAOlOrkG
CUacuHbw75K28iKSMaXw4HbcNv2qiXy//uZHImGXDv71Ul1rXx1HrQ0BZhZAjOu1LYJxXUDUIqx+
U59UkbIJopIKwDeJTdYKz6I/OTRQH7euwgrJvJnKhu8epH4LilzYFsVuw0Of/h9nSmRtKIntTlnK
vMB69SCr+DSyZso2dz6XVa7DJKGMTf/W/Qcooz3iWVx+utxCnzt+C2cKdTa/varURfQPM1TJveWa
3cCAmjytqomOg+TrQPEhpIN02qtQwqVCj1Of3s1UGF8ATLloHjDPh1NOIe+c5Peb+c4kO7LLk5oz
+VUrhsuiag+/JasbvBw1wZhKKXtHzrUu0joLnCae9BRGcke21v+kFnddNJl62Pxu5Q1LCWRwkhZU
B8fMfZ9SMInOdOms0NHTE2Ji0d0g3WW3nLtGSxmrnqgAM+LJqfFuwbAOqI7xe8opFP+46T88I14N
ejCUTCP93dyuJh0sdTG1lDmvlAJ41wPt61G5qk0FEe+rlQfxwNI9u1E7MmUv2tff83lRjm7UJtpb
eQt01Dtjfe9UB3Mn6Usq4gX3K/8/2m7E6K8BSnLxPWZNXsVGV8J785wC3TurG9n+LWbJdM8GIbZP
H9LtZEgGkPYv/XA/mK4AePPLB8FEQp5hwWRSE26uoLAW59vllRRmxFFVHTFnexymp6gDzF/Y5Ygf
+IwRHtBdjHotKiC3FmmzmQ+mXPlWLohEQN2LXWRyNOCKKmq5QQIdx551Z7eyxavcJoGERt2ukNcy
oGfA3B+aEvW9gzlPOQTuaFHFVcFl9RDAt9uuXQ+qnQAazLVF2N/44vERtuFyqHucJJ164Md2m7lp
g2SHxVN9c1QWpk/HvvNnFV/yVvNbdAx/DPTGsbeHWAcujeInfhIa4Qor2rFpBmMH5ILz6bi7hApC
UzBjkTsFh6Jy3dpvmuNJxLzaaD03Gb4m/Q9nvodPePQQoZuQMk1GToXgp2aKDf73RmcTJHcB+tYl
wHPnDkIWq1UYjTft/11GbCCCyvXoJ19foolfgsc2oX/6TPy7XZRXtudCnoZTgIhTWPca1p3dGNWx
WBkm0foLOcy54RCnoiaXKXacU5yPYFFoKaIhr+9OQDkSHukbNzZA98kL4eFr8Dw+2yXdDKpu2QjU
d5Cm9e4f8cf8sFQcOWdsoZXCDOVRrXPqHnxN1t/Q2dwaVOr51hhvwdfO9YNO1jBtIw+6CTmMEKZw
Ec2036YGqtm9lDN1mFF9sJAdNcm/eJXSHTVlidC564gcEiIWBsVNDHEdNwTddnZkI7CAee7Cyt5u
595YP2QN7QBU6QB+xBLt/9kpCVqmHOdFrH9jAgEoyE5pZb5o/cPS+rKfbUivj+m5+Cg0794rDVz+
3wOvlHEcyLvgvyuxZ9oItu3DNTSRbYyEUDkD7+zqbggJuo2MsUtIheANJB4QTvXVLD0Hq3RX42u9
FQMhbng88uxNfWLABM0bveAtYkCgWUtEDT/oBwzF9pxjXJb5z7l8rIu5VqQHUNiuEfoEbo76mVQ7
Y1L5hw8cbwyjNDrXLO3i/ecIJ9qOt8bix0xs45U13jt1KKpgU07wOIRCl4EL11XH5uDICWZ4761E
CPHY8wXUaecpEYawqDp9xm7bIx7tLAuaMQl2piGaU07jZTPsLTooP1s+u7ilimTxUDg2nOnpTP1x
4bC/Zy7FhnKO1qGmTOj1LsrT1ZG2k/3V4iluIeeHVBWvnCaBMLvkAIUXmkyLidCHReEdneSgRHst
x11nuw8PlJaQSAyCx53nff9iAdSeSEdvnSL0H1HVJ8Gs00LEJBwM3JQDTgd9y60Qk6f21C+G/lG0
RhqobjBYhwLv0h2zZPX4Lo8WcjyU56/rQMHIpD1+nLUD/hh33sVmJnU9mdHmIcpfc7Sei9ye81hl
Amcb8rAIUWqau5P0Bgtd26TzRxDGZkqb4N9RG4Hx8wFRn7jP/EfCZsg0Mn69Pr7AS5dIlZ828/K+
E0LiPMMyy3JP7i4KDoC4wVm0+NSXa/DpR24n43McfKyfcD+B/+hAJflmkkTL/PMbrNAjHFLwPAp5
ah4sSAKDnf58gLLBFxDg5ACDLVwBqKXG3fq6MSNeoFea4sFP+SkqWi5kb/Fy6VEl0kayPvbbFmvy
OngfM6/Paj2RhjacAnpIiKdP9LiG/3IxegmxgS1OQ+0cLLZ8gZDKBfccBBjtpSX/gUbMrmy1OL7N
ZIwC658FcGzKgs86YhI24+t1mxNIpw0fUymDtr9iczaHEgq3NniuEnwjIsJOD5c7F8x9dL3IWFBD
c1LwmiXGsKwFabs5tIvZLSp6XLxieskBF4PMxEHeWzf8H+zr1ZHVU8mfwUi/s/BAYXKeR4+BHdkc
0Zn3SiIiobuDMPPg2hCSxIC65b0qKsN5zXXGyrq3bCXr63xViqCn382wa81Mg5vPPHtumjtu80Q5
p+a/ooNEdiv/vhp8erRbWcMoJl4+/6LkbMAGJtSaU0jXwsKuIBIcJP92CNn+7mmj5+Yg8Uq9yFO9
IVATZUi+3Xj2LnhbdMhbpOz8AWMZRvqwKKrk/TI66CuvbrTsRc6b79UQV0KjX7gr34FIaHXrlZC/
n2rtU+E4cU0c0Ndyh1PudPdP+bUNzXJl/msxo0aLzlRavVc1SOV2/Ng+UH49T1i64/ViHB5DU3uP
vsa2OtD0iYmpy8eXMTNhKMmLfK7eRiR/zBWyzcBS1GCUCp8+KmZOiv2jNdzCnl89rQznSkBzG+g6
R7/Lmhug3fEK+YcjsChxZ6jq2jehwOK6NRv2SWj2RNzuHAhL6ivf/C6glBHe8vd6qR5bi/FLiEfY
e+EWa0tLyOA08cbpU4jJjbNM5s+CcQbkhyEEU6giAfBHL8jaroaQlQPDtjKGYvSvy0jgpGOjHQuR
tYvWTxctpysHUJ7CE2mhA18v+ylGyPYauAUj1PnCoSrA7+7kdhZBL6UELb7cO3eYI9i3JHGqRCgc
lkOcczWlSLDl4GwLaezIGpwu9btDz6Jd7qs/qBHKo8LIOKUclE/1XVKy6WbkPZuSJpmRYKnBDxfs
c4gAGZQWcTtdjue3OlGYO49cvMSiUJp9C+aYIVaOOsHoyvjlq8e102n+DTfIFRV6AU3xQGuIo3Fs
BGoPsdj7zj6cHDeOAgmQpwa/GHZY8z3ifv0hc1BG21Z9nQTlnEW02bUWM/Q8ma1xVZl1Da1DqnvY
A09wasgObj834EM3AlC9f9A5gaguuse5NFcntIaTMG7k2zGwQ+g+lhzIXWw9YhhyPCrFC5VQBtqw
uNyY+j7XCPBcq6cP7LQmRoG6rqnF0MmlfudTUPt8v82RgtIpkxO+1ezUNkAlM1TYrhAebgt3iYvj
n9tPavYU9dvltmqfIuLuvuRDkBZdoRuLRxbZksrlUQmcFc7moVYaFoX+5Xd9P7pyBMSNHsxXbavO
4wWL+JlU0NA2fYv37pf4nEsnA4XXg9hK1Zv19ufgZiUsuBnOAG9xipW4bVBtGSW1CBc8OUc3BOOb
5Zs+fiH8bpzuhKvHa8sdjTNMz9zQWeim9e62HfWET/pcVQ6b2mQpHJ6ryMlKuOLkqpxxc6VDAUvz
lVK7OKamh9VtDoZANtpbDKnD6uaqrxyJtAQNr2+uMptBuTZI905iXdkSblDoy80vm0dpoDZVVeeQ
APibzEB1WtdZjowqnx+GsZu7YRNkntorQBdTQ65to7Ftqx05harfsoR5jWYquNl3KV4JPuZ/yCb7
gFICp2UJzKIi7q5JSriq/yhB8jFosYoy0c91KXXCvyeRjL447qrvhe+u/FZ6hDuT3A9R74iK6mmN
Ykuux7ZOdR3wSZKqwnyXxM1NokzHzaAoXuks5Enu1AjiGd82KdmdWKkFug4rwmsXe/u5fyh3vCwN
oTsK26r/uQyKqCVrO0fnh2cmUpp5qIu0dnK7L6uM4Lll//sMj+0SH/zEnb4tsTOe2PeGpFaBTfzO
PHwoSXGKiEdnLY9v4K/AZRXiTYw460hRM5I11XGCvu6DQvyhS/lI1NKiYDsHf+bmef9bREhs6eQU
CoQvOH4nvAwPZz3POofONO9AxBC6K2J5PmdvpZW3SHNRaXu8z8AnTTWhcEX2yRQYxTl+N5rDP5wq
CJbObqIHBztKA58bNa1us++ULJQ7YROdTHc1c6HMUDIAT2EiPUTTEVPUIS2PIsk755Ec1VFrNWZV
I4YS6dfLnHHWKq6HsjlDSHGOnUBv9c7edRIpwGMd3Q7duh7E1tGTuq6Lo4Da+MbUoTVs6xzV3Fn5
AlXWNmAiLR0V7kxOerGOVHmqRJyn1y9JLUSQ060VzSgWVSQlTiVhgPBauTfLplK+b84N47W//8v1
0MiNOFGsH274DVt2G7Gyr+2OUdfdgNPvOTNSfACI9Jq77qZLxCtKYK4HLb+eFRagEJr/DlYPhF2b
72IQ6OvA4L44ASvc0AyiN+ESwNnc8S785C8T/1sYsvNBCNBpuuSNTbJWGnEnvxwDtqttC3U93dre
6hzTkq74Bz5KCV+h7PXFEGz+xJsF6ycDyjOSMXuJVsIoTo9Q0xgte8FXBOKCzfrNn3TFT8UGxBH7
fGi9BPnO4TO16sceAXnlXUomcbru7m36gbKFkaBGwlQhYZxmfJpUhWINDfmV8eyU4ZAQvu6wqL2l
YGXrxn4Tn9tIu/ViSJc0aw9pAW+eGvcL5+UR1foEPJe4MNCZ4Yg6P9nNiaGZw5xuGdiKjEXmWIDb
YEqLCqPiMeEDV5douMEmBQzGEMPYp3Y2CH4N6h+QLVV9NWW+O1brZgMzBXQz9kzCBbepnGYiOXio
pXegVgaPpfU0LiPB0P0oOpv1uYEubsPXFRlzEMTz5XWt0HW4raesnNo5MvwsNutX5jQr+H0Qr2CG
80c7lnT9PRHPbgZeNmr+caoEtXZRoIORJqGUkMknVnouxcSHL5jWIBTM674+n3vLRJhRgdgSDpWa
JicVh0gFIRWSl1FQGvuJIAyiALU9OUibHAmoD7nb6YimZ5uvSXgYIs3J7db3d/oxGKdGASlFpU9V
ti6t2GwXoEkgovBhsAUls35/FwuBMIgzAelAHkx84DnEcWWL0e1dCpsGlKTLGqqRn5/tZzEReFmu
SNFaDc9jG5i8UkdGxk1OY+a02uLEG9iB1oUaA+U4GRPuU5UhflxNGb36Xmn7Ta6mJw2vjP9Wmqei
PAS5Z+Gc8CgIvios3qwCp03JmcQ0XreuK9DO8XpB1LPle5+SY439BJXLuBpyV2BpvOlhSShf/MvT
AQkNQGzXNPYMt060JWpos29hvqyOfP5Eg6cZRzFTb7nzQacx9OOKls1VfzfAncE+Xf9TQyUpVaaO
wScNHBZuip47q7aiyZ98EpNFfMbRUdV1Zv0GbWbR2pwg8Yaoa4viV8C/QDArThtU5M/hvVAEju+O
Dti9iMpBn8a9ksK5vTcBy3mmaJS3MW+xVk9JYiW1wbvz1FiXmWsS2Kbl/Y45w93FVq7AZV8hTL8i
CJN9SqUiSOPPwl/Wjx7vmBYSqqjOK34NqdglGGkwm6sWKw7ZpklkaIUQRt2t7O/6JKVEwsZ+0bjV
93tertaCpyaDGcEU+j/KMG+hNqjI+WQB/bB9OLJeN1Xoot6MTaFE2piO3VffOq1mc6hXfiqFEhvY
D+f65HXNdlBuUm83LpFLqZv5IBF01hHpGW/kzInHtr5QYphwWPCQMFFjp6WL59m9so6xSq/tpMoM
b7tAhJzEZ218dTBmno6Iib4mC9bMVzUrCx6V244YNzzJLY+U8eExJNL0FDM6bMyKI4pDOZ8ITTw+
F4P0UlDj+AWX2uR4e0TCkaB4PhyAoLluMMBPQBUJin3bV/isW0QaHCrAeBfwJAVNtRrYT/yJutxP
g5pZPqCb+m9hx7W8m/BD58AdTlKD4aJmG6NJkUo5GGjdjye7eB+szM92oVRekrtFG1uk+X0Dtc6b
Ls/W8Iht/fN38Px3gb8JnqT0JrdRcFrZRlPP3eThB0vjqZtoEsm/u4/O8WO80TSjXYqiMhrqni7N
jT6ybEqzahSTOKWNTuPwRPq3TPC+Gs+y9R/bJksWYk0nQYVdBupehPU9LvoWDBfTUBzvGMb1uidt
RtmXKHmjL74G8NnDmi77y005PbsCM0xaytazNqum+JHtr/K6h8M6ZxxIIPvTUi7NdNQVJHqRnMNF
ObsfpWtAYgHssnmOS+G3Lh1Va4awgs5E/2DLUWUaXu8TBPp0k0jCWIUTRYai54sLB3pUIJ/wU7DM
hUm6FLj+eba0lRLSbXIw/L+0S+Q2YwgdtMallw0LRXLyz4amrMMDPExMMJB67NF0iHvwv+933dG7
sEqKJg7ploN+3JNWIddNtX75cH9eMHeq4u5/N22F72QgX0zJSI03CN4gPPvkwn85gF1dB38IcCjm
h3K6SCx1bgBZQ84rE/yOxqowxF1xpexU/iT1cnjoInwIjw+dheGrZlxIOQsKoCJ5D3aGKRkonMge
TCsyJiK/kE521PsR+p+o7JvWwAmqGGdTVAsAbZMXiVJ0QG5wI5OC6cDw1P141hlVAks7KCu5Z3O0
Y/Ffanv2ooqIPA1bAD2yjJ8nJbQtSOXmMxu6+waxyqG+iI3JiR8x3XA0YYFvFZapfBz1enHx5Naq
Hkcn8xM+3h24zoSaRNIhNLOVDDtW80xX5HLrcHA+oUeNESAZgxcMPypenIxTmOeOUK/Nohr0sCij
ZkbbeBM9GfUAp0LQxgSvqvj9FPjLqqivr7twwBUQ3MdVnUVMvOj5lrGvfHEn6iNR9djiKB1Cc3UJ
N9ITm/LiilGcaRKvrzsj381AJqa4kUFCdV3oD6PEx7SFZgt37mM5p35X3PglGm+KhuZRiTss98zN
hWEIdSyZIU6IGAlPBy+0q9rTp0BnwKrgucmckYGsaTI3E07Yi/+Leuu/PwIbsE1uTuaMCmUy73W5
eyFJSJngokffo6ya5nvSmwO2Eh/pEmi9ZGctr5c75u9lqDbwlLJZqJ77xdSnWgV04WrglJRHV2Ay
QeAN4aAAeT6VHf1QH/sthJQtlEyhn7DO5jBzP0l8DCdTgxD3PimiCU7VqQGthnNBZbkN6I/RXw0m
+fnVLO+4hS65CJa+u/D2ZR0kuiSRzdzjqEyWQ2AADAyivnJIURmQs0Y+/fInKnOfr5NiTtQmi3Wg
o+D/TiY7/kH1DTR3xa+QnMJCS+k06znrB5lV0BNpiWOG/saRrxRyz82XBFwzgy1TquPpYsaMh1es
g2OFEqT4TpADnnXs2MsYm0mbJQICZY6goUrKH9lSzxaFr6qGPfpYu/eVymE4vG6Uju/WvzAuoYT8
MNGj9mFtHqclcjClZg2gKRQEA4I3ibusN6y2l9aF5VapM4Im/b263ef4PHLABkbbwbrE6MvRILba
vsyqWpb3bz2BuPp/3OihjY9RC4B+dxnqHIxuCjikCizo8A95bDqRND/jP7pEUMn1HT3LR5ydd57w
qJrwU5zH1vZ8cAc45Ve8fyyk4tP6VLd8+KdA/l7Rw5lHAhHrNfz2eUIKQ1aIwJLG7Jr2S+oht1kw
fF1sPhMPdu9T7JgSrBDXkboK0oYlGLxa3wQcct80oWK9ysiQEOhr5zStMw+FVsg7+RQBNc12k4tB
833/ZGPYyuXRjIZU2QmyWQKIO539AXhqXyo/XDQqmeUOzTg92PIq5xvMNLhyuUsFELaUr+cVsm7N
GMU8uzkq0DBCY0BzmWzmMTmBzgg+O6zFKmYpIeFiMGOFlexm39sXcW/QyIpFLq/10N1gorJUoBIX
2xIPOUb6X3Io4rLf77xP+q7aZelKquN7vl4BrSjVqOP7uL4i9d1iqlKSe8qrqXl+SrgCazqdvE2x
MNhK9U9M7o/RUvSzk6sub+06yWTxwHz7VooYgkKMbv2/qH8wOvuGw6oRQjtWWCrHH7ZPGxlgtuwa
MVF47NU2wtKzgsg9Rq+RbvIrUeewwaYNuD63avJIgDU9XEf5lcjikepXwy8+Y6b/CV3wal9M7uWI
MF4wkeRYOeOwwc7CYjs73AeDocJZf9GjGpV2/hFvANfV6gtGJ2G6iKntnbe2LCWPw1W318t4NGLv
YX6RYaUdN1AtkHejEJrxtEgLWeXNuif56p2LbFWDEuOj0ZUuaX11x+HLo8tHaDEozD2jxnh7Zo8U
w55LW1+ddUEEa6QI1Yu7/0naNNkgVpy4seAhFu3Hjn/kmlTsUqfgeo8xIlh1ehpSh0qNb4hdh+MM
aAISZT61WVkRfqjqgrlx0qLcper3pSwqWB1N8iYSdNHeaggLVd0Rouw5QlmB9ISpOSC4ROqu0Esz
qFcDQ15c6mli+UukumRDunba9/IOfD9adAnFZ8bnrZIcWlFpqHwTEe8soU9C6jI6iGyBCjot8Bu1
T8YwtjkMm/BnRLSgInruNyzHLTmDSV9wGc4QWt04vH4LiXcABbZnyG4I3/syzpeN8CVTJ6Enhdqo
cE+Z29z+AcjZDxfoIXxTxPGutiRS7cLpEjVXpr9XD3lCYpEv4G6dMtuk4yLXjM95WqVE59BRJeNC
lvS9PMin7GyrA7ENCmfVkNZDId8Vfz6ZUEOZnS3/BNPjgejyw+RzkZHWPlXBcVXNgkKYDuJ7i/3H
dvtCm8fLUjNVP8UPi0VlkHgFOQsXeh8EzhOZSWPNOF6koA8D4ElF79OrH8iQCc+ItkEqSGeNS/P/
bFxPTlZFGQiTW2DUvIa+FysTLx5ZCRictc3a3B9JfCMd4zuD17Gn3miU1qoi7uuLHEgzR1NIt/ei
bw1qL8tHIVMn0XtaTKYnJeMDC1km+91WBFlJTmWZPxbdkhpFh6Q6nsLBFxNZahOjK6znln02boMx
ZmgEFQyqO26sJ1TqwepGM2lFVf6bynqxEIGzIckfdq1Tr+V1MlhkMAuceyqp3PuuIcLCts5Iagzz
4jvdR/6rObV4kd1HfYrQygydilHYoSFUh1jPMMwdV2FGDpFERDR2gjWtgOgTQM6/qJwB8eX/SSSP
jK4rtnTvTA8AW9+I1vpQRPrAaMGIyjd8K96/IunBreGsY3HxUNmIiI/I9akP/yajCf6ZEz0JSb0Y
JPiMtUUkaGdxlrKzghty/KbAlcWzdaKZtZoACypbfzTyDCjVd3a61f5HgV8gq+eJGeYXNkVU/d6C
ijtMHQmzEJ1Nc8bMw9g7jBDiUbNx+Yeei5YuxKdUgAFbxS7q2sNJzK1KU9jWIdpVy0H/3U722mtx
AjoiivjKBljiYN52roSlHJDa23LAANiQaSKer+fQ3arcLXy97NV2TNnVqit4TBxKzsolrSZG0+ay
36jukUinUXIm8MfRLUhd/XXNOrOO3CcWNMnvLnkweY1PfD0joE2SzG3XvKRM0cYuRFPWzf/GOPzp
2nVe3UGC4OmWIPDQFOo3CEI6Mpb2Kq67ULyIEnTZ1x52t82JXT+tVyD+YsKbWu46oXfEfVGMLNwK
wHnMVJYC+CxnvhNwWZtSkG8h/G+G5eaRYgJS7Q1703ORyifaicbubzVglhLa0Jqi29hNI0xb6MHM
95Ztlz2OuOHZ8XjWPkvWL4KHVobt0K/rCB+rkGaESEkVXyJMk3drpkI4G5xWaLw8DyXObf4GCkd+
3IPhteCZ8TDm5h/88QT4ottT4nvug6aPvM3a9SliFZFj0fhpJUF1XLYEX6kVKY9tJDXLRNAQAfBz
yVTBBVSgf6WWrlUATJJ1AlwO+D7XxmkroZ9xWZgL9RUGlp4ioKnjoW6IxWIJFEVbXmlLKi3P5ilU
oS+KmFnphoQtDXuR/x25TEw7f3d9x1SzbeDmCS+rZGIo2p3ZjUJY77ruKFdDU7QBZAimctYXeVzv
tnht/ucD9oc5p8qjpbqnpGAblrT2ix8DsiZcxNZ0LuqA3XknqQMdBBFnPx0gm3J4cZfN7yex293f
P+4sxH1R3oustKc8t0uPJ80I23uD9Za/dWD7UNnE06sfCtD+3ZUODB8qBydqKjscR8pY5Q11gabn
EbOtQdkyRjg34SkcnXK974yjIzzAyNCN/KgL+n6hEShu+s4Qy65Pyp/VcnacfKeeEPWHwOGMYWID
Dmkj7k0/3OD9icMnCfFEpFr67BTos/1keI5bG5oD31DlofZ/nyUcSeQ3OtSUt9D0ZwyUqJAF0MqR
cUwAr39hC1ZQXCs035G2Sk6MOMv2hxblyWBgHlpr4AAmcr7pprDsYdvRPyk2uLrOy4OM+I8ggk28
dceVIayvCQ0Z5OU98AKv2bejdfvOXcRPQohqlHmjaxwQsIB3QeaY7b85oQWvpKDIOQ9HtyP9MN3j
noBxrunwtn6suSo/seFTVx7RR7D8YQG+Ol4hIWNXJk/F+q+w80LDeUGBhwj1WFZvIwJ1jhqNtLXe
n+4xsGM/S71Q5QhUS3S26WgALhCH+6aSZhBUAjnMFs/13X4d4MK2jom6FK9P8YWjEB48v8S/pBYc
hHzV1dS7RXSS0HmhA3E1Qp5jf9SH2NjdcSoMJp0V+Q7JLmayGiNgmRxl/GMimuTsn72B8zov2dzx
ixmzlNuoy0Az18y/2QtG4vxvivAtgCVxI6aTRT2LB8yWP+BIwFYT1OaLqqZs9leDgCHxMAqcg+nv
JEHKFqj2d0usXOmdmvYfr3Z69NFs5HSw7Xytdz6ahYq7bknmH0y5u1avvENjhCTHu/LHgtpypPer
HETqvFLA/+3SNV9pLVsHpdkq0rEokJgktqkW1qfIYPuqffAuaHYe0OnzBERg4Wv6chKKPv+AAeYo
VoWcmjU8fNESbTs/yRR4BjZ1T2ws6nqhqtvWrcIBgl5LnLpCYL5e/sJpzpsPOYvqyIu1c9TN4bBu
J3vrYCGy67ueZzgZVAceVrImdIVSfwINyxJMt5KyOROIHF2ExLAGQJd4QT0mhhTTL1oaEX4aIw1Y
xqwFAtnmd7Rt78pIzW9QjhqfIOx34awLu/m+IuDumrXAZ22wvcv+b7FAif46GyLm7yAeElKpfiFs
VgW1ojYm6WaVKQgcNwrNmpqHv/9yRbEZAGam66xWfTF4CmdwqUbKEuN8TD2q+YDrlAFbJJzdlJWZ
jyneF84sZw626pPhRKrwnaSt1EmU8WgZmDINrgmlYBNk3OutH1yEs9uRLl89Z6VnCZPjJW+pWiUY
yAiPmiWM9ChaPxG9tpHVcOwH/ia4lDbdRiIbd/10eDztEImkjbdYSRY6TQZc5Oc0z4sMe0cL4YRw
tKfj/o4xn3Aixxqp8MGcp+KZozhtuFS+hL1aRfPAZtO7uNN5RhwyDSnGbVtm45zZZXizSx/wnBfA
tWU728CFVpnJJOOPd0EdQlQLw09bM/t6/6+O+J+WE4iUdLuR0bXEg6L+0Q/pgX0gCfTduoG/Lj1u
wvsz1+xFcyiO5i5tpxSFAr8yOuPS6T9TS5jbN5pttuiDi8zdVOES7Fskt7UrZOaIy3rmUK54dWXi
weqo06JAE6Gv/WS4DP5a7DId7QJUTU6/hiYvyoKjSXUV46/Dd4SSjWCtAUxbaz5rDnDvmvhHdQ2y
5em+M4kh5SQPqfQuRa+OkF8pL4uWOBlI648KDMk93IR6TFX6FMnqTZaClgImJ2CV2n3YLaSN3A8u
IgGxUmVVRN6NoM9/e9mYpG2TUx6CeahusUIBougyZCoupy0n6xJ/imUNUjU+59ETwdkKYFutxxYC
YWQZx2RGpY6xlhIaXHwrhlwnLNi7PHVaROnYYJE8CI1Py5+W+qqeHacYJo6OMxHcEVuwKqvIO/1H
F8y3RPi/gMcdbMvwUtwE0dIIfDR/x8fayzL43zF10/eNcJw+yjdiGRbT3cUWZ6gMYYTLUP+1OySc
//1aOiXiZ+41U/goeovsRsDHUKddKwWXLT/KZVeriUD4wgxF9aHAcck/K91enfXtb3FIMGk+OQJr
OkcQw7kK/NuumEGNY17fF8inYWkOiN1qa+cSevnHF8RsYqo1joRTRCC2AOVBFNIkRY0G/1pHS1od
sd0y6sInm/O1OijaBJDOkD5SuYgqq4cqh8Slk3ldsRO8Js9h9U8KkKxv4px9cJploBHcfWi0Su/m
nw1eD+8JcfIoIehopvIOZo91N+0l6e+rEda16gxnam426yWWIyOKTXj4SM2sKYJmDObjoxUhUNPK
Px5EqdOEz0aCfBrulNsX3YAI0TWQo3ssyDjRWcC8lhbsZZ9zCbA6bllvdu12OI6V+jArTOxL2xHv
PB2y7WM/FK8za7DvtKd4nn0G1p2JQgaGfGu7gszhZmQq+NrnK3DDxcbO/NcPve0CGLwmmxHNu0G4
vQ1EDEwgmg9uCr7WlO2tcRF3nqPVDH2SVClVp8bof7mjUOE47hy0VWwAJzXwurVCCvZ3JVNujWUY
YVypQGnIDRyAdSHRP+EkMP1J0mpdjCGVedu5XKvsQobkgk/fNEmPTp/aqiWc5jYIZnnLsPBuARGf
kp2USfLH6pUyDS5dRB+Ka0Ml9G6rA/fIktWCd27KYuLZUv4R6yX85rBx8fxSjNIw3NNj8w5JDRAU
ZE4CmwVezvPkOaXNVdzOq989JuXCMuWzrCIamjrMHxgMsAJJYvA7WDg+Jk972LyYlehFVYdfEGQK
2j3KD8OCml2XOtMW5204PYC6b1NjcOQPTtjsd84Bfy0EWeNNYNrFdp5ZOqltsQh1klcicg7gNqAz
moRtIvQL3aU6Tz1JZhMslKzqXkFP8OCJY/+CMM8BWyLrM3Bw93KuKeR7Tt/Wrc8bSjXV/WXyJaar
23cAztdN+9lr8sibt+BUvgGylXyDX+7M5+0Yz2BfDQKlAyaFAysfVDwP1WyX4R4pd9Ukpu9pN2DF
cNY/hIowqPdqntTT9XVX9wxtAItdkfl9iqlzdwYaA9l+8sAj22izSnceWzlN+DvHj+deUS8MNeKR
6+3pXSnKTsi6tO6OOkdBww25C7Kj/nI8poFOhledWm4sWkLVpvqISAk2E/b4gwua4MhY1pQAy4IW
1Cz4V3SFFJvbIQUnfcUtP4ptsRH5WGP4Q7Vk91QAQr6hM2o34onrtvdLvpRZoDgQUhBDCS4Bw8rD
HWxWIC0r8C0UPD2jn7YL9/ZfyaSSXB2sm+a0RRybUDrwESvkse/79PcWdd3Tk1f9NdtIHGkBR3cq
7yHCiZXMB/M66d3QyipMRudzRQJ5fTm3abeLoL6eDX6e5pJYcNh3UHS93WN8/P67W4hY7caxguQw
7+8RehZcyxsWJdD7rcLAz+OuLUEW3hQNlY6oH455OAdOAUvDfSX1s1KQjfUjqhfJkT84rpp0lFvL
maR+5juDn2fdg7OpFM1n0jYw0jCr/9k0t3j4+J5hcaw67e5O8OwDAzLgt2fKcPUOQiWCLhzS70We
xmoRsWZqDoI4rR4QUJoDvPDwfzyeaLjoPyBm4l5x27WJsUQz2WT/K0BSHUdqEAzpXnaH4B3N7srz
7hJq7nVwZuGsYRQpHj/YeQwphs1u6VVh1NJNgX73ePgRJNG41QsDvVfrVA++f7UYyaQ3mLTuRFNR
3b33FO650s12X1IPDra3qnfv8XWB1KwG+0YJUidYrPfRahMeBydYYI2k9bRvTgAZCMwEE/TGqQV1
eqIuJnFwS2AKCGgzG55XMZ8ejTJaCTykeoptNYzNgec/o9IgyWRv0bQYFzkSqa7XGhrXN9RWSdL/
WB5aR0UOcYI6DDI+Lvl9fty87tZPcKr3tlhLQqrgb3N7wqr+vXmEi+SRKAJLetu/ND+NdTPuhLIi
SC9Zg/84JMR66f3J7q1ctOAnmNcDxMQ7QAEQWVm3xJnZ31jtVhxjUMBRB6V9NZc9HSrtBaryiYRc
+D0Z9CAT9PMiG7oeItvtCWRWsfGZ2dkQEUuWNrC4UgTK8cJF96GgmRBh5UE5VIn/vvyPSBcWtNA3
P/h7eRUGV7jeS5i+loHoAnhSiuKNfLtHYHOcciQikEwVVeomzgGi97cJuv4QyQO5NGFsaGHjh59j
7eCEhZC8lTAviA+g40XDUaNICUQPVzGKbjQUYl+Ufri2piekviWXbHXXwvs72yUkIe8GRuK096OO
OmsE2tn+cOgmCr2G2LRHcE696VF9SM5rQSJJUuvP29JJTbquAh+HxTDh1sfnRv5FZCCd8WAXkoPT
QGoEaF1mEjTKGsKlA/QyT1sVP+vl/sO5MJdTHs9k3baOz65YmL453eT42IX4Hn3wvzcArhklug81
JddGEBL5gcNzr0KpQuQe9CKbQ5+KNqidLdpEl9tnu7UuE726+hFSeiXOUbNWwLODU5EP47PgFBb4
rzDy21ywRiPXN25IZtekkCCgzW4I3Qs31P0rIe+0MPGZMAxn7YpBp9wgdbkrum1vYWXxct9nSXV9
5HJX6XchiYHP35Wl0Jag0h+B/GFe+HnpOAOGKsXFXqm6Jc9CdsLtS4FsnSLnXQBcMdEycbMat2Cd
lSKLyLpcYPD7iZ1lB6N9dRvbfAsjirJiP+mDmRbl3oA8tfQVwmnoOctm8J/mZFApImSG4Air2oPL
4orixIKgEQJKPX+K+qXGPZLvJ2j99lccY1QPL+p3UrIut9IM2vkMPtPiT6sQ+Rd57PfAp0dcsQHC
/NJGakn/eGzMNbInOJLHlsd7MCg9QIxs3K9qVQMw0n84JvjVGpTsnVAaUhXilmNKLWjoaTAncTiC
p8GkGiqlJBJhWoCKufqJb/6FnH4jWxUrdUZwXiHhJ7dJWMow/UzPkV6dNU+c3qInE4ugNjTKdWT4
qVR8fYULU0xlj5VvlgF5Y+MSIxwqerWUQiqbhty/4NvYJlOzfPAobHIHiRZuQV31C7mmyGZ7ejkM
jE6xXaZW4TZwwi4JDaMzE3luZOnghEK6rRnzF598+7jDeK41ZDZ2x2Lq/HDLtO/yzva0+DMxNlKs
dMB+SSIGx5kxuTP9i73isqs80Q6ijU6peU/F6NS9riqJHBgzQ6dVlg6IGR4N25T3+oDSvwlNVJ/6
f7YIO4t7UuAOUtu+PAN2+/2nNocWkuFbR3M3IWyfxH5E2kVuO696sAFU+/ujxjBMS7vTSCfFlPN9
HYEhVDux1xFpoPFqsqtR6hS5rInyCe1H2vBxfV/gUUfh9jN+GxWA9ReqVg4viJjCtV7zi9bLN84a
858LwmOYL/CCkXanKqvfVAJyLVsWvgq+EtPYEInL9UttozzM+QUkhD6rgs8JA4ttuBGRNga7Tzxz
Ytp9agbfcJLwZRS+fcDONE9nR+4+GvVJcYsEvzP34KwBBlgaXY9xGCQf79lwo46k4Ue4LbQTFCzh
A/Wr+YFvNS51o+1g8zgfpdJk/FUGSLjGn0Mi6OOm/tw+N/0SnwSG8NeG72auujj2tumWUl77v3Yl
uquvVlwy9zKEUb/PIZwsiJTmBxC6OHrqq+rjVs/wyI3W40CgE4fTy+hwMWIploRv0ZMYww7ByzJy
UVr7Xzlf9A+O3rUoaY6zJ7j60QTs/H8dbsHgTa834Y1dAeGkKn+fRIHsH+KJOBWs3vt2oMiBS8Eq
UROH3SKm4QqdV5XIMNtJ2Ku8WT0qb6mRjmhJrHHjCa6H7cNA8ucOF3TQa6p+HoG465Fy8QCTlUA7
VIHr1R5sxUit8H2dzVeu5V2h7Cq0k0dBd5gf8IUhiX1zlSvb5NFZbK3A44Qq8B6AK4dEufxnejfM
ymU2cE0GD5L6GEx3+m2zyLgjsfBPGTp4DUtCszTs2q4JE6omx0KKXwUOGGmrln+cZnD9gwsgl0Ow
62m/MOtKR4dk5VIKBvyJuULX1kIlCGw19DLk96tMd1F7y2ydzOMkzkeBZoqo9+cQUszNEDGxQpKV
XkQY1LiQuTuOALccRcVLFktnhKkIB2NAwXYV1TucpzW5UjLPrT58lHTwtGE25owXXbwrDgvB0Xgy
t1mwmr58KEiVMM4iaiWxN2PCQNOCRaMu3T3V/2wS1FJ8+XfD42HnkK2C14VwfII/EMpy0q0BIodb
xkrZkfT3oq+eIdle8XeHOseUFVVnSG2KIPwSDJFNZvDxDfnCmw4vLnDeoYD5u4UoN4mtYp0Dmn5G
nqHeS7GQlurTHDCzVsWOgGxCbJc/ADajtXKgZZtGiKAdsT98jrucit8dwLGI3TkqA4LILVQBf1kA
cIi4g2xwfO/tLG3jyYr4d5ErytIgZxDT6nEZyE6zqU2iybbG8IoSPkZ5Qs2hSOB3bKx83j42qQ4I
sfP7qbG030Xn8P0ino7OhupxpNn47b0EsxXhWuCckaQFbnTc02M2ehmQALYX3D3qfsnruphcoUk6
3rcww/iJMCBQMal8moHjFxChp2BqsLP1c1tPLefC5ZxUL9Lrcz0zY7V2oxwbXblljU398owqAIxL
M9yp4zIsZSdj1HrjeDpdihZfAQ+g+6w70f6/x3JhmckD6aMx8oBiupbR9cOaJtQ6qmUtiYK7sYWG
ze+1wYvWSuUcF6Y3JN7z8CUZu00wv/VC7k80sJiJIKGb+msy40Ex1PtHT1sQSIA4e5DAFoBtsoPW
ejVSMme1ohi0QL9IgdwGKF+ZUupdqaBkSSDscW5PUhlv/59N5wORxW6bqhX90UJ6+ia8p35YQCdv
EE/NTV8FBs7pumBzPVlCFxGeVG97eUPXtsoyxUFUWf+mXChvGwB5hE43G2wb5+bA4fenQygASBXY
ZEf2QivQkCPr6tX8jAJFYjaEb86Wrq+PfkY2MCCJvlS523ki2GHhqczkpP/OCcdJVpcfdC+fQBsp
XsLM0PrB7Y4NAxmt/ejSBkGHcu5Q1shfUrQ/wfLq+HeU95T7KmeJHildkaFgRBw2cq9bF/U9yoA1
gUFxlpZ67jCX+yNleiI+25BUxhdfLXMwfxo8Y+YrDvGV9BzGTopVHbed6FoI9BzFHtIQH0xdqUIq
XwiLT0/3fVG/6N+PorrhkyRjhwnY1tFgqaVMTp+ibMMNeb9TFP14xdz4/qaYzg36mpc8qaN8s3FF
u42uNFqHhUBZuLUHWVrTaT1RJcz6/mzV1O5OGaGkiux1SIcontT2Yu/8RXXS4iLw02/fnh++Lutn
tScPJ7HQ3SZ2zdjxHFc8Svg18fNoUR9FCEIfhhm1ZapP5YOHgXmbSK4e8jh6zxo7kyIOhyQwyZ+K
MHJTHwjWbI4N0/aSYyw1euKx6ZNDGPuUrr2HkvsvY4Ptwj4OOMnETXdHSJ3pngeuganB01K37NCE
ip0Ec/z+NnZ7+3YOMAsRXOBw848oqS8zqFYVNcdtkIMucfNhhHaCQ/smfvCSL/vZ3Pz7trzS3bGe
UxypsfM1LVxadAB2LZ5a4344L+St/LznHM/ORvzDZkLmszPG3I3b1ORDc7Brg8le3u1zrKvLIiUr
PApI1LGg2GALuQFbGyK9Lk4x5LB6MepnbZok6FLEsJ7yFCH0qiNdHK8mthW3v/9yNx409KP+ZeXt
a3epEEfU8lQzsrcwKlREAt3heTYm7FJZF/nTXDKUQBLai8pe1k6f5Mtebnn+cPj7r0S+NjcHeIiP
kyJ54iccgPf8sFwwXg82Eo/1VoUgTsj1VXxccEo8bStVvS2xE/nkhmoDXiRkQSmrnOxJU3K74w0p
6i2DRITcixPuS5opC/BUzHtlg9sXOabH3v68P8e/tEZQ3QHodL5tCKG2RdGB6W3DQVnXWaCZqkdx
dRcg4FA9poaBluT556RcEtGfZDw2kn9dQu7fQR8qww/6oIxB6gHK1RvK+uexyoer9szK0to5mFbH
8u6cbi+zYtKDs/NynKjCqimJc4AXnqA37sSsaW3Y52cTeTJWGgjAXx0cz8ChHIYQQhfI5Ul5w5RT
+om2EsMC9U0EeOQjYtoT6Y7bduDNYDP7wcN5Gdk+oVhteMQ5zeP0j5YmBMpWpeWHFmYDm48eusvT
ey/+sXWyHnuDeBxUgqbHgEm+wuu+1KYmS3zPDB9llC6g++5GuG4yPdSNUXak0n6wZU8eiEq5AHWA
h3Lr6VXNGAs29hCLG5t76vLdSsfNJ0Ebp7Jn11H14FBvaV3yDe8Nma4wu+rZISZSs8OeJxIqkeep
ZqfWjBrP1pk/IQFi5r6TDco8WqJa93onfFeZs1RKmYwWW2+HZSNTfhsZFLGFVwJI38wxxA6os46r
zlmqUVSmBIR1ts2YQo4v0te41WzghpQEzTFoClq0LIdX/iY+XU6Rzh4AYvjxSyXHMqXi6YANHiiI
61JtnMYVzGl8QM9B9Bl+I8OS6xCJ2PgAC2RI2q5drQgpHpUBKbMWm0Mt0WMj2Jxnsq/iVaXd9FG+
JnCowHKxPtx4EhyUGRCRmmFDsDj1Rx1D86SJwKHAdTG0pT3qwc5yJ3h1UJQ5tGvAcrW9PNwIjtKZ
Y4pT6FulNtsvRGNp3vyfoGcMRH5Hr4Yv+npZoL5ko+ze6fDu0AK2N6+MmjDwsrg25nhjWIWyGqhe
JzcabGGmQQ1NAgoQrsGRZoMOPePwPb+libmtxXBpfB1KrNl4vfAWmcBaIqx0CrdAT7C9WscqkKka
vfHX+4AXwQTH86JUdltBgg9ZBY5yWQYbXGK6A+Szaq4zcGXWLyEM7/81UYRbDHo67mpeXcvY2pNS
W1Ndhq8BpbGEou2RPuJIVU0EeJou+JFZFwn0Lyr72u2atSyNobEPApOwVMEAlWQoRMc22WMj4qiu
DVL6YY0YIDl92M80VgCtQdQsLKiMBqypSPTKGlbyu3jyZZaHnBjvJJ3IDpBQu2x83913Dxs8YDyp
QNduLWnQg4j2tYfau8T1k+xb9U9txRF0kCIU6/3NeWdO177BiPWh4VBLKiDHwUOWquBB5+1PbJCE
BwSSbvX5wAZHcuQ05BqfcL3XpXBGERAY9Vac6Nss0cRnrjHvESm3nSWPjViF1PaSxamXfMOiF8Hx
f4iF+SuPFGfPyX4WWYz9SWg6ETlquNNRbYo9cRENHyv8m1ddR1qxkxY4WLTn9o7Ip6326zgnwrsJ
iU/d7leSpE2IBtvXxA2nDQx8U63a+nMo0iGsKXm9JZW9IGW8QgFErcxScBkuirLV3HgF3wALKi6N
1bl7YCDV6UcuveB5YzU4Va0YkLHSiS+D2Jzh2mE9IRgILkX8IbmuzjRJPD0ln2Ha31cGzc1hTqJp
RHvTgTEBX2YLtINsR1b9886VRPH9flt6XCAuqKLjJm+8qPjBjeS1O82sDJ5ynl5dnb7UuwvX5Jr7
No1jPJp05g2tZBAFnl5EsNiMOZEd/zC+UZsEgaRp6ruR1SWVQYILyb9JxiGU66fC0svy711BlntX
ZhvJU3Gkr/dCjLSiN1JwrYaNv1D5sAI+feUvqHJ+4/cUBKxIdeb1oFR8NZgfZkKMa+IuK4tUizz0
FAl7wRXr77FowGSw7hMxx6dlWymjHOXEkIBhk5tITimqD7XAr82WJq2t6MuNySCzTD3zD30LZ3t0
9B9ozocZapvB8ExizbcsZODIzhsFNpxLapZYxZ5qu9Bh0XDLzC9ItEefaakuM9/StC12heo0u7t4
MU56jpPnlcMI+MERA/UUFyl5th6b4G8yb4B46NJE7IPnnODDu2i7ysOQ/HcTeQ5iN6H4xnadsliV
QRGfEfwWZmxvNUoyHZrD0ulIiwzViPLxs7TMsRx++QhN6i/fMD2olanGgaYRZdPDrJ6fXrLTYWQq
x4dSgCmGOqNwToPaIUfvBwn/sxeESvSWFLdKDYfkwf8vRR7FPe/TllkQC+z3QcDDeThEAVCQ78BE
ZdATEzaquP5UPwTUUqva7Lvc/m2Tw30gbKP/W5LJl2SjTTfyWnLb2xPbW6muCBXo34LspUxbXfTx
k22lDcgj3QHXnAOHC5WwduZ3TpVngv+YcwG+RwqcSxne6GOAmXIwInpgd0RvN2JT+qppaR3tBIk1
H0E1nKaXUFSTZJh+ZpvOxNdc8Ed6fcan6mw5tWvTwgAIpm/w5uQSYMzi+2J9Yo41KRfo5pclvf0D
W+Zm/oI9zQhzCKQ7lZRkyfJPinUxhjALr9IYG3wftWZx/B3Z9gl6v6LoYPwB1iERMV4w9h+YKZ8z
cbLsx6nCwiuRDeIXhA1CbcMWNvL8EdlfHhK2/hYCPhXSvvODmDs7IxnndkMjj1kv8UglvFIwVn6s
5VnEhr+wp16R0gCiKkOJH8utqBarxRWxtkKjAVcYdu0dMV1LXocfepkLFiscU/8noSxt7tz26Oqk
fP6oe+NIornqqjigb1dpXzRVfKGuLjBKSvJkHPLFM847J3FGalynFV0pFDrvf7wY20RrLLq+tSKe
cnTK6Pmwsafv2uc9+i+gkAOknja5eVQHVJBbCDH+XkouppR661UseGy0msjde68keS9UnjU7BuVy
/bTZNKD22L5s5Ma7bHPJIpWzedqlmwmmAtB3YnfPy4jwE3GCyjwaCDhM8aviw7vHgepVEf4BuLf+
8A63qjDj8WO9tuuNicVVVSXksmT77ba1j8888vN6/7+6JboQePUfGBX+QJ64f0V7hokQ9u9wsrKL
wgoAplRysYNrzao9td7k8X1wACz1+xS+udojQm2eQOgPw1F/MXthMNKGmX8iS7V0/T3EOXBJIKf5
Q3B/BaEkeJyhwiR5RAPdNiOsd3bXmfJd1LeEXDJCYwkEevXnsI0Od60cWck1dZp5MG+K3hA/EUu8
tHduEnuC7iFbu+j+ABmyKJbXM7Ek07itfq+xpqjpWOpHfafOSxXEGlThyH3rHj0hKH6X3CsaSn7+
BAAecKBiCNLRdZJMMWo+2vNHCL3eFXzM4Hd6D1eJGBFKr/n/cNKejP5gj3A4MjVBWSk8pVJlsqjD
PStutWmZgvqBEfbk1/egchTYogx5tYbtb6S5/VVT0ZeCOG56IkJ5yaN65tWH3XzAepFsTVQWOovX
YkVP6RIXX4Otq0ynu9qqP3iIUSbnKXgdvQ8OAymK9yR3/Bu/MhhxsE2nrE4hR2I54gYslG/kfItI
lmuJxJaRvR6Fn/ecNE6CJqcszlCDpKc6oh/Mwsu4E3M91wZ+MomrrBkLQLPKokRSoIBvoKq5S/MO
L06SH1IcJt3jYj/v1K/Ups2Bfxl8QPxy8wzpL5JqrV6R+U/d9E/T9RFfo47rg9HOoyxYXVYI/ahS
3rIqvh1/uCzihgqtPEmbAdfHyvnaybSd7kBrPQrZNA+Cav1BRajuue3wF8Unp+W1pIwAIhyJeU/B
jTPDfe/EmTqo0KE9JFPeDMB/OiorfT/4n1VE81x9X9gutW4WoETrL+1OYfd/B66H7/x5ZO9wPpNj
Q+WgCh8l6FlfsWyOCDKjGGblaQqsvaQCFBjS4uK9bxSYwg2hP6EJTh/clrSq6SQ4AkbkKHRHUNRW
k5ydUzuv9BcmTte6MMXKfBJd1g9xxZc4IZ3UBe/fbsQspcAw3TyLnHEyBopp9eIpjNNQ+d+UR/63
rd+152y2KFtFj4DVutMvUxMGishxEvmVxmlyFX3IBUDuWmJHZVLT3JTCtGlwWGRPy6bXx6fb1pcv
HwiO2fU/JT/0HQm28dLUNVsphl8b4zhwnvzBEy9vKS5QuCE+tlaMEiwXTMQDRHR9RuZ3GL6IiprZ
2man7HIZZujvQUG0k0aqnV40zdIj12QxscTIXw9/oDK/FfPqCGBlTXthF/rllN3rwnE0OdSatLPz
193QsgWWkZPKNb+8TvJVXUc6l+7PYAuIUSvRTovpt5ix5niO4ajFrewDIPmYsEKmh++XWqlF9FF8
C4vKznylxoi0qJ2G6aAbrzQH4HTVFr3PqSSsPJUgYI5dDSio1q9UgChYMYXSOiF451qicz2D1+Yn
ug7GfatbLP9o48prioXqX/OI9aHGatVFveMVij3RuIgsWzstnFK3Yv+2vdGAloLygYsnGnKcwLv8
HE7K3EwYka9EZgdbhnk3TvsigPIurAsCy7+eZUK73UbxfmfQsiWa7q0uD1iIzHnk/Kw+Mnnbg1yK
d6tQwJ+CQjCMuAb1f0Gb9M9CxMECIC+wpCT0F72dT0UgTm4SrIvI7guleWYc8FuuxVs/hLQE5O1P
roA82rSFshOCwoKOrWFTKomGA8rQHURTLvzHkIhZhu0/ZyqZ+Hve+bmUFxLLg7ed3R27hrGh+5rX
vYy0jCGcVTEN1YwpdMjE72DIe5HOxM78WIVR162o2USCYX0PHWMyDozdlW2Iwtnt5J16wQRDeczB
lmOYp+MUwA7Ww1ILtmO0RxHvAPWKhfIJCtT7cb9jK1QsM6csQNptQaRIwP04Qn+aDSOlrvOjIzZE
47uAm4QDgw1vPw1lF+MeX+qJyoJ0B7JE3Hr9/gu6RDA/eQkOLrly54a6G+MqwS7g7ZNUx9w5Enx2
j80ndi6rhXXenW30i/m4XeLuoEKwL1MOOPvi4fGaCiqOm+hw4iIT4YImwHTDOmdcqwJO0DpahrV/
cegpUI0ucltXgdLfYdATyUD0RezVreTJoc7kKiZZt8Ljt4u1poebpW6cOvthvpPCm+zKUWDtPD80
J0Y7ciUD8Kqf3seyO/4u4AtBwpr3oHwEaTnKJE58O783FKTLBeGCJLeFERv/VYUxzYI1MRPb3hmz
+65/TlIdJGcYKfqxYNtIMf1vpTDoSvxKeFYrW9OCdHh5HPi04Rc2x+U+KvYsiVhn9+Wh1m+A5mIq
bEgsZWczp9KO/ajqqaxdEPA/aDoZpeQxme/fvnVLLn85lnoS9I8FpocD2ebVGpM41BMTYQYyV14x
S9gpWFhO3cjCxG/6z32P1rBTNTqkuZh2p+ima0+QdEQYzPLH1dcCwbOAjD4FQFRlgbtEjGwRS/UY
1ZmWgA9onrT5O4UJJl/IKSM2Ua5hUXmuazCgy7fOtfVBVGkEwKqPrNflLCbU61sEjyprA4URflH8
pk0pP0gE/uzNDPPT68/EqWOu5XFlrDa9a0andzQEvr2uh96Hs/BZM/DhVivUDC9J4hsiWgq9/Jju
IGNDhkXFkqzgBC7fMszj4SNir9XN64Aq1EJTW6Wx+Qg+vYYl/PIEGzwdW183Tl0dIcluOD1NBN/K
d6vITmncKVAn4FJOm5J0uJ/sWvMeYk9zd3T5tRxPNSosfrQsqnje7V909rekYA8cy1Tzu2aQbL9y
tNaL8YZ9P5Qe1NmspyTITiC87EiguLYs/Ls9WGMt8t+E++hWjkSONrOi5aCaQ44ctyzk2m5txAU4
SXqzrct6jDJzn3dyxDJWXcRMJIml+seoetaXVQvpGLhV5x9bZZjqBiBIwxZCJlrQVCWDoEPDwv4Y
RkrGLObcMMT1WOQdeDU4dK7UWl9wojQKWSVEUwRd0GHn/5v7vzsjD6Mut0zPAgm7o5G80oC8n8dU
UR5HIZ0JzyUm16TdpCRuofECxhSbO95thR6npvErSEychnKyYa5f8PWB2/updh0GzCiPR1pyQlL9
u8Yf1/K8Cel3npkQmD4tU4eN9FMhlExW5eu0Aj5beX9ruBSYlpgcRFrZen1MoO0xnPHjOruEbtaK
KwU63w9FO4YY6cSJWecO0Pku6x1UIsbXA1Om1xEK1j5pNnwYiTsqt+RMhDbO8OvxEoitXgFd1cH1
Nk5gk1hhW/+ZAizekLjwKDPvsLbt1O2Qu92RHEm2FW3Wu4S8YjONQ4knjdVnNKtGQzNaCHcahGHM
G0tQtDicwSoVqtaw0e0DjEMgWg7cEZxhlSXidVTXts4c1LtMnAQ9ln9TyOUHUCvEbwGsjIXm+6z+
E+H9vpd8u8bpFnXVINDmzgShqxsp/9CgNLu5/6gtfTL87F3xT1bMSwEXlBe4hm//oMibAgHk2jZM
tXwU3WwRhbqvT6kIZbA2/9b+/93Tr2ub76bKYVDNrNT6mGmVRXy50M0RGwLE17D8exhaGW1pndFA
YLG9OAly+UP/GuLPcMyKqEEcSS8lQj9kSmo8Eyh4TxYvGYJDdEwotq768lhFNy3TLiroWzrS3vSg
i2Z0PpukLOsncD1OcvLIOxtSWNOoBFLf8IvqQmihAU7ikVH0RyR70VOcbmhbrUNC3Dm6Wz9jAQHa
4oqygIdw8Xjg5ZvX/gsuWE0gYRwUvNoR1Esb3WwSvfrro0triuNSsb6/8reEaf47sDhU8uYGI8/Q
ZpGUwK5gfe7IVa+IIS6t6ORe0iS9UrVxnFItaiqBREQMX9vodnweuno5oV+QKOL9lS/yjcYUerSM
RYf54YFokFtufB1+tFaT3tu5qsRqJsl706t/QyDHwku1WITnIl3ABXqne1mvKuIFCDPPg/T7IEyI
sivO4yBL7ugNu6eZ0bp1lUFjbuGSxW5zoUwUOXWiX1bCHxcdVf5gHd2zxIjW3aZXMBGF04DNDO6K
ozHpmZ2+61zU88Svz0k+aPW0gvD8ITcFDQPLQ8jKNRl6vY8gKYibnRieoTptnq427yxNc2U2Zm3W
vc8LIUwKzt6D6RsMN2G8F2CO82Veg2IjTjNyjB0sTMF6oPtUqTZ3QJvZUYCqPea0Us+2DqG+uuik
MpqsTMDuPfd4wcSs6jbaC/DaBtqfPz9c45kSX5CWrrNLSiknp4bHSees3nWggcLH10V7YYgLccUm
+ILZDfzWCCQch5nlpHqYHCP7C1AJ88qw/ylKVlkwFEZFpnPCaKbgE0nqydEoF6Y4aebvWdDqU9qK
mIdYGTpXFOzjTaUGPH6IcZLG0SoJbpou9inslO7y/eQ/mOFZ3Ic3iZLKAHuITLv0aaVYlBj3OwrI
PqwgzxZWM2jrmV2ZGhNOCYpwKpbtPibOgDl4tFvVltChseZnpzjMoQ7caUbsMtpShVsSVPbqSG+6
UuC/PDGC7RB2HUNlN3KCN69D2cSknlypp50+gKwaCDQI9Fq7NR4EI2S0d9xLwDYTv0hR8AMgMSt0
01SININ/1oiRIZAfUGiFD+3TlyJvTyr3HStdgNySVKhqH7OjRM6SO4irC9ryKxZixuy2ioei0Q7B
WsD9S0jhj7Luzy+84lHM80S32vujCpJtRrRctJ9bj6Ck+awYXTVmG/wJaBGxKj/cA+0tc+eNNmHU
xPsu3JJi4wttP59ycH9PLCwQh4qZfUo0QdeK7epCAT80gwxTCeNPU5kvrQc7ZuzsrPwU7/mqDg2o
1mLOq1tPZ1kOavhEnTTG7Ekju93ZAaeiQ+LK2cgT81yo1ExdxOvqh6KlrGijjfdccq/iC5cG5+4V
tOkeaVbTQOb5auTHu1iDjky0UyRKVK3iatkJr61t7NTcrdVgQimTbliC1fBXDHNcGuf4xdcmB8li
QAqumI+6IRxKgHPzJXMt6Mfd6woXCM2YPf4tkD74nxF2J7sphpCfKkvPZRYfbBBR5tiLO1APL2t1
SrtbKEehBq2d98TuutgLWt2bIy8O1pOmkzTh9Tv1NcXN/GmLJwgoEhY1p4I+I0sEoHQsPEziSDnu
L3i9aMzD2eZfc5SuGjUhuxN/64SJXW5m94DOMdTLY5bjeyWe+k1AEua0jEMOGImERrz46f0xmF4n
pGAzQ7se5viLOkN8TT5QmgO8nVC3JvB2D9orQru8RKoFOcIfu8080MhOk9A6EPGQSKY4KmN28Idb
CLlK+sYQ57iQP5x/UCuDQFxXgdlNGZ0VA+viI+yt714dAVN36YVdSGQ0x+1huUMoCfqZuO1WsBcb
1pEcK+o/m+4F2v4UcBbfepFyxs2iUIqoCj+Utgdf8Cl+XCTfF1/eWw98Re4JJznbwEpFLI7Bdow2
13RIseAF71EdBHij0jH93Z6fiVEKjn015PIauCTqExAQp9MFYLgDHuNypBa0MmtFISHfEV/498b7
v11PLHqfMgCrJ9t9akhCrpMz2O9dX+L/oJB+PHtd1iNANUFxO60Nh2E21RBlOr0X7IJM6naqLAAo
2adldPDP7iQReX3Y18xibJdN637X9THkv7EbBq6Jw1snAJCKHqANDTLzchch50aj/Qo3wSGwq0nO
lDiF1vwHW93dggRCw5104Y3Uueuoi2dEtwCqrdPG0ey24IJ0T1lLNT197PLcmR86XKM2+TPENUgm
NahiS8uef6uHglz1lqtKwCJksDOTlrZe4mcRwJ9UFH/+R6Ny5PH/fvuTge7YjyHb6YAmfyxmtHd8
K4LLvkRZqNnRHqjPQZzEQdAtl85EP/QWNNqIl0OGhvMslYTacpqH/gIIJoevscwy3+UvE0Rg4a/w
9Lp+T1/sdW936hs81n+OjSS2zsv7IY/v16uLXeJOHlKURwJKkFTkbnawjekrjZfQcc+f+ba8Izzy
eTuFUTzm+UDZng4dlcHFWATzdj2K5gLet1RIoHaoAu40etr+V+Lo7h4mON6Uy/Wv9lcRZkUgJ3Ys
COZSgmFKuzqDdkiYgJ4hh1aRALZYkdtKgaXuao689j5G6ikeFhZ3+hTW8jVVbFI2JMBE0i/dQfjv
sN8L8NZx7lzXQxd14zDxe5/vF2Gasip1RPYBIEhQpMkKy4A4Kh8UQ8zJd9/hVScDp/7ibLCHhUiG
u1Ig452ihBJP9ymzPQltbW9J5RlNZEZZN8ezGOSdEhz1CjU8SXo7SJvZaVvpGE36gCIcvHPvj3i+
21NtnN4O9Y+tXXyPb4n9jVyIu59rnWYFW+y34tyI6DMgfIplmkhdwunTOGj3KYr+o5/9IL2JtrCH
MsXjFPVE0L6heYlJJYxj1rBi00Ywfu6ewgEy5xqTqjefjwqxziq8HVzC4pkh+0tT9hneMw+4nMCB
hv8hSlyi05qpyUz0aaC5VAw0V58+qW1vrQWbpwxySZ6ixE5MQDrYLjnNELGxMlreXL/tYn+uv8OV
/AGyYSaPuuEZ0rXgGW6v9bCBlkJW035BMZEQ0O+jTWA6m+SMUoDQEdErR4/nRitAI/sCTnv5tfWS
HzKa0yw/Tntl4bFt6WqOFWIegFOJLCeFsB6BJlkS8jCQbmh5+tiiq0qDEowS0mUsMq8xrNMv4gsF
6E2cfjcT9MUcw9d9uZlnRDy1cfkKYda3JzkGGdO/X1Z/xbdfT+2HMXf059AcmMhUxdQYu+xgFrA+
jMe2JIJStIlNYAuhlwqc25bDxGy1T299/qy8ADswVaGdO0V/R5KZJ47huYF0BxnEaYXTROj78o2R
baW9ARixJiN7qesT8DQMGoiYKnB+vHt+Jc34sFxqeelzNqQTJgnBW+XxxowNfdy3WqMvTPWTRQ/X
lis8IatT9i+/vCLo3sfjiKytcDIF1uLu4zPh1EBsCdPCjrR/uKrQvTJEU9NT/ELMeR8MmYA5MF7f
p5jd262nUeiP8PvFpEbunuL4+8uuw6vvh4qIu5+iaRk30g6a04VtHM6SNcwvsPUfQqSX+96RlST0
HpuCAQT68MG8e58tWMEYYFvDcYp8AidxRf+sd0YBWFIpjHhYY7Q+ICiYNkRmpFT64pqNfsGA+jET
EKqYklLXzSz+iwg9jG4uRdeE2Ld1DZGViT+qvdxhG8PGNorHPCCCEVjNYAV8znq4MNYgGlbHY1O4
9zcTswNTU/56VwjRPak9iNBK3/Dgy6gpzrz+coBPcapty9iTAMszXyJ8F+krMuSUiYnmfcvCYQwb
mMEATC6gstoU1L9SaaSgsyliMDgV42/6SDg9mmc5qZ3ueLe7kwuzyXv7aYOVF/HTzkpZKa3Rya9G
Z25ucVSWXsjwifXd/yAMe566itsPKP6vuroYfiCTSHagPickCgUlFHe7jputHUcGpGnIKu4uZ8Ec
vIwadW5qShRMA7Z6PWXezx3lquYDoB1Uy3OWqvdmbwYlmU7WZnRvsePdZNrbin48glzrkrK/iKvZ
7bx7PplVHWRRMzxQtROKLiOKTIyZgDsISLRpfRE6nLmMZ+8A3Rbe7m4L1+LwExgP87LfWNyZOe67
Bb/Xmw/Mr1Iay1WVqZ+/L3M2rQdC6NEQ4RP1EYY1Z8A7FsxthHUqZO5WS09HI1ZIUuYLQenL99fl
pYQO0AAPAGutpLHh2sWI4bp1DiHSRvT8s2/8bSnVrEPhC4E9Jc5DU6e4Z4Wzul8FeQ/+WlyqJhls
N43cvwN8eX9v1YOjKfd4q+ETi1BNIFRYJjqZgdo3bIEAC//dP3kp/Hn3ZlzigQSVrQWLzZMQkHCQ
534HaQ1fOw1rp+jf1dC52nyVeI78SL7N1tVhaTNJy9WvybMgaoIYstBoJrUuvUvQu9xbOWyA9PL5
qq3JzflhCwQQw7ez3BSvg7R+XHcVheySaheMR0vvv7RG/1sL2ezTRDZ1Kx9gpuh0QEvf1EE/tMHQ
0dihktpbzcFqTrkLV4+tdrdooQlZA1jcnU2AFWWRy3JXwp4ltHEokn/kV0N/kT9SqrMKpjEwGT9r
SAK5KSpnQJQ0BmbaiUt4xNDzCbXzzQ8i8ij+w/FgwsvAagctm+ZUW6cN5DdTXZvSvMFWoYI5UTxd
j7L8+qJ4iOHndz1Tyayy8oiLQs0OGlbhpnFgrD/nzAsCPK3D3VtMbwV8ti2leBmR5yKht1xpgXP5
A9BDt23wWGQSie+CBz5KKKs/CFQv53JU2nO5VsCufx7pvwHO4Dn49DLVs1kGu35ywt0xiZKxeMVB
MebOIine4/SLJroY+oPHRspBqSGSRsT7vM4b58DEnnuhpsXW9PzqwLorxdP9cZAct+xmnYe1fyfb
/vg4wYLoS4DTVEq7k0WunkDBvfyZhhbGMsi7UH5DC7FMOmb2DJsPqbDUnkeDX1EJifUHO3QJuKSQ
eMFiPA9bV8PgO0t5vlwmG7Ean2h/iQ1x2OQ3+FLhE7e8VVjYcjWhkFRIW1uUsMW/5qXZQFumhatt
66HKiahEeETdsOG3CSSSyk800DMq/DQSmWd6mnTjLiWLvlr2gtaB9iBOjFW1twwRsyMP9cNG3Z/S
c3BYW8oop67gsY8OySrlg43kGBshc5DD/88GN/rNGLmtRlMU/4zuw7HqwcIh4EOxbV9AQpEEQZIU
32eKFl9nLgX3MZOUlBpxWiz0eq9dY6zs2CgGPg0DpOaPCrvaDxwRF9zWQRRP7NKg8XrijOU+Grak
eGqB+Y+B+t/0sNSZTRO4evVYUAL/90GLjLcnjVvDi6d67GrBkFT1aKOo7jhka9SfFRn0bFs6knkM
df52GPItodCJpxVMUp0MKFzwUrRcKmwAjDvUroySGk9h+jDzxV1mzCxvMKbVTDNBOIGTLgHc7BAj
Vq6mcboN6K0RvXW2v9o56bqrzsRQZmus/D8HTRemKJzPcvUJQhbBs8vdFpnawaZsJaJxVjNfoJAN
HDGJHHEH6Qbve1w2WPOoCIAhbnOHdoEBFquqB2YpZTxWDmmj6G/ORQtFoGxmPd3vr5xj2zS8hcgj
lnR8wOqpCSv3csvxjrXExtroZIG4NqmvB53BrsdcX+urSAQCVVBgUULr/sDkw1EvzzRXSfJXVocc
E0yQIEdTDws6hdN7jzi6L4YB/nVNkC/N60dHz6aaRR7f0NclyPYGSdi8Xy8+p9jWNoA+vm7HxN72
9HbY+5yRi7qVyk2K2l5q1qbPZ0UERjJZxUstX72ceumrXWL7eY9i3rpROn2Cuf4nP8ccN5Y5W9qD
oF5Tdxb/tOn2HuA6esuUMrT2if32p7Ts3g8uUpVuGhjHUHgio54zreyoOJMyEtGDMRxRavx9za5F
5FpcYuRAwuK3vwgdf5KXKIrpTikVhx4ZhFU3irXb6tIyb7uIQW7WUrZmAHijxXmyCN6ZcHTT3pLA
A/BLKiRevBeo2tjudbZq7M2lrtZaoWMmEvQJZ9fbyb3nt/F4sNydPwI94U1KYJQs9fVIvLFsGVxd
eqVX2l6uB1am0dQGbnn/YgTn0NMCyKx8Iax7q07mgE60q3VTkZSU0tVi3P1AAhfZtQsVSQ01y4Kj
4MqIJhfXE6GwxwYldM5xrHiQ0Qb/UeBbN1z1c7F4SI8NtyixyqN8kG85aZoMGLTxEqFWW28d8GoH
5oOLGb4ndT/GLxWaOvLvudkX+VGHBmY+RvTpsSGrM5QMXuXe1jSJx1qM+cdpDq+MducQKgzklpIa
3cSMH9KLD2nyE+Dx3Q9RDzzemP7bvqjW8SVz3leCa0V3Uyrw6JXnng/QJybyby9eKh7R5A2JDHkq
EMW7zt9Amq4Ry/HNtwkLsV5/OIDshR2MstV7/p6M1h+CaobG5rieRCvT4vHU0OcUZPLXJFWZgNZt
ohsTdC+sfvKnq8/+bsDfCNF7967jnmWY+2qY6zsUcT+lQhDFHXdJpe4PERMCWTQDWYLlJv8OJF8d
oRSlbc6tEV7OMw7xjhHzapoSOmUlkpymhPnlXaLVZdaEKzkWKcMr+ihe3tsNiUh4eo0VkLF78sOo
1TC8MFKMuAUtTEUiFB+c8SD6uixjKO/JjqoukA7QkgUvjU/TUzK4+QTTokhQ+EjmY7/+i6dXH3Ns
2ZWNOCZP57z4+8XbFT+Y/StueXXiiryka3jM0LATYwUZk2cn6IM6K6Mbxzz4EvgjKS2UHisgetRD
tOjxZmO/DoebnXl2ANIM5U1JsUw2J0qncj3OlFblsNnLlJ3VwYBM4GONqHAWpYR0ElSrwQaxWFGD
xEeQHV5lTlbTn+Bq93D97hdeCTwDC/RT8oM80N7e9KXISuqH5tV6IaCsqMtQb+UBYBdo95SX8cNi
6L0YUkm2Ier8Lz1GgMJP9MExoHJ2NylN1g+4tMMi2X2qLXsRZXfR1SWrt9Ix4RcsPK1ieZskDh9Y
IQdJOfM5v7GESDV2Bv7KHDg9qzHMYyXLg6YKRI35qB3UNhnuQJmaTXXdTFeujZiBUaPnoj7Cle5c
Cd7ku+7iWKcfpDlmydWs7K5GMDus3dhibvT3qBdNdlXEA3s6FffskOxKh+0ThomplIde0Y18kibA
juIU1X/sVdbr/K8ErsDKZy/AzW+v6/i9/CefSQjcuzvFkhXPxCHCKgWANLEMNd/2JEERXbdOVOo3
M3Qc9bz1rY770fxqsndi2y3PZ8zRtV8S1R15EYzg2E1tDDaiCM/1c3FIW3edqzxFc2EPnhf3tp0Y
x+C2W9bCjoR9Nj1paUsMDdTCs7cEcxwkEa8RcMYkMsZErDB+iV0FeFwx69buV9+U3MMr3D8UOmjU
5BNlHam9YTRDmN4JUMZR30vPBLJ/7Kf7BvX420dzjGV0t+cWm4xA3inh4OxE/afhE4jGgMEDtC3g
SOet1SsFdtuiFd//U4NbTq6D4kC31aeihNNaXdNfLbprePt20JDGpeXIp1yaNTinXPpHrWleO+I8
NLI3QARP+8CFJ5RI5fzjmTk3WhZhpb+CR6bbrSmpMV3MFZMxR7J6nPOKnClp1j7WhH9QUdLx71Fv
KSrrxNEawdRcMf1aFmxDhIMIvrBY2GviF5FOrX6cgs6BgElwFBJUsCoBFus0l2Yyg0de2/umcOAF
tI7VuGBolZptWOB1mXmmii9IQO8JiNsm9KGUqMpy1UXW+O2N/GjT/WJoETF9G+4POyIrRRQixwP2
L/kpxWZ2TsQPTUOQ2LH2YUZgPYDJ8DGiibQ3eDFEfM1VTeIaXK7snx8k6z5NURf3KKZt2IfESvRy
6hVAjM3uJ8Tog0PNnWNTbFJOPc8DqNhJGJsHcRWNgDB2tIl3r9UPqlEF5UXZwRRiRopDit630YL8
+aOOWh4BtezQsLGPio+0AeJTW/w6mfIfovTRNW+ZPYdGGu3Wzp8En4Hhpep5fYs8lb7xEzj96ZAL
0jaFjuHWUbFmSczeP5zerHlhZboWEbyDcJnEU5HgAp274bnm2tQOAzXlcAi8POQnlM6P4KUyAALn
+9b5YgQGRhhmyJHZJXVhmtFU1k1Cpxt5EQrxAv5t937XOsrdV3ZNyxi/T0/xJWtHwxuH2iB86ddA
3bBNy+tDFcdyBhnEFJ1VBQ/nxAnLb8eNwjxDwelXDEg4hmnGUqHBM99wYMxLaJuphmhxzcBdASV1
jH/PDLTxjpoS4oeDkvhgR0qYQo/a3HYdkNSHvbp1w5PRj7JWkCdFb7wxVJlHCg8hF8ksDhSE2USM
BSI2yM5xbtzXFPg6nOJ3RuyCzuo07g2tiJHllhNIPX0i9fIUZlAikIT2Jt35K2C/yGNE358Fy/8D
V4og4OzGHBBdF+rb7B2OtfXRATEnhSjHyzGYR7aZPaCwgo9OaAYxzAxD2b0NYNs9Oz05Oa1V/Or+
QSkLt8SUNmlp0pdMlTShkCTQAAa6DHq47WKQQsyJFqQore3OwddwxZFT408VR2V1JSHDcNWeFvLX
mJ9Gu8jpurD/Y3he44ykT7CKCzPYpr2eSBgcFeWp69qiB7pSmmULE/rytYY4FtRMvdmiTjRth+cY
rmOSDRUp64rrA8m4fAsOIv2qVlatX+XdMVcn4gDg6YKSmqambkSLb/Q23VuStA99EpgDwEpTSI8V
WA/1204skuYWmBjBMZfFLoLzewAdv8eQGeYCCaIff/z2KdcY+u/8EkTAnjad/e6SX+PCLX9g12vA
G9/R0dS8P6mGvRTULyQSFtzqI4rejTBcV2h3GKIpxa5YC5g05NVxbk5Lt0Wrk+M2qRilC90YZ/lm
CLn4ojDdzsrqLcsggT4+KDQ5KfOlncIRrS/xmJCH3AwMSSOrQeilK1m/nNvrO09Yu+T9Bkzrn+N1
XOd+35T/qfQrqTMAb7Thw9mLIwoAoFo0M0PcZfWC4uMmW8tEUsJ71Hiw1K0cZLJAewrQ8xi44Ygq
3yCqGJC5vYSs3AkeV5j3mLD1NUpzLXKxYTr1+hkH87fvPKxoV1NAG/kRtSS5igF9n5ZnPNI0WtqQ
Wacj/G8PltGe0y/wQwMdh6Iy+aFpDddVT7CczH1mU5bo9TtsjoMEiIO0tgrQqgzBDvry3iFBtaC1
+m7CfE1bW4aYWjU1vVkwiO7l+ZaFAgBmpzbal22s4UrfZPaqs3dpTIaNpuuDww9ylegxo/TugqDy
90bYfSiDqEfv28+K0tyD1d6jdHisCqan28iseEUG52hHmXl0VocedKKpL7TPd+h5kvLwupzKbDse
iCTsu5/WZIW9zqJ3oCm06b88n4b+AlDwVZhGmOtTTV5vleCGL5YWBXxhRKVBiWIEBn+QJYUNYMA5
Yq9haWCXc6Q72jYaT6FNAPPcwumhpxlc0QhrIOq86dVuinDvWS4Q7YFPqR7n+VkK+kOgDCyVCDf+
w87KV0Zx8S8gDpMheXGNPm625+fC3Hdjf2s9ef7Zn0fCAbRdcyBQSswMQZ798w3iTSxVyXxpxn/x
iggRDFccAJQsv6w5LnjIOx425ruis87cihGw+aJqCGyhx6MkPITx5s6bol6EypxcOmSv8vBL6S44
6lm2epIrjugbWTA3fv0cU42nibzwnpz89/H68ZZ0PRdFoatsafoFDK5hNd2n93duluEHyl/E0a6Q
vWdUOsmlTrx472coAPZp39qw8jh5XYAXKaKg6i6H5ehK00OUTwuV4G+dxR0vJ088ISJPDWB/nEme
1m7k7U9Nhr9Ao4BzDWWJ0n2JQ4YdoPaOYnbtasMAQ3EzL3LYU0a9JjZyLRWSQYStmNDXQ3IPOTFC
bHoeBMRIU5rCcF+dmEgLaJh53eFt879H6+CWPHhpKebWqd0cGATaWR5YzaNRn95336VdJKrwGH1P
kB0GRZWVBAaqCFPI3j07imZUHZH9cmcwCK3jMFuF2twFXci5nvHYifxQ8sGMnb9s6QLnJ0GtnYwK
hWu0be3i0fUor6MetCcllpm6GSZQueZ1et+0LwtP07YjNga3LrSxu3hCS4o7ak0cvE1AhBXKma9/
/Iu3LArBYSmzGd9tuvjAwzE7p4PZtFpabUgFTv7BnApdUS+X6dyMYRpREdqgVFBKA3x4XCG5emvb
4kydLU0A0GI4CGDZn0il5m37UQkdgR2aoaH0tQJh0GUVjDOBtZODN+rmZfKB+b8oU89Z8/KhhxgN
Te80Wl3vRGfl+PbMFpLZgcemrzDc5OhZ0+th3zD/yLTn8NpWz4RPfeJUNRu4t7iDdDhWmHSKpQBr
VA0RF/tjALHWZciNBbAN2vlDeNf+nhz22MYPDWTxOouw13TJ8HKgRFiPlDF4Fy7ezvtRysf7C8HT
UcHGQZE0X0UHzsMRciNSJ2K73XAPLStnSI6LOWDgQj1yLKUkg37jxcpcqG2OzfL3yRIeCmTcnQsg
wNroHWgSbXSe6yQUHNozeDt56pf6KHtXpoi1bmVSsehmbfyNI9u4TYyz2KVTHtEOil93/demyGK4
F+CUMczoDMMsiBK4nxpRuX1jTFM4J4kFnB7R5ewi0W0sZaIWxueOo296NdB1k/+kxuqc+UlqKyWc
PVqu1oJiNTUmlWy5UgpVNsjZk2/ge88qrKji9xjaNoPWTCxg8NY5MIrnlpBFh6gKhrdfPaOsc0X9
jPJhY8OGLRoBRRVBJMlWMIernLuo5S2zhiirp6ntqhEG0ztr1Eo89kRmvq3Zm/bT/d1/3qOxFGCe
JNukdImqqif47O+09xuFIZPVfpqHsn7x6tqSMhdmXO7IVy1QZWfeoUfKkk8KDhCfigaccUY1LHW4
hOTZxE5ik8Ow7NiY9joDOYzml+0dIW6zGURkeC0jALGX9AN5TIKJg6iX+oEE0y1w2GM5bnO8YHxE
6fKDXYkSmh7+s3lxgXMMV8SC+VGE6hRtHF1UTEOgzWf4J0vVpKuCfLYhISyYNU/cMsosHVAlN/AJ
aHjG+mqkOZyiCqigEG7wIlisWgqoXvnk6Yrpw8gkVbkKkNvk7CeBEldyLzyO1AJC4NSXka5i24JW
G3s9TqL8YI+mQoi5N7PjytdvF/PSRIyLacPKbbLYf77PHj5QuMHIovHEAMj4+uJvk2UPuPyOK2c4
alAh2XqK3z1Z1NjGOrD0rqKh43j4ym3Q+KJaMk1XEmpPKPKSFoqyT5Sm5Pl7DzAvkmVtDIDQIMFi
7IKPnktkedKlqgUW1kTC2n2DkMyi9bYQVMg/RcGU4aYfEIclV6aWi29VTTB46X10BHm09gX5pe8F
EwRLfkUM9PYN7jViQv9k6jp7V78M3KPSzedowbYgeuhIJLXus/pvi4RVVjC1alUSxtdILDY3rt/D
m0uGoq1IaXLEkSIkEa/5PVzRA0zxAfM4NaDR959lhb56nV+eH3D0vE+iQq/aaGVCD0TBnOMRHaoT
Im9D70nRQDFIOXLCG5Jr2equLZGM/quUIA8dLXmhadXIE+zgJWtM2EuyqXPtOMnqbzXuxHIWiJ85
x9Hv4mdk1jLmpAqlwGT+RpAAzJu78mrmNFn29D4xjT6FK2E0CAXX0um+uJ3QwWytHteseFoBlzSj
0xFHqOqb4Gn7Ko6haJbKOzvIv/Cnb507YWJfod5S+JCaYb1YR0AFuk7ZndCJOljImhUzwCrx1V7G
S4YtSomg56Uu14pBygdlw/IprzyhT828vWdQEEF6JVbMix0cHZv3nDEUueBNKEKrXZbeGBSteK+U
K2P3HACdXucjwBrGSf+JXZKox21gCPbBZLG6xEyZpasvsXcS4Q6gzLHIwamzg2Z4dMtqeR7DeL4b
pzmWYQVYSwBH352r4Bvjgblc2r/N3uhQwShC3NnmtT4XK+vSUKzhUS5FHyhaJoIN5lTX6oX2jJBf
p+MXlaT0cwO0FkGAU1Ta1eiofXgwJ4K8byip3kD6+JCenmd41xc3pFquVVEMNpggJ4bG0yGFsz1y
JPsIcl8P7l2VGebtJR+x4QX534v+VUs/9h0AGWyswjGGpn7JL9Ghoib6eS/5JQltXRn0uXaE3RIp
MLW0tAmRB1foZMhqm1aRerWnQXiVAmCoDBCBZfxhpSs7yrgsL4vHSH+8G45urhcv0HtY0fSjNBVm
Nmsr7kcotXj2dK+iqHYLVJBRhQGjfIF49YDEViW6agiEvIA6eLm9JMCtAdhVmV61dKvgdck4XfAN
/h8qpJIUufEDng/LQrc4pyRsgVR5EQ+9rco0GSAB7T65MfV68jEJc87juQ1aYCFlwVo9ZS3dy8QZ
gIBLxYMoknbEF/cvgtXMsR3/v9oBTiKzlaoOnFmIJE+PfSaC/KW3GYPioiYLJTP3Sw5yI8qitGVL
57Lh1iBGAoTR0i0QxiXkUisAUg4ngOxU8DNHu30F3Do0wncD+ujK8XOTv6/KMSM6soO5To2UP98f
Q697U5DAw8d6cxEss629nIibg+QT9uYL3HDSlbi8npFjKgBUkBnPzykNis9q6BgVxgQcPImXxBiu
SC5gBeHO0wjuXvqYXwos7C+K/KpwQ4v7qEwQ4brZtbdS476o0l4rl5+NyRyUUb+XGtjnVJB9Lc3z
q7/7yjr4ObpBhjVQn5DJcPq+uGUdcBVTbp2wCH0H0viEFsqk3ooocJ77ydOCO1V85u7o41ikIv8B
NXNzG//LnAvWfb+aExA8McQ68QGbRsBfH8/HcxeqMLuM9g5MEdiiVD8I+g2+cDvrSYrUXWM88Szk
GanowrVNBM3D3vz4JysWPFzmUMWfD9lGKeyWQgIpP+JG31Yt4a0Z+98lMb/oW6S2IIJw/otB8Cwu
jUPfuHAwLY4BhFBdSAbR4u6Pkh1oa2XxXdlWIpdcDBsiIhwU4rR4UQ2xW9IKK4BstS8NgZKl7qZE
gDW8fma5LUPAafs6hN4c2Z2ANYhxw+w7YiVV985noV2paomj1Sk88gr/v5zsb6H4j+yAOoECG2n0
OhTILep8EK9eFchU8OlsJfY3Uw5GvSyoAeo1RoCYVS19haLA03krtdHxAXyFPw8+J8UzPwKPGXFx
VJUirKnRKtkIVP0O9QCsgTrYQfGTe19Nl3mvV9fTCTCkabMkp5ljmNgnbMK4jMuuXkPwKfwVoBy3
veiXlJadAyoOigoJxxXMWR36Ra84rt3UnIEecdNtEHw4p6JqzE+y1Q/LTcinialGVJbT/8GQwNmc
LyCW21Yy7MpDiGYNAvUlE71dOnt8/8rcBwIZ+b5W2o9q7fnI6f2uM2WSQ4JbdguRkH+SmyS4Nvht
g/Zv0nvJf26mEQ6SR5rm9aFSrFrn79VhE8gXwcOgOqjWDsEKedu1oWvxkBK8pt38S3Rxot0JB+DP
iKb4zgdLQfx6kUkIADYc9DnqeVwosA/xEs8ay1Y1uWhE3nTtgUkm0765+xYMLLv2xJWCE1MO1mJb
zs8E2PRPYTdYtS03Q9Sp74gfqyRlhpZ0tLq3HZFIc6UPis/qW2fL0W72dJuBu60wddsbPXvhQtfh
ynYf7J5jDl+J7ItwsWcDJcI/toUdHhYefVhozav3LJMJS8wdoFO3TjQq9H+dmZmaWT1z7ddv2Ji4
Xr8Y+mecbo0BGNFW7Zkun0rfPAfiYKeEg0i70nMxcKh7tpI87F0zLGthzPe4fBbL4fPBjWLd4+6f
zjlqwUCvbXqGyiUprNQeLHvBGT2gy95sz8BUm20B7OFXgqL65S4iDdSY/7TDK2UoXbBPp/mXRS/n
m85SSEQAvUVH+0+/8jdWMNZJLxAVckso9vq0Whkele2CiX9nEg8DF6/ApyImRL8jfxsNSwlesydv
a7Us54LSnrbvPtiJV/pypVVwgaYitFGEczCtmwq5Kh5yj4xJ0iYrF33hkPF6NDiHEaYfcdvrUFHP
XvgSZts14ITnN7Wt9Y+HGx0feEbpoJArjZkubnKLRSACG77N5lhPE3obBeHLJdWG4v4CMEvt06BI
rKrCUasiNralkRV23Kyv9x8SRAdbYryFhzGWjU9+PO85aq9vdAY2T0c4NEHVd2O2jTdtoqzqYvyV
eWyys8CtzT9loN9Yzkx+SoS3qnT00Ys24FiTBrdYTVEEIHNHY33fVgtmXWPZlGODJRGTXSJLECZy
uwmRI0uS+awYH1ArvRzl2G3j6RziL7/43bn6FuY6CEzrv0VblDEzTuGQBAop33l1pcKACYhlb2GY
R/BeqQPQax93f409JuZL1KfY7avZr9RMrAMg6RN/RGQRU88vEFLWfJUNbxIITgtWv++ob4iC4jSn
p6AIEKnBHl6fJG4eUezZVW3eNGjuEJfa8lgcpPJKnF+joIzjY/d9xORW/GSzUwMmAMle/unN93i9
wPQuv1AbjJUKFVodAadKmv5+69ObkSGl+u9pEZ0eL/oqJD9JaWseR6iUMyXa7kiA3jkYndHU9mnM
ov3zHF0qp0LB0gsiS0taysQHHlebGoBQj8/D99wlwbEN4l97OtC8GXR0r7jC2bre+P2+2VnJYstk
4LU1veaMdCPEqpb1UgpYRtHfnqPB+A0fyDrh7qxa+kSsBEd3dCtp6YGnGMMiyFQ6wtZP9Xp0FkXA
f7EAOAnNUfIy+01BK/cK3nHAk1vpyCbpH12gKRB8O93S0boyCsmgOP2FGUtve6SVr+sdznjoZoQR
aOV3IOznn3nZxszwn9ykoohvkOs4Wsr7rM5zLi5mM1R3ak5Ms6R/OFeBXuoxMzfulPdgvBX/YlDf
KPreKaqZ2WcWde64m0QQ8IcDqE6Zda3BCWdYyGvG3xERV19Qn2rIkDHjbYPpvk/BE6l00fdgTQvD
jAnBmItui6PeouPdQqORW/xIYwIPVYMdMfa7AENSRKqomDJzMAsJXX+CLKb0b63ReamK5Q8uFPn2
eW5ykOMwt3EhS3/kZgADpdZI22Q16zkPvCBqW+sqktDpUOT8vpO5tQaAi+7zwO7a8L491K6O1ff5
bYXrmyOBDTXcdKHS35x/L8/x1pE1jR0lXsKf5eh5uQzeDH8v5GhGOajvjeA+h1ms2oQemL1XzBki
QuGWVFKiljWW0zqTsrIB7AsI8+WixCj3uityTDyPhxJwrBQNuSyx+m/F4PP6wDoNzcZgkeNqAG+Y
sxwNMGK1VwdIWiMRK2FSYtzGdxKu7FgXNfYQd8f2s9old3frb1/ebp4xW4UsPMejjFYe9Sw9cwX8
OVQUWqQ7vNUMXfygQrUP6VnNHTdfvEQ/NMSVMWZwq7IfuanSxEs8odjrFjsG1AD2EqbigptkEXj0
xcJaIPpnv5uXOVIg7KEaj2ZD66j8/tUfrTLNActk7PrWJ4auD4qoiAm6HAsCAcNYPxr2rZpDcYg9
Yr/q7JdhAuu83H8DSVqdrXOiwZVxjnWY2eNZHW1opkX1T9YytxvYFMty2NEGBr0jWDXCr7ePKzbP
lIFCBO/6CwsPKBMBlFotfDejICNjCzy1CqCZP776Nw/ZODKUgNtP63hS9SA1Yogm2wvwprRWT7jB
kVcLmZUkwFpUMOyZclkbwrDTJHACQRdP8mx9GHnQeXgJRwfUeLpKYbSL5O9h+GNtGjr/aSG0bGwT
BJey20AfqXETWC77um7+s68rP200e6w5tx7Qby6YSKKWondKSinpKe7Y99DEYDYdnuzomeBj8ow3
BvNew2saFEoYTzK3EmDA7xNdpvvorOruyiX9Ds4/Jn+lrYiwnGqH7Vs53Wn841fSg66gEB2mxFSk
sM8Gy1C1z5RpbxmntyfpW/hKoOWqSEaxvNdHvYkDQQ1llIbNOBxjfSYvLcoOOqBAqLPDJWSeSReV
3FjMQBjsWrSTY5sK9qLlP81a3PoZ/4/cf2fkyAZ6PmxIS9OI0PBwdGJu7rqSd1mk6j7KkPUejIWc
SAF6XLlTxjVrSPwM7GdS839samSDmp6m5o/D160Tpfy1RwOYYwKFPPKOtrPc1xjNMHI5LLcOu3YS
DED9+W7h49vlQAHLtaRoAaNccWjgjsLZMgHOprwRaVeM7e/y/z29SuEiZev3oCWNYSOnLz+Yrw5Y
J49dtmMVOJ4mOkQqPmvvpy0Qqzu1287avS++IiRdZ1D2YmPi4RTu88F/1BCWnv/1B7tgH1muqWZ8
XNuns9NAcyYM4rdTb+BGaB4sDNxeApPpCTDJZC9TuQITJoCaPC6hjQwD18f5T8f7h2owE6qyDm4T
ivJ/zzeATcMvv4VICArW1gZjijsNowJ/UeTC0SQSDGl16GskuKM8c5VQv01620hL+wn7N3aRo5BE
36zBQzLd/y3nGfa74rny5dAbz8SOfhobchre3jjgNCB8erbqmwLbAVHl7fKXEtd6hIF8JXrK2FGA
Goi/91N0asiqg3rEJwXCw5d+NJ7EnJO4LTUo7IZiNlgwHxMoQNkbOJd8JVFh8dmk9DqZ2FgKeZpY
mUwd4ldX+KJdDdERCv43qeua1OAGo+dynzccf0NLqumcZdNEZN8UutDR5xSMr0Q0qzAxgtO1cYhL
WWHB3H9DzAMON/uFol1ScVdiqcbHW32cCaJTzN6FBxBL7E2QMqvzXVYRDSF+Ss8tvfI6BfqDWTaJ
I0gBLna7TdYVIqBmY+EPOfCx5IA9fhA4NIWU5dRtWjBUijKrKt+dXKP8HZ0L+35yT3+M3e1WWkne
/Tvq7Ne99jONNwBoJdDGHTvo3jUqYt8g4qM3PCyuC+aRa5bZW/7+c/0TfwFV9m3SxfHC+2Y7upKI
4WiAw8624Kd6UPfPffLwafV5ANCmgMETvB60we5H/HGJuWVN8sGsTVOjxCMRZGwxn5aBEFEr9RaM
yW4gzDuRxCwesMIQM6bE+X+itfE+X4ESY68y0JEB4VnG5GqbQVarN3gkaYmfApmSt9+3iU8XJdLH
BOs7A/PXufBVb6NjEt0qgFUJQJFOeQZCRUtW41bHsLwqKWnogxaJ+g784Xh1GC7Y0xHULx95AFfq
Qw8NCizhMwrO4z0D/TLnKOAYohU799a/SHN+7CID1mYbcvgBmNK1Vlf14To81yjDqpD6a8L4GE1l
Agtkw6iUuz+f5g9LoHl3k9TeSXqboeSl+uV88TzjcT217Rqk9QGeNMJ+wFBnVH2e/BPau9/C6F8V
0Yn00h3D2N/dzt1EVIsyWfCGVmz3jj+8iHiJaJ9bC4HXR/0gRiGxzTME4x1yrjRM0N4Ie7ro9HLs
5U2/ylWwI7UlloLjgIwUGasNTz5KupFea84Sh4GJlyc6W6BIoqOGRXlfTgxrydid4dIHVzNFnu5C
XlIDRdpKlrQEOscMyf/y9a+jdOGpgsfAN5sjiE19146I6GJ/I6G7IVNFn3xU1y3XSolgZMnScn5d
0qrymAQkXZ9qfPTqgMaFotRZptrDnY1WkwtbRdKJPu5PudhsTKt6wDoRiU8LKkmfuG0SMU2MFZZ4
YhEfA039mbfftIuuPJ0NU6e9YeRO5/v1cvD/EoO71HCidxLAQkf74Tl7eni1LuCsfv802CflxO2K
o9dJUAtqXwYysVqOktuHPbiD67F8iB+zoFOXtbrHqIWeaix2XTh4s9rlkBHEOcASgxCkkMo1irIS
aIe+kQZjzDa0h8kqMcus2P/Mqnuo/4g1vAXAsOm18NOX3mn1o7Byw7MzVDw9miY/r143wL8ovPuT
Z8PxHcB2tCRGt/NeFGUkjxvlzlmpUFs4w9uiqPyP9hfzEomTYRQCp/oaWXA2CvElGxRs4TgTmzHP
Sp5MaHmPcsH+11Wmtsf6bcUJT755/V8SoL3r9bAtngJA1wi5G1diCov79t9gCh7Em+qjHXIY1eaF
lv+TUEI2oB/G24bYu7KZVdh8GdogMY7uDFZV7YCI7Kx3ltUODoI9jHy63DTHnWcfZBdfHQoYvzYA
6mQsTXjr8R1icYoTBXRcceGY9BLdk+zbmhQAOegT3flqfEHHBsB2wb/2akPGmaOY9Udn3RJAvvCn
eRbdvZ5adDyJ369ZwTgFNDApUY8+WhNdKr+ndd9wsAqpQXgImV31BewqYJS4ul0KdMDuV6szIoBH
KsZlq1KPYp5nT278dxRe1NB2MftFkZArCU3YFdpHg9B70lqDTQH19naElqKv+wo4mb/4NHkXsbBT
peE5qzsBXyWrpOlLR0/gNFTim+HFKtT10leGb6puHTlTPZU25cgGLfRE3stRMHE3TlOtJnad6g7z
ywHlMs1UfYC2WiBlECdKoOT8wvrgsyhTZY+4+be+0diY/ONevYnOyv8yPZLhYzxVF3Y1cl9aAOnn
xDe4iCrdMn4wx/rCJppGO/BCf/guGdSH+ErdS8FumZ/UNN4cFQEg+G98zMflqmHSXBZC+l2XJO8t
u0NesSHmlfEPMUlBFtPVW5JX5gVLOXNlrRxPNFCAMtSX5lC45b3V8x1+XSfXcmjycy9HaYldDFzw
SaaqXYYNeJi8YlYsmtXmbikJtMz3hnsStTzD3Zqd+7l0dVodZU18FVs6V4900YfaL7JZiUBv11bT
fF9J6ZDsZBRmgcgXEgB6RNWE2ooCGm2haCHRPiSrWbhlM5y3cL0DcGkMIoe9/zcdH5zM5BmvA8iK
ZePiWykcqIGWQEPdH/Sda3P3Ww4x7PnO9FhPCwivPNXbVLfu/4ZTAqnfEcUUIb6AGvD27OPKKHCa
s0r5W2rq1RGk9hxLlC3ggFXe9w611VhBZMIIz+ZzvB9zBQOXlx5MF36ZCOuRvdLytprZZm4ZgRQn
HueGFC7+MRrytx556kJXfLLRSmXw7kJsOo0lMo0UogPqi8CNJuQPQoMh/P3/l1fJW+WQWk6xtNTr
Jh3t7+B6Zm10cmksQtYbmMrcxQFhB2wwZXtby0k+BW4oE2u1ZV03JdcWUiudOLd09GeXdazegCAO
YBGpi0YBj1dI/ieWmQEBX6wbqrLGdvnFz0qO87UDHuUQbqRY1Lp+l2fNx7tLECRnIrbOLyJcqQql
VN7qxPgRzp9Y6ircr75ZSUul13ocdfgJbTo9QSQOfEM7CY+N127bkepH633PZ8ZR8k/+I/hAyQc5
YHxSAepoVAjlkJMuDyjSsrk6fsFaQNc1E9mjwytGprj+BxSDI6tmMHAcHUYsN56Q4vgH9WmCCPh9
aqPuBcYZm369yHhMPLKcM8r16fVp7Ms2RxfxjNZUXXPwM27AlVvLC+5a0P3ALvipvCGJEIv0ggZe
2446T+oFZRjW8qbVzmyBCMgaFXaSIFG/zE2srwtC7wJt+mQ00O4q6b6SQfjlK3SIomu8BXWhi9J9
vg8i+OMOaeyoG6Abkpw3uYPUStnwtXjZSSydGr45x10Q7ZPfkRes5Qw7mMWoWbWh0eTygwOdfpQl
FJ5TNuE5MQXeXd+XKtoRf+Ne8Hk9Uj5T6X3QtDA8o6iCsEiVlqssfAPmiMevWIer8l29B8clAW4V
n8rfIuRv5QxAFGvdDRnKb8lfZzJ5VEiOu8I8NjHPCV/uzQIi+60D+Q/bPzbOu41cV4LhP+bLz9xn
thHLPk250bhPinrOnVmGZ+eWzXhOIBL5MptoCUBAyPfCS9FNKAWwImbRhCNJqcE261ROKBQH1ai4
WAxFJ1jm8vAoy3KfalKV/aaJ4nKfhv2HR2H0uSbBngvditPA7/1TzuStaud1xc5QKvDdgw+MjaOF
1yh7t2UBYB7UqKFscNblk6rJnwUqfGIrMESSC1MZ0n4dOgkHNZArfkj6aVB0XbkXOfT8oBRTWWB3
rS38xMCW+LmcvpvTf5o86wNHQ5QUAL3w66Em0aPglBVaZ8xp9/7zBf+QYrjc7+9+bFo8wWzRVmk/
cFNzUbWX+g/le5kr9WOjLQ5KwJds1ZyYNSPMf1znqQdU/KJaX6mZZugRldXetsgJ02RdGENMk5RG
n5DTCVpb69YEADoq9VsUPvg9Y3R4KX7O3AfchqJvoywrvxFbiHznX8MSHVfNFChVaqP7jZlLdOJ3
UyWbDLQiD4aURTIHKd6o+ceGsusqUtslR6ZT0Vc8Pq7MpZgZoZaxfdGPh/JQP5ycx7/is/3A/Hgq
S5o8Bg3untKCZaG6jXweqbKWzFpK0ht1G/+vWgjWjg++ZvmJEuTALlE36rH+5LHW3Ctg9T3r15bu
lCGCbyv+oIcTqMEH5iysGvBEQNCvIraB2kkGaW3oJgWiY8QARAHn3yDp0JjH0LguAjPTy7J62rar
bSgZujaU6vnfV+eLOD/YMR4PejTzqy9A+8IsUMe+4BMkCG+BrUM25CBZZJ6GiZsrL6KR/SRhoQgD
LynX59IDdxhJNXYRosWc7pNJYSqSVK6Kq3KZ3N+nOEU3sfmjvG2rPQ8asXLL242ykY/WVl9gQ7BW
xXZa2XkBNdR90QkJIA3mq9E+f1NFipkUmeGEInBz7reCJ02MynWe0ggTAUWV02KVR4gpIlbwq6OR
vYvzZTdvmAERQ10M0nsQQ46gk3vJjz3xXk2eygHS1lsHVIUsRNQHeYXtcoCR87VCbDp2IZKIe4ph
vtYcA4A/iTcdRuAXpwqg1zr6WnwMTdGh3LqGaxWm0XhbfPnDFJozgGlMqwS+cMnGMhfbSZl9G/OX
KxbJRr1vSBLKa62NjHj01yxHa7RtbOuCuIXIBkUKlLtB/KTvM7VuGtaqKWtJtjOdMv9z/jJoiYU7
lPUWbTTh1FgaoWXsmkm+8ZJY1QohGvTg6j9u1FrfnBtogO9Y9cq3Q2jFF5gcjuhSbotI2Qn78NV/
kESoiUwsKSnKoTu4HhAxdQdOjmrKPzu6bJhyBNfzYAaeypn14qVw55nk99MW6t5aWJICAGQRgnjt
q5s+LbZz9bAA497W8g/tEqcVBCyS/yfKs0yEKJgTHdrt0V2+t3oTJLMI6/+R0DMJejTN+dYgXtdA
QFhwQSBiRRRGA5CvVAeuk1CXqiXRMo49QXuniWBFLgGdyeQ2ElQNq5cfJO/CIJLGFAuPNcrAkfLo
TvT5WgIZp76R8WJ81GMiyqi412+ygas8/wmkbPmbh+XbVu25k2YUvdpywyyt0z3AXFaHfE7G30P8
ikOp0L0Mu6/zIDS25aYJscI/n1fg9fOlRwoUVNlO5i61DTgLdYcqZiQ4cqGTpLSaUMyFWtJvT3Hk
4ANfNwQxZZq4czcXEVRSeKZidBr8ie8df34hogFjSy7D/M67pnaO+EEZuMF+1/mQ3G8rRrQ7f0Ja
VbtsE3gGfQDWVxUJurWwBv77FiUDXMnBhR7D5U39kKeRCvsT94Pcg+CDzA3q6Ak6+g1mx5AJr9wm
BIZUJWfH1zDvhDa/Q+zL23O77/VBTB38pvyYtxsx7vnFXsYK9tQPUJ6gEcPv7yCIkmyNtUs/YVW7
1ekTzFZxcKWdNJUAZDv4cmcDpQPDsRCUoZNd7lVn8n66VnevjfemCeR9U67ObRzAdq0K2M1MaueK
lyBuGS+PUFPE8D9Rm4Ez8wiNQwgX/MJtyXAVmriW/NjN4o4vSUQaqhQWIJoMJlPYopoynCEqdRa2
HiIgRQJiL05yaWNB3rxrf8JRAj6xiSUqfDsSAMHYEW8Jhy0YsqjsJ8cvU1mO1w+kWP6ZOQ7TP382
jgnC7OsfdsRAD7cqCF2WlSVBAhPd0HLKQS7bBz6VQJyR3yBDptsvm+uZSHERUGYa3f/x1E7reFYJ
7QAkrt2qJ0MnXR7VJtc/0s+24b2AumKdNf95McSaT/+/dv/ZhCR1g5bk7t9uR5oUOfMLBq2sQRet
c3NXUUK1Y8iNzez7DWySUpkorDqES/w2cg3MXocPQwSVptV25kbrAHwFaORg3KtR/smNmO2ab12q
X02mWRXTpt10sSjAvVWEpr3OcxA3RwzrJlRpD22OdUptrkpglYtSGhJ355Jcp1xTI/bQ42hOJHC6
hfK2MZ8jK5tc4VWV8lwUDmGOaal0cGhlV8TbmVUDjzQJxLWAwEaSRz0wdoEuN+zbuc93jqsPG7ow
d/yJPE1qgirkdISRdtCgEWVAupQOI9/I6TpyKaJXnQf1utASK2ChjaRhkdzXntMpePEtU9mSagKv
YGPrwv5Mv+PHHXjQ1e7/EFRc51gzW6HHG8o7vKqh1TCzYbPuObXArAY/3f2/R/iEkJ3p7wc5DGWP
RHgMnjfTK9BmbbBaCSvlIAN9e2o8o03i2jkHBQqv1yq21jQyv69qqgd/kth+futJan2hQhyN5ujs
Jq5uG470pdh6/yVSCbVPFMyPxDs7P0L7bj4g15+IYquV5bqdVh9pexQEJteBmh0qHHHDiKa6eCWw
gImEiuoUi1Yo2k/zO1jzZn1InW7apHz9cEd+PptY2o0NsqywLa/bV0pFsjHiHzXtxGvf8qtUpN+t
yaKdiIM+x+JJhV4Ofykt+XxXMHRBiHKMy2cu2guDKTDbkuU9iUi0NwNFHJ/WgLFuygwVMKXkSzmi
tgK7llwTpb4LvrNg4JYcqEU71H2XEAupWVGwxO04X+ieXq69KY6ijdBACN79Vmdx9qslw/e0iMAv
Q5sTtT3RbNMdNQ5/cX72v80eb4jSG22e5hCTDzXBVE5C55VVzNONvYFLrkC80w+PSANoaqxp5O/c
NaN8Qgtbk2GzycpHaSjkKcid4r9leQUmFNot/DqpMD/3aGnk9UmKNU6FZWathbwcnI0M27IS3Lie
HQvAv8qyzMgTAmj9DPw6cqCmHM6MhJKwFwA4sWWzKme86OZs77UB2KJV4gRas/zCTX2ufW6bI3YX
Od62BkpvvN7ikkrTyV2Etz+A7WgJ9sGv0iRwX412b5HkLmfMV7B3oVZYFcL+eaPL5tIFHtczEXBC
bdEfVx9SW29AyJ2phRRD95LhHenj3a5f1Y5pm5UH44qeA1hd/rsvL7pegqTiUGY0vvUbgx6Ce1QN
zP0oKETV/4gI1zmZRh9BMWzo8HTYP8TTRI6Hq1Pb+gYopydaUcDnAr6hjI/Pt9lAZS2D0uyrq4S+
om0W1D8gPZyv8a4rWsYCPSSF/2Nel2z9oqsFvMu6mN8D6EsO7lIrB3Tvk/jURoOYHftCMbLrYt6m
ZowTf6vE3KfGqL7Xou7WKryjZTH84d6RIpRfyJTbMib0fwKHqg95m2s6s76jTz2xVnX7gOIhKHw/
9OyCF9QzMxmeR9EXu18aZUwANEHyw37Oxo0BiI/34HxDgOtOIvL9jpPXC53xt16CnA4jWU0Nj9Ue
V38WBLHypcSZl/d1TP/Mz6WGs1GyPclvFk9W/Yqs341dX6Ibds565BMYIXpsYJaTZxn7TVM660Bj
eRW58PVAxkpnJlge2n1ZZDtxa/JX/cyBa015lVU4H5ESuARRdVU2KFxcLteRD/5lXWG4r4tU0xKi
sa3LZMAehcmUz01FpMJIa8lmnpWIc9vHxblXMZ20AQ1lSDhY3dPMNCltupqRsS52tlo7paLX99q0
KchNSlKWKeZawTl7iUFcgFQqYYinFjjzxB6bJKpy+dsdPZ3hP6eokM4gyBVpKywB5cZ4WYkpz1pI
2lxl4WGTyKc+qox9ooHrcHtRRyjwXDm6tMdy4Cw6ql/MxEnFePMNxweRxUKFJ2gAiobiTmB3Ao7+
yoY4iW0XL4iDjrSrufFA1jtDQ7nIQZPcESnDrOLkg49rrYBVqyfOOGWtTuhpsJV+BPSyewao6DyN
+uSuYvPEZTcV2EAQiNEjvahZnJYcaWW5IQ6EVRl5Mudv7okHGIIoogKmJOaFi/PlQbahzJD7S9Mo
LuT+MTW7vqFd52rBzvfNZwz2S3fY48TB0Wuz2G+1fcZV7hoDuTKNSFLuol1MsF7Oa/J678YQ7UrY
Voj1AhTgE/uDzUdy4VSHJs0pXW1IfGPXpom412f8nQNsn0tS0Mq8MSsAxIQDWc3vx5/Y4Cuu3LpW
00Sr7PeDnoAisyPWUfUAoAR+oT3D6osPoA3ZisfMGBPhjTfvh79JlyJqQP6JJgzzGkJF8RMY6S8v
Tjj/FqAj2oMgZLqn6m9W5EWIskMuqzaZJ93gd7fwZB9rTmmUFLuiVFCQHfVD5KddWERyyOZZFq2u
vnElnKUURQxmbwjSs85818PDA5pEuXicWSSX7DOKJkszJk6tfako/3AJAtTo1R1F2fI8GfNsYKj0
KF4TGSJoW27AMkqahjS7d/x5yMujFi4SsEJlx/7igzZztuwYyeh6ay9Cuna2yXgg3bC9SMXhGf6b
NK2UeyQgi7xTZaKSkwr2rsZgiGQ8cnzgCztSI+lUKqHBuZz134ldyaVcrY0j8Md6CvozdUOeS6mV
ep5VIxM7CVOCuGuRVaYDTlZxni9MpZKvDXmgFvbVELhZ2wurdBinAgu8VzWbRvTdVqfKq/I1op2o
unalezUK7ooqIalXXAMTRqzVX1l2DiBZc3TJ/TBUODvdgn3iXqcprFpLZ71pxZN+TgBw2mvMErDT
RbiZGJ+PZVKVhjqfr/SbOptzG2af6BDR8c97TSNuLjxDB5S+u+oAep+6ic++TVaEi35TS/h2fRJn
EHDuuIFJzLBA28XZIXq03odM329tamfsSE89wgv1YeFC1OC+fCqIF1zcD3JT9bhO8dTOuv8FW3IS
zqZ19PGcaygCvC0SanOHiUeTzN5YM6+0RQiT0it0hjLd3gxvbTe0roHFpR4aS3WknuMSIoGDsuyx
xq95qHA4tbfYOgEKFOfCqKZsPuFvAH1Dj6IOHmgxCdUVaiZOWeMsfByiWWocTyfxRsqHiyujmiGb
qzOlZ/Z5quWNCwvJdD3BYG5ESj1m+rPWQChMuQ6jv4zH//ZnjGBNfmj55TSnWu6QEBuW4/wGEaPg
Ysp/yqTxBTHmrWCpe3nNYQ/mDpZLijITRSLIZS0h3wl8Ykg5AcqefmWABqg22DnB5rKJ2SbSQm8R
f30KdqlvSyoXUhtveXIuGh9xAq+M18tNN/HV+DxkwyNwtrO6cQPPERq/vC0CgYhGoH7Mc8ar2qvB
+RMu/Zq+Y2ULsF648MBN2jlEjuDZGvw7k8tmiqlEC/DB5TWzQmZdVigAHiIfDTOdpmtHlygGrnU1
SKZdcxRmEtb5ebsTaYMxkCQeSlE+/g1A0U9uRHM5URCZ4Rmj392HXCIvrjZNqPxPGH4YqvTdPKQ9
oyFljHgQkeyIh9aHr/w/7h922iBBFTQkWBAoaEOmFwHIPnaFdi9IxNTC4W2pWjGOXRh1GXT9/yl9
Lpi4nYhwClAVKIQtHWdMlByc9UknjKYjZtWBzlk/XFCLgkEarcyvdKHdZEmKnAqJ0L3rN/jyxaIY
JO69kuo3LYiMjPBIbc/QCV190zRMVBRQUShGqFrTBJBGOsbIegJ0iRwVER4EbR8KyZI5GHGN02v6
N4HOfSKmDGVPR12+G9ZRCBDOyrckqGaAPJdwbf0KvWiaAhO3lpW9FEV0tUhmA0yaCB9AxwdZCY1H
JVYCC97E8xtvfLY8orBgILbGEG95evoF1dDmVmzk88zEsr/5Q1gbxCYfy04J6R3wpgFlBK1pTBqK
dEJbNpTx1S0ojacx3s5MBFomzX0qXqVB1M84tp+PDUbu2a8I6RRdbTdQv2i4JE1BEQC00T/IDfWj
HsG/aZBOimBsNfHnnHjEecdgVLyVsG+ZhOcptZ+frKH+jMb0SnqI+by2tttyAe+01W/mLZLmkGFB
vF9hdt7FcdaDaMyZiSxTphDdFPZzGz9ASI4cSnzdv7ujZTGZOrtRa7q2+fVpIeyRN1n8td5NpiIL
l8MEx6gACELitF+QVlokGmR7VCti+oUhN6gv44hFmkhqSZUun1Aqmnrm8ftZ6OQspg5dAmNpREPq
vX69JBMMGFEvQN+Pp0sgdX1miC09tXb/qSX+k38MlUpl9i8mxoOmJMpVaAxOYV5O+woAeckafi4j
E5mlz3qdcKRAb985b7gyrCZ8igBcjprRJkD15qiS+MaS4xSbd0/B5cK9sJAO5dEEofLO6n6wTPDe
eyuqu6GIL0Deu4oYe46nHVUMEWbIjwRkIcn29lC120ei9pc6refprj667KbYNrJ8uDiVT2cc2rkj
37eqr3bxY30tZu+f/0FejGKea1OWhcdTpYiBv0/r4u5dWU/3TfGxwSLU+r57f9HdlbCaSBAoYFPj
dLjbus1EMVHpjcEagNMQrcaJbs1hm4vGNAg2zceB4NqtEFaM8k4ls+b2vaxQM5hnT9ogz3wb0+b2
5ZqRt5YLXENkz6aT5g94c3Ls1XD7J89xXlIEBoDl1saXHLbVj8sZPTnWYa+mec5zVJ6XfVwyFYtD
j9Vq4y4ypxHngOA0zgCSniEX2b5c2ZHJN8lqxPHJza1GYVMaEYjk5kQhWb2IjXsXEt2PBfBE5rVb
6dysGzTjTxpHmWMS1QufjepmqrqGjadKBjzr54Rmi5lmbbB3/xliTDKaWrYui9jBaGdSc5TY011J
b1m2SH0xric9lEHzBCNIagURUP4qUx5Sajhy0KaksWEMbejKq0V5nCqB11qwxmwE8zqevAKBb3xT
Aq48MTE/CsPjhR8s/xBsweg+F5b+9UgwwfZAZSehUlfCKFfAPKsQiB2XSjaQO5+L0EFWzCnLRPuh
Zpx2MoOpkMb5qIhHbdJOpMuqlvMpOW8jOKjQ3Gc0gNAUaqrNcrAdS9I9jtVu3zU+C3qPHAg2dIsl
Zld3fvSXltxFQZGokIL/Azwj7WtMUiYyK5svZD0wGCfPlUTkRltyyZ1kHK1PSIXXo2f9/Uu8ZtQQ
pTscUIMy/fTlEKa+UpZUnYfkmBsN52PiRelQ4mv3Crix/d2MWF4WdtTk7P/SZ0TDDi2v4JwJmrex
PEQylbzaNg/LSlzU+I9aaLatdlXpkD2CkqIMLdyE2NibV3IKBoCpHCUws8UvDbVqjgL4/8rQk0jB
cB42bMgmkEIW60S9z35OR+ubECbw0VfT5EmI60yx3wlUc7jVHFrREOTqx0c957C6cfxA0NPLCCCu
eA+GP1KerIHW2GCALDx6a/D2qOQ98EDeYgUeCxI/ufjskMNw15pWEMG9iHnVtnRCGDImPG9icvUC
Z0NbjR3AskFqalRQ2zOQHEcszYcEGaiO7fYdrgZMUWSPZqf1QQaU/CB7fIwkGn2Jsf8w+XIH1J4W
k2FPtjyOh5Ut5RBnZahmCN4Bx1xibP60f/n7wvkLU3a/zlKRf/j9PanIZq+3AAXop4JDskjQSSfp
hJYxUPUEZmoxjepnMZUp2bPJnnTM9oQ1ok+3wzsxpEv/TE6kvkGkNpOr9YxX6YOsKILROL3Sq/cW
EeSOkpZ8PFmBQttMloOLyKB6A/45ShU7oeGc1pSpzud2mOKhyngaYxpGk0pGFTmPX9aF6gIMP9DX
7WcMeIahP7DZof1Sf27w09lbnYms3nDRMkrNJU81GKpUAHd5AFf8iORAXXj6zudSro2BBzSYRJSh
2GeeDht7uBknOUweStEXML+jqIgVf+0fTtRqvC4vd6uc+r5DW6eppswx2LRpoHuFBngRfRB6tkM9
kuVzQcBayJt8ffAAQmfRz8ww12JUG8TFAy9dq6fZQRd34EcqaHJA9bIOwKmcl26xDwEKiI1bgiUT
eE3SRNtAlD/GCQ8PJJM5WE3kJJDJTa3lAw12OVUXlH8oHtj7qcg4ANgdchtawNmDv/8tBwspXf0V
8336EgYDb4HUzVWiP8RPuDlH6tFYN+eR2kjbotsiXPBOWSDYtttoEq9rbDXG1KEaaW60d+xyqpL1
ZVm2kPTkazqo2IRQ6iI+2t2HlmUfS2W6iBTRzQcHdg2MA9w/i4UXiPJwj6T1qS7RszGYPWisPxMX
7illAnxR4JicOhTPXMmgulj4XLwGwG09HzvF6ml66ztOdepmcJl9mShJTa9XG/nUyhyEBgFmEvxa
J/6A3uscWbj4AZoTx8sDJrIdZgxp4CGARiBFynMjyCCDaUarVF3JVfUhLvPUPvyw5mikOIz+OC9V
pg00YsOaVHfpZyn4/sqJ7NN0vgYO+Y0R/NQfxFn7GcicB0MLlIwqP7yZCBeGs5kB3wkape8md1qf
nWNCdHdMSSb5qi5VWVSCC13lalf3lIBEcwg8cG6OvzjZzBQmry2rX+AaiI4JJ80T1rZPjDeCyYF0
9FrSXM5yuRBJ/s9sWKjgMnoEAMCjXfY4IgwL3PxQLPV09rNy32QW7vJbT3In/Bx0qou5W0ZBkYHb
qGgqwZz00sXuZ4WSVOrdxPW1Tqzxgzdt8A5AwTtZHKyI1iaIvg4cbRRRhK9bNSk2JJ3iXLDwDn41
beqVzTpWAR+bv8HagLUXzdHNvq595tr5mQwcdWwCqC4HlXRkA0vEp5N4mFKrV0UseIkuzOMGSaC5
wcNX9qNV1TRv7BtmIlaV1LHSiK5AeAuVrKw6DvkPDTZq074f+xDZ56riafNK1auyChbjC4VkcVeq
NldemIgU9iyneJvdnB+ybBM7ljo9lluW0U2jSVBpA4pTpTnwc/ky5vy/odi6c5IqoxxYfBq/5ryX
MHz9vM6PnMp3u/rPxwaqkR+cEiSYypt8T6eZ7W9dvfMuux9fWijcvs/GrShMxFdCIv1rEIPMzwnK
RMpjmamNtf4+LFpfyYFxRZK/ov+665cCkSoZ2Mta9PQXX/3wwItSI8QIItC5RaPJR4oY2SqsU8Hj
YyQXxIxWg+IDrleoC8+3VSsGJnq19xplKc0Qv1h74Wq8NM9vlH54A9QPk27WcnhB4cyBc1ZmiuNf
VdJ+mK4ytSnMJSv+Mji7FakuXf669jDVZ0/gIY1RJjN6g6jywiLFVuaAXZucQmfqgZKXBNCPqTwr
mUhFvRwe8O/f3XfjtG5mPweqqv3Kn+TklCgS4b3JH35clv+JZvAhDxLygN0fzgRQJKIXu4BBoKXg
BOHlPnN1evti0MDQkMhhf7q1Lw5Sr5aXVg8eRaIGVUZb50y0DqolVStHygMgtZ1pwqhuw1NopiSc
F6TOZF4g90uhe4okL55aysN+UHX7z6+s5VqN+y0Mby0WloI2bjclhH0/6Dt6znarNGeWdhblO7iw
2i5Gby3bDgxZsn9HWIXDgmzLJE85aKAnPF+PrFlUAXQuCI+RVvrRb4YAAjPUWIkuZXsAGuD6Sy8e
y8fHHj4glIWGdsWcAn0vxpJJf7wzX9xfnUXiwOgBLtMtPPeJD2QULd88qOFtlcenGx4fNVAScSF4
yoLPd03tiZuFy/MOTODnsDr3+MtCA1nU5+8P/6U9fKGwv7DXqvsqHq4tndBD2Rzx9RIDOJwZypdV
1DnjhV7gzt449xUV+y1JE2oyulfKGajEqLPSAyZwOcmfv04xzixtEFVlmdn1zIjN29SHzGbLlhWX
eO1EB6EY6uv4S9G7nx3GDo3EM9BfRg3rj3Xw0iySXh2KmwAJnx0tMmw3EKVhHu3XLZdgdtSK+s7a
+VfBsnZRXYq+pxcCOi8CEU0SGVjdb3Zmwg2Tf2tutddeTenNmCnt1HdJfhF0VsvIEsR4dwbP/qXP
9tH6OLOUMZBazUs7Fils/1iuYERh3r/Zr+lPDNq8Bd7vI9X7jwAT4K/o37V7UdnItyzORDnubqrs
kbvoZQatFWzlMjjlqMjbjSZERML4TVXMyYUJeB9Ge0WTzYVZ2/2GW7AQyYMRi35yhawS4WABjAm4
8SnDCh2iD8ZdIYxDPUunSnJLHh7LyC08lxHgVtpI5gQRMu3NHPE+gsXhx/8FM8qAnQGC+5nShSsX
iKGICOP9hDeecBxwSr3NHWWti9aXxP7eqHB7BV3c1BMi/WoNaF7KUEAeVu571UjmmiwZ9OE6q/B/
RLl95+uyFRaeTU6LO7apKawif3+E/bB5SuxqpKjR4boApr5MsfSnWayZQFeLu1bJBlDH4HXxoLpg
AzAzl00attyFQ4BDlz1ishFh/65KkTGFWOv/StoQecMEiZQrC6fW3X4SgQ7wPvh2/pafaL9bH6vM
Z6D6kluH3FVyqbZ1d+md/iicTVtpMrSSWT3c7NFIMZL6Jq9UTkfRbR3yQK5UYKV+CW42nNrzNIuz
qmadq8kJ1kEJgTMJMRbXLnJMPWkDpW7ZItcobZJS+8907TKh1tB98dHRo8j2W6rmTZmNX4oE+6Be
uyeMyeDWdS/dpwjQBeP65DqN38D0yiZd4M/W6nDQwIknqqHqqQfEIgt6dZ8qfz0ZG6+/mUz6lSSz
KKjYAA0ikYUoBOuVNDAVQMUO7JAN7SxtOidBczCP4kvHyHOoeyKDMTllYKCL3CwJTSjt1UMhU5Kk
h5yWdVh1BHdF9UTLg6XtHiXRT4GwQEZHUte9Z6KnnsSaBDRn+Zfwe2iWU+YqV9of7G4UtUh69x9B
me0NFsWzmX9qo7bwBZhjSEyWGWa5KfT7H6CsO/82t3KSust1bUk01knOxcFYBRj1oOFMqKm42XHR
GBh9TZwlMkks/yY9DT50qZvadmcLMNcmTaJvlA6H88v+FyUblUJiAJcb9e7dsh/oY4axTjobvhnJ
qkx6mtwNVtiYHsC63A+ZPHhFgmCKf1S/ipEKaVHSc+suHwuYkd3kbvAQ1yLDrHKTXUEmfCetUaVY
WbqOXTSPPUW5ixTKx1S0Hwx3ZaIcSBgF5dsKJnBS7GoAJibdAHQzM7QKmYYFS3CBByOg+BYqfvsO
W9RXD3o/ZPICBZd1/T/7gN9SBYQFcMz54J0lnZBQvQph8VjRcQVwK5bSPx0XJCPn3s7RY0x5duCt
2wAECDhHkkkh51WjCtKQ8p3zbttt7mUlk1Sxc7ITQX2/D9uGMiR8d0Y6dqt0v0FOGeFGUTKk0JF9
vSgPqiu8q67d+uqYtIFFQMJviv9UVmFYjlMzZbIvUm6tJ4hZ6hs2lQPAplXHoTJqldHER9HEzMkw
mp/ig8ySZo9kOq+4tyaiF3uIFLRRP7WnHQl+0uF2jDf9B0o9jK7L23B0WvgEFiMnrcBcgHMOz4pm
yx20+e4vvlUHzvuob4LOQ5qbPzYqk0ExiOqxQLHKueeQH5xlgNdsOSfVkJKlxY0JP+ynICWuimpo
pjc0yG3oj+e9WCXCoV6k2zluxC/xTmezXoe+VydqffYzxrRNDFyZtQkCVZjZDVwwu7RAOmlazd2D
T9jYuZ8e/2JNf+tOP4ty6mn7baG5Ul8CU2souvU2eyiP3+pyEG0cIoREZ9HwELJibvetaHyk6X9m
AV9sIX/nSI71SYP1+TR6/sgvFy7TJlmVYaYlvnbt5mSWlve97ej0EETHKEnME+n3KO7ejecngr8H
snMcy9vc/oiRhCKOyWL25eJSEHXLsXbWeRM9wIEj3+3i8QVpKFxTyq6+WlkET4wXe0XNpLMCBRjN
AzZbq1MALHeQjmurhhdd5VWG6P0Pg78jQhVI4JPcQwe271HjElSYkhU/m3+f49m78khrwD9x5PFp
JrHwFSu861MR9ZBbmrPxsvMdIL79HUnv2xjSYHjg4ZQK79DWcXDZcU/bpfc8KGyHoMFJBdb1MPDX
NNMKiRYoFdq8QMrU4vPPUlXw4mF/IhPKKaobGmZLEPd83lCembW29caOmOKBlL8GzZXgFvdVZzse
WF6De/VTyFsmiIx6Hje/aAGJx9aPEE6MoK79cwCtwC0RI8jAJ4R9sr1/QQdABzT7U5yWAIVPqpNT
6zqCmEfyUY96VJ4O8K2kOsxi9bBhlGJJIvQjyXvKZOL8nZPunFm0F5UVOUC25AD2TWKrO+RgCAFI
92HAgvz6BhRMLIkXGjZJrQcVW0JEMBEByeY8unDrLYgGdREyEeeZv/v2ZBNPmG7hxpUVndCgFvLx
cbSYbKD98+SGMl21NuFKuQPs8lW6hiqSXhqqFXclzm/VlH7OT8kBoYhphF9g22aXx1MAzbNRV33+
licDsHE/r+Hy9PMcr59of8Le7sPwqnabDyjB8Itf8a39G6yuTLp1v9HwHYlCw0qdkrYk60XOVYQ3
Hmo+Va+Lm6MbyyEt7B080898y9aRgrH8FuudSltetC+RNaDQPh72arpNcmKetFrMC+7mVo5gHNHZ
YrQ+qdSwnga6P24UVBbNvxw4yT2oJp4FDB3hi+4ADXvL+Tx/5V1MSk/afzccn/ny9NhHPpV0Iwdc
+mP7YzZZnbZbiE54/uJCW63rHucOiwITjkgcJl0P7QJgWMSvkQzVAAQNTdLnvKeUYzIHwzCKnhi7
gBSJngfcBr7sbFBAHH5OlhgzjXshYD6V+WcPQQi81BrkuyQNjCpBHxJ3Vc61OKkgddTE9sY/dWw4
eaNeNvzWB3ptThTLgO4FTDrMDZLKSJwbNuYa7aef1B3WchAzZSEE67+UlFP4ZNaegjMq47+rmuuK
ydz54V9FjDs43fKfmnheMGvTxg55C91PZ+hPdAkc76Ms8u8vMXWeA+pu0AutBkgFxScGeaPFfo/O
WYZ820JGR3BlQaV/zB9Fo6NuOUWDcg32f2cXSr4gZuejEaGWM/xnkT7bphrBF2den9LGLmniYAVX
sY7Z8SzDPABzR/+7dIzqPurhdTVaG6v4aBYCP9Dw+vs4WUm0qVO1pIoyEwuDuSeEkW4FmvDgi0SO
tMJQmft6leMO81lG4aVvWPWalAR5gDqcLRBcv2VMMPMaTJmd2XzG9xjsfkTogwe+vRUBhuwX+A04
OAKrQJMrrhBOM9KqoID5/pxhQJ7WDC366QwgYRfKbczgmjuAOgUVjVaxC4qsHNtu3SWxDdzMojxa
vSIqBz/7FxiD4tHv1NtfC37h3wHbJZAzW4xfh49rM+jihwaHASSNNMX0Mersvany52aV0HNg+lcR
g0RHpHLZOF/7J4Zdxx+fy/6VGvGNw4jl+t5zRvIpbJGboFkCaAEsNn1cije3XpLSv5DnhLUGRjlS
U7VRtTzKGLgE0VDPLfT8c+aRsvD8vP9IYIlyjorjqC1C5xzwQfsneHudgNWxaWs9uIWoPolhwmYA
Uu8cEa76kLXSZXrcgmVrWOyihCcN4uMRZ+zcyd0sZX1kOertCya9d+Vt0HGdv+4DGm+2Yu5Ujopv
1ASM400yu/lQnVJumAAjZ15VBgmnFUsfC/jlLzRbMH/RQF0n/v6YyIlVZw97x1I3tH5bD0SkCBjB
ao7PcwYtXhpYOCeowAlXAapu/ncH7goeUeIHzCqgoVKs9XqV/ODTwuD53U9944PPLTFlf1XqpRT2
U7bOJzP0At0r1SGH+UJzC9I10EtDLQK0MRMG+k6rgIB4y+Drgz5nnwaLAlGMoFJlaG69PPzplNVI
KL3xt4iYXHPjWU62jklmQxuK+xBMpLBiRfVknnmsrF+wqPMgSXMFlvIS8I/i+PnLbWSJp8t8CGSj
R4MbYd2tv5RxwKD4bGoN0Q3VwkLKYPUrhKAPUp0goL8GBw6wEu82QGNcMUHDDw25qLfgz0WnAH2N
P+K0JmrXoTF7McO/0wXxaG1nN6vE3Oqduz8/fei4DFbLAdbSR3hZZEMC+IqCCNg6VLHQLR3pGAl4
XJ1pda7t6kNP9d873lOikfbZ9MzPTuNtX4jeixc2RvGFFy8Nv9b+6jjahl8BYe9c/Xjso3yIM8AL
W56ra9aCfUyFcBt2IoEHLuhy8+u4suCzNfgM12epV4WNqkK3d3fynReMJ94xg23rMlfvLbH3BK5k
8TuAej363kJe8fsexLLWH4M/W5YzeeatI70087kGQ+a1E1uFzLyZ1IyXpQMFtECej5ykTFhMAasr
Bdb1M20BaAPdbGMYRMYlbHvCOmF1OaF/tvZyIZUqVf8f1LS59KeVi7cObAgvSdRmnsLYZwJzOVqU
VAD6dJ0yFlGkRM+KhdRCCktI1D1QWsNaSoIbDUI3OUFHrfhX1D+IUHYz1lnXyDvI4HxOB+JcYM2f
ltAAX98Ixle0flN2sg0MpBGcVwTn31fHltaLJlitvnBEayFFOnLZc6tSU58W88eUZDAeaXQ5whwl
3Ph4Ij3Uhire05L+EabmVqFcqgcBEuXgOHndJPztBdabHCR+o+Wj/u1bOk9QIQ/8VyYcC0uUejpz
gNBADFiudJXBnlEIMcLOFfZbEUpcR9MRSo9dKXbqMutEZGppRWQaRu0zc/G2hXWZHEjyjH4svriF
CQ+5/saap3XeBbL2jZURhDeVaTTeC6M9kalxakOxHvNSpbw2ncOqfqcJ7oRH8H0nady7a7alEfB2
TPcC1zGEm7IT4Nd4jEYR9NxsW2yXA/bTsNf5iQ0IdKiONLaVQgtWRi3SsaR2kDr0SMG9Ce7sFQQT
XLPYn+mqN3XHXzq0DHTHgsX6BNbCg6q91yfBNokeuy+7SvXz6J4nqfpxm17zAQv3sqfp4fnalOeG
BEKBJNvfnEhXJtZlFBxOmqSkP8b6ubQlrsrw7GoDGx2k6wvey4QQBj52y7JNaYwHCDqxAyIwd8dw
x6jUDU7ydf5xhZCyhrB2RzGXZsV0B4/6RGMr+oLNhktmtip0Xg8PzkK0SaWF9re5cmoijbo/xpnx
pKXMnckvA8ElAa9+pws2ypcCn8cOHj9CEAevucsR/nVhd9+LoSj2aHWj/uikUZOnStVP6+N/NBNS
oY8aP33DAau/7VLx9+CT+JvYYa9KZM04GtC9iQF9UyBBRPQ7kkUtj/CRaJFzSmB6vS5Im/xnokG0
+yZk2sMBoAwiDBtowUEI2Rfk2uTtgEBFK1QvE7J2L1U669ohcBcT4+tbi2AsSkh7uBoUKkNIY3v9
Zh6oytiLdUtHFTwziXoWG4dhzr6ePFqKVqCAaBtDsIJgMPaGDsSl+g0aixCJrxTJQ6lULCLzQ3J2
3qVYAKXkxLkj2hH6c0qfKKYBwWwDzfmgVlFY3r7CMQESdY6neNLD+WpmSeZjmeaLmaBv+l5KwMLc
ZHveJ9hThwqMvVKxCpIJfiwADBjzkq984LK8qUUaqyiRO0+sN3hC2BZJo2KYGicEstZZa4hw/8Hn
N/7OeBbYLPeEsaSHKQS0k1DG5kxvgZQ9P39pPVh95Ua568EvbwZ7KQ6rZdDbwaWubvw3hJrcdMK1
XPkGnqbRvdpIj23+7L5XvFHot6IYApNiN8wAdBIR7Bbf1jApSkzmTWO4YcWMbYVdF7H41ZGOG9an
sw5b7Id2bgFiMKfetxZX5tAXpTVwu+azu+KVwfLA/Z41f0r4q4xRnXevebvk95fBg8jRHSUXhDnR
CgzEfcF46ZtuU3C8B93U/SMsjIdv1nuFG81wIAvwC0EqBv1MJZPnbw68SdJRHd7whp+AEu9hm8aF
aHnTqHEGptur3d62xWT8LweCZb38icJavNk7t3xkMnI30kQWcLLrzbxesxNtIaZVVXx+AUr9cr2n
xR7MmyK0KYiLUe8Jz8a2LVHgaonB+HMioiU6bjPv+9aresIE323/E5bemOR6gTddVHt7Si90Ch/i
ucCnad4Y60NeN2NBGCYSatLsQ2eKNFQ5wKhL45e0fF5yzYama1KuwWTiKJ8hcYANcyrC3h59MDKO
8BplmeKRzAZMG91P568RRSnkCDrPsCLrECCvG4//qTEhK45AjRnDuk9IxzaEdXyvK5bZsfmrt7iV
NzoBaSWGz0U5RhG603vBoLFye6LTyG6wmnvferhjjHoGh+74TVmG4/7bI/2vt4+qXkPSMx8KcDCV
DM1KPfE4epcGm+kfURvqMO9MlakCBa3YNWPaTJqdy80j/HSWtLP22a20vLNo2XfEDF6i1f0qB3Ho
B6GNqho7Gh2IAaQPe9+x4+uyZ+DAfm6I+MbW5Mpm5YTAq+i/ObnESnJgOoFY3oujemH1aporEyG6
lHZR1P9Ctg9hrXDzwhN+POOoGPnGFm072a7+y26ElxlUizZOsUn7S8IPK9Hk89hqRQ9cl1LX3drS
3UhShnv08lQt+V0BBS+S2xPJtsUv6wKcCCJ+vhwZWs8e3KhvRLCtFZF6RYRlJ9Gs2vzkG32fY2TD
f4sYoCOVznw//kGFyKp9eyLSoJ/9h7Gc3FSP8ZbDEz5OxVnObfFXtrEthxKrrYsJVkKVO/pLyVgh
lsY2W2cQ7OH4IJV+frZ1JkTaP75GAL9ugO+5v5itNpv9oTYT3ofgi5A38261ae/mKwOHco6FhVDw
2icHVB4iQCByMtMh53OB1zanaOZVToTyHul+UDft3nF0hWiX+TrCcGlaMcaunMea8fbM1Vo+0npW
Wofc+WRzziqFSp0vYGIa3IWdq96CeFHhH2AR8Fz8IP1TWpcO0iaDlTw5sb0oKT9c8ldobtkF42xA
slF1HYmfl2XDuRUagCSS3hltkAss7ZI6vRkt3qX4pGnr+VevEh/213SWJGfpjuDsRXLW7SraTxCJ
eMJwqhenR+fXlCkkIPPuvRTLCjOqQbOlo4cVeQ1X7LoVJoMmo/BLlwmISS15rg1zvh+gzerb0gTW
3magdNlsCJmkWDT1sR/en5g03XpOLxLZog3G1FOQltSg+vmYiDuWlfefzgiab5wET7GKKehS+bIz
ep5rbCYh6cqNoMtclh0x9fM8jYKiwXyLkLPKIZrSWcdU2YMEend5Pp1S8EoZKh4dU6iG4RvlW2sU
6Ueq9w0qw9O9YOFI5DLUjicWZhZJnr+vcV/7Cuc3y2yzRE3H2A3R8DjMffktkpyeQn3W9zPcMt77
5vjPurR6IJhBaxAtq9sHIp84o/xyAzBY33P7rsfLbepJv0SZbMXFzSZd+yHXx1RHqnHvmMMoI9Xt
sw+TOQSjcK1MhEIu6qoyYwAGQqEQ15gX2i4UMsP1Gj3tBU55Mun3ueOQS/UHBC9VuYJ9itSLJ/7v
4yLted4hVsQeIJG7jl8yF06eCiQZM8uJMCRi/fwFfTAEGmNw6ux0sxKk1WnsAlOpGz4y2IU1wdNK
xgWqsHplNZ9TyXlWFeE3srpuJ9G73U2GPFvBNKNJw+Kb1yDkKvWpApFuHw1oKvvMC58cbMaVB1Zt
9hr3gTWM5XEZQcCDWolUjEMLlzEQLDV3xZlgzZmDWIWWPYh48k5K90cPRiA70/+1Zs1bWkCPIqCT
6/S/C2Vnan2KxvAbgcLfkHmLKEoyAPgmtdoCjZJpkWBSlVS2OAqvehQVmfGqIHWho+1E2xzUjku6
i4rnjTika0J+YlPPgLAHRqWgL3V65qupt7evbrAFIKOngrq3qEmyT9NKCMSFiwLMBH66Bpv4PCdw
kOs9bwJ/WLlR9+OGaQWmaz8bjdHIylnRMNrVtkdb2yJVIN+32UOTk90Of5jSvK8oBeNDywlUPWah
2GoFxRwEOtW9DhtWlmMEsyUhfVMMhbNu42vDSY2ZWwDydgdSFoJhES7ZkAbqUbYFPMtiM6bmX0xp
wNmHMBSq9SQETW/UJXXJ4KBhwTbkH95jNJa01XiQLCZhXI6WIJW6DVj1ypKqdYNZpPC+w4aoN7I/
tkKT1TKcz6LRzSCvUIOp3sXV/r+rElxM4dDVJXVus+8cR87STfFkYPGGVU57h3j2JfEBqKqy6/+x
vnjtlkuJ59NjzjMe+ITAu0gF2c6jeN6jI5iaw7shc7AcNqiLnUMIwDa9UWJhZZRi1OvIap5he51C
6yHZLktFvR6IEoLgMd3Olw4uARv8uZZ5uuGByelcfV9SU9LRxkLaDXxeVQqRUgwJtummIieVa9Ws
9cICuq85rMs6lviRK01XBakqvB2ws7avrz5XUZrU3glPYTgJmulwqwpvDiAVM3wOyQsD8y7IhCSY
n2FCA56J1Rbe9Xq/SEh05cFtHNPdN88wrwLmPQtD9JVsl1Jbo+5Rc8FDxq6JkOClER3ewuE5CcaF
YjEogV8o70+9mR1H8UWR0iUc3k7XDQdDmbj0KG/ML0VqhhkjpL/GwW8RQqsGfN+oF7Kr6ldotYH9
CIbXhqhFb8o1bO5oaXYYF/yYuxSlo5iQZuOuRYXtFbqRWnHkbpzlcD+CbM/7vl+EQt/u0IX4ThOf
ED+IxnzN2yfp5DIn3ZlW/6RmbjHlKvYUMZQ/6cAUB4FYMLZ5tckVVU8ieI0abCY2qo8s9Dh1hMOM
YsGNExnBUzwWeSwmyZavaNmT0p/Le8K2xfDwLTvKL1HBZ7W5xSOXoMV/EXFrmVw+CoAcbABBc3lB
gQuxqv1b27+xIS6kjoeL+kPJre0TMZnOWtv8ZFJ5kBvU/xEPtgzTpLZ6juZQ1OMJBcHRk4gIQJbj
ZXhD8maVF6YK106RjzkgrhkNQacgN8GB/NdlOA2OjU51xQaAewB4EnJ0P5gN6ALkcT+CqMZoJCzu
cV/x8Ya+cePuequVFQehhtlG2eixVr38ifUr4QU4fLUJsEYDir3xjYOrbjplw6sYlXE8OIyYlqFH
LMwG9WoXxditU8CR9k4G2dOfviu+aFqKGymwcs6zF1hoCIHKaxukQSUlEN76HOFhlDmvFPxJiznH
SFvqU8R4LclxW6AiVhL3UrWb10KUpEziQtYXalWxEmJOnXv7PDCqmQt08cpalJF/Xrojn5cYc+SW
v4ENMeDnr0ztpltO0e7IAGer/YtZB/aLAj5+cVPBjNZwn00x+rNLTMVfpiWXTrsAQBVlm0dGc6V/
UTNDCc1nv4qC38qen5wuvw7lshQvWKHgvshcjZF8If0JGyxZQfSrK9/58GpTdEg1f9hkn4zmEiDw
272l7sQc0DGVgwpFQOZigFFH3STPbZ5R1+eBd5s+d+WSMdE/zIMqDt/DmuMuNlJ2hM5epEnWydSt
50Md5HSGHxtfAh4CMHDpZdxTWVQq2BC5vwuScG05lt2dWZa/RXjEnL4AaAnZMjylX2BRcXP0gJ63
2bsXo3s3GkalTrnl0PqyKcV8dcMoscuodnEEE3NSUNNpPFUd5Z56l5L9vk6KRYTiOVwujIhFW/v7
zN0Q0bk6YLqMYN2Vymg+lCMtd8n0lWoBxK24EOGodGClMkywhV6hcTbkqhwmE3lJROGB5pCAcrzu
viVUo/55YdyCaK33HD2pBwvCSBxdG7g7prWa7TOIEFBVShvq1ef/uHvxBDNqQfLRbwK/OEmoTLGC
PcgjO7iFvXbfCsskbN0ZMmQ7YAOpxHgQE2Rbc0lik6Djl7r2WQx7jdQPq+FJrr4tjOK0eG0/ywXI
a9ISHYcJ9sLB+GlH6nKGJbgevHYK376GlHRArvywujOdHideRHK6UOASW05u1mEwx2byiJRj+shj
v8k3ox53Xt+2rKnNaGtsBnexo+tHNTb253Y/u6LHpHSOZ6iE6DMLVrsfXAYR/wL2ijzQfEmGxihY
UhHwlcE9wfyCUPq37eAcDuX7iDI0GgyyIYKiCm7BxHkhikJQE0lfwd/HwtA/DbRxIA7qaQteeuEf
2XeUb9DkFz6QT9E+dxOnThze9++e1qncpQvmOliz81yn9syo6ATF7kRgHgkTS5EhWaeYvQePJzIm
Vhsfyiz4M+5igQHIl5pBz9T0dOrdzlXhpELYEEpw9vwTIdP2GY/B/PKsAfVY4SocVRIl4SozzRXk
UCzq6O9MAuw1RnfL/LEwLxcwhpDONoz+UgGj7OjT4L+fFXlvyiRzhNM0t0CvfsL22DOtqMSHlaZ4
kj7w832xWbj5Day9VPlwElO1UtyhEaDP1FU2L2PALJ8hm0GOTZFYyIWuyYFxC/kO9ctEFl8v9/eZ
PQj43P0E0MBopTMBN8VKJotd8O+KWkHQumCZshgh2p6SYlwaVC+O+NeiBKmUzmdFehl+W3sl5ysq
OlTGwMKMdfYpQ+yDu30QPYLCahDpwtRpu0DrKo8DB1oYSXU2YvHwLPsM04PtU8qNeauDFlaf5FsT
7fej5IP1NthU8b9YBG8FssdA594HYIKwyD40lPE1nyLSIiWoyzYOeQW2gsTcjbzFxFys1dX7UU2P
TawTO0qIlrCFW9AbSpm0o24uKNok5YLsee4+fum0GN1BovuOAJqVAGpJtEd8l3FCgsuVtbKAcp6R
rJtoDHuBy1THnjAYFTjmZOHjiLLUFrFor4YE8sG8oUZgoxZo+9nZlzt96D/oqYdJE1JGm2F+0sDS
M0IXObHv1J8UTQiwi3F5DSxsn/e7eOgwBuWmAYysNRB9lpeIoXFVc4pKYQaIzLoR8N/zNCYZkaMZ
1q4GIAsIvcbAJU/A/wkSKuYoBgpwGjXV3XGEZ6RJ8MO14kufmZSM5lyXF1OqgZq4YqkF6VK2QH+b
ENPsdTVL1/UH2De3+9M0YjYYQXN5LGNO5JUSWrxXRQzXC9ligLLx/skZ42WKoF1b+SO028GMBMO7
S7FvztDwXiR4oUNhATQCZATiNYONJlIHMk5nxjrNY/iBhWZVN+kisbACiP1aQcTbQn+etcHAGJ3R
KckoGr5+IWoVEN4JbVI5iml9+A/9QLOjoZ6wFEPNpyC+JgckjWHT9n7gbwGOLeYtVJ1/3nHHyUG3
QtlHFqFawWxhiKUeeUeqf0cvrRdLNOFRLkCmgBLTUwnwPvrMZSIuOo+jdvagO+r0Wg8Ji/2KL7Xk
9UAsxEUWsQJkYyHXBuZhPNW+RETY9Pr4qNOyr6z7Gky7cpK0fr4da/BjlcwrwqUDR3NrfTA/Q8of
u1qSFrEUx8mfVwp6yXIaxI37MTri63lkrxtSWrLdCMWutwipFTlMX5LGxB8EUmj57BUruP5SEVDY
KFWi+dmpycb0hYW6J0fS8xApgqY6C5HhqtRZGbsICSizSQgfEab8Pw2JAMRladEXOazGEM7inAxt
0vjfgtQGCOoiJnSr0gUnCJ26u3AyvN0z5/BJzgqfYxumyG5uDgsLu5RdESl7knGYJ1el1Qhvmbo+
rXl0P0R8ZFlpAjygVaxwyEUAqKLplrufzgL2xMfIV5Nlz8QAdEM0PA0Z9sxIGNZL9YukmrVN+oRL
rw9OnmIpWOYxgkq6OzkMnPf58wZhpiDtQlwr4BUDrKOnXrLMZs6GIrr4zc8vq9HAw2BjNuaqEo8l
lEiXcBoFAhS+EkG7aP66I5T+xTIGofGsvFt2yhNEi2lWJatoSRz7Bv8DjwXFbfRjoi5yFEnXl37E
jGbk7a/6m6UxRkiOkKh66UFgPSVE5lQ/zuIh9aMnCZq7i2x4Yu9gCJ5iA/C9VbcJhS5d4ZZfJ8Y/
0CuzaXWfX+InbO7WBsfEcq2uayOLg8ePcmnd41rpjt7OjMQ5ojdx5b4Fas682r3Bp81jIxd0m59Y
XeEELRHvUEUaOF7jy8p1gPswY1Ngm2IWrqB+LU9c+hAj048pOtMx3NXP0tYyBjPR3OG4I2b1IVyG
d1FflWtZ890lNaMNojMWl+BdXRfgqkKvxi8nIovZYZtNzSD1XVldCveMhfGLojLC+4msA9i+WcN8
CLyy0oAoI7AfR6mwPhzkHbKHDOyuC9+dJi4ucvdnKtnGJ+9fd7ZyX7yzFnr1zpYTiYLrVrMETK8Q
/F8D7SCWHZcASNkRgvx40mVBzs1yDWQOZCSy+10T5YHJgIwILpVw43TPVzNe+U4SxjC4oxbC7+3f
Qz0dFvePt/y2GH+0gSG7FWWPjsD/9MqDgdLspiZkf3v04LLvMtqnpgwrnc80U6V4yjJEZu8w4jiu
+WrcPMXrlrNTHCYY2tkIuEh7RrbYLd2x7C4hQ+Bo2BY9iuRfliD0dWMpaX6fSCubH/dyKxKzeRVt
7rEEtHkjxmgdxpy1W4xl9q1fp8tqtvJDeKhOlhIVJa3XAvJFI5t4uBFWrBvdVb34qhmxhta78Nuq
D1H1INpJ0kbsCZ8+DbgXJ5Ix0kNek9Og/baRJFohD1vO7oUL1IMklr59rR8++vRnXcAqQY5xFM3M
jKJTAIbdMOD06HCHrmg/zEh9e5hga1afs7Iebht4NDCdYbJxXT6+5vnOEeWvE1pU+z34sRmL0Zqd
WJgBKUxRBqIrSeJx/J5ZHvgbB/uB6GY9OfrZTJZCwSD+dvixVS5CVI8JoajPRbrXUaYEd3XoC5k2
bZPNy3fEyF0b8fsv7XET1tARTc01eqG+6DfuSj65hwvBNMAOSpUWP+2KNWe0v2vaZAF2HSXj+cr1
WqGTElJqLFd/mhqovbvwz0HHoaWr6KlhT8m7C/blxk/JzY5ppMeZIy1ErVP6wpd1G//StvFvqbax
CEmyW/WyVeqaQ/BfG0J+NznRzjnOpxUiA7yd1cOkx2V+95kARGdPOqvzavMsSTjilWxCFD4fd0cW
Z/qbEv+AD8kexCBKqCmLbToi7JLjIoKrynWkizMEAzJZ1kGZiZegyZUxc1qCouMzy0X1uMcJfBBm
YYLEfi39T8xHuaEqxLKZnsapQEWZWbbk7nMbkrT0GFVq1d8LtG81f5MZMDrdYR2cJTQFvmEyfljJ
yt+3w0QZeQxaU8gG2sJr03MF63BAoCG24bnnr9o7gCiH/4ALwpVyVxswDJzrif8SFopufzcgFX99
m+pq1i0zUm9LpA0zrqJi0yzsZDrADKj/rQ2N6ThlegEPkfDfuG0UzaKCe9FvYDrOH/lF4kxQrMQ2
IkjgNzyEtY97jXtQ+meKiHuDujWbmTeAdbKRm6wWLZvv/gu/cJim2KHrRLCGzjXJ8aYRrp2i+Hwk
0gprUQ+9m2BYR+qSnyTe+rtPwMEy9noJAKJrjdLfuD75Q0nc/ugX4VmhQTufacKC5HU7eyZ8gbHE
k/MDVegZ0sB62zw9wyJHJ2AExa88YdP/lnoMq2WImPi+dl/mq7HAbfCnB+Lix3uQyIi//iu2C2gF
d6hylZz8quEtC71IR/3ZbpLVr3royAAB+HqGJnPpXvjgDie9J7I4RXEwfjb+Zlt/zAFsJzBkccZB
rTDweMkJJShrb+XLRBedJYrznvjeqG0oDErCVFddZWC9/SPaNsLn2iF2NKzd552Pw0I6gPM8A5FN
MvUIrm7epf6CkrG4fIttDzx9O1CEp1y6a3W9qVoKFyG6vhGr6FB+88/vOy71keIwG1WqxBJEEy2/
kKKo3bO597lduiV42GyxP2MpcbII9mXlDC10cG8SWCbrUS0MyQeCdW74VZk/BJWqueJBxfK/G0QK
5ochooRSORxx7sWfogWK7ZgawxjKANjfDLvaH3klebFNTeD0qGMv6vvJRf5GAbNeeomYtXw0qU4r
hYeslbkCxpaWlKohVYcSy0F8OD1OODsywUlNSVnIm/8YnUwrQBfnUOGcRbit6wATVRFaLyk1zFJf
k/yYWee7frSpBGC6UtDE6UzXutoHnD3nllTexGyXsgcQcBnuBwx0vfo+DF3bolIlU+pnTPn4QIeL
vP4YCT55M36ZvW/pTiH0rpM2/iiICc058NV5fnx2E1ygCpIT/HBjsOrRs2vLuHaZmrrB/CHSFhR/
+QylhNdZSXZ75L+BXO6o4p3q0jq5fjuCmTp+dpNUyC24ANSOOqXb9xv+v1VYmB9NlcGDlpAg3VdK
r6+bi/OMVBiWYWPlNCCS8woEgNY3I5B3dEZEeJxdL2BBHhW/rN4PwXTTTMPAigJpG8fazZJg8OBh
L4eRgL5CgjPTCS/KQfBU2R9m6Xdzrq8BGpgkQijkVVhoiFv0Xm//R0/HO2sGrs/Zn2J4qhSKxn4O
zwTtNnXoxBGjxBfKZQeY1lcuwaTYYzv+HTkiVbWcnZR+CrZ17ZdgiC2Wg7bhvZs7Y98rHm+tH+QS
YRmyera/g04pOunBxk48DUDNyVxcJbqQHzQ/ZmBSuBPD5+vzyIBIp9D7XuSb1KOFHiATAlc3dDDl
XW7kjeFklI9p4r5KINyrjKZEtCb9Psg7sjbVrmdxvXmDKk2uKVsHN6bpof/UAyJupMiJ8uzzJ76I
T2Vl0e3pIwe0rha3H385WffclCovJG0cOlf93TLeSwuzfqPf84z1yL4Y4DVTXxOvT7AnVbsswvrg
zRspTLh9rtm8N03dLrfe+tw0YTbHkPqKey6syDdrugEjZHU5FNUtnWtirc/xnnOf1vnZ3gJfiei2
rU/fxO7/nWbDr3Pj6DaDHUWg7xoUOvVC4sfekAV9Gpxs8fwDdTFMJft3DMhM3Km5eAT0QzeZtFeL
GBuEiwVMK/C6sbj5cELyRbEIHBwxuq99y9ZiLy4gV+Xh/klW3eaauYJE27NA6Qn73EOAjNwuESen
Bnt6N6O/tO+ruzTLSkYnEYiXiNfTNHJJpfqwBNB11ylhxfySSLE+uMAPRXI0YjBjUjiXmqCTrILG
WSjoBpXqGa36wu/lE2MgQtrhDwm7ey3ndlgGbfJTaOT30w1jkqi6mtzqvO6XoERGDmr79NqFa7vT
8l4L2EsxdVveYXlCaSQoFLhOfjF6OewaM3nprS8p5JPh2cbqKyat+LhZWgPVSLmvx4peRFzKgDfv
FgYz6rWCn5x583DTgs1K87aLkhOGsJ3ooVYJkbo70HAER9pTRdAUNf6xKE5FGOgj1Gv5DI1SH0dN
6kaVXV7NA5Wnl4l7Fp0hXk8P/tHjFNuXokRQnUcUanl6Sf6zcH223dnwcc8CewgiilXnBVygAdzI
1lDob5QPvcIeCwv6IuvjdnaDG8IN1Yn2j/n/tXjmEyuPTfLoezGfoFEaTgSA6u25k0Az+N0oBo3M
YnR9oyAq7joOp3oFFgl1GWzXLW8cBxh0/h20AY5Gz12ik/kKzwOaMEeIkNMeL9oh6tu8aGABIXJK
Mubc0Sje96KgFm/kU1HvFcKMUzy5W4uEEr4KumF34Wz+kl8E+XWCbN1R1L6A5bnZ/tj7IQ2hoEII
T1BcxONZH50WyhXQanRxjIuXrZ4IghwMZmIY/weNJbYtJ9/5g5BeW0rQfv9v3TRtZlpaf0U3QYmo
zQwlCgqEbtr2fx2/xFcziLRc6wex1bRskSWJA+xeDQQ9OPhQtyj/0LyWKKUl93Syw0ZfzYxUrp8D
8rcRr5kfo03TPH1jNlkSP7W8dbgyFc6DAnzAjOw3DX1no56prlp9p1P5dtD0CvfNJaGYOMeaPLqg
MvGL5tIuhbi8H5ojYMvQwa8hDqRwOseJHa96XbTbM67NCvCP4NAcg1yc739JzOecKIK3zmwhcxwK
HqGElYcTmoZp6Thq2hQNz1Z/tNOWBx/aPZjYBgl90c4+kYSUzcBnkVTHRDZfg29t7757ACZud6a2
DY3fr/SRRdi3Y2y8RRVVqZZe2mou94VqjzABSVjNrVL+eL9ZHcYxdCNR4B33rGGAr1bQ6d2IXNTk
jjG2JW5N13B3U7+JJjHEvFJyBp/IAh3gGa9Inf7HhUZY6tJUoFwRXwATlqSazB0780zpWhGdr2JK
6+vG7WKRpUek+6NyTVi6t4qFJaX42rLRm0mfMf0uSC/zxl/pS4BxkurEwvC8tBgr1daIvd+9qJ3h
XJS4BR0o1Hbyo7aaCqfzSJPr17ZVwlyOy9kQUsTagsN2ARaPk+63lfgpOgBomIGsYThi1rre6M9R
XoraQ0MQHu6XAT7ux2K9cDTtriM5qHZu+Lx+WuK5VXQkU5jmZtwuh2ZJTxLpL3aeY0OnykFUyue+
/s70fmwOwCu4CYqaK+r3IwZSoPiqFp1m9ExqBZRg85IGpAWqVNQisVT5td8M/VXWtuyfpRvXgJOI
gRs1/VNgpxCIsOIadcWS62w3rE9Hrj0MLxXw4IqpijE96ZgcpNzykHUc7Oiw6Dp6YfkQFZNrgPSZ
NKm2CbJwsGSbVlxh0ioansf89abB7KcVjBZ+/QipN9VM5pyewYhZ3wsFNnE4U4HIa/Pb/+JttBKR
SwlAMHncbZGlsaSZu1LqddOTaSjT5ShaZQOT/ObVsm7hu1qOpDj6At7NLVkrWexMVmcCFAdkxz6U
GLLyOpvxuV3MWvdgycDmLerUTNxGBYpzOiU0mCiYdRcLeFDHlOw36vCZL54JJc70770DSkWEEUHV
bBk/A+phH9qr9PNpnIiBSREEsn14YM3iMtnENnHbMOGKsKEvPwijsbVSznq2xcVBdYojtnDVYHmY
fjt1YTm3Y9UyVTpdPz/gDb2YXBsPEiBdmOObebKCZ/+l6iNC46mEm72NmNFtV7jrIJkIvBQOaswE
ecBH9jlvRh3CFXElMy31rGrVFbW8VMJK3YCk5A+eHq+ielLHnCdopUyLsZ1oExv/OcP3+ZUiKZMD
iggLYZ/ced7t2GBtDekRXYZF5/4/aVYeo8IkVR714+Odyik4HISxl9lebZABu1MbqI/16RUvY/lp
B3kKy4XPvg9TNpMNvFA1WEmSf+RiBgPhoB9O2kSRcFabwdAMQsPKrgZkxv3KrvDEzqU4rkjole0J
RX20SS/xNi0ZUH/Rikb6iPJfjANxIZR9DSckAbAOlyUJvJE9ZAAu3YKItAxxZQLvHmfEWSdcei6w
AVzWxwVsUAfeikjj7Ehz7T4BB9SMUMpRHtD39Jv8YSgUuprALR3t+NBFbBfpx471JSaGtjat0xif
YIodzCQ+dUm7NSLbEh+FeKCj3zOY5cahVI0amsMLk7Pvd9YwGuqMdHYSIhvOPfUOInI2Vc/WWyxg
vc3q79QOhkNCFanvwSxTRyRixEiUqGRGFwXAXdVREQZCWorChAWTQjtRWkKi43rYKl0wSAYo3scv
G7NT7wpMTy4fibJKWzqEhtgZHHJH/YTsKdOEDVE9UpJWdRV/QrrcDDlEry1PRJ32P+BNxlGwBOn+
Dgi5+y8Bt5wtsV+Q2YdnIkkTcEY1k3XyiYbSDp1UqY3xLXCDLrOcPKJEdyYvs8CKEc2CHCm8vLkN
ageK1ur9PUL847hGijiTKrOsQoDT/REsQYmg9ODErSqU2FOIg3vZyvjCNdhisC1olHY3OgPJn9zL
dY8RdgwDhiKCUTZFmXltMXaDhBQ8QLQxx2Jl9EMoBLunDTA/4XoiIaQWEmcOo39gZL1a8PTslEyR
ILWziuAQPN4CTfJaVk+KFGf8ZS2658PQN78darfSl9BwP6cGwtTfUixzxxsGDQLfICACWm/+Eka1
D6n0nO9+soGSK1OtheRYCfrHur0Mscr5CZ3ckzKlnJ6SkHY0Z48W/IMpRORSs6MhQMeOk/nrj+Ll
4aBr1pKQb17wBHnvmHZrjtl/2GYTk8ywrrqza2SMiLDt8zafOzkjKAUEB1zC2ZrOBSGOh6VtfC+X
FOlQLfPKagMQs8x5nbXhh7JPNF58hvOLltEyq4n/SBpbxiOUNsTPes31kk5h/Ng5TGcAaRsqGSvv
mNQnB6xcgLFi/og8QsOP2rPqjZDzt8OwqrEFwJ+2Ctsq0CGs8HtPE00JyrugltpQS2NnVSZawM6S
DJdpqTKbwiEB9v8qDebebHaqZ/p7KR4GnwsjUOPYAAdvHE81dL3nIWwFhCPiNx0eFidt9/PXBf9b
uy6C4faLZQnrCJJRftB/lFsNCPVP2XCkAO+WIMvnNSbud+QYvePV1KmrmKB+s+gmsoLxaaeJtre5
BTBkQSS2ttk+4hNe6AGu4sOwMMuG+kIRpSSU+E/rESzjXBZSbO9eiPJ5BlHEx9VJtD7z8Aaant/a
+08ihY/6jrqJG32dUPCbr8HmQG8AVXwrkqkrm+3ZJf4A3MbP3GKgxYby9Li+J86NfZ+Dw/DWPQ8J
QI6MAQA4odky9S0XMhWNmw1EfRnXPOwkxtsbTLwzLWgnKGIifmi4jbVOCPfc2KzRPc4mr7PaNQMK
dwpkuyBa/bZRksiU/1SqFgqnsMmjxgxrThkkS+S+b51NuBAAG9cuI05k2fS/411mXRyxPjXknVV+
IkrVArkXVsU9r3pktahIGcC+B9vKxPWVg9FHvXLQ2Gq/ed+p1ztI7CHsoEAuK8/ivd+3fun7s9AD
z/3F7+/D1R++W0v3lOjYcsd2KoSBM5bUvlg2vqksZxcZVriIEDGxf8agGyvhEIBnCvS4MRHE+fY1
UggFkqwKnAYl76Glo9hoLb8FyZ7a+satsnX4YzRBq2FCZOkh6sqa+j631vAph7A5hKRJGsS6pWuT
zDwZD6WigHHcJUkyFGBLu/fbE2uccwLKoMCRuqUO4G+iMpfQ2PF5uSBFpdR+fBo0RL+3vh3JUX5p
MZBluBSJNPGnSJiPh919pelWrzKWWU3267OkMQnzs+CFwnz9IshOIKlgiGy5Rlvy61P4DtCh9mto
pK7om7WK8batOgjMdaaQhXl+FGxt85iuSjBLO1iByME1HIzENWp7sjJ8pn54UP9Ox6r3FmkKN5zT
Sw8iaSA8CFg8w2jpp79mOHc5X2MkSGxI3Jepb8czHKDEh0dtfVNfNpcwey0Cx2T+qMzf0WnR2kQm
YGsoUzgHHZ/lgcrZZ2238MgjNy907B/kTXhCyXXpN8K8MFvJyXZ9eX9fjlUqUiUhMhK+fPzYaSz0
djjVn+Mha+dBIkgg6Trxx8IyH6JO5+8751zjTtUktzfOu/yf78hqQyZ3DAhqmgEg0D1IMsclDkVr
MrWe03kRE564xAxr5JisZQ4eNfz2td5Z3jDM0Sjf0QBwpJvDu2PXqTykKBPOiGbQF3Xm/09L8V4D
FqyX4KIx9r4Sebkn6c8L6pyf1YOm93JWYDo95Wwz+vCyW4pLTUG48CwwgDgQ+OzKziLxQ7yZNp0L
mkZxnF9MtZYQXvxjEbCByI927u4Wrh1hqgvbMFuDe2yxLPPAvMSumn72JgQKT5VDV4KAfc0BfoBW
JU8htHvedvTrCPzTd51nxxYWEogn2DzqZiVVAOjFeQ3E2RqPI+iggCNeHrEu/IQI4h2C/QNu2TO/
+5D2aI8EkYqFvqbP6Y937ghMvD+U7+6ka3Ni0y4jr+cxgJDdb79FvwH/KnMCNV0NHqwhj3dF0uKU
Cnvk4ns6StqFVdxFQa3se+7tJ9CTrRhBjwTU55tJ2GMJPLFh0o+IHUPMQPib2btb0Vmvw0L34pGX
tEBlDYOAqrM453XPWkseuheYta7lhkla5n7zt6VOx9i9mMcXaZJECliTF5kLrxwdm79/uBp6tLGK
IJMCFt8ifadkT4ByUQO65wQMrOwWTuubySfhSQgcVjciSXNOb7IWGQOhwV+b6Nph22qamxupTQY/
NUo1ClEtNbNfz+iOlLlZlPPW/UQNr9VV0vb9yJGIdupjGeQTqspLfEpM09iJhrBIsm3HdqSdYQcl
M3FRn2EFe26BSCjoJMaYPHEFHLFRDAU5bDop0hA6HOa/RvBir7ZKiIvlA7jWXt8btEswo/2Xx1pc
HnTK3rV6VcL+cwCcInb9BW3ZK3xFRgkj3xIMKbZAVox23zsXjzyTdimKT6iWdvuAYmTEoiKjoMQK
iJ+nx+w+HOtBtdGJtrKN+dW58jWOyqYl1+UX1MhTHay4ZTq8TnnQjw6hG+LqMzDVWs0FIibNSOes
umDna9IQxzEaMe1aZ11forfPV6Z6R10ea6do8Rnjtu6yKnddN3MYMTEocI0dAb3ZEOu2ETIz7Ymj
3OpqkEdfYb4vcZP/UGr6G/1vKAFGY2jU1im12W+mCpZCoW9B244/jq7tM9fBJRq4ywo1mRdLLAsI
0wHGwuzOcmgHY3rWUpCBr0vq50NK6GkHO+p7W+Kh+QQcA/h1m/BrJKQksBSexuOoEFUpsXNX1kPk
RBQTZBkeOJfx1JVTK+FjL7YArCkFjA7vE/6aQLV9kPtbKMlIq5dTZenA7apW/CkbI8Di1YrVJFze
tvdx4Od5eK8ecZc23kat8GDguvUxx+J8yo5XNbIc1cWfkzRKC+Q/BhAjHECFachQvPJf0JLyqAvn
b3qIG4+2oHFv46NM8BXjLhsmOXXP1Tf5kuD/tUewdqPlJ/5+gHfxE30cShhaLtmDX01KiQgzPgYv
cRosPHaTMFKCuZVX2J40q5oamOgT88TWnKe6XaAHR+bYOx+iLskiuYNbm59tp+ZlUg4hZBiNF2Zs
TYqMcpOX6QzfG3zkCSVVUfX99TIL4vKSi/x+IAMbm6GARQz7fe396eFzjffFrxgQoL91PWJEcd6F
2EZxt+LK7eOUj95EgcUM/GGrWbXH2ooeWAH+s7Cr8rzJjRKxvIL2NpiKRhk0DAEntn0K5soZWbA0
gZ53tTasK697FGsSdTwJxGiVWcDfkV7KVWwPwIgiq06O5Ug5mvEyG3Yw7nbV19DXUmkyv5btu7Mo
NiYjMQwOjad46FVo/kWPY+Rbcz9AGBlgoFzf50M88LjA6faqbapHAdFUBJA3JPMp1JB3hlLOFjmE
oZm8ogoheHWQvNFa5Hlr3aayZW2S6C49X1UnKN96zrQGgIQPpv/uysCEEsSYylhzCiFreGdwLE/x
zKiSSmvGW34pc6ylLqkCiMV+DN82iwQ0mwdcnlUa4YJ7bGus/RTm21EWeA6khvt7XHcIHTfeepve
5jX6swTw1xBeEXLC5avsRwT6KT8PaGZujTQsKViHSGRDpEnY6ZKnNEpCsjBkkPk1pi1FzOVMtZyi
RiZneRFv1LwLjswmcYa02WAVAwDKLwMgfioWiqsLtJVYJ/PwENoeArir6eZ9jChOFUnwz1pU3GJX
xiUbAS1Ci1Cs+/AOH0f+cvk0kTuIJVB3HO5xsPFgWX/xTpD8hVbmOArlqodt9U/2RXZU6ENVe+en
jImvSd0RM0raJ+vxDACSuJESSbo1L5ZzU7lER6KYofBDrmD9S4UnuodwV5rnvqegJE4pe4CRZ1H5
V80+dega/zWshvpXKsKDAEPcb6/4sbATduV2fdDm6Ye1MOL75znYqcOO9E1U0dZOG8kSxLFfIK65
EQpNG8jiOT7VndlyrcoX8e+ur7MlzqDmARaL6+Y0X8n+QstJ593UFgBV1LlGbKvJAna9MaLPaFHt
oW1uFRN58Y9o/7BAQf4s/La4zQj8xuBdQyfDuOKOUYLXJil12XVRSDq+UEQ4cjWAvFb8GOYvsNys
QJTMlHb8hJpfg9RVEFlo7m+VkGBjA4yg9okagPuNpVeXAwB+J8ySxUH/7nWrIxdWY3RciX/V7St0
0bQdsl/Za04C+P/4esLUQhn6NXr6cMOIhl8zbD6upnxhxqZN0UueyZd6NlhxW+ptoMY3vplu/NWq
YqBdaf3hVA0GS/qLYFqp2aRt/9bJaPYXSyisPfBgqn8SSRqN15q/Z9mD+FTzz+3zbjU/7A8R3NTO
xtD+NGn5Q6xTTbgqxQutAepnhl7vQzxREr1Wsp47zyj9YtfabGNvicndjwTaf7zJbkj6jgEExGJT
KTYEPGKCRFnc8AUEm3ykJftJm4kPrCpn7kL65o2m53+QN0EdbzUsVVKmkGLNINxo3D1paRnt1+fs
pSM4CxpXU0S4RziBoEXJlGGyBD/XEBeSJtLXQutyaUwZiGYkMNkpIwl9g2oC9TWCf1GUYxe3v9dQ
kfiDD9OU61gL2vh+OjE+U7WvKrGYIystXLAw7pxpQDSuv3u8DKJL/Vuryv8ayZzO363HpDyoL8ej
DE/9XUm2/D8Uzn2lDlItqjJCqReARMsTzqB6i3ZSY/RbBZEnuklLpB8UVU0hXadJTTGy2DsnNMdA
gY7rNvGCroVRYOK8O3HC8Qrt6A1tRHUfaoiNYDwVCPdgDeQ8YV62dBgwhCFVHEEqjUw4jn3Jk9D4
RKeMqMHGmnD04rl7xbxt2T6g+o+ltvTC5ZUnCGIM+WYsB9HYwfZSySBm/ANss6Iz2s1alkb1Li0j
pyIUUyrKG4JuVRkpPxRMYABi1CeOqgYa5c0LX7rfv/Hp6n5GhKsDw20LsmTvCTwnHwlcJVo7hhfd
MLsMElKg6xrYHtSIG7/FtiNpYeUerOXAKOgUQx2UCOSqvc+jaQotBg7PKtfFyIWx5mu/WiVs0sz6
lmZGxHfOxLVyILYPAxWLBGiyXWY2cxO3z0FGWrH2Q906A/F/JKyE+hvqKw3VtTdtAf2gyWBe4Lp6
cI81OF/EWjwrQ8oj+HflQymCi5emQFxXJG/5/BD+0JJzJG7EjiaHT0FeQqMoT7i+HLF+5SDpCTyt
EqaxoY1pvdumHpPBsyPWQb98Be1c9nae7+WYETU0U7I6p1PjnlFme1/vBjCNvxSzk06DMUJsg4JH
ITY9+r1u9kJ66HL4+b/0eIJ33mr1u3c8coDH+etp0uTjHt4g/jYPBBUjQZvawKPDLBojZzia1FW/
Vs61KGVtcnzc33trL22LcortR6pfpFNuZUEq+KBOwlC4adYViVdeHGUaWZwCjJyNYoNydglbobmH
JjWdXIk5+3Re/aznaW9qb1H5vI/fA94yc2nfc7qzT7dh1scZxwVKMD/ht5RXVghtats0hkNnsQZ1
xYwxQ86+mLaVkdwNVwTpCIb5j2OExGZsKU7SV4KxF+0TOzJ7uT0V/PZp6s7T8F5qGOHn/K6hzuXm
BKOE90iG6XjsytwV+Zm1f9FIjOq/GsNq6QTNO7q+nLWcgjU8RISiqQjl41Q2hslTfhEoDxDvOd8W
PAgx5pAPhANGLqXYBS7QR4Fd5nGl2ryZsL+OfW5Fnxh+CuEoJZ5U/p6LyQZCGmysSgXBPipFzSJS
Sgx99O4D1w5mkz2ePP3CWSTZXBaD06Chnr+G3lZA0g+5VZKiN97ZQsWfNjkyq9jmMBnj5XvkoaX2
iV9x6jnXN8/RCLgd2/yVaTgYwhLysy/UL1U8hIdi4KMWdPeFSHCZJvO1qtQ94nOYyTJEHe6BQX2v
HzY+dijpYLVss7YTU3YWj05SdAY8BrtoE8yhDqOSE2xvAHLGwGTYMd3vhB/v60coaKZ//j2KJC6P
ZqwcFkE1o9D8Zt/7N0c5SpRYsAOIerp1KdzIhrtR4frafkmYVY+1yyr5Co5EOJlPJCC+/DV0hIEH
sOFog/9/FBu++b2M1+NkuhntnAgVLEyRJpsAQT+QYH79QZdlOtQi6Twzww195imx7Oj8CLsREh/o
0HkuNr6yFeED1R36C7LFVkRcSL9AYMVWiQm1T25K4ETEmkp1dMv0Ipu5lMv/gs9ALWBPl0QylDJl
Kb/Ls9q0GnZwpVTwKQIXQWx9nfyxUQdhzrEbxi71Dg1EP+iclOPX4bABBXf2N1BF4pDWKqLXTqlN
zVXjujq+5Ws+euw8md6Uz6gRKlNz4yjlko/WMMIX04SR3tXePsLn8iYQqOvOXqyQ2vc9dPyjDHOQ
kLzV84DHh2DNu7yNQo/6Un7jIuaQxDYQ872mkLssQk6w2NMdWPrh3v2QRLJnbPiMttEii13pP5w4
7844TpIk4TmUdwMF9JGnHsrBdUkAS85DrHZf0dvL6VMlozSch7gwqSNX9UdH/bnKCeHrEJYK+2Xn
Qoo1gnRfHi0EyGj5KR7vz9fLpP7PTtgyHB5XCiCe+IBHq0Ib8vZGPxNsZVR21V5GHy1VaoETD/tC
AYUEy6WXSXvUhQ0U0rgRfxMQGoqKOY3Swh3brsBhMSH8ZeJ2tANGEjYJRqfQXReEVodNgt0+UpWz
3eAnqjWqRHB4PQuIrUH5r/F39u0hKx1te8i++9A33hY3Xr0uSVlayTFnETaGLDhFI1KixSR9O/ri
v1HXncOpaZaIRTqFFKx1ZjrDEeXgcTj7yeH/+W/bixTQnpl5vM/PUSTRXYcVHDv1A5kA6ZDpJ0V1
LVaC0gIMZHUg1At4f/tujalmZgP8vPIHMMN1jna6ETSQD4KB3nZTv/5e1hwU72P/qaLCe/iiGs1x
jw70W9du/cYsjpRAyy82HqSsKxfU4xsKvNncDLtbWb1YtcTFJKntUne/ao+x5EpYoQn512C/1Ies
uz5ihB0RR6i48P83CEhJxV/HcEmePDwwp4DCIJgXuNLCtHzNCmL+6thBsQZDPalgAxHdoIScUe+K
5dTO4W8XacA4m3P2UFguzDt8hUpDaYWUYFfLKczE3iH88odoiBh2HKkjQ6fP2OwxSkg+xjUN9kjg
jtvnZEVIRqhs+T8We43JdgXHFJWDXTzcZTRgAy3aF3kqIPdHlqpB9CV8n8j2HU67X6tc0oV3O0fA
1nkSnP3Ap9940oXbA62PVtuDUkcLj+UW6U47/E79du1ImrHq3LPoAIzZWJ6OYSo2Se/NfVAtq1o/
pp3JBTQ7iXb6PPx+nnGFW0LDCHohFakVfeCf44WJm/E4GaCCfvzwrM3Cfydk1BxXm8ewMsAeYcnr
bjdvpxE/84HDANckc8rywgnvd04CW39Q7BHYsmSLsd8Mvb91J7ZLPqqDQqxsJkwDmRzb2UUCGCmY
i9p99moSTHglDsp72Px8xM19NjHjiqS6YbxsjHYNCMEU+ykVOZlz78AQmbPCMq/jGuf379PlYhGa
U3oMviUPtH0qZKGhJr8QYf2CRsT7O/G6ziZKxTvOKhbqETbzUS/rjQ04U6I4odCGUZcQwpCMjpI9
dwALFEu/EwpiY8+1+hAEcu2eyVzts3A3zR7gjmW2oLrNp3tnBMLkmyj5WvgKGuLPDC1vMCDP+xle
JDvhaVIzcPYv2nXbKMvG1RjZ/3A/qmTgY0IS+ozjCyzb86I6jb2x6AXyhr6goGXmrMyql0fyhxkn
LSXHKUpGpvtbm1T/yERMop0ouW1No0+rE56HdQoYauRsRIeNMlRzOhqqe3aZ4p+ZVX54U8YkngON
pVxfkmY3ea5EUKKQmJ8d/tRHCD/9KvJpsaUjofntBnVlemuVU7q0oBj2G0hcXZ/sHg+0Gy7Phm1Q
gvGNBRz1S8kSm2MTVmMpot4JlMfXwdgA9qz8Mv0xJcV1OOEkvn1kpVARjGZLDFf0WA2rONTWiJ4z
F4xOZRsg+o7xKhSd5WBq+knSpLVD9XcAy3wNHxXqzhWmIKRTKkHeKEZGq8h9UpJSVDf5Pgrq147H
lHq0iYRdgAoMSftCmOApXbu2pfXB03ceaCDKnvTNNBfXfAISXHFjjOxOzsk/UxKcAo19TuEA3BFP
RwwXabtiJZYIsrkQv//cQ2uZg8e4KbP+tEBDJUR2pDQPZHCOcduKpBGrtTa02p31KpYc0pVTaTj7
w5p1tj5T88qMsyIDPCbQDUUNrFFKwHtExPj1DKmCfoednQeu7HHMWio0CC6uXh44D6VxJrf8iA++
Fhs8+6j5TsbMFXMyxEpgP/tVN0R40gq37Ly+HOVTCGaQQ8wqoaZEjT8QmyjBWZvsAaoGCPdJdHun
mXhdbeWeRZBUTHkEmu/rxoezPI+6INb64EerOwZ1ScLs79ATG4qTUJz944A2EuxAHbxYjokI9yH2
QR5lI1AyZrZKgCp67xopIFjCsbWBZiYg4hfueUTYnSJrQNPeK4mwT1WDfNsttNWvLxvBiC7IMxa0
N+4tqtdFzl+OdSFFywwrjuBTecEtFYfK3Nd1kOAZfPXD3MWcPBQP5QG0r6lYql04FAN0Obr3gnFC
U1yxfpiznP1FfFEQv3mvcdmd4oRDnAgiqkidF2iVp8LOovdFQOa/24e1rgkUVrHRVVZw20NUcQWk
guBVmTnFa7AeYINNTafx8IM4bY80j4Ibgomq05nA3+GmLCKC7aYm0oosWKdX9NVDh0YAJFRQS9SF
O+k8DmTtChJq7ZUHCYCZAUKWC+6RwpJ3l4u+Pd5JFhiFV1UsglDKaQrPXaclyj2uvIhvgZeQLMno
XlrDpzeKPwJ7w6eOKxKocZ346wid9BtRUTocupX9fdPTGSgA+PrLWcO5n38VfwWYvqUs5yqLWXS3
gtqBTU+SXVnSCHtLblUV+54IhylY/VfUW5GXEPLw0ncBBX8O2JFsyEs5idfDeM+xX6AzD71oVBFB
6yQLu7fxnbw0RyPza+0ZnIDvSZR+RbjKiuSFpidHTHW+zDwFQbyhx84yMCkGKL/h2QrYhhGqYwXu
3pVZ05LSHZXvJ04nYnwi+mcloZ9ifq9uzA0xX2yNedp4LCzxiQsBe6pPSmr2j1WB6c9GsCM9Hkow
SqLj9c+yGSKE7s4HUKkK+Q89sj3XuN3z1aSpXuIVwk3/FpyylrjAfYifIseaPFYWd5ESW6/7US0w
Mz1aizGTsGaIkdtwZITjQJfCTb80uDWBwT6xb+7vjY8SDPWi9r28rngBYXCqOu5oaQljadNEtkTg
9ny6dTZvRxGiEkFcRtU20WAZLTVP5dVgp+GpsM04loVEGhRq09+NQ17uMYoWL+oyCFcF6/gEFKp8
md6AUWS6meCABeH3W7rC7H49mISJqtzAeMcUoqZFlm9Za91KjrYfRESLa9667VoC0cp2LPpaZybD
mF6cnKazXmKwGhFPBs/YB8VuIirwyMewCtj6zDoyAnbhQxa+w2+nKAjVf6iKfTngh5nvnFxKrlOB
djTpS7tRYMn8qAWU2LHR7oVI/mFsMKPhTsMWss43yaedOST/Gt0AxVrM3HmkxnOIjXu3Sl/fqAYZ
Nrs2sC27H06yNzWNj6Y0bgJ01D1L/0CZl4OvX21DRWJY1E6gNezJVAE8ZTCoKCqn7kI8WF+Pw00d
4/ew1BSzptjdBhN3m97kTmYdyv8rhZYnTLTn3umamXqAxO78LUobVzuaBkhz4uEI8HDSGlmzyG0B
zmp9tjOGZotQfAQmlN/jpr7xdDcck8M5IZKvTbW+N7VEBbzmSrM21slxnguiaT72LjxWetYzI+m/
wPl6E/O0LMJ2ficoZSRRcz4JNnqteNDJ6BbPBfgsDhgFN8xfU/B/IeEr3QPNwSAwJ0wLMSrXB6In
OOYKB0idrwbF+NKG/CawfpkbxwH8JTp/Umnq/IT61x/YByeHaQ9hnK0cZ2wQ0rz9R6botOU+dq0M
Fj3WgpZdULA8EREpANOGSDhWeBK/uUKyFc8H3fYRvzEdhj8kMOlyu6q39LFr9PDs9TdzPlrY63/N
G1ihHNXc4dkbaeywmKpLzvyx0g0BS94C3lQN7lPIMBrw+FJ1KAFh77BidnKLYBHqu6onSN92dHj/
rZDAwlvY3qwcTXAfAKwlBru/oUAJK0HlB05EJZiYaIRY1nu4hcDRngIFGc/lq3zLCwiaYbjypjz3
EAdnfKLpLt3Xji5GUloCIHUkl0aXGr2SHRICqFeio90UHQOq1iQMTWpm3jhwYZZPHwITkru1JV1R
hH2JT4c0fljktKNHrGG1RWY/MXMHhdg3jzMbAn4gWdjma5X9iJ/ZX3eEHKJfb7prRfsolESbLdjc
Opyu4enH93b4yCCDh7/RI/N6uxeXC1zbwuaW17iqZpq3vKJhU36Bxrqh9jA8bkPcX0WGTjkQGh7j
zJPvHbsgp/iTEOYBB1LWLQKCxleeLDdgfFpjO7WbQqz73CK1tJS3IykV8rLVBcaiNBKAs1zdG15G
H+OYMvyV5qLGOD6Lg2H9FamujhoXgBlbjrOnglXtzwnFNwQnZD+MLZuG6lnu8hBoyqSEGeeHR2/x
Wl5C8POR43TCrwVPnRJY9wyoV/zrv8WJd0atC/T67kwvIk4wrmHxiNnZzLRWf/sPJHnJH5Ue5NhU
r3UcS8cRl9zBiqz0Br39yYjWk5zUL8JvIPto4lU2n04Zu3tx3UDpWgRwEmkjTWbBOWPPcpxn74sJ
i1rg+95Yus3dPEwktTpQy3Ub43ONCvfN5Qjd8X4PdTqhA5wPjf6bKabMjSarUdh7gUmhn46+S/Ra
7WBwgf8XgD1v/pXLa9f5ubxeOg3C4i3diQ/B+DTbtLXXabMUkzJhLPFJ+dgy3iXhrmFJhU8hXB/7
f4u0B5df/07X0b8o0FIKEyy/t3QSLHwStxonSQX2qGy3C5mK6Ks5Mc8mM/8NmPFs1dJNw8vwMG3p
+z1hFlXNJABad5UJcMu9vVCD1SMZ4XWu5eStAYPhyM3eN/qEup7lmAFZQ/qcf4w9//kiqxU+qeWY
6vuiX8iW5tZCxVWD8DZSlFKUO1mL57KivFKmbP4yzj7XJ3dZf67ED/2CaXPK/4ce940UpclR5ZID
hY5dHc8Z4l9Vji3hbOOfGewDXo7YigKxtpgBkPXFkY/YH9CT+ds17nMxuHaNneW9PqvlG0hxSUaw
zFFvhDcGgXZaTNIz2QVY+BzBcDaLBWQwHrSXxhVAiRTO/m0NJf+uT3rgD5RX4CeGHu2E78jdcxob
Q44NSdSOK4p9EQi7GwpC94RBDjlyMqnHxMffNOe2ceWpnJh3mk7Lk/v9oJa7Xf7g3iWnVsvtfq5p
Qc70zzutJTxt6m72GAib5ooigIdffw4SmCeqF4qkrzSuj2vP5laCjrL1kwtq/B+HEUVx7kPfuRG8
RuoXnhBB/eKDngH8amjpyiDSnx5AeGOwHZ9kKW9Hxj4u1tQQiNBhMs9jctH7TgDEv3Df5S8nvJBe
EDQDgNyCz0sSL/UgoBaiu5URHCHLdwlBZxgvks6AegZ9wDkIOm/+cd+Ojo4OrkxWfM2X7BNShTV5
VThVS/ssjKPbrj/7dJjS8JIRWtMwWOSFVOPOfTq3yx87vkFZQ9xPk+parsW065QLLMwb48qXr3/l
HV1NQ9OLOsS5mFv4APeO6m2klbmk1/+790Uxq2Yh6iuxGa9mPVo9bIH99rb9iH973ceHneWvbzFd
ddqnWZUf07n9ROOGakNpj6hcKUNQFyY3nHVR+HoRc+k0i6IfeOUeHjkJjdwTaY23rnUOegoLnx67
TA/HGnVEvhbzjXBRbCbS3g3WkxcwZq76xjqV2i4FC4sPD8cXK9uyV1QCJA/xg3W09rNvSe2iE0CO
fQth4/rf7Hnwn/tel7hMtibFEmbSpL5VnVhzDkfR1sWphYGMBSpW0W5jDGZQ6jWAO40cRttjqOIC
GaIeWl1N+uVI0TzYRoQHBMEnV04COmN9cPz5erxPbhBgKqoryXlKBBytEbVPO/Ab5nXvh+dkUBRl
t8EqY938/HHFi4x+QP48Vw+Dse05hSs8exEYbFj53O15E+B+xKoewW59XE30lRy1hNs5RcJwBkTO
VmBBJbD8SV9p4wwmB3GiL910AF2+8R+M5xJUO/pWoxpIRo5FhzQH7PiaNyyC2hQWSAC0WOiK0fei
1+VN9Tf1z+M0L1hJMwN78r/RRzzs6c1OnlHT1liry+x5lbjOjwgdNh5Umz4ldTQ/3zBh47NWIDv0
f9WA89b25lDgr4LEaf19X2EPNRXfMu3kiYJedJqBB113k6GddaHtT01Lk5ZfyG6FYDIu7DlOq76Q
mZwm+cscuVo5Auhem5M837Ody0hDiMh/K6abe/bq6lMeN4UYm8ERKryVhSeaxVcDZfBOc0kC0O7B
VLxoV8iJqCB5daEWjqR2uKaYbtxV2yO+QlsA1r6UosbyfS9WRPN23SoFrBaG408fWD7kXCRjObu2
jgl7jo9PJWYIaWV+TyL5YLtELi0kNdpSF+RsSSrefPuRELQlotXlj7U0uzIoW7b8OkiqomgY4Tkj
vLevuwDGKyb1Jksf3ukFMwztcQkxwA3J4ZxIerMtL9ANr6sbSR1xLGXtN+z/esyjAas8SeZr01Ap
2vqTWt3Jid3R96dJwcO8ywf9QgD3Aw+IE0F0W0hT/VG53uAgSZW8gkMGd+73+GmEL3IWeP3W2lBi
KW7UA/KyToGt63Hg1/cQpSYMppHTjqaQUtR5CM75utT2vLQ1nOUCu4uYnRQOUvA7lyAKf2bvghsl
mXa8RJTkY6zdHEm+pyVHAY424BC23QTkpWkCG24AlAXrweR3ovayZk2hS8lR9OaejMFuNZF53WoS
YnGZNxZmJ24yzkY9D53SC/sloQFpVUqOQAZefZ8qHhUCv4W2h8CX+CfLIeg3E8olJor4f84+aD25
/Mk3KkOmBHxH2bYwVO4jp8EXFsMoPT0J/NmZ6w9oLfXQZSgqc1vhw+/yjaRSf/W8BFaHtr7Ifbwr
xd0NMq5k20lcxntv9qXSMey8W05Y4RO4kYNDmXpfWkXoO1Mmt5LkabTjxETzbMZcuSPJOt0EpiRZ
dOiu+uahxl7YKSkN65QfgW244gmjDeOA08fybsVnD89jy5j5rDqYhOvXzB8pM2LqIA2u3XnzZpMP
CrMnZdNoL44x5SL0kwZid3BkqLT+WAYR4pygdTwW9fN+QZXg0wRwdsffF90WFjeU3N6zba3ldomN
1bOIK/6HZ1ZF1eaexYCmV6JNSXN3CmIkfPCkzhqbDKlJwmPKER1lsAFDGsI++o70x7juLkX8V1ZJ
iwwbaPy7PPQYBbX60zLVT4iFlam/j/oDbQ2w19C1CLH4V2QZ9hhw1zYvpOpRl/uOFn/OxVkhrfmB
H4SQK4Fd0zHAXU5G6dyQ50hORdOsiTaQW3TrD3bznlbUaHDOxTAvr4RNdMX1A3AaAJHi8SpSoLpK
iiiMJIu9ohSkXc197sFVYuFze1B103wQXPhpuNreuw4xkeDoGMaGSL+KePjCSDEBQzhNjQpABsSJ
P27n0mkV9x0G4V2rpARmK/Df2zlVNMDzSqCIr0sbtEups16jDDM1vcSF1xy4WdZOsW6Hf/C3leT4
LXlE4KvxUdOPyQ17dz/6bVUD9RS4uGjrmpVZUvSf3hbV3K2QduR7fvf3uDtQul6jQefj+++Ajm71
fK6jHVBiyTV1zpGBqac0VZhqz9dh6dyHIvkEU9MNeFJ5xBWtH4OZkEpVZcmgaYkUoBxkfUbcs0yR
XKkBbQrkY+47lSgOwb+jgOc69dUqAanrG1X4zDIndNQB8jUktcyv4wo46Jw8ubFyR7oy+lBeMkX0
izw5sw/DfdTC9wOx3EKVvrfy0NzpHWCAhfaIAF9PTFek/mV2X+r5cOF9DAQbk5ZekSxAv0ANSWZH
cf9m9+5o6ykTQfjHwXwBLxQLiXrdfv/VkyukLgvcReJlnuZdGhZOrX4erv05RuxF8eXOZnqCuKxm
NBZQlg5ieDGC50PoZLl6CakgAKqQGZNlJngyRGHFSyBfYUBe4bRa7bKgdpT3zXK1g/nMfKYJdmPt
vB9NpJ3faLuSx9zmkAcYfkDilqftSMvLzmGpuCY3JgbGMQbPKQ65d988v9lceYN4PkHeZoQ+b667
BdQh0BsCLNUC80cH0/H8MltAujOZjhV3CUgjwXkT55ztArzmUTFWbG9goc/azRAZnJXHf3JDrcEu
PjoQI2RW1SI/pTQudKZ/z/quC9ZoIAlvyfGZO6qdhaQlkFAT35I8tenU+kq8EWm/tC4D54dmMxxs
jzjdyKkQ5nM/Y7h2s+b0w4/p0etKxbHYhloQvM6I1Fahfds53abd1upWUpqN9a83gHaLPyNr28wY
NcJ/nb6wkYUiqompBnXXldKD7w5iMpVY5ACd7EfbBdwkw1snGJ+lP0wuO1AukL9s+6gc4UGPh8A3
j+mMbQW/klE6mk6kG8D45Z+ulHed1fTmGY7qwRSyHrjnhmufo5UtiNOSNTfaZzzOjhgOlhE2WdRY
6KA9nM5it60N+DbgPbK3UHHpIQhYnW0h23IfASseRM8ajQRvemO8DXuRPLKzTdxf0hSqHx+ombhM
cPTJ18dDzHECraQSj/cNAnGsl/WhR0eWdt5TL9MOfjBveFmjRH+TzzAohE2yoQMy0Fdj4H6MF6Fp
y4F0/4g/cokMhKDFiRhG7Px6T90wQKzeYNqlND6eqjMJV0pZCGv4x1KI0rz+8jFpgZLytijgwg+c
m3L4rpUvQgssa/UIk2jT6k8q45Zj6fXX9AnTxLKKiYaKxo88m6rcpp2V+AUXp6H1afO5w1rql5qd
FklzPY6EbhRe7fFTTIJaxAVYFqKi8tTcwLCdj/HRWGdQqMq0qqVsVUlynoRG9dZITfDSo/4xvzM9
RwU8vLoyMd+1fBGzoCT9nyGEw5npu+UO6rVrqNxHO6hQjtc/JHGIV72cB1f6mgaiges7rOE/8GKR
O2ZpgmmY4//aDfH/6JZbTwKsmqpDn7B9dfYz9Iic+elhOM9jRtjdVbBjSIblVNzV7x2xFk4KlO1d
+NR/V25Kn8PBamRrFdGjgEheVWyPcE3tg4+yetsA/T7xKenIKQXYxWB2UBm9JQa0Lnre1GSh6igc
aOtCEWALvZJQbxMb/QUaLcNIjG0ptBrbzYHvpLZqdLws43akI82v4D7XiuOZwhiAudpvf+1PVz9M
nHKdc3OdmT/hpwGR60Iq+dUegFh7aNyDjvDQI4vWSTmtfRSLbVIVaq5XG2W56xpMe7sI4PJhmk8C
7YvtLFx/Yh4gJNBnrSAMaDoJHqRjB7yrnDzNXnZqKMvXZY+nFqzxZ/GdRICo4WBXr/M33Pv7BeXK
4NYqoZy+xmIamqQp/GL0o8MFp/97dap5Nk6kPH8PS9Cqzu3FWgPhq1+BOxZ+IB/zWwtC9oAjfZo8
zYjfg81i70GoqhnuplyAQzG8n4DHm5AmBYOxb8Q26stYq2+hpsXcGHcrUnndP/YV19BaFDPo/jNP
8tW7tJCqfGkujHCr3a9tytW1TdsRPby7DeCMdJRM0B9mUjePK8tdL6Qgm6s0OrVe0W0fIorqzyCo
d0MUaSqB/sYlN0Abu1pD8Nq3Emc7+c8shoLPmiChI17G0MKp0YjZPFqdArkjkleRdHwWKnjgVCv6
QEAA5/WJET1giHOs664PZAsVkU2q/tGu9uR/DAh3P0oRsQYwKQ32EljsQOe2d+BfgFa/S3jDwZeb
Fz2hmwOhPHTmEBea3MotaYoNx0pfClydh8Vb+P8vUbjPhjgoLGc7AL8fi4MiwvZkAb1788Cnp0OQ
mL5USxURHkAkYx8EN9nYRYgsafclvm+EO5odnpRQqe42/QFKl8nBvhtDKKOsXwpjS1GeeEbDr8Cl
KQ/H+2IHqjoxuxrLEjq7grDJSfQxTamQG+Vade8pM75n7nKidbwC2HICjCyj0jPxZxM2u2rjoZnx
rHWvOUaZEW/PYJCbIrXJJcj2K6/STnBzyAUDIufoGmvk9RWS7+kU5kXGemIKj8CJxtMMDzKM5KIu
LuoqobLrCd2Twmuws1UvjWLU1oBjiA4cRyXrgFHARGEKlCUWXIV5y/sZyO6QuzlMwpqDwF3cAwjl
zCGVo/ZzIDhjNrBVmoWX1Zcv1u9JAkrJop3dc/h8+ZURNuWoZctYtlcFhJTPVb5HOjA4oiPsoWn0
+yIkdDSuk8cDDejCex5z7Zn8rakU1YBDKTqWeNmKAPmLZZqfigDwnKcB56W97D+FeZvZzdP1UKdC
hI0P6Z5+xUqEY+ag9Z7+Ww1RzEtjI4KbKTHeEMuKfdnEfaelgvKtfd3hOdKLO2wMRp3GhoVdzWX5
UOSrcjQCAD6eTKY0Bx9AQYfvjZnW+NFDpORacH3g0pTqx/jRqhXFnaVVhPfsLdcx5pvQ5ZZnFtCF
XPYEu0E/hkNa8FCiS5MXCXPzywOWlWaDTBT8EIAGBwzVcLVSyNmnzVa1eXqqUTUWydYaVKOGA4uk
r20WLndQ8ENLg8v23Fqahd1ycnZHcgV/He4B0TH+tmY3oLEQ6RLrHJxrXAQnjNs630eWgdrEKVoB
SEVpRtEo7pk4nzqEVEvqTMp2j2NVcd7eu1q0kmYlFytiSkUbEy2Fxiltwsfz0JonFkZOf4OADXjU
hTTaTU4FZVxzRqkuT8B2aNSQx+qUCX/4qTSmaUcUUjXbrZfxqo6xjRYOHroOtjKU2H2BJHRhfer9
z9mth2LNzLy8FBrmwkEv4Wzn0h06ZKNv1BgWKLo38KLtN70aIyJynITwPGP7SStEZ6KiyILUP+st
09pTudyTYTcWXuD6C278sZ0jNEitbIqNxilGSBOcRpvY/N0HSynituy6misgef7HNOt7WSMQS8kd
DFhALeoUqRulgVrElmx6PyAE8jyQUd9AQHmT9rOnuFedKPs7lz+W8wGOOp87/UD0+I2aLALUAvtg
1VvACTf1IkYq2WuHUL7FNse8fzO4zEU3/OwpsnJQJsLLjEDyhjzMqmXmBzAplZd7AInBAXhaq5SJ
LfoXmFgDRHC64YCFRgyNJAMHoIGjfcO+D7/Vs9iMfG76QgvcykRJgcSS/4VLy96mNAaU/LRWoNIs
mDY+u3L2BtI14KUGLWCg+yWRJgce0YS8PYxV/r1z9uOU7SixeIK+e1nOLiHQqK/z+YPhv4MF9EjD
4Yr8ROyW6mcotvG+Cq1m5LHwSCB1zvjHZ7keJbnwEzMdeihJVo+y8U7X4t0sGxjmpjf1hxvw0xJ+
uBYGh1OZp6Xgpc4wX4AQetZVIUdxX/O+UJeoi4qfWDPRR3vQqqGtqmFowGxbSp/RjpIPyPlqhfO3
hcSQzO4KHf8tl6I0pnX/wPPhOOqn4swwceIps0eBA7JG4nYEoKfL+ZSTBt+u4mguQnOxU/NmmYVj
num+3Hralnk4O+lr+ooTjkj8nQQWCGRHi0Zit/5Y2vBc/O8qUO44H4/7nerGx4YnA0MdKLPZLiK9
FRt3i0VyFBy2EWUhcgtiL2mgVZeJ4HTLTVNA3Vz4rK2+zc7mTLUZ4//si4pdn8/sGMKEmmpABsrN
xABfAmJL8MY59rhSbsF4K7ZAG8Yax8VHDHszNgYKKnsXw4F382FpOs8nPtqJ0WtWV4OaZN6J5Ik2
YgyJrHOW3ExUWsTds5/vn78eoHqfZeQkVEvghAHYuqzr5AKrt1L/7HbIcn7/DtkcWY5RCfMZSyux
ZE1qyahYYibqyYbkSh2XXYaT3W6gEqB5mD0BWx+VmU37v00kuuBwaNs5wvAB4OVXAmZjj4VdCIRF
sW5esajeX2bUqXsJvrJaynM8JSPPKiy5ATKC3aTnIB9fNrzBVu8K3vIoyGwVbXkb6hu3SZdnqa3w
fpermICiTHI3E566ED5CZm0FOt9bGelXLAPtUCdsjt6AqjMILM7hKwmgSlWypF4wB3bZ4tCRCU/m
riMs66P1q4TPm/YQ6aaCyAahzsz/dDR3J8+c5u+7COQkjxG7X7ZGi7LxOHg1cIiBToqceNmD++Uo
aEicMVz1xYB8cdrHvaBSfTEgoPmFx6K1AhGxpcm1LFDIg055Vu0543e1ejYMG9agmcyXmguYWvR7
tgkFYuG5UWsm5i0/3JDbZKw9M7t4BFZoPHpXPSxwEvPg+TvtYEixKkOFNUE3PSPJ4SK9C7ZNjEWW
veNyPtphcdO9EeW11LYywvJGfJnEKWl0R9RmcqdthTFAREqt18ErUaAqFZ4wuGuAsc+/V1nNpebU
+NbXcHnDQ3xTJlkgz4YErE4Yz6qAFG7sIyds2bj/DOCg6dJDWbhqIrqeMWwig0kNvjViUJZaASYZ
oWH+QUd4zCk/RHkqz5gVRYD6RZ/qW5m0voXkv+gwDqN1DeuZ9dO/yAY6iQWOKiZK7ng3VmN3BVQY
+KOZUkw9AtAwDU71jghmPfJcwrESxhecBtXczsMH330VFMN+UWqg1RLZQGIWRaGNJ7e0WJX9Z2Wq
obgaMLAVaKbJv4Eecjra2LYuB6iravLbS6Xs5+aW4LgDlrIMRGkQzIr2HDp49xTyL+VUVHq6d+/e
1L1TseeMMal57Hkkdq973XOkqYovWnFFf1y0VZXdzg3hS+vC7M4wATD8oSws3v7UKfdioiMgHC4b
9XvzoGvZ3wG/RxfZ2x49YQSmtcyzJZEOm+NvGdySkFINT43ff181nB11HTy4/vRlNqw4OUio26xV
Jk0oiec5UOkCQr9lx3smS+lvjVxZt1En1hdB14R9f20rmz8VM1cPpIG/KUX0oo/GwC36oG+G3PL2
IFZnDb2MJhmqqDXY/3WKOJ4Ps1K7yDBezEF7Jkcv1bOAJ+J72ivi0fT9ZrokcmlpTHcXMdPrC/YA
q7sJKQWOHfR909Ila+6fm1LChn+WJZf0J/QsgJUijRue3LiKS83RrEB+D3PUEXRkBkM/G57fHwr/
eVNtIdXMjFep5ihM0BLw+qdNJSDwGVHDVTJzG3/+uCPfMmONN2J8ZGUl7gJD7EjXRtXm213hXG1K
L+pdTi29iUKMLG5NP9zetXnmGZcvE/Cy7hGaENLE7OvnBDrBAzhJY4NaMC5pEEgscFrdvLSGouvM
RS7CXPVxqIgNq4c9TpxXce3i17Cr+EMk5Xso6vYapvsWERXJtE9LsmKRKmN8PDNMjrVqyqbu2C7e
ss7BwTHVcrEtMRnQfcerT7arWPgKHic03NXitcIQcGfZUzHqwjwp0xOHqHs8AlWMvCU/ApNdifQm
Wy0PLIqaJqg0ZZwEkn7VPHrXiq1Q9v2Dr4NlCzL3BB8WWzVkW9jGwxQpc3DaOJp/rBx7xxvEKZM5
5XaiJzNNtteV3y/xRfV3Ko6GfHpEp4me6rX9OYMpEZ5usJ1tYIkio981wMILVouFhyuYX9VA4MHl
q8s9T9/GWsMIqTBSVXc2sI8cIgi/X24l8pFZH2zTayMuW9VYSPPSVCzjI+PVaJcDUiAxayqC3p6O
qntI82zXsa/vq1i8AOPN7jJJKZUxJquQaojsR01/7w9w6LriXGarrRPDayyxVbdF4ozrekXN+2sJ
dTboDVhCbuSQxCHsLqp6ulFPoTSW8nxl3m23rL3bQ7yiek6TtTlNHicIQBdAj8kKHSk83qVb5NOx
3WFRiuxA90OTwLP1uQw0VsLQXHrMjXgfreKSFjv5nbKMRpKxw/ABiay1R0kkQg4yzeP90DmheSTw
mjzYOML4Vsyv9aMg2gMDH8KHr4ggrEAj57dCs5AwvROFPtJkaRfE0EBmbfnaH1/it3khXw0q6etZ
d91pMMzwaN5NWSHopPYlDAai9TCH38c+z6zCXZ4fQzOprhzrx1K1MMMaJu6U8VMB7GvUmhYalvjw
i3Ur1WK6J0XyTNFlKDgvDvB6iFfxCtCMoP2S1pe6QC7dGhUbFQNB18OyzqnbMS5gVfybz46Q0bYo
oeWU2PHFwfvkxi13/DcYnz6zi44xPe9dFAk0USEzxil9ruUPTZuPgIdOfbUANJOwql2qG2cir9ef
ePgONXjd2frFscJSKlda8LTVJWCUZ1WrbQLbBSdJfWI0S+ru4DJ5G+Iwt/krzD6nTUi57dia91q6
Jage9QkiVLHHeh+ReAr1/tnNQc3k3xt7BuyNyTHyiGW+jpWBhjKaJI+C0apfwcsLQttqjoNgagTu
cVkxLlQWcyFTRGASI0/iWs1Uzhi5Vw/B0s523WeTnuwatbyM56cd2HEGwMcKB3/u9cnYyivsfTLw
FACGgMTgiHEqt8bLMVMxSTt97BIKf3cLReCwothcrTkxNQuyx1B8QVM9EVkUbBuZ1Lr9/BPmRNUB
CUH8Pszf5Fg+gFszzOZjQ2dFQ7SO9EFzJu5CC71Vho+N9BRzeDEsyexN+JY2vhsM6zgRNHsklNyI
oxAFyobb6MW1aKjNoy7jOia+CvEtQVFsEZ5Fjq2rJPsMOug0H1Wll+CpQEPfwAO8DVUGjjuyDloR
UbLNtVo6Rz03LeO2v2IJO3YN1tke6ciiRk5QSfn3bAf/q8hubDD/oA6UNw1LMK+dD4ojTsap5yvH
gtcU0TJMgGe8jmY9ZGhsWiTIPIQC4AbiNCRxvcGk/vwKTrH0ac8lQPlAjFUQ+L63lau3idLe1Xvp
zxpvjmjjcjeAUDxITnguSXi5+REwjrCa0gDLPVukJprbw46tURzLju0iNg+Qcahrz/IEEAxiKhar
9EM8OSjMLsn51BdtrYYIdcTc/eE4dbHHUaG2vr6B5GCmzbFJPh3XxaXsLZMIuLcm159OOAsbpBj4
YAWDmPxVDqNDvwZfV6Tsrc+YoWx8RwQU6Gp7In5vq56lwwjmcM0MkQoC2aHH5sC00HU8k1HaT/54
2oDLBnJYY3Pz8DzGpqhO9A5OAp1vHNx60eKScUNYd/odSNIQWEljhLtcHTm7WetpOR+GVApUovFg
eKkfR3n7BUiOtiN7u/kkdWEkSoE+3bDTtax63O8Eu+S6zhn64YYT42UKp7QP6bCYccV9HnsCYAZT
44rmHXVGBvCP8vhqtCeOXTfFUF7vgMEx5JHVlDC6pDMARmJ+jfy2CsB8OASTIsiYYoqFJc1mTlTs
7ry82L08TgCYtYIwbfbS+zSQHAqfuQooR79JncHH7sv2wPQb2zfIFT+G1NHgApcCoMdnDnty/GZR
bwlxcNnptQOhprfGjG6GAbn2TvvqjUMpzthzaI9k1G2okSQS3orf8YA1aocXamrZUjQ+VKE+H8kt
Iyz10sUwBq3jAVgdbbtJMI/OUE96HmY7ojQ7f0WFEvrK3sTSC/gcKJdb8f+5aGqJAtFFY59UJDSG
NffIR70v9ieil/9U49edlgWmTRvhq3rJeQhnR4gjjy+YkVKqLerxatl6skGhSiwOd0+6bYLRBXst
Xr9cxrLGi8+Q9XE/IH4msq+q+rlgJgf0vUWrSdzy2ucN4SgTnGnhGIE+ujTVVWTKQ6avH2sS8stX
pnkrLrFzd5/U/27lzOQPHpMZqhP1L+B4Vhr25Mi7F/i7Ch/NbHBuLBti1I8Y+94k4/KLnKqqLNnn
UplW/JIPvtBj3A9Jd9bmF/RA2CHvRAHjDwpnbXeF2XN6z1xDhcq5Bhc9tV5bM+No5elbHzENWKVX
a+feU3SP3OnAg1ilsiWpzcVHy/HimvK9b+234Tm0SpmaTkDEkHjxjp3ROLNR+Ot8NRmpLlpO3ZJQ
Jwe7D0gCWnAdD8ZA6FRKkDn0tPcX+im7+eC/Ny63VC8m5mICMM5SIid4ZsiwhDLGKUC9FtQYWkWS
WfBZyPDtfWpOr9rROJqsNEvRX06oRKdw5SB1N9HsQJhA6meYhfqa7XjJOX9ow/kzpCBbo54/8Ou2
/5U4KvHC7QdzTPIe0+m+SbWFfFt3QrnfxJrMfHmfapNzHN/346ShhjI/8u0HUuP3wtBLNbuKCVrI
OgTtKyx5IbnG77tDHdFD4hqVn0LudhWPQ+uc4azSTAsol5JnjuOKGF8fbzGOoapMztJQvIPa61xI
x4uruk+kslkxgJVw/QHlrafteMloFB6Lnd6PO+VFgS/9u9hHmlx9M80vaMsjkSKV/lOUsMZr26Lv
SSC8fDvCuWEuGAt5cxy+yzhMb3bYY/huwe2/u2Eb4UGnBf/4AL4tQpKt6owfvRxYm//2ip4/r24K
9XN3JdxCkg1foGW4l4Q/bvwsWHkBW/7Na/3HNnUJQAl7zYyMQbQ1fOgdRTMBhqjKZSfPZ/1851iN
g7z9yh+gvz1hsnO1oaacLyMcVHOBpu744rvhhBWiavCrMBfxYrBobaEYdLhcjArYNd+rcxRCO+jx
LaSWNavjw5h5nNKVuqEQrVxapdh0EXtb+dwprFFwuJVjWv1eupysChJnWrCHFmWmLh9KvAmswHe4
w/Ogg8TJ3lB3e6G3Kyv+sCPYVPFDuxCvOMsEkoBS7s/Yhe6OYw0v9YslpZM+roIyQREYbfS9Y9fw
JbwU0dgxIJAgT0GFoI27c8svW3yraDfsKn+ZXIDmeFNIlMLDwvmaVz/DvsxmsaVRGNY4hiR8qJsU
w15TUxbVCRGfPvjfHyQ7Z+JilSNuFCB+DEghg7hB4qRnFzpKnIQnLAwP/zunddZQOQbEPHrzo/nF
ZwCqyCPQOe+HDztXidivSwm9LdGRlfW4HMsX/HNdiK2czsiwKuGFnQj9Ihf+2MEdSM0R/1k8TgBe
zTcQ75HUeafbLqg85EePVtRlgaoWHPD12iDTyL8oHctNMpEeWDa9f9ZMUwPGt+75HdrofxFhRmlV
ZwnRL7uPVFivVTBvr7spGOplqdt63E3tbm1Vt7frqot3CReL+e4VlQWFD761THOrz5F0uRDKhE07
b2L/MnqlC+5q81UePEdBCcuj5OsSVKqb0ng1HQV8Pgf2PC7grbSmIs+bEL2brnKEa/DQRDm4uqnd
idHH+PLwRzvf8urPPa/aB+klcM4Oeo69zL47MU70F/zN359qE4tpyKMsAnGgJuUjTtU8NgMUXoyz
kuEHU8WN2uH//51n4Up7+ivti7tudAbbUfyS+RkPWRZOnMQJ2CnRb3smIBYPOaCerObpL0CEHTbw
wc+JaCADNm4nO8UHsBT/hxr78zdd5A+DpWVPScuoQS73oNo0xqb64ejKmiG8rcI/qDQd5PMLugtG
8wD5rg4OYmuQiqZAAI8dgug/Ofgv4ytIelSRbQI4kPWJpqCdOXX2A6H4Esbg+zwQG0909bcrsMgw
+XZ61trxjfDCBSmQXmSPDlGvdyQKCs+oA/BefXfAImuxcrG/VIY0fAR7UBQ8h9/hPetVKrXsiLRT
9NrshPNCPpr1pkj6qwKIVRIVqctSgDKG9G8/8ElXFjNg7A+xBIev6DtLVWCRjVv208MxY+ElZuYG
G79v+7p5oJAEcRa1yUtXOOdM7hcDsy8xeh/S9Zle3NgbWLxq8jiQiQhtQMGbWCuHEeLMAcwgNwCj
wOJKjoncAySruGiAKGMZ9ByS+XhVK41gosSieghRZETkLv/zFhV6R6z7bGStVgXJ0+qUxGXBFhHu
rM0XlMxUArWKcPiDzYF5BnHxNNdErdWHZIRtPQ399PtGCEMvb9HYP3OHpEI96DA0OWWAEHTet0/v
RKchDJP5gzw0l21iqOifKe8KoYpIULJZPVcXFACDY06KW/YuD35Fkf78jhe9Bbs0VO6VIfIuaTuH
ftAQiInV8BKITG+ysXgos3D7m0q3Z+Vb+EGLH/psVgg1vHobU8CeKWos182taV6GEIkbA1A8kNcQ
9WKOjyETAwQEynkzzQ9Z87U+YWhQ3NcgpDxbDP7YBWLfuvBAMjzEbD10OXFtX3QQt0YRrt2OJa2q
tORXPkxpU8SScN/JB+mwLmQG7++Mob5w8v5rM88IIPcIsSOd8GIFoY3l/oJkt8q5Tt1/W2H0I+fy
RjghkBmQPFzXFkZ9ebaaFdEej6wxn/qLeAwyKDBWVIL4aZTUY6ng1bhkqKb3b6trGHS7CtUHMS1D
WCJ/Qq5CXIDkHhZc81MmPCwZwaZUq7fszKNWFd4M2pLKrn2zT+4MaYZUFsng9II+Hc4iWoh4k0+l
m3HLP/fhzbnx4bTcojv56M05npgYcnt7C0vQgc6Itw1VISc2znjEvlo63IbKl6CXL71R2OyjmDfZ
JuoHZfNI5BM9sthRhA6x8mnK295A4jTGiHaq4Rjq1kzndA2uH8Ryo0BBkbbWU6iYRlMPXXbsfdkF
DsK4gm7fljgrs+X5Q76pYy36uCXDX7Nj31+/F77xUbC0rFEyQRh+/maXplEOlN2o/GrJ3pmUISK1
gRQu4AMpS4AxdvCqRLIOSQxsdURp2E+sGgOEW8FXFVswiaJ4hsycPTbP/9rRYlauWdxmJ9FdBLSY
HX/P+RF5LhVaXq7yTztT6Qloct8sm5hQfr9ogU3bBMNQwU78uxT3508uchVeM6kVUxlu+AW9jkAC
sCXaksElbM/+DDNOASAkcbNjq6zM8iEEBcK85aXC5ttcymepqSJzrZK08o1e4lmQaGZ/oVxgtSMT
Ay12mRuQs0s55kspWwROQz9bH2wUY6Bcq35G1zkoc80mNpq8UlFB+dM6Bi+Xl9dxzWM3Ndm1WuUm
WW1/zF0MZoi7vOQEu+6Z1s0DKNJZ3kjzIhNNb6OeSYjMDxtU/AUsYsI6xVYvWx9Omg/kMSyfTbM7
kqcL73NkmfCNR8fPJN4DoFXilwC2N6s1m12Ylm6VuJI8yhN5AuuscrjjqhGm0arl/KkoSqpiuZOf
jmo/F0Swg0KuMmY6VKzCBSMmkW9/7HsV7RvBEyR05I+6k8ThDB4F0XUOqaHpRQQpgDNCkGrCQYw+
1SpbYBmw6OicF756rpkb6ST4m38OACJ9DbUG8xo6ruWl6M6xyZ5PMUTxc3JXxiphk+UGHoKve/ej
aUJOOCpL0cpMxcX6jgLMdpt4yf4hljpfynmbTIR/URI3bDUmssrZepM/et2zvVHOt+X9sXsrl+uK
YNplVR0h8jVkXE4gmPYMo2N9eDAvazrc2OaEeAlnUM/DxSnuVYC2oo8UbD+Mr3TUn9XiQMdDLq5h
g6YWfJd3UmB2OnFn9vm2WXpJucVSKDP3HuZU3tIKxCZKn0ZTdJxu4WzEuDO2eK9FrXDqD1DVUGfi
WTU2nuJNXkDfrT7dVN/7W003i+dgb2xhs/4t7LiQFF3ovX/SNhM9ozjmTBvIrfDl/VMt2oHrJUVC
rUjYij9pwWgB5jP/wgriNCg4GYZ4THGY0vsYyrYypRJ4679Ldv/VjOzwBFLSaQU5I5KIvRAALWwX
nhstfbIR0V5hIrKggjZ/p/0iG1JIX51LmMMFS5+EWC8cJj4adWq9AKXTy+W3uuIFJTKIEGUSL7VY
ke0kQ5jf/neD5EQ7ouqRLYZsqJm3vWmBmF1wb2u3wBphRGFX5L/ByGTvtYtfNAplm/qWVQvMHvBi
YZDEox37ofrxOF2IydvF/rlsksDznbLvJ806Uzw4iOgvKnS/8Z30BpN5bd2ks9E3sFaP6CuthJE6
4tCzSa4blQw5WbrFwYHEZwHqficpSbjpJBr03sEPz3FmSd48lScRiHAnvshslPMv5D6phIPrte5Y
ExxYZekNWZGuq7MzuCvTWcqrHcmgHavVeVuATiHP0beqvdxOEmLdq4+3MSHQCzL8VyfJwzE4PRCR
aTUv/JTGWbq0MtLtRbTanJN1KITt41oYLC89ex3ANSNdpNlLQbAd5gvuSdYxAV9VxICG1yO13oca
wfvRPt2TDb0+Vb4kyp7AjScX5V7m1OjsXIhx5dmfi6DXvteK9SiSHqA1dUm51Gk0BcgAxs6mxAoc
ZyRqy13l33+3SqTbW1VydvsEjGFPpFDAF5t7+CiPPocMWHkkvkx9F/CuEkFsXV1WYLztscSf7ZLY
rKSv3QYhaVX/gXgd1gi2QKbxWqvg3OEjBJMsmNGEjYq6ildXz92ehCWME2js/PXrI6uf+y1iQp25
KwrklzMjnJsMI6wpaTc/y8Aom9k3WVKL4KPUY8TEcWoFbTwWDwZEJFsDm2X0vbjesneFStOFp7d3
Yohn+R4YLpRGBaMtXn1fjsEWN41HsQJ+21NGD1JW9IqmTZqV1X0RRGbVp+hPTmCzwxfaacVKk6Cs
YcoUIjMJB0E1Gn2hpPGE9ImVw2LtjvIL0IJqA49a4ltwtvilWmn1d7xCKZYG1xjC36v4CbSTHmWq
YJjxFD4b7+CgCOW8K/0Wg5/VMZMtpBcA+YQ3cWvVblm2aWmjsAn5tX3GcT6+6jm0j4niku9ZEM1P
vaDtUs9rvosXdseKutazy7iBORsYC8o/d5k+6cheuQYTobxX6KkeJTnig2DO/VALU9nZg7ilz1xj
VGPp7uQqxRcsuvCGsaILCZCgcNY9Y3/dNP79LdNUiNG3EOKwujMndwu6Yc9+zdEB+m8v5wWedyi/
DGWEhyu2uDuh6wKU10i8zrhHJRujNjhxclhaAtY9DxRBn5jPh1dqbOzugM0y2X8etE6BUaxdCksx
TlOpRz4MmjJE3Eac0jxm9kj0QaGaNUBs4C0qnWHYy9ZdhNsl9I7rvsnw+KVJi+om7gMGueGy7fo0
KlcsgNQV3pnFjToJgf2yBYMdQAoLS/854OfsLcoyXDIpXeD00PrSPmLd012C3CtrupbTMv2GunXL
TWDujYp6+pNfErw0ApSoMZFZXDGS3WiVXpJ+IRcYnsDEwcO5VOmXMzNmvmjRU3POTooZAFJ9jhwo
ZF6rOFZ3knpUy7PafZsNq2td2C78H7+zMPJhFxHszuuSg6nIGbQjqMkMMYjp7TaYLEEQaBAY26TC
XATpuqxR2Z1vVqRfx4YkH4EEMasb+Kqn4tP1eQNCiBhGbiCEn+0Yqal3A/ajwsn9oeHqekvv8z+M
JOA23i/StlD67QX2q1X94T+ipThANmVX/5C631wWs1cIiKZLtq29aKclBB3EjcrooDnqI8GY1Qpc
Vlp9mNkD1DsrpyVEvagg+Jl6jUeMHYgaF8zUjbO8tNgsTsCLGPcvkE68fwlywyK5hqPyD8Qtp3Qu
iSV01SIYa5wlM6wxIsjyFHcpdGas5XjbNbOEXQ4gu/WatBM8YmF9IiFfqxo59F/7tTjhMOJoNzal
PQ/zsaT5gplrYYu/AtLuVuK8jht8OM6pRS2Yf4WyXSEMfETjrsgeHCRnRQkH0oYLZb0+vBEkuXZG
cRV0Z4NTGhzcdoldo74x9VfRyvgy4GVK/XodYtxWK6r9GF4jbkq0tXEskPj50Zk+4fSVeSIvbh5Y
XggXZTLZrNpR5tnT0UVwNoH488OEZmijRN7O7jYWTbkyoD4dNd7RjgnGQqPrDOK+xwcrFPcVTkVd
RJcMvLZ+lFOETN1iW/yHHjsexGcpdPcQglD9zJfgkYkbwdjEJT9WicFrF5AbMBM5xn/skefeDaW0
6QxYfbVtGXFnOaO6VqmQ9kY7iv+cML3AC7WJfPrI5s3joAemm1wlWcnbCUjrqQxq7snFJm9zU2+w
mnIxjj9ByxW47KQrQON3gWIinMuFWtzhjJVTSBQao0pl4un5gKAkavw7Xk7a3dtp5WpkXpSzUDEL
XLmb8UJzLKTIPYv1ipyg5QGEgk6PkXv+hKrgpxbn65G9POv8eYSiCzEGD08lX/b9Lv2gYoIz8STh
5vcUAXp8x2O413+EqxlWO6WyHaz4PUG89OQ3Qp1nwiF/blst5E2RNvBc09WApq1wRoOHm93zGQ0V
45/6wdtLDUkbV4NPioohcRg8HkrPIX4DRWjUoIAkrRyu9t6QPQxguSJ6h11bYHi3STWfmIAc0Jrw
OdAnIsItGICc4abGuWQbCwNxNvK1kP3gtdTCF24o9PVrMpyBZGLH1JKOW1vYWsna97DuaLRgGbLx
loSwRwxVUAduM5+Cin2V5ieAk56FftGj/8nNkd0WncvtoYmMjMEjBUim6MIwR1xdpFrTYRGInSTU
3xXUM5IzON1ah10+PV8UoTTslyFBz1VRg8//UTPAgiVkB/qw1mASA4gtWLvHd4quUMLqbkTA1uxz
3NQ+ixROXCZYh9DFGtTXZVCoNjmPmw08Ly4zeSAxUyyC0I81nXosQJ2T2SRYx96xrVWPq2Nqyf9l
yyWZ6KE65ktbVjDFy84vgHqE1YA23UglIhZPA4ATyD4ZGbqJkd5AkqdurpaJ6tO1fILeItm+0+Ia
3eGPO2xt+w5zlMs639VoaO4fQy6ezOZp3dcN0j+5UHPcvi4WM4y1BSRzwz8G+YK8+44W7zLR1KFQ
TqWmfBnedLEOR6SPi/NfvX0bbZEedHyBeKYdT41quoM0iyDxusTo/P4lRZoiWilevujjxOGN2dT4
y681f9KRsvy/CFWRuENZxD+kSZ9T2lvsdICnR6QcKYBdJHaliB6QY7fpX2p7vKi6IYzeJVtYq3HG
kpYVI66r6m0YQkoidUc1lqryVxf34PTOm5cvL5BWMN488mj5SH7Ag80/Cnf0kml0xOMgOz+B/twT
n8Ul70TuyBp/3Cpp0uMGAoK3neEz1L1PmIaswHTx4Z/8nnOgwA/qNzHd9G9k217RnyzNJHR+49bj
KPgKy/PQQGcOVFQWJ+rTfgX1Rwx2UNjryQIx5AoaIcU0QwS7YyHDaqRoIhdl2E4VFHjHsiGt4U+F
To/Dha/wtpNkrFcsuj6qjwwUXgDY4X2DVF8LT6LFzt1GXKIJ3+OtV2vodJmbFnbYmEbbreWGB046
Lb+bNiadOo0DHR2WFNEsnJp6ZM3pGCJdo5RuyS7OwL99uCbmJjOZYKpRVdTsBix/02PG189wWT5k
cTRW3FiCCSf3U8m9R4PlD5I+yzW7jlK6HczdCsUsBULBFg5cnyWY35QeTx8u8z6geEnEC9sanjve
Ofr72O+QwmVca2cRfajGFVtX4vSLzGe6xz+jgj4TEhPRpAPH7g6UTYQo7mjMGXfV1G0VMi/G1JnJ
TA+m2Wd4wycDnuVq8Gn8EkkyIGq2xHfx4ImFQVTIn/3/UxS9Df4EvWwejrEOWKo2fAqogLaTDGM6
Xjs2cEOsBg6t/K0ii1A+u2vYics1AjihnCiTYRIo8AC101ZIj8Qg2Jo5NaDboifWr+PCUWOmD3Ck
Tej1KjyNtqdSnUcQ6Wmj3Lcle+yhDLVo7oSxAV6+voTeG0Jmi6qIh5mqQWo75uUfSJ/tkEThe9gY
NEjQsEU3PG+bsPphBBkb25K7dFPceKXF++HCPt1uF68VeG6OfiRy1z1WUzwgLIEBg+hSR6mIatG5
ohKf0w7NNMnxfxrGKevETwvErHfa0a8X07iBgMNZqMCLOfN8X0ooXKCRV1nXtdCVZr/ShdZUwefI
oUHCI/01CRWASV60kajXJmE4zHPuU2cLuPZxBHNgHiqOfZDwJWQbyGQLxP/sZcD+VMkaXddoBpJ7
+QVpMJzvOa6kC7M9hIjl9N5cyM+vtBamK8+y4ULCiyOTWs9WpkrkQmp9AfxxrLm9r3GoXwbZK9Yr
RvyPqdJZ//FYoqlTed/mvIJzA1qg4snaBWUx+Jy8hvIXMbsmGS7jk25XqtMNtljHkWPcHUU52X9K
a8O/jEJBcQB8iHK8O/fmMtfOiIBXw6WhefEQHpUXqKlQSUmwPhwlbcApgnoSCIrO/QnR9DbDjqLo
mSnesvMl1gfOk0RPjR5Mc0nJ3B82aRdwU1WlpcUMaxogCed1EsegDQKZkKDo5zz5Hzm7fVx8IQFp
ALxZwreQEo1Q1AtvbXr2bqfuoDsRrLsyEkEP2JNX7IJ84wzgbJHtlSxBpoVorCkj9r2btgQgKPT8
VU1/cgoZ3EwIhFSdu0iODBiFgVGpT2TxrwLOoIC9VOZT3Oil4KDzAVMNmVulDewBnvp6U0JCZXI6
PhXgZdA92Ju4YdkPOakeDAQ6hA0CQSwFeyhPLhPaWCyWkZOjbW4yLdGgkGEeKtvAuDmQdFmr6hVL
dql5ak/KCEfDJHkB5lJi0HxE9kj8nUflu3XoRDwtSvI/KDunpZFgvQmAoODn0wwp9asLWsG+aYP+
BJcyZY8Fde560phb+ARLVyzfs63/RZeqjoOsUeEZPk+2vnMLuqc4LxCr2frafc8/fi3K9hNxZxC2
f75qROKXQ59qne6unsgM36LAotGfHVxZnXphxeQP1h5qO3kAC32/bLgni2ZAfTijJZZb1m4qhTJU
7eZXOREDC/Vsj9vXLwb6Tbvjs3eJbBqoqwz52KFqcinXq8lTBpGaPfTJy0jETNiAYO5rf4DCKW6C
xOCXe+7vTJ09c33IxeLcfUaVO263VTkJRDV2RQb/PCTKflzBB/J2TnSUrf3HPoHzaxfqQlGcCzaH
INFwOlzfLPWkD54JwG6akY6/coyM5f9MHFkMlNLLw1n5zkEyVABuZJYHcPHOjeW9eeSv+EcCLf4f
R/hYIbMvR9QFw7QEnBUmLfug4V0MON2dEOvBiCGNhHp+6TPUdjKn/RrH5gaXLM/7YKFCsrsawtSU
TGUxkD/X/PuECkWVgw2nFH6j+9n1yOhletsW6TyerMKom2jzWzCXCefjrFL+BpShTsv1/wHekRpX
8qLsHvNULXtUZhFQVJhztSRhAs02Y9mxa+gaqjLNDviOZccC3JC2rzVTpxqQPVg46aNlfhAGqnhr
LJWxz6YazUWq+q0qwtQK40MXGrE/eGwc7CCv4l/m6r/gVaqQvVkjzpzgRcXcGIMcU0GpC91J0yiC
2p4K4PH0PXDIIFbn3WT4ufB70/fPHU/SaL3z4mF7fdsv4vSPEwmdJ2ncKREGsy0bk83l2Jzz7SAN
z6Xvcyy0EJUKln3eddqTdqkJ3qsx43MdJ2qrakO3hnbfymbqLwo6hsc4abq+bjp1usQFdYklk/8V
LL0zwggAEqgfs3wavf0LrxgqaiKqS7gcdLIJzLXoOW8TruZ3fkp4pROWJaVCDGsg/N01W+jxEvwy
N1+PHg0/PdVjbKLPxwHt1GeIGU6FOMfJUy7roxYfChyoXUh/roO0FyLNlpYzPEBo1yEB0caqxehf
rF0fWGf0ChEpVn4JDYXSsQjfd8aNG2syQvDji7XISXr0Aocb+6FX4AtBK3oAxC2L3X/xDdZ11goM
rYPmpt3qs3g86UPktJimvTdZevsA5s0JKIC4RFFymqXiEMVp4S62XlbbSVMxPwZ3mXKAktIhoEeI
9PcJ3isInl5rjmjqFsVTSiYk3oHpvGSM/AlHkfDVU/BtdT+1WvSS76s6HiYe5CrQrQR15nzfIi+0
5s/6aHkkZvjGLzajDZHCbBZtDaq6PEDaGxjVh/jjcyU3PDp6yX5prpG6sl/VaSCU9ITHYFfoNf8y
6p8o771uRRu9NzsHSi49+Qn+w275xJ1NzO1NE2cb7d2bMomtCCA5HG6tqllMWWGCQnmTLqW8qNrA
GrIgO5ttqnaWzTEob7Em1mF6BfDMaE4i4ae4ZBM4DvfBqtMXs+e4bDT5W9l3AYis0fyhOTWBtnqo
F+k2TfTmlEl2mgpwUtZxTM/RlDrYWd1Qo4nX2LpgG9yJ3wZAOuBqRMkIiHReRv2vLIFz1Tb0lUA/
aI2POTfdvN7vNVQ7EwAYp7hPNyFkYCe00AesXU7/vNObejuZ2TQF9TN8d1c8JZQ9CngOBTh3B4wB
cRUOL5C7ESueciKAc0NjwhyqyDt0dCLrJG7xeHJqtGBUxEvctXg7VKH7MwO7bJD9c6/LPWKWlvZI
CJ3UGhZF3ZCYSUCBqMw+85DfKmNy0eE1G3g22RCc++1jtAovrXRi0yEV23xddLrORqlnj5CDtP7a
spbbC9C/fw5fea06AvfzO5WhC7Kgo19d8bm5f2x1YViSlGIvIKcBEpy7IvXjivkt5EgWqx0X33VN
5X/l0MVF127VAxqYDEpQmyZjivjIHkuqInSQ6V1f++Th/rE6WTsLLwBRYSXzsqeFY3Y8kug46CUJ
TSq+zxIGydAsDvh6nw6kUIFZthGN5fqS8KM3bLcJeuMZSWVrTstm9mXgIOXlbTteRqCzggRRfb4X
kb46JKBo/2uuubhQQpsi6rrcY0qDSCuKusL4xPySBQk5lXjfhS/nB1cXHHtkbAz1YOJnV3iRKYYC
Ck6OdzuW6/LGa8BavVF8/0nI1P7VycYuN/0FqxsiZGc+9IDYhjKFM590ItNv7uXw0/TKkeYzntqu
uwIy/NrDOyOzOS5AwZgC1EgjcV4BzREeebFWZs595PFBC1CIFoP+f35HMnLuM27Y2Olcj9y70Q3B
p1YDDHTHypVhP/zt8JSQctLez44khDPbIQp6agMcjX4pMu5kNWULFjNWW0rv+CgJ7wPus92DtoDP
7ICCGaD3/sLKXOWi0TjCyjh6U2r6QnLMhnsXrU5B1WBjEJdBzlGoh/KOBJK8b6t+QSdmVYNLnlo0
vUNkxsh8HqoBEBBNtN2Gz84LIcUB3RrKTN/TEEY8rP1ZXMftAUyIXwE6mVgY9gx8wb+QILfIQlnJ
2ckL4lFE/Lq/9dcRZPMwRzjH6XJC3G5gcub1aDyyrGP97aQg01iNyjjQeVXUhcFux3NmJQVbFNC9
nGADYSukvM277xOBd/t/uN99P1wQ7yoBg/GOLNsZM3JZ5P5PG2xU0U/+DGNEkACDt/VJznM9NCVe
X8M10X61yzmV2IEIQRP3AemM1Bk/Pb4lJVbV42YfUNYLU8DzJSbjmUWLyiMmh4BRFl1Wnkk8etRH
OMvV76+n+us4OLtKlvLEnb3Z0LlrGNNdWDBoQENTHAa9kS0zhr76qIVMYH/9OxTfJSp3mxireR23
q1af9ufCFBueO84ZnGWKN8nSnCUc70S5Qs4x0slMGE2EseOMInAcS6KGiVKbB2ov7uWDYyKgpnj7
eZDUzbarMeqx2ufVZn09mDQbz4YODz9RQZM2tPJb8o41r1pJvP/Hxsj2ho+L1PBUS0ZGaY0b8irK
+w8sAqO9Pi4JzliBn/a2V1Dl6pVeGDRqZ8BC6X1u7KX/k3q6sPzBXUyMrFkIHjJdKPk5Pexr1ZrQ
tmoRgbh2dpfyjZ7olaJbVUJpgZpLzAg94IZgWfa18vxyTyOuzr7riCk7G0IOxXLqXcAmjvj3F8zw
qv0H6dH3/Izsf5VoeWBiwRygbORFDZwOCUS4X3HoTX8glStelKcjTfXlIMVdvSZ38i8qDlcIKj56
Wt04x4CyZcUbW1EZ/8Cyh5qORO+dv3YDsYMdRGFwryqNR013HllP/Lr2S1aUqBGZj5b4DcwwdWDJ
u7ROcF091E6cZ/09FCwG9YO3jR09E0c8u8nC9DGJaCIEwByaeLXmu6Lshi0TWsASzYg8B1thsNLN
mmKuPsqefkUsl6Bvg25S0yex3NeB+/gjcTthcrCGzHb0UZjaSwsyOQkRRUlOoZVoVs+TijbG5RED
442jiqp9cRcHI2QBVxeT850bNGXUiw5mjWsh8n0LIWDwOhqsLB7mF45xqUfEiNUyNq3EgiDY/a9J
gXJ8F6kJ4kID7YwcEuaH3JejP3kBTmBrzfa93iotsOyJ5LzxHqY2bc5XIyWyLrjnJUux1RzrYBJv
4PLFBiVMYR+ivDFx6AJJDYNZnh/uhMkC+sHk3+HRn5rG4XKNVGbbdhquCpt5tgLhF/0fJQvtsCyF
CxJWJT7uSyaMApqsfEaqfbIGUSMkH3S0S08zGAzyE8YsUbhLjiRyXetGsg6FDDzfUIq+mO1uCSsg
bmGnxXExyyVquZpBJiA8yQ4VoFuFe7R/QHMRsYBWBLJsuFvSdcgMf3qn//KMB6KtZbzcmQoLV0XV
rXeZ7wkQDk6u6geVsTkAznaHAEWasMzOSG9NlMNAYxbA+bwdvEVU/C3GoJJs+ZekQ0c7Zq55krC5
7izeCbkqNFnGAl8vGzNyUQ7bU7Kto/Q98T7uww6cXs8cEIc295q1ubLFwpzvjj5uc9HJ3xKlqIjc
Y0mD+o/e1OFG0cRJsa0g4UsD9DXJLg8y49GklkHvuq8S5yUJ7dxxaLFvr0pqOvlntReZL5SAYJ9b
tNn+dXPt7Z8hF0JDUJGusbffds0vXxumXTFyNy3DzHOZ3AK59E1LGUVEXwp96Ly7TeCcHtLdYnCw
zW0yxiTZxGT1fXskqk+SmejDJy7F37+QJ1QQTJHOIMoPHEbnKQZHN6jTGrP0Dy/k0ypo6s9/Cnvp
IgLjsanX8689SNwaTCaw8c4tWwwZZMYVFOauPwsKZEMSXTnqV1FXbd0B9shwJ9TzSUXc0+EXi6Ad
3e3u2I3fgy309/2PJavui2kbj4egq0s5OiepyEy3yOZcgU2LVNrecLirrU5TnjXFLQTgAN0k9hj+
tpjM6CksS6KS5yCPjCWg1dmWmzABk86GZjz9Pw/7UEFVm6j5U0mV/7IjdlCK2aMyK/l0AuZm8Liq
ne1Y7mQ2ZPLGHctHepIuNvv4cS2ioieTuG/Tgbtl0jbY7PWIseoly0OL+RSprjS281foUn3BmS10
XNGPE2tgObI082CCdgy08Wjs2BiK7nluKhy7A9mgpoHDmy0oCdsATul8JnscJ6vL1AeEpvUx/fiX
usP5wRx+p/ExTxip0TK1MqqIFGbWiMe9rkDV6txmPdlrLJgvh5ZbngoJaJOhzO1Utl2kZT3sgw05
s6GyyrzeqQV/nVUey5wjgcxsE6dyGMvTolld/h8kYuU+4rYKW1dfs0IH38BnIERTdw1cjLzv3b7M
JyS6eJQyr8h0py1ylNm8St3nFWqeGYS5Yd6Belz3t5ypvhvYXK/PZgTQ8KFpD29aR2h+pumqTZOJ
Z7mAcK9cqtZhZCWuIhJvn8xr0ikAfYUXn+910BSa+eYt4cTR1zo1Lk10y9rXK0Nhr3ZMeeTEfHfp
bnpRieKS2pBoktWtPeqdVMdEXCF+QNoMN6sDHP9NoNGeLcTOt+oIvQz355wEVjyGS/Qn3CQKovmf
JTcpObsI3e01CXuMM5FB3Xooe4Ok6eT71tayUpWz8TN6h/SxlB2l9qjAKNtufMuOFsfUa1DTxYZw
y2bgwt5xGq+34mfx4j3Fe/ffXR0qPe4YSEdC5U2kp9Y+tLF3K5CcVumyZOm7GS6wYl6aHo9WvH85
HtWnvYM7aMV8ledY2mH4Nq4jB6u3Pli0RgRY8En0LIq4JkSxFLV81u+9emwfQUfXlbWIuvB06V4t
hWyZKCxtwGCSTmOLH6uXN+IGJuumauh1XCVFaPh4H33oHFOgIoctLf8hdUfTxjEPCDasuUMzsPJA
3vDKDZ6wQjUPtuYQDk6qfCnDZnolOTeneiULtwB2sJjmB8Js7pnG5a2b+vS5Sr17aL5kt6E/I6K1
9/k/RozNZsdkMhEv4nW0TPsZhk/8BI/4SZ3lvmgJDj4KnCZPD6/YTsw9uz1b117HYxOlTXrYt4cT
BitsPPhCG5QaoPBIeaDDNooFcvwkQ07SnHwlN0U/H9rjqx01RGy3rCQ7gO4l6akMU/S9XA6k4MKY
KdLI+oiImdCHpnKxOM9O0JtaKnEFXKiSN7CUh7R1rnQnab++JMppwG8M2KEgDTKlS492wuMuEtp7
NlkXT759PAvSEWiDXQHC+o53O+tCLugPVmFMEmMZh0y8FQyqQzdg3QAqPigJ+kWDvkgDDxU1ntx7
gR3eOwbhvAt1rUP3FB6RpZNMFgEZsj8f8jk5HSxuN6aCeQBj0OWDTm7W87drgla4Jpkv12FUjWPn
XFaR9vRyPMlmsz04GFoKYUv7NvXUH1lWxwcEQUSEmzEEwaxH86/3YKw+jkOUdHDPzqYm1lw6Sgkw
nPPuJk+gRGq8zNYPbUylqYMvSDYB8WXFypIzQ6F6IzhgkiD+InIv6cKSqQcoFsW47SA8GRz0tWqT
8S1BJQWHwAFKqyL2CYOwHVkxoyNJwsUoiAUNUf6ftCZ6ezthTCPTt3LOdHL3XthOquUDlo3L+KsG
Y4MmQDE/QWvLAaiXgdNhcv6S9xvQbYkV2MCos0zceApIVbRvzlR/az6XPA0yV9xgtuoDv1r3fch/
plQsN97+jR0TkzRQqP/a9wYtAFy9vrNVd4LH7ofW0WcVQTlThb3AIH0jnz+J0kyx0QgpMycJUU1p
FW/fFGYX3zVBn0dWreScwSt+vFQ0M0shh7Tj7IxAmmO25uekdZpsOmkQ2gV9jkc1A9T39wOjFREJ
QCIN4yNZqlsP4XtUOh4q7j2HDJYyPJNOHW3nzIXN41zDezlfISmhOkuh8KcYcsHbJ4tMUXAyLZI8
Y7LVOxAcDpGG6ij4ohOdzybekGbnF+YczJZ+XwNZ4PIKhnPTfIgt40yg8pNWSiMxpqd9uKFFRlAt
2esoj4XIeA3ZLiR2ACwleMqWDDm+AF+CJrsYtRqEdxrmPZODMJNxrqVWvR7pjJP/RhUyfkwUjFsF
26krMcALBSspEBFfE/Z7xyMicvI5/BqHv8f5p7Xi05CX8oY8ZJpsuQ7aY1A8j5WaE4n/9jqQpJul
14nJ/5HPYeQBPVDxtPNmfdUPgfGQVBcQ72BEcUjwHxixSOUwdIehrniSNVptbBjnd5WKPRs4lSPh
a9w7ocBAhNIagb26KCfwY4c5UG+NBOm2QxlhRU8KIFORh1UyeDOmUrapHQAPHYX6JOGvd5K1Nq88
3k4R+d4XQSQJeh5iCn4PuKa2tmOqe/LAN0pGhFQloO9SP2MIpFo7VplPAOmb4naYNR3bcOKHTYel
VbnsCjmNdqh9+CWJNvk1sJV4XET5JzgBre9WgXk87AynRCaWfgEz9ijW8s2TJLxykPLLGtKWpyri
a6skzdCyc+niLfTvl7TT3a8+z420Z8GUqMh0Kd6zfCfdhvIG4G3SbMBqvKh4mHgLmuJk85FYqtYq
bSQc90MtMDIxqsqd07P3z+URy49m6p7tiJ36Lyzh3+tVno2GaOHObnyBHetY4kTxOMhI3wOklOVz
lmKaSkaCjkTaLxzexopch2jYEX1Byp9bcWE2E+cmWHc0Ey0DjsCw5K+b4ek5/1h/RrhcxnoTzm7B
db4QafoO05FhKA2AHU23SpcZt5Qr/MGEDioDAbsBVp/EqbpIKgu98IOA9E5OKF7QXplO+BdKGpAQ
7XiUSjUDF+pvRpcHBeS/qVMx5jkCTZ1jPtE10f+WwEfXvpQR6VxPzJHYNaVgWTKC1yA9p0LC9htD
GMzcy2jTqFhJ+cUO4fBapBS97L8uHmPMVtq80t9VRKG+Xma8dmlUwlkHpdNqLgbAxjMdH5XXcT9s
G67cYh0mR1jeKVhMB6D0tPx/uIjXMEd4Su+6nYLWVN6j0GLr1nQVSq9g/hC1BjdE4alGskaPplsk
ZsoaABN8gC+uoV5qhJ7kVJ8mJr1s3fpfHnSOVSWXf7S5Xz0pFXyyYP4KTLh6mxsz9r8StfmbK99L
a+/USZODnoSS3a1Rr3tl6KOEWvKFTyKQLLqMBoU6TOFCmQ75C2DPTX5M+a9raThiS81xgWj2mxHO
MeqqPVYhWhEr1TY2uvsomIIc4ednWwIE1Pjs/oE6nZQFDsPX40qDj61OYBEq8q+HWa1YUJJIgWIM
/TXX62mRBlyyr8Nh1efTtheypPN9N9JSOvXNBRsB267hByq9c8n0cpj5DXspq/94z/Bgoqqp7js4
jejbTQSUNlsBwGzCMAvmDl86O86IiIHmVFZcHHTp2oKABYhQvc7fDoDZNd2KyTOCNb5DzoYZBw6i
K2suqukM67D5CY7PVZvp2HTxKyDBhQCN4j4JGoi/TNlP+T0UKOy4UdWLeFp58e0Rbbowaz/R2hlE
c7uRbZR2qmOOG4yPpf8GTsy7YoHiy/i8DAvPwejUFoTUpKUKMj1/qSxPAfxymplN8okuVaQAVFDB
DLgH8Iq+FgvqLI2bm0KuT74Ia8ODtaxCXueg+QNgVEYR8Jw7MdwrJfyME83xUh5qlOgGdv2q5rKC
wX2iNVR/3JQ4bWkRqhbiLw5jtqk5Vxl3QsjWriu7IpQyC/tDd7Z8pQe3YcJ/Td103HAG24E5jsiH
CZvPWep1SNXChpux1a74ISXaUtWTs0vdmflEsHucjo46ULpzYrLGKERVCWWmmpy/swlXwdEB2VuN
ljAhux8eNnFU8cwMPYjRjBeT+2Ag4pU/XEMzhtgUd1IB4gHxumJDWb2KE8nj4D+2vS22RMLGwE1u
FmxzH2ryUyZz0qxwiS2NBKxHAG1DBijeE6vA6gRBd5KIAClPI9KEJPIWwqyO2BIj1F9lNfkAs6fS
VsmF7Mv/N9JSgM81rBwFS6iDsCF3FFQK1EWOIAUf4+AUjS1ErVUywVF2HPOj0V0o4d+61HCw6JZt
9beIKCdIA6k/3K5/IKwt8WWoK0i8fZHIjvFPTg3O8rteJykwdEMXy7xLv2WmHD0C35STDdlXzpY2
tg0OV1VKEFcXUOZzacwD3XZGbO6kFaYhgIv6jXwrNhqpfZs9sL0v9XEm4HfwLSumsXV+MiysQOiT
i0yCBxZtppAGfcsD6uk2beCO9oBYKpJWBC+gSzE44Q88M8rRHuSt3V8TcPpBmaTMppmrFR8/r7hg
MtL4FDuQLzZJfu7rJfzvDugae/EHoSKS8MCHS5rdC1pjOoeTWsRWDaGaYB+U4f50DTB9cTHh5q5h
9CriGQXtyb0BqoIeghPfoVYRmGMzbVqaPJzv0vXx0pkQkxqoweEEjiqYXl+MxacrPY7o258jaDhQ
jMhUXnlewq9hv8yyalNduYu/7Lm2ORfoCsm3gWGbd13C+kP9cQQ67ctWPy1J6oOjOi6Qaz2yzeVa
6P25qlyqBGTaOl5ovjP6GFS0D3kB8EQpp3xySsSfZwCqkV6Ll+gC51hJZKyyZh5EOHu4hRXL6jiS
CZA5B/qEe+/SNqv4SVcDS0bJ9PjteEK6eFQ3n02VypFEqHvOlf8gz09sFsgDimWIisi4cH1MGldX
OOqghHRO22SLUtqIkl6CO8KwzZkpvJhKzgT+rcghBhD+ddauvOZqnOaKSNK+zqoWBxk5pSyOXAxs
HSx5lU0N6bLlvxOpoRE7iA4Ydt6KTLdfp/3PhDL++YsU9WWtdewsyHZkpS7F9FB4jH1nm89GuYQl
wyimv/rOnprcTSQieOGWGyFXLRL6CTjR39cnwlZH3FDRKJhG2s3hZMVc4rnXhvpT0yA/ng6NdWGf
Fuia3LcfDVZEtWpzNKiuOLkMRqYqL+7qPA82vy53yLwBnYQ4YJOOqt/JlVlcaT2vEXTr/JdvimOu
qk4pc7mzBbRb5z0Fd/ylVStzRRke98wAdzS3MizWjNhutvZVD7DPHcggoDW6LvKCUt/xxx8rMjOp
eHfEXbdQJ/pnU88JxMeBpx+QHvyjVs8R1tldunHFzwo1OTZThZ16jK4KW4NiJ4xtVcs35NnlFGzG
2uW0X4LtwYhiHx512rCzgbSOhbDLO7IeTImNCXdLcKfTrOeu+h24kGODp7wA2pqXOrCL7j9uBvm4
tQvOa+yuLP0CxCdEK0AhCeWOjHJckZvM26g8e6NzbgGdZ52aXmx7PuGhBNN6rUQawxFxPOZoCBeV
rHYCvIn07JEh5uwrlD1AXk7Dv7kRLQMSqAYWc4LYGpXC7c91iEXrMBrY+qsFpr5ee+v2P29zBajK
40YucKcXDNeBXmvmYuw9ymZ1ySYFdGpsYHQXwXsfUF0l4vgvOBnW/04NeHg7VfUM8aV/4hhUFrx5
BOqdqUS7Ig55PrzyG5LGYRt3N8TsGWpms17JkXcTBj59bdZ0FPfTee/uTSYoVRaC2/fNjun5UlHk
EsNEqibKpv8fj2en6Qan1EyC3ZxpWuf2vAQxk0JjptVY3PhCOHdx7EGrZwI3PCP5jTmIc0a3OD71
BY4r5R3x7mBdo7S/i93u7/zfNyogfMUsOgespYVekQVBoZBA1knRsvimj4utBuNAIlllFOp1dmY7
bgMwrHPPfzXCRDk+5wiZU1aOYpcrNceedFqkZmthOaVWHPQNz/j0mDV1FrWFCAJxtd2P82GSJOya
bOPxfinxtkSAgELLlPoom+J/vlu93i7lLmiJPQHwzC+Ml3VVgkOX+7u4NJOG19nWhmGSSlQM11Ap
5FlO+jVWQTTF/4xdUGuSEyW3GUTPlFbjX+YfgrHAu7s/bqP1HN6jGhDH+Mk2SrhgwtCf0Wqxeh5v
P3dPSCUDrrz3OVtQqKrEd+Px5/BjmFsfbpHkGVi1IuzUuLRf52Bmm9EZVjsPUQTlkahv1bdC8j0r
u3sxwJlte7dp+d90lplS43LiaTEE0/+nOfY4ii+X93tgFzsR/qUef0S4iPU4PAFWEebG6aOrMJgD
C3/94H3fuVhY4Qvw6AMFOpUGb7X3ntnONtLVkvyXmSzXkJBmUsLR5DnIbmZ+OnymXq1G6NoLItas
n/+VQGWQo4zSMW/r5r7E7m4JTKXnqdH4/jV7XCNmhlS/JAbpSuBz1YEd3oBgZOILwc48zivsZiZq
ZbEoiabbUh4w+2YgLiZMYIthK1ViVlMvzqqP6Umtloqghyv+WtfE5ApLpelmebxTCnJgw2t3mBgB
sKmiicgdcIs/lIMt1RbQO3w1ynMw+EBadO1jba00ZugXdGl2K96wJDvJbnN3OapiJWnbO3vErtN4
+fZ591zwJErwSNYHD1Ah0PBUYCGfSGF3Ut/mM/Eh6/dO8xo7J/cahtaiNyJzuqcQ3ZjvANXkXvhN
bF+p/Gutak0OKjlsik+fVwgaeyt4P7doOcqWuGTDCvi5P6eVxm6FS/CheGgdqYnEkk2jmB+cAPwc
qb+9ZMH+QDNr0V6ECCI3gBkRpvpIEFcPjtbAMwvr7bpb7/HlwNMgmIEUSuzsPRxIZbdap+PUKXn5
IJnl5b6QrAhCAjwCgH/6XpHWGcpbAjkJui6mbnCOPrTdGTdUea3cBeK+hZIBQKOhlwk+KaJJFW5h
eOtR/XGeCTzw+xAzBkehxBeU3wGKhiQkfu0IjL4pbcbfL1z3X0aEYCPNO0vdbzO8zn6LrVlmUjM8
Yst1eWTaWu5XFiPl9EBgyvXvNisdKMM9UZAufEiTxK4CSaI0iXzFDDFj+PjWP4tJn2mTzTojVJ+S
eOXb69PLfDKdyu5x00ZnPVZvQFQ9igLQCaefD85AYZRWym+kILb754Ad5JT1A05d3h1AvUrQVy1U
TkJSOJuueoa82esMOOlOuA+TEve1N9HBAOE+GfSskBN+s3Z6YhNAwYqREW5pT40QOlFAw2eMRlqT
AtsApTvNY/DRx6FxZoSDfYbJ1F5Vq++TjUe5tRIWakMqj5z20eVBoMvOJAemHKJl8vJ8eAr9KMlF
0vvw47yz5qXqzzTMT5TPSYSpHED2gVqbdg4p/eLq/i1vu80PbZgoXr6TPrkzXvrz6mS//cQ+O1Yg
QGFfO6wzg0m1sO+gKQ29GYYQ/DRhbKfYsp4nYPEYDbPW4/Jo9Jnibdu+L9GVHFHpqfD6bDicDM2I
Pl2lIR3P1lmxBqFFhUo4qe5WIixhVdY8Idy+WoB0SU6+e5Ym7mrUTccfnY14l7aPOSf5jQMqqyZh
R/zOeeCasqf7M7CHwTdqJcvr1M3L0n0viiFew747ME9oIs2zLSQc9Wnrq93vcCigYQr3NX6c917Y
dxGO03Ld4bMueTi4j2ktbawDJ1+bI0LsMRX1vXo7f2iTNPmDl9ZpgAjm8rylyz/jF4epvpm+pxp+
tFt8Gj/mLgAR/BZIq4BF9oB1E75OUVQuW6srkbuIBxFkwfhrhNyEdQrFaBWH1Vn2sXZAPnoRKAxN
j6u7W1/NXVrY/4hfDP1VP7f+L9MU0GY21fdAWQo7SbW/J4QZtSKYawmruCpBrrhUlC0/4mz9Gw2j
FshnjVweG7k0qXBxj9KvYbevNYIfGsAWBr9UpWXMzVrgr0+oywJb611zgWEYmowilJrQIZ4WEYJs
mgAiBvrXZOI0KF8aausu/LKPkp837wkVUGkV9hahEs1Xh2ARJYg932rBPGhBI2olTOTsor5Uv+gd
KV3A0K77h8iOaw0kEzXw0lY5t81TJKF6xqXXCWjl7KeCWAt7IQOo1irSGP6hd2Ehh89fkpSmZaLF
Iq2mnUG4xv4c74tFcPGlGXWo6xgqBG0mTEeDfxz3yvmCwQQIfstkAiBuWiZX7M9lOAvY8sJXcQjr
MepoBQ35Fw8/wMH4itDqIy6O8DoQjWPLKKArk/FuK0FueGWaxLRqFlXi1kd0vleu0TsISQf8cpr+
1ROPe3ww3r1G4piLVsY0NkA0g6QrKZM47X1ktUNjpn2pY5smvPkCM560GBv5vxHVbxch0hn7BNqH
aBXFlPDGv9kN4Y3cCdzyttHpn/retVoURhE9pcUegaKQOOeo+ghuL7+J0rqtxrr+Qm0CWtCUj6kv
U+mpJMPEDA4lwWLxkpAd0jkSjiNQPpPe0n+JOe6nK//U2mR5jtmj6P4MZ4uCdPbAWG2cU/1rXFCg
UyGOmFn7x+9UEObRQfiK2y4ktGTRVTC4v/G9DT2NWKEmLhp6HLe4zjN/KmUhalWgS50dSbQVtIuT
+jQnKgNqn0IJfEnZ0wqA5cZGiiGVbUNlb/UE03sE95pw6obFa/74nJ8aT+tJSQvJNWjUJfUvWWc0
wVZEo4kt+FrsEumA14x+04GBqj4TMzP4R0FS+OrRreHhXIKoJh9hwAqxTeIcopwa2PKRgfJG5nZj
ihH8f0WBEg2hBj2rJI3uN3eX93ikuV6oXR5BJNmRCujTDn4s/L2Ov43qSPZUrGZcujOa/AuCIwbT
1Ce5JI4DGewEATHo6ALTJSZizR6/3MFhghURAjXLtl9ZPgIgCDZMsgyzYCU0DnHgmS2kOu+d8azY
5Hi8aZDCKSW2bGSSyAseOo//PCBGOqWQf8OOshtyxpD1i47Dhm4/UCKe7uIXIL/VY53jaVuOrsQ1
CI7f+7htiSFsv7au/f7zJhpKORA7+xFeetL9eT5+Kl3B58GP8kc2eUWIHd3VL4OV7U1YDTmpIwM+
+Bs0fZsj9RjQXKpJMNrRfJV7GUFEwyz394Dw6ee3hEaJGVNeGdkq/jeVPBp+6Z5uST+pQz+zLJZi
NqIbaxT+3WoO/zoBeg08Gfn7E8IMNKMMwrvOqbVu2F9eusx/EaRIaWjfF/KqNE4djtE8mn9xw6IZ
XyRBMUmQSLkdEidOJg30vEPM3zjFqol+8s+gpPeQWDow17PnZi8K6OoqBkdz600qX7n1XmCEdMg1
yyO8Cw9OYjrIBnqh+97Sq10RxWnZShX0wKiPoBcdlBogOIsevoIKGjFndyy6BkkxkA25kVkO47qu
SSstX3xEpBKfvhVuxvUd8EfNSiK6XPJN3861tObhxeHykOo9CqpL4AsCbZEzd6t0dOAnnqe0LnJO
gEHvMmUpxJHMVLUs5U9fQkgkSfNDiX6cyIzWLXEnu+5SRjujAR0o4jN0wJxwMl1GCMVVfMuCgyE8
6/btuN+Ys422pAKDQVF6st/n6bgRoYwalnw2EUbD1hEKLvXEi1xmZNoIj+6/TegWD151r8iLYgNZ
XmfEBiiO0ats9REoSBxvBOdOQwScw29DCmksOH0GYwPcABopamNtURYJ5H2iYFPR7mIZDhIq6pNG
sl/Wk5WFW+obz+z3qMKnM0asNuXyxwW57TJfDCpSPShaqktwFpS/8Acj6k6L2UmKOK4/+5aKqiYD
mm19rEHbN4DbwcUDdmnJ61lgLkhUF7CqY4IYp89vlcSdV8UrCyq2Z4VFqYoTvX0bpkBvYLHWiZYQ
WKkQJJJ2+13heORphUaO7xNUOCUunYYQ9BKfp4494hKymbstLeB2sqnuxj0B3F47YhGaLtnUTKuU
0tEPTJLmQl1CEvlVLl/vVr54ZAYFSY8ZV1b0ReN2Gnbzrus3GEjc45CKt/DzSL2nTyb0tWV27EuE
8B+8QIiLZSW4lGIUyUUa8UuihqTdNNWItdH6MFhTsMo+2ZAOtqa1L9ApKLawiP1D0PiQB+lItQQB
JQF2EJYYYY/uNSrTu77JVmsgus5c9hIlhEsewCgaVsZZgqookWYhlOlNEL5a4u1obriY1kU1WCB5
SxpMR/vSfxnWyE2yEhYV1J4RCuE1TZVZCk34BUqmxUcnS9rqW/qxr9QIX9MAep0+3OJ7+RMacBeB
mBHxg3REJ0CbApPCak0caDWknH855KbYb+eI9xjDbt318gr59fRcLythYylBqMffGhvytrxFqV0/
79ZyFhGwlnuO/edQH2hdvHauyA+pwOcL/SG3IA/bRjpSZ7Q+6aPD8SAyXWken29J3VEkqMvevLRX
0fG8y7HYOTlmFSZl1W6SntxqFN/bGH5a/KDCA9aLFhOYHd7m6cQ16piGf27SjBspmpQlNCkMjOFt
rXGtQU5rwC9zBYQjVcAQOXRBCHHXflZm92Y0GRWTWoyPL8eMeQJgUPzs3Wnw4rEH1L8zLm+uPHsp
PhhjaFZy+RNW2WmDDXWhfdm04vkIodYEkteUI8nukOjFzlci1YFJjZ9quxevIWjnBa5lDsmJOceg
SLAM3RGGwdK8SdiWhSl+4bvIPpB2cDTg362NdddsEjo08FMeS1VQC/FwrR3tyEWkGuhWabMZFEXm
125UlL2VRJOPoCLwJsd+q+/4XdllSX6A5QlBndlMFywwsOLkVPcghPPY3bVXaSX7salIuvHj0ILj
br3o7mlHd/ieu+5d0H9Z/r1v1qx67vwZnlo6/RKxkOQETMwXOLmgaTIMzpf2VWjwRAPmALDrLhLi
M/Y/O6vjan5bNp68X+bP1wUSlnXThhWDZA2C65gSpZSrhPUWf5ETIh3PfEgGujtP7W67knjyZhV5
uXYxtFU1jilH57at6KV9rrJub+D6/NB5oxqmystaAmpm+iQrriyZnM3Bze0u5omMRR07gb9G6Qbx
P6oGgQhS0IfEHX1tATcdHFG+/rTxZrYS8A7VMCxtxL7qPecBCchfb83qTSEGe3S5VIHKQg82uBA5
Vr5Uqvq3Dn7Nr0qObomUiAdRpVWRR3gr581ZtC4p48LZ91dER/QuL9zAg962mOftOk0htc3jdMKe
ByyaBH2izqYehdRMO2SH4eG8IgtLJGqdbmkS+SpH4aEwelbRmADJcYqFZ+TUKLQKdex54t0Se2P2
4Voizrma2Iz2Q3Oadw8K+fHCm4+T/oRd79BIa3+OBpVMW8OFJFNX0nPziOziNyFFwzkKxf9hKTS4
lEVL9gwufV1NesPgelqPQUeGxxifOdqDpOLk+3AFMenuNkSWtEMiTwVk8Oi6ehRcn/2d2HnJdFs8
vP5SNmCWOwa+6EwSEr8x/7Q2A8lryDOzJa6vdSaBMSJGySc1aM9VXABgEPnvMToUg++T+GXISPAZ
knxd6zHl/IIai7pUHZf3drOhEbiD6n6/2Dug0D+DoBY2MrKtXrDKt8DF7/s0j/xIOYQYSEgbrhGh
QfA02K1+pUK6q7rj4ap+U2SVeDhtM+XfsT4blWQ8a28DzHN5ZfAnAFoY/DziktJnDORjqABfnntF
vbdEisLkQ3Wacrr4OuHwxCe1LE7PStWO8NImwAIZ5hZNt7pBFvluY1KtNPRZ9hbwxF2XylSqIQEI
byMhG7F8z5WxBsnqlmQFOm9DPlh4nmf5UKAVeL+QnhbULEnP2tGfC5+5H+CI97TzUTbWECCVlqPO
Q54y7ujyDQFt5P/xAwVnf+lFiN+W8fCwDRLAMtCCFLN5Si4ynzOfaBSvGaO3sgErxl9zRFGuwhrh
gc2n35Yw3km4RpgbZqafz+eedeCnol0NMAVLarbctyI8i1xnDNVOTHgCtOOsnw3Ry82I082ImC3l
HGDS6V4ILUnMuWFPJ1RVjEUMEZtdpcexz/7d3vyq8ZtyYPKZB1VfB4hBSMcewkRAgyry56XxabiB
lk0Pd7dmY9jLA4zg30WDsuawTI7+Y8nHo/0WEl9h7+0ExaBDUqAuI1cdiDUkyOQcwpXm7k5hukSM
pfTIP+7SZpXww4IMMCGhbQK+/+RF5eU5N3VY7cjIl0Kjku+8VH8Xi6kXgLWQnJd7jEbxpeVAT+o0
NiNqu6Brc9WLUyrrSE4ThVzr8x+lnWjnQICW41qx5wn77K33aWzVKJ6G6uVZrMJFkgohGuN40mYL
Rm+lPlZonLYXV74Bt/YUrZJceSw7p0MLuzDO5YAaTmyj3YgJSpVt0pmfmlgi2AytrJuDylq/qgNz
J5ALbYDi1PFiOh7vx274utjRJtitEzcB3g71c876BJWsrUfeIJF9uAqKFw9SjIA441QpZJBpcFIY
j3WRVkQCitR00RJesOgWxh0Abi+Oua+xY67Nbv7rkRcwji5exL1aulLc/UImXvTtAnq/U4MiksaW
VNVGZNIS7PaJGRxpzeVrpLoQEj4SJb3CwQOah3Ge6q0tQ2A2z3z011KgeBFR1hpTx2I+dt07/4Ho
0HPqTkL0hxPsL6IB/7NNEMxbXhvzo6eh5FBCcAZJjFWoE/eT628pjYSpbUZSbsz6hKdZjCRj/tCk
PlmoxcpsK79JbJ6F4kNI+pskUIcDSCGQp3uxL9PUi/nOH86Hska9y087Bkcq+kswqeA4hC2b/KHy
CA97AJOI7Pph1iFFeKVcDy/jz97R0IKAGYrk4hMzdYygGSYH+nk0xorZdkOeMkdM6bl0JzRcWgy6
xSqxtkZ/f/U5sdt8r1G3tIq+CWAq/XYsCwoEOS8i7bvdDWrozR0HIqxFp92Wy/36i1Rb7/8XZyoO
F8Ca8wrrxbMHmZL1Ejd7SUSseQkvEOX1nlgTA9r4pMPFjXMZPZyygWZcpKhpQQQa2JNgGloWC44m
BMKHe5RNMJX71sg0OJcjW1BEs8Rv6YUz+9tH8SXRNU/DXYl+yLGZsFMfZoMr2WuGrCfmoQec44ye
q/I/475hW42fam0RA4OMbo2FziU0nTnMVHYTkPK/02d8Mc6XDIy98+hb69aG295WwoPLYu32clrw
i5AMMy4pHfC8Q00IBoVMTT/3km74aGjBTptYn6NY4t1NXf+cyTXvucMCkpKE6TRF8PXUtjHTHiXD
9WGT98nKod/P8q06utlRPIt6t2WlKz+CiZ75JcvxuF/jKJcxWMgzlbZkcXMeEg1nDzBZLkyvzCJ9
nMLKWNen6mQBYrmfxVNnsNaGQPWd4SSffy3IIlQOJiVgmrqF8JlJEerqbGob6AE94P8kkuF63MwK
2wy+hN070I25CKP9QWV2jRYyDnfGNZ2OQAunNdjIRRsRhxQUvnZogqDRn+TfAvLD7tSA9DvBwVsq
dd9ilw9Im8gxFJXD/RT8ctCqsVHFzLA6B1/D7Y11+z9b47yE0LtBSWKsKloOBwNkSlAiz5Kdwnca
X21V1QAcRhgql5/lyGvd8S+8S3ICvq4kDoyiGwUyhEBpaMJT4TPeomnb64dnitgOHAbPUbAHfM7Q
gSy4aCOc8U7GAsOL1PW96Q8igSnbFIF5VxbHvN/DLopa+fTpn9ycl73uOIEn7V4ncMl+U1QeF0C+
pCTDsPT73ils0gLBpfKxjsUgsBP7L7CVgLt2qB3ChD95sKfuXFioRosXCa4JeqHz2XI5T9RIc7bl
FexsnWPpqRtM/9rMyHHZyR+QEkebd1Nju6sb8AFclR78cqHdQZeE5Is8kpdzxfnPZP3m1S7Zxtc9
OEIDY9Lu0+wq9pX80uHRrN1lKWKdburzdCAjjZqOvMz5U6clMx5sLj8v9RqwXKXs+4l8AwCKFu58
XGqP8lxraDaMR7QEcpcD3HUzatvScBBSBsbeoky94wWLW4cD+wWh+U3VY92DEbcRCk7BKaSlYIJf
UIJI3YEv5ZIGMvuu/iNx9oE+74U4dn2DFYeAxa0dp0QxSvRsZgjLnxDItYR+U/3S+Y6beE0673PR
yOhhYyo2Xm6H+NrZ5uXCD74TzJ76ycejLRvk65xeVXBPruGP0lT7vq4gZKjgGR+cMMHcvVnpPzDw
ojPThxx1+8c49cRkCZJz1xVaQEw+9che0H3xERLRGP8G4VP8m3aJiJBwqa4uitjkIgqysZeO+r1b
UXoYQ+ULh9Cl3dewcB7wlv9A6ZB2cOPOijsLt7tTNscIgqhOwKne1aXzDYespDMhVeCT+XYVr1l/
H2T0NkpQowRA3QB2dx5CR2BIs4mDmcgwY1Mk60bpqEq5DwNA27LJl+0UkEL8w1nbAsvrSGJ5TMbT
kNQRKhy9agE/QlnRSW1M+PT1V8dfH9lvBY7Ld9yi3Pob19wYKl9vKTBrdTMe9ynX3OZ5uH2WYzMo
TEEoY/dfHx20oj+YsK2ysl3MuQrVpG763EafyYmroBVdMgAQwGrp2vPeP9gHOKSpJ10iErfwHplV
4c3eTeRm01y7gp7sfB7/bGOJxjgFCoo1RAI0bu1Ii1HcvEUiyyR1DmoOvZ1oIiafTvbi6ttjmjMk
W9Q7Lm+BBRhHDgx6OfJUMOChsq40rnXqNy6avdzTLGfvaFrZPlFWyvvGJISsjBLxk3cgeZGjgCGm
1n6YZrEDQhYDCyNytrKSfBoPKjgQ/YPq68qj2wVt2rR8kz3d4GM1gcZXBsdN5qv6TzAeg6fjFPya
XnnU6xqesvPjhPWMuZSoZ5f0LlIKGZs2S5y/CU1nuu5lOppgkXo9tCTwC6RRwjVGTtMxb+tEroDd
PvyQcfRvB8C2+MyhbOj1ZejgHMLafx3AMam57Wnb1y6soENNHe0irP5S3sBz72ZBpDi7lh4QKcsq
10LpTesIfnMpbYrT7FLssibv1ZUGD16ernrT64BgiEgFSeFoz7MkxFpmtfGGtr7TRIRaxhT+D3qg
qbwvUfDhCyivUxE1e2BgZB3Wm4A2M83SjZL/0iUnVbtEV/ZV+Iw1q3rTYWLGgoPKkBzhpjfUP3A1
7ER4Ya0eMA7XGwmThDCpgjeSEKNnfbaLO/pPgHXM0+2ztsC+gNBFcoWeUZejQ2Tdc0IaNIJ6qApi
UdhuAegRCBlYHTYMc5n4q6NaDeRyrvWPx7kxX+1ZrSLuWf+gQ9vBBmk7qnXDO/gSAFIJ/EZZqD5P
UtUq5RScBIR/grxtjHwvKDHJG32S0RS19WV1njFtoGuE2jW0FM0XLCGQYpwIPnjt6QL5zqJeM0k+
KuXNqY92j2n120juaxXtijY3GHYY9nWETc+RPJGVOsOTK9GZEHvQH7GijOYOm+EzhP66tDhopTKV
b/xpQN9EdufhUyBlRCKj6XP8oteuxcxFL9yMSlThS7x1ubSZe0WbKoQ3kqtzx3avHpiUwc1t943G
yrDAnWyigNxPLrUFEYp9jcsb5QzmxOb+L0iKVDvyRJRNhUotLwkYjp4RBKwCyBmWLcXAW8yXykdP
jWvsGZjb8c+LCdt7C0qGTewg1kPWrX26vCK5YRM+fFOf/LpX4+DEex+N6ZA5XKxx+xwSRRhuavgX
uCKLZdWR78jPb2sENO00XhscA2Aj+H4OyFicCwxO35j/yGv0Ggqwq3Hh/YqNqdn3/L8Dc01qoK+W
lYsJhjN0J4eW05U+v6hBy5nOVczNqRDvpMUvB+ONifUe+elmUNeiU7+cTlG7mJVlIXWF/bNY0HzQ
ChLpaTHvSdLyBqYzt5Jf3Vywe/TFcsP/8Eg3Jutdr1WLxl20+RSgI4JNtlKmb4PKJn+3ThGnVpc5
ElCLefKe1hEMWFYdc0Xtu+Ri5HCEkdrH2e+d9DLGyRO90tZDPWblszc0BHwHXo6BqCgFPLKYwS3E
QjE0XrsTMRIdspLP0PVUAXunO3150SNLox+T5ZTqb3l/voCL5rYD1OQL3tQ8JORdE3P2JU9398xw
SHdRV9Xsc5oL9gXL33HkH6pTpVpe15YssBOxRNJdQ0SUbYWJa9s+AIWlI9wiwhdtSAnIniTzv/rB
HdSyKnG9uhAY1GHJjKJj3cuWRsPW63zUcx8zYLAQTq81a05hEvWo8sjg5gdf6MZN+N3L9OXETlBB
e9oerFGkE01J5illvMzmgISi52/3HsJ0rukPSS5pxjrxV7dhtPoogzH7UeZXg/HHRblbJoqMSr8I
IpGkYmA/sUHwgJbuk5ANVIx4yEFVMWMiyw2INbIOaPJZjSpjHwXJyWUlxrDTN/28kh6PITb98H1m
3ibITE2WJZ9oqPCjhytrfFgVwHZDg70N8A6Tfwfkl/Qx6x2JQj16M+3weXXHvPVsRRycNUWb3ZNZ
UQko4VbU+GStrnQHCiM9JzNQUkZSJdnEntrHga4dtE1E150L8GI0Ma2yTYgDqkVdXmUH3x1MnkA1
iZEs53jCSnCeUL+teZwVK6+xH98TdooWYvlTGYvOagHc0cANmvIZG/LzGUXABcMka6IHWiJTcgNx
4zwhdf56iUmnn0CXni28+ACMyc6yWVgzKGz1QSbInGC3IbKfrf5OrfiRMCnr/vXWtIN36/rARj12
6bXt00sea6XtAZ3Q1gZsjTwKUQDjsQc871JPk5mVJh1xs8s6O+N8FgWa3EFfMVxeZhVq5FQxycnn
mluSabIPEpgjKtWdT7DaZ3+FAtQagzomw7T9e5iz8H4DlQauvtgFyO8GibchBNbM28HY16J+GT+Z
4cGIZaoN8Jf9E3DREqjzolCvIRcDDR+IY8gbf3BLaW+cPN3BllkGLch7252KhNm1SWP0cDRsuWSR
b131+/CbWtNgrtbQiTFTwkPR/m39sbz0pKc1BmaGisnbUhAqPHcGz9L3oBeSCrrZ3phH8Oc3sL5y
v230xWk3NK48nxvCEt5fJ8Cr99f+RilnYlWHbMPr+Ts5xhKP4dgymZJ1k3aJdcMPmYSzBNbwONOC
b7XSGMnnAZ3uRY20rS8ugTcLKK/Tyioflnf4yF5/0a+B2JrItoVQBHl+B6UQsxAnYXdsb/UepTci
/evN7sruYeJyzJFdpi9EGAg+6iG27mRo8J4eQosDZ4/1MzRQ1nQqRVS31VG7aLgyZyLlvU9xFxNj
HYtUA7MGX+fxV0NHGxmTyHHFAMxCm4elQWsjd7/R7nY3SIO1QHT2KjEsKePr8lzr94yEMSQUKKGD
+jIBrUU1Brdh8XabWZeLs4nzz1pyoCjvUI/RDwzJjd995/sU5/h6NNBqaSjYk+sud+oKWkXIhiyo
0zAlFvUcIEdGkg7cubvTWAR7na7mO26N+LzP+JcS9grfKs6ddaOYDeBw52rpQd9RzLOK8adI5u8E
CwRwlXOidHSGNyxrYQqd5Uu7Ku6398Rp54RP2EgBtHIOWPHb59QwrJeLu2uBaYffnQA84ZcjI6/8
XiIdvvni+F/wpWEov/KFKW7GU1r9JL9X9GzusOQDfok/yoenRRSqNGLpcMD0CS/ILnC76nNqOAdG
/pNrflRx7tI72/LSGKsS4jmo/kqvucUZc/Lh96l0HrLXpJNHZ3XWgonOreIVqN4EhQKoFz+B30Ls
IL4VvwJMSN7AKjclb0OCNJtJuTJ9HYFnxlWKvuca1XUHqnKyl5KJA2RMQDwXNBrAwkLbDNLW4cic
mdwl1KHbxIdgZRjVTuWTLjC6kzmMXFx63jF9Mt+oUMfndbtHvZ5XyevSuZyVtblEtof5VwaXDi57
GxOqVX/6FxT09F+FgWheDPeP9Mv2EaKtyv6Fvi2wnlTDMhrM1B/j9wXzMhYAXzoEOwDbcbUfndBb
kahSpjVQhO7s1gfVBA/j4KCkD0xNXsnBQjaRoVZPZmoUqb698D6RRS/frz4K1yr6Vue1JoHSzXxt
5tLTW9n8fsXyUTeM3BMLX5/2rdm2ijJ2e+SKLvPw3IYtHnXude3eAM74QUJTXHxLSFWcGmAF10F3
wHFjl+Rjaa0bXXwwScTkkUa4Pc4veglZ/vFsF2E9/KXOVs4Mg1C6Rg1j0VLqex5ssq3allTMuE96
Er5F7eVfGfnRmPbIamkdKL3B8FRTLdvYCWwCxbvTs89qB/gQ0c9azIPC0WsfbCtQTbV/kHNC6OUr
USimDIYAeZLj8rhvIJSSWCKrQX1YrYhVm+rBTAAdYlZH0KMNSDN1aNoYYkOtG1KZm3K/31Micw+L
wrqj3RPiNDhcuAD5+aiEkC9+zMjCjx4CqP7vjfCDOgXEsMY5XFUMSxt0nZG0AeBa1hGcv8e/1+0X
FX+Weztz+lD6+B1OAET+1UUb9RUK5vBsdxo9jJXRWf5GKu1Kub93rcFaMPKk+kJmn/HJXi1JFljP
KQ5Ge4bNcbdErX5Bw4XA+NxQK1ff+I81W+KGsX2ozGvxbEaaKxD1sSeN24S7pAxk2QDusdhUeotw
evBbNLxp2qDs2i8Ab1IBBylYQmgzUyO8Jd1vGE4APOHXDCtA+H3eNwpUQQY94eMTmCEucglqPLAE
MtN+kvIDZODjaIwZResXPheyRpjBwyEIl1eK9lY5JkDmVTA72z1/frDPfVyRius0GWRFx72D7m5D
cDrnP6qmhKOrgIMSPGKRn0sd2sUaxU0fJqcSWll5NvFZ94mGV/fGphYZFmvAxYmzrrNfi+2sqQlu
GVBPup3TkygMK4PnZQ31kOEAzQlpbYKPI7kxgBTiHWkzpAHgMWmG9GuGxJ5MjXECFu7y6yUoUSht
KP0kFUTVGyZ1P3QGc77d4/9b2q5RHZvW9t+cOCsCb8PUTAddjE/LcqdilRt/Nk03uBS2suc8y6QD
XHGWrvL4p0IMZeQFYzP4JTFTF4ZL0dYPANtuIpiv7LlIqMYZi0UWMg99oRBgWQNHeVY6ktB53kr4
npR107//y9HZB//PjgZwZ+caSvQI2BFPMnErCl8bSPvk3CPR3F4FhcvVOecc0xlVgnihJFc5hw5B
Ne7zj6OtQ7+7WfKavZZQ69GEHXbWzCc5R8TIbbs8pXx1Fg/q+qSEbKGSuWO7bIOkcdoPHh+3cHy/
a5N43Qib7a9znDjXi1LkrisC8zlP4uWuOkk1jrsneqIj6spwJSFNAo8mLfWUIrFBdxeSDppXahg0
Ork6IV8RyeqDAVmrRqUr5S8DAjbH0X5ltx4KNEBJs+vijVYKzc4L5AXoe4LY5Wdj6d7Z0wL0gw5H
KJa9C8NmS+W/Y9dznPUuyf0JGCab0Q66hAxWj0Q7DJHvEctVdQjsPcabXNJE+gX9J4VkyILSQjfW
XlmuThJPRELm7BvNhcZK58PTlyqpTh57hAA4ZrciR8aDdGSsN0ZjqhtK5WlfP0xPVNQPM4hrS4jE
TLgGF0cFlmkeIjnaohgxtDPm5SncFXw0tcQI4GFXYzhyOn0e2Fnm3qLiQwDJzkVvd7y0msaGCAqU
fAl0gqhCbjpyqMTt2PeP1026do1H9vAE8SryKdKd0GLwS4EZt5bhqytMz9/8iTvK6v4+OySZ9vhw
B4Ju9gm+THDT9b/jU6QW2zpbd2v3Gwbgcxo3Z5kp91XeVWeVS0TDJf05yk/0XI+BRk8tU+SFbp3+
yoitjN/DVI1c4Qt4gIPaT0YDjPNc8Yim1FebOTIMPEnzobvaU1W9LcibVFSWYfEVnxbNYNZ3nEp1
acnrtwFK8ogXlRTy9q27zDb3D8p4vsDeOVdLW8sT+IdRmUxk2O+zSkLuOO8BhzeO0c6XzUSj0pSR
AqsmoP6E6LLHnqfGFdFJWHrGuIQmjDDN6It9j0N3NhRCpzp3olPAu08qkIZ85fUVdKUm3EW/n6qg
4Df29KhJcAL5UdPheEVWnDLV5ELQQRgRjawYzqS3h5v2bEmi+vMj8NnhNJgxm1d/RKwiolqc5XmI
MBynKRQ+FLyyi3sBhWwUM9BXwE7SLgxQRFyMZOqSijcfh5PxzcE6Viezqiu2tNsYI2dy1ovDKKMq
MBDO9p9bvfIqcafjSzJFUmLekSzc+wlgzUB1rF08jTTKDbTJM3kJeFRE20IQEpl/Nlvm794FZSrL
zmVHXC0aWIM8MCkb5Cr29JzcwuUmWhAnEpQlWxS7VXE8uvcv82/LmEA/j57LuWZlCuBtCwKmpryE
lL7avSJ+jXq5T8ivPBzC3105XGKI1bG+eD8fV5UnkT+zHayEIho9YJ20mYfyO9i3VCpAEMuj+/du
T26ifC2v2tp7cjMH8Pztk8WbPCb5n+nahnYBOe+kphO1HS9k6n02hQ01R55w2I9jYWz6GeOA4pa7
q2n+MIk4QNZLljm6SP5xjgRWR2Oaowdo5/iKA91DP3OhfJn0RWAS3wQThL+W7NuveG30j5fx1kNl
NCxSixwQMDopG0Lbuf2qDsUqYcI+ucVrZVIpg1AQbJU2camjbrOXh2c35ZNr5C4y/tIIKd3SLIu4
WHfN0EC7itJK5FvpC4QTrzd7gnO6mvp5YpMEvXgu5ysJC3/cgU59mXSIFhAuWmSUHsVzg3qOVO3r
u5o8cfMRdVsvbbDAvybn9yXz5Kp7Q1AAFqXsaexGhKXUaK3Dg70qcV+GuGxZybyoHg8oMa2oBeE0
KMwAdrXbAUzn70FyJYogFCmWrLRPqmM1kTigyQ7lnCEbvkoPDzUtwKhi2krmFbAQXWZBhln4hc1j
/Ky5jNzmVXIIF0m+RtmLy0a/spwu3Zh+3HtN+aFlYqcHQeR0Wirfw80tdHeH2CrtQtVs9Rc8+KPV
UEr4x5d62uhjrDy6oVE1NONU3+UK5oDUd8DvEvpJXsjRgSQwRaZsAyhP66/ENtmFL+ATHmm9TYjE
zPK1kYfa9+fpAWIRvT9JhxrWtaoYA6fHREemXeZp0/lYuFGs68AS0gH4V2Oai/pqVACvoAPtbyBf
9JHKAUqJY7+5WU/En59uagGBfAv+X014ispbMA/o04W9LZAvS//ZNY8EbQDknxg9wuRF+bMrOq3B
roja29S9fFm/knHuJ22gXRjOWH94730VyD/JNivOjUy3jA0dJgMLW7YMjwbIMsLR5KkyHdgiiqQV
eKdukb9d7RyzNWd+QZDVkPomiD4YhyOToDSEhq0aHlqjanM9sYp/J4MkIncGZxziLLH3TxlEIdPT
TGBsprWxtFjr1dk2Sna+Hqia7W3bE/uZiq0avBM4JYO8ezrUsDio9/mg+45nevoV7sAA9wJlqEYR
GoQI3fYwLNIlXI4igq59kFbKcBbE1vK/rITbUEiSjQvbWVt1hAujz7HVzqZNa8UxB3jvW9VhXGdI
11aqLuhjU3mT1zHTc1b+Mnxivbk/aXS87uv+23A7zInPCW+pCVkWLs7wxE/9NNcDpS1h+ynZGNI6
Ue1HL63hTkcRYSm2t2R0t8wgZg8WavS7T890msHXDNqgwdNJZ3NsUt4iUKGEUBIdUD3gIlmqYKS+
Kgq4B4a2dCm2KjcYLxcdMok6PnLbe7qKQGauJe+nyrnzdbNCQ5gOS2TLUGR3+9GCymuiBvqoHCvK
zHehyUFTqhypVA2pzAcsDZftiVLwIehEZYHd6MSRgHegWd6Y2NXUA4PsabP1+hHUJPe2Mn4QWSIf
9DZKowOv4qy8AaDVNOkjc0gsPfkpWC1v9keRdSi4GK5AYLaphP/Ilb9LX1dBL6j84mjFMM0o488L
9DYYK3D1fw0Wog3SCvwYnrU7bUojBR7rwkxdjMBUewKjg1KFX+hZExnYoH27+Zz3qtF/XCVUvDRq
3tVKJNtz7W99rn0X/lxEWXpNWUfnLhV1n2p9F9zImmxYELkXA8XOnssj+x8Nb0wr4uwXMVDMysZx
P4htBczQ1EQ86q3TmyFM0jInySQAMGbQdmpF0Kz9qTkKMcMCtS5ZXzOBK1cCTWUWgZQ7cYkK2a0T
JwBwg5eLRXB/CrZT/PFQS4HNX/+2n90KlQ2qCj06nklTerlEtLu/dbKk5lccCdzQ7SUeWoBubDJw
O+Pxxa/uiytZg/b4BpybC0XXVYNbbG7kKZTWjP2EC7kr4rt94cn5xlHN9kfuQOpcz3rZIQtI31l5
SFUWoTh969ZtUv2nA7tGGdRZrahJZs/DExv5ywgtPu1NzdnzZOaKb9JDssS2LjaFIHIRECPiFZZV
R428qhe6PqTHei9mh3vUsOuEYgHhsL9hOtqZwc94GIStFzwc7CZNluBrvSGU0jUsMh34+aDhFeMP
9vqqCM/9APr16pSZH0whZQm+o1ObEUDE9T7NfJtF10bXjOTKLhFlv54IejffD6yj7+fQ1tKbw+ug
mQYIpIQC14bDfYKXLzkh+V89BD2w+H00qvG9wOyjC2BJ2lRro1YH1OCr2Hf/PqSRnysrLlUxlTNo
YU3B91XuFtwze6nr65Aki+ETOsrXXdq9FUUgw/LDtvwCItaGl1IBv9i0Eg4Y2NQuJkGIeVLJ20Ul
zLU6rmxudTqUurYnU+87nqJATcRma+cRCj4XRvA6jJCiwsDixnPiSg7k9CTbBWsrEi/N4yC02D/p
y1k9LVlD5RFH39bcoYqKxN/HFEnoWIGCCiQ/9bOCFRFZ+CIbyBNxNUAQp3prE5U4XLjWKXHtr6k2
YaR5qVpJvXDCdx6FKdKHrtjx+Zbw78bzvjRlKmEjdR2EAjF7JECD0p2UBsnz2wn28ICsbrJ7LLeG
Di6de0+sWXVROY8ALE0ixxXu4Y64i7KxMVsphFh8dqOhHoWmJByw7vzWxMYXBIjfUKO8VdzeXc+F
KEoq0r1bbW9MM2VC6c/Cp3L1oHnU4xWVvT2KgILue3UNLIfVWzJhOyKcRxecezgHisRBs+0ft0mC
eelsSM5MDrcMhAFWpw+lH73qHAqXhnlm9wxAvbbaPJidFbh8ngAG9ZOSo/PIgWp5fRYndfoJZFvB
4K6q3OXLNTexO0D991O8bZrUIxqC54pYop/Kg4/RVo639ylPZTEk9mLMG36zY9yMyyolEqtqnBiQ
N2SG1lXz5pXzM+TjbnaGmlfjeaVeuA7uCyEWj4JUYPcuUPZcUMdl+KBnnEckFxsP7n+uCG7I8Ds+
6RxpbpqJ47M8jmfbhc6viQj/14l7FT23jVsclK2yWDc9FdQZ9v1pm6i8gYAOnEzyVyGr2xTOCKOD
xYN39owVAe7AqOyNMs9OQHp10bKkDhEy3YS5tmEwloHIzgYfNZwoSfdA2V47Gke4p8QFbf8ur6jp
Q6O+5bTSEObqeUyMlmXAmETFfqiGJzBEwdzOdKTOw7u5VdoeaTs4kWiA8JqgqMiPleUoSVT6Nl60
veksXHteTcLgO4XprCiHG/LXPt7nnQIzSxEhOGWk5fHZYSYMb0pMLoPL1+wv2+X8flD0SugjLiD7
iEXDc1mOCKnZht8p526z/8AVO9Nv6Olq7vFXgCgQzfpQ3rkDF89gNMF42o7UMonEyM3hVC2sW0yU
CQHWtUCSuFQeAih16Kks3HNgeKqGf9rIL/tRSe6Xs8MiCyFcqxkCUdPvelBC1DtU+s4yFFLFbUko
d33SmheYRXVRL0dW0KMf4hZu0k7ROhTgCxHX39PwBQoLUoVeCy+tU6Y4oTKrhU2S3eZxFuHDHKQF
SthnGgWM79LZOKa639UU5KX4BCPA+fFbHze0O1lgp/ENlxyQOnZXT2IDKuagQtpJjBYpRE4ykgoM
PtAWTQoX6NaYXDkpeo06RSUo3BMelwC4/GidEAAjxrSUFEjT1OR2drFbkaMcEpxdRvnfAS7wshWy
0l9h83erYU4RCkgU2y7XIs0ist2KlMtovl7+gYy5ArkS4U5eT2crXEEylwbyswGU6geH36p407q3
au/dCyGPhRr+zwPwOgKu2v1NDEzXTHgDKMJuf3EwHCMX7ymlPTnjvRdbOwPfz3yvLOHu0k7CBGXz
1gKd5xSoshOW4PcnbkWJu8LjK4ATkrAfAN9EXEFB7xsXnJCVTN32SCmnPULiUCTVOf0AkjlaufLo
q0DhF9npAD5iLGJdYMWCPNNKPmX+9HQDnf+ytIcDYcX72dXAzSliNzzfI3QlAofaqbUK6x7dQPk4
wUDeNbLy0bj8wzcGyG2iypDHLGJ9qPhR91VWl6qHw7Zc6gywmmFmnD/4GbqukuyC7kupJcTDoxH8
kXfFaVUhJmXq88N9Tu+LZhAmvIKxz2Oi0kER9XQP9owH0ieN8zhvYEVY08CfIMrpOuw3r5pgYC1e
ISHzs8VV7ZbWvPZehvDsvmofrXfDbX7k5h/zn8wLc64DwYSl+6en0ytgSpbj2pEn36rXgigKWuVp
xkWuA+98SgBEEbBvKyx3kRnVrJd2rhmv2OBfd4PXVYnhhKIP4e79fyCmS+g7E22jDDBVZBnsLTvX
YGexc46WQaHFQ9ECy5D91kNt04rw4G6z7KLQeW7ip08eMIUZKZDW+GxlMaf/YOP5mbtScVUjR1p2
2YWRm9Y+HoQv6nzQ7tBv0K8gqLEzsRSkkfaWWE2MpK+1YNaQ5BY2vaQs0TgdsI9QBL8YKd47kOw1
mvnsNjOJ38citsYG8hsd4YmE9liRbXZChtV6ivjrHpMD39pyQngG4C4VSiY31EFfaRYEVTL11Ewh
2r7EkNsTZKX/JOYr71MgaylVxwBhFfomotUErJX20pY6yTNOeKEfrI75+FmuGFT0PnW9Y9pBVX+9
a2WqjspbLn0cCVoQZ3K2ZY6U4n/t37MShXqnrFXdrRk3cdyAJ0OAxXQysw7Lw6RC03y+GhLgNA2C
eiYbzApoEm7Es6GpX29+vzuCA+pWTK0zweKmBY9cUHLdcdM3sTknw+7Bk7vuW2OZAUk2BqdEmBYQ
1QynrAmpSiufoWVo6kE/erENb2r11saMq6K812ebyI1so9trXG023BMJpTviWr+N8qWQi4cMhzBw
BDbwG9p+NRHcYlcRyd8YlvnfLVjUGaJtS2equpp4FA/lWhBfrx1fOdCouCR3sDSvNwtQZq5vQ7dG
FGxA/Ilo3UoRvvh/HiFbBKsDIqdJSWLxYfy/K56uSqgPYaFTb0KXNaLdCSb4BOwjTzTaqbbQqfcC
PhLtoV+yhE1uHDOCMpKHiZw/XXLzWesu1DUNn0vDXTTfIrisE6CokZXxYDqEqeJaJTlR1xwL15oG
IskOgqU4gPEiWhgCcrK+uv6Z/t1i6izq6quZ3g/vPzlG/AkJ0cuojz+nqhyQBM98wFnjIN4dd5xZ
Pbq11d593OR3KcrZHfDcfzc0/cxAQbmrinZEQwZmAGs4AuldMS5KKq82DazLc1KxzSiNAasBlvFJ
xS21e1EV9BN1iE2l6156G2M/Dmhep88g9APSDTUnkSZl1FMYAk6st+1Kj2hcdXUpjQKGzI/Cag+R
GXoj2N5IMhW/zUGwLXgmeJVGnVwHVecNmmBFq4GEsrgGAk/xaUhU/WwKpsgVBzCAo2wlyaNML/U3
h8f5SJgihQZZh0lI60SVo/lPEChiauoB47D/vDBTg1r5euoCnQoP9Iv9aXuwcR6aWjbKTrXg8RMi
629JFG+0x1olJk5MWve7ynmcbkaNrh3k/4aYsKzqYjrMV/W0AxwkuUmQCo6S7UmC/+aIE90mmLGX
/zeesktD+pyWnjFm5OYRZSy46IJCBkihZ0ONVTD58WYbMlQRGjuFDJBxb8MaBlHb9qD1H/lTIkEU
ho01KSq6Fhb7H/LAB+bYWlXNYi38dqoO+nDzXzLo8LKCvwGNQfn7yfcB9LZDlQLPSSo2nvvlqZF8
fRRInmQrh1JXZ6K1DT+HUCyEs27fnB896MiHIBrZ1sRGupbytREQMXqIUz4NQvWzzuatHUI7P3RK
5W2x6B1zW6ngZPagdpLQX2HHxN7vf+5gVr9OdudgE/g/OgvkygyB8BZfe8gVrQk9XkKItUPZHlre
r6uPjW5GniPUsKVSuarb1Q9kDzpIhddzLfVdq/HRNsFwggxbZ7gC8kPo2uhSJEJqtHcyO1m0WeEA
NUVGONZFO51FxRDHRlZzGHLVYkFHpCK4dMlX69fX2byTtqdn6z9NqlA4i0QbalRp6+TezJJnqIrf
yCfCNl6nYExflefXY86E2eonX8SsUYbs6dM9ddR4MGyOgTWw6bFIat+DU1l69wiwQTbJFQs6SssT
EHinxfhyRTNh7HcmXbpOw7/XX0khez25OBgun5sf79U83cWgES0v/jYOWw9MveHKIpJL7JKK1QV7
CKjr4INWZ6/1H5jShhccHy7fy46Ysv435pDq/2P4ayJCbY/Xf6xLS/kL2k+qgC4PY8Be+R8cwP4v
qEiIJudcfTwyWrT77G48uzCoup/Ys3oYVtPEfRKt2HqWdPH9ZID+4gQJX6/iwaBthFXN+GZdFaGH
WZsoAx2N4FIebFEmZYuX5jJeMxl1Y1+xTaIrN6sr9QkV1d3Zv0c1EdZxI6HQDcBlRBfn3+j/31mk
mSaHcUIAUDcS/NmLJMQcjbiteXLry+lWxjoT8kEMzk+1vUrUl2r0QQ1LYiJeYgIzhPTGZzwlOyWb
zjDrdWhXm1gQtRtC5a2laIxbxxiqZXO7C/s7RPjr8rxkkoYfloL7qpZO4uvUSTY4LAihPGYM0Uco
6A6p85dOrkrcU5H3KtCdoe8LfzECaRjWZFkmGX2MmoS6PbQ1i/cENYraCts2U0IsNbRp654YHEFU
5ZRJ1OKzCFsJZZHn6OEpfjNdyRxLkRbQVgdiOjNS4vdpNaZmbV9Lwb5PVuKwRFoKxJMz/QJ/1XLV
13TO7oCut72gI7CORz0FSbJsKGGi2Ool7PQXJ0dM2npb6gZpmbcQl3aOEE/FHDb7x4zJgp9dIn5U
91f214lS+Ew5ljPude3cPJOHFx56SEBNoUdvHLqbe8BlUyWAFKeQM6w6sjzCJxixBQl9/TboNwYn
YctRPQP8pilkvYa2gh6jMe7Y0x025n2rIQAotCmDCl+fgRZ+CHuvPzrEsGzsMDJlsZPwz2hufcoQ
UszVOBIkdjk1NXSHzeDYRaSZ8QnAKXQ/z+XcUsALDym4hexGeD6mG+z1C97LlgqNlW/y89BoOHTL
ht9zvJNrU4xFC8G1XxbeT97cyHZGf/7bM4Xb6io4JDXuWhUBxlGzrAz2LXdij4N/PObonC4+cYvI
ypXuJAd6P0z3debJtU1f7tYmLsemOPTbVDxbzEr9qjvUW+vvtW+jmWmotdE+GpmPcIsKOvwLWLrA
LW8UX/WBLz/mgP3DtefyIa6zgvEngIJj0Qu/9yue27+GUmCwn2BdE5i3Hdo/vsD9sq3VNUzdYAq2
1xzTabXEPNUE8wYTgjsrbGk3S54iHYgo9WElle/paYBir4MSXV6CrJLHgytPB5YGJacBR9W5uzOy
dv8jyruK0GDNsjOT5K5YrtI84Tb9wV46Ied8xVKU+becLvcjRtjthMdrjleYoyOdi/tOAcQWyYLU
PnJ8IFKkdKcuIUY9eFz7KM+7ztJumUs2ULrn4RyFnP3T0Gwjj8NH+wBzJJTKHQMIhXG9HAbO6Tly
hctI1mhUVM+nkp/o27+fuRnVe/bBM8zEW8ZQAMyfdZe6KZd5J1qkQ4VmsA+shhJwX9CDCRC41Qzj
6gJPIuP7P98nTcwVxRjT+M139etSt1sJw2XCSUnXxY+BDKE09rvbo9qWxlAa6u5yfN1FYove6TIG
zUyGjK2JeyBUMwgr8YRzgTTtfeUbwjv1HQMYnOf5c247aC6yVWYCGpOy4Ut1aRGs+F/HlljYJqWd
9gqKZZWFM1VW0V1rqQi+ON42A8NPl9P8dAA5tfA4tY5syCljdQN4RZP+UOgAtxNXtrAW3SPSSWNV
l77y0u71BQSUxfLvbzeYvlS49/1lJPTnGTnbIGDwi1WGIOxLZvuRKI15LpRlENeJspyB9+ffTTld
SrHKwpyZ86SKJlGvymvonP7rR7yd5pNLc3pEa6IGT7kI1IFL9f0fXhKphr7YHz6rmxxmx3SZwXof
Zf63rm7V4H9CDpi2tnJOmakdUa8pAemoM/s7JWR/NUdxh0TEU3viMxSq4r3a+h0Ddb1urSqVKTrT
BNnsV8aNTm7W0pPUwrm5z4F3CPmYUm0BU1NX+OTJ3LZ+1KX3srME7JhPjXB5n0PeDtAQ8YeS7w5p
i6Yr7texeRQ4j3AmPABhd4L+ZJbE0TbA4ZDOfF1Sr6W+wurbYahHQ5WmRJ3j+e0c8TfhmcYSVi4q
S6Hxe99Sag3ZA27NclVDW1krggO33lAOlEP3iExiPDAtnSLIl4iREg0wONNHv6VEPNKOWmoYtzlE
OzbM3suric/E21w7Kb5XPpRW0zEkRUduDNsuVLj/0dsTLgnll5Z9crvSl6Hlt1HDk3Dyp1CpK1Ib
dHN630YKV0gitTI58T8SCg1+V2tZm5S/NYHB9HjzIRWKAYzJY7vjO9+aK3SwS34+NEOVyu0k8RAU
MWK2+F1LVS3QD669VH/Uish71PqHLnUZqDYzcjcFovld7gp0AD0B680u1iZVYmXVy2OzWHjO71+4
B7/K/I9e5bMp/5cFk9k+Fe8J1AhQpYJ6aJlTB1cnIqHaQPMd+a3+ezCHk3e1MvV6vAMOA8VHjf+m
Gw1/QKweJkPofH4pIliFkYMKg7QXD70fdd3vqbCbyyOpUMg3hgH9aurl8jCgV2hwtbvh9GucnMHX
uqUrBzkckXRb7MkrwcqoGqg1L8j3tRbo44HXGxXesEyE/n82LfP7yzBsQAHAPKW1Psz+HS6z6Ugl
K40pDJjqPdJv8gWt7FA5WmmzvNydrG9BUJ1R6VfMVWu2CQI+ZYhm9OqTYODgcTGpkN6YgmEM5BUo
W4faiRiHq71kdFUeAvDqAfK3i4onOtuEKlCNSLQrFDz5UrXLa3f1oGVTdbAQdl4rO4IFBBnjME59
e54sVKDw6I7nI6ly86pXW2e2mVHUzqMh7dRyyfJ6g1lwGzyrfws/4Np04NAJ2Fjbn+Bw2joIrJls
pFPMz/S5vF7btBxeFvmHACR4C5UE8dK0iZuLfLt55b83JK5OMROoOMlT6gVN+s4PEfv4p2LpEGCi
hZqTZisW9Wq2s6BGr8gcaqRVLBnzLlQMt8oRhN6LzS42DNhZH/UW1032gC6I+x9xjdfkaMXJ/Mvv
VPSgYLRW2onzj7vQd0zEbkuyLsjWFLf6EAyI80kEI5i1jTiYU9QJwmecbtKCkGdXA89Mn/Emj2Qd
k0nB0PFj6JRVRvI5m/IXDkeKSfPWQtFqFDj8W8F+tu8o9Jom/xC5X581FwPFpiQ+2u7JQEoztr55
Fskc7HgmYXw61BYgbo4XLer/4JvaV4s2mOOeacuzYu01yHVVqdSA1ksslik3OY+TsSVN9/+FRWCl
/6BNqnsp9RxL90r3wG2h0BXt9i+FVx2XbMhvh8enZJV+PCBtzZQNxGccMoohQVcBlFQtylhw0vSf
ORaajy2SLjOScc1UftOzxS+qym5qz2lVy3h2lCcfFkQWncsmTSenGqBPwj7489qsvwz6FFHPkNER
7x2IAkumIfU9w3XLK1OKXDqg4449gKakm8sP6G0dmDr1sFyeSFGMxLoskoV3b7YWg55j4j0rSpTE
iQoPuiHjxr2oZQRZNqyYgbM0UduLmY/f+/JbjDNP20hAA1rJTKRrMYv2cuE6Ai59eGoY4xrzNUCF
Y2+/djR4jnZlEVbuw2SP7y2/wJjAWl6BcofKRInU/p7SHzt73BbqkEYNwnYm2wqtINXjoAoXPDje
sGMduTwDiPD2bisw3nAxzV4hjwaKR7VeIP2syHVeVIMZQjJn9UbF/+9sF2XakFWSDMUa1XzoIrLt
+ZEMPn7/YXi0Pdyxm9NCNmva6dysXKpdA4ga2F7FmZUQ5U7h1jMrc0eX0xL7wJdmIlg4b04SOz48
shZ/WTRc/Id1sXMRJ4nOYnX7HwwnCzF3o3xWyHIlEq4i5UE7UCFXv4yLH4JDqLJaSPzC92HlbyUd
wbpJ2UBt30NyShr/JDV4YtbkkQ1V4Lz+2hBD3qpt2ZNmn4qEPLplcfMFdPmnOoTG0ccSqZzCrqj1
9azSawgDu0CdwUQYfrh0hOTGUfNrXyYh2Rzs/Jq28VCiyyYkyb69sH2zvWphtHPnJDIExewrNtzY
k5VikyyXqrmq595pdyik7fg85X5NZP+1cev7oDnFAzE/5Q+DNf4YqN9FWX829O/Wikdry3X5CxsD
lGtbH23UUie2AZ7dAY2y1JPt2fVqJmui66Mj8Qy6adDkdqIkr7yGhgpLMYlHMU4zeKui6Tqm0XD8
cgH9FNQBxq1paGLBii8Gx4XZlfBRBjVcblO8VhGG7zeJueVRSYva1H3bmB0O5kEebqxklwWXaHM6
JVBj7AL3CT/4CXDXq55+IrZ7UQBLJQmuCdSfrbf2Mmx5SmVLm1G3qEerWtf7W5bJDj4WB0KxnrG7
+llnFi36NMQoXcUNDmn7FSnfMoS7pFAXf9JHUr6kqlufM68Ltwi1fD+j6wqx3aS9d84cwKd8V4po
oi+LFEJt9MIZC4HlXy/JwYBco4nc2Bqp1siMN7hRYMrM3Ey2Bh/NGTBOmyFwuOIki6zj2OLVlMz/
AsqU+jL7dYQ2wXy6Fh5nB5aXEj1Jue2jUsdzSITYaRCBQvrxzRGX4c1zjh5jLfwRi/Mrz6NJ54Oc
afvVlC3nvYEqoV/XTMIeO/or5IwutISMf9ZfVk/BC59QZh3aszu2VXHm3YDKu0oeDcam6kJyAwsQ
+x3w/GGd7WvWlZjK0eiNl9r8UJKPX1/guBqECV6ZA9ZNNh/GmksO6IbFWEiAVLLjxRDnhOeTxKfJ
r/74DUMOacCV/1/qkZElelUZzTAdlKhRjYbSlo+f/GxJKphm4WW0/3OL58wtbLFeFFXq22kXHg0Z
ZzVDG3/SUm61MY4t6t9hg5IUd2R4oYOUwEstvM3dq25IZlhPmLzizLJ/toPERKTgX3A3h2PEie6n
U57tPT65Fp+ErvJAPkFjrjsoCQJHZgWcWi7LISNUv/u8nFackVcu/SAnrnd/WEceaQliR9BGWj2B
GQ9LTsB1ZIZgK0Il0aBHiFjRSQDIyHyU0Zde+eeqKzHas/Ha8lAbb3dsm5wJZk4+y6/7D5wVp8b/
RUR5z0x0Ouy5pOvSdcK0dD1MTv843EKCYlPsUup2gCblqBtvFoykEO1JM6eevOKQPaPfKxU2af9d
l+czl3iFy9tkfHoeaTRca3unz5wMZA5YPUKGu/h3KVvkvj4GjcObdPxgHFLcldfbhd6LZKqqhvLx
xr+XSj8TAIIh5rkwOpY88BilNpDmf0Iq8hMYcli50N7oRczasXttGOYKMcBv3wtiNjt2IuRftcDh
5iCB8q4sfdco1lcX1ADvU7jpwtFDiiGqvRV2ESE83fc0qXl2hWCa8QGjmxw7lt2Xnb+bXv6Jkf+z
d3x61hBvSM+0orqt2OB4r/Rwxx8zyL9ngSzcciJO7I0ViaIlfGw3Uxr/6YMQ54LDyMzdFE7bowN+
rmw3lxmicgW67276rj52w5ldpTKWvj8AmrhkFaRB8T04FgVcBof0GVY+xDgDjTvr33YFfjiEofpp
CAUvvQpY4viLKvnCYct9BL31So4Y5t4WzKFqD+SeJwoVHiG6TM3DHAM7NIAoxKvm7CdC3MxY0UXq
ubojmTd0xVOGgCt2fUcbMVrpMX5JrM/5G6StvGiZiju3f1St2JVM38Kjx5/Z7Ph/NgmpB8AEmzX+
YEM+R3DzR5cWJL0bBrM3SmsQrnPL+OniWZIdRMlkWjZ/GzaXh6WOYn0Lsl0JNhQh00FsoslCg7/Z
/EWoPE7JQYiMH2w2J7Zmm1OP8kH0JP//jMA+1WB6nkYn/JxfuQ+LR+Sul9bh2Bg+cj7FJsP4gW6n
5I4RBCIVn63g2OmP2Pa6UwuCr5h/rN0fqpofzaaxdZYrzkVUEh7KBIW+DiXLG5DTfmJOv8Njh4BJ
ZxzIHP72zIYiAnfq5V1IU7FuAPHnbBJL/DCvI6pNBmzOkWsckOIjx+Pmka1+oLvXTlwzcwvGfK+X
Rmm8L4hQ5rXQPrx3XDExmxu8bkYh4ojzV/Qm/L2tX72P+XviI6d2oGyYBpwToK0tMzROouGWdQhC
WatdWSbgY20/lKUaT2f+50mxFVqvq6wTa4qv0jI57wagi4GGYaMg8ajQqT/y8cHnvwE6o0SduP28
r9F57Cy/lczNAdAZs4LXMY7ihr39ylDe3q8wH7FBHUlf66l1nUicbSnizSP3IIFgDfXug7YvUgRm
LLB7/zBkgiH0vC5IBLJTkTUcC+nt1i16ZW3Mvn3m5Iiv5Zu0g4zdWAVv/quRD5/Ex4sD/90cRes0
bUOyBcVeTsP36B0KgiOsPY+X09uHVrIueNb0qWqoPLzWhi6GbszB8aTIdQqMZuqCtdDWS0i+o//x
PQ776hu7WWOtCAFtSoKa72qnKgLLh64Mblvv8flJ2MkHX6+g4w9S2f4AR7SGwYHSj2nawz7Y/AGa
7U2Giu24wY9vRT5PeK37Lx1krsM9Psa7p/y/a2pVj0MF6pQDB+zs3+DLwGS8bV4pGuHb644Ppz7B
qx3aaTc9cEe44MxwDWWd5jaQ9HakIzPwvYEP3X0ecjRj/6VGqvs9xNP1XUXBXRyRIg19/jArDy8G
3uice8whdnq87QiVbV7tYBkM7NVp1YuHZb+XXKTVtcvQ2t9W7d/S4eaj0DujcHoAA4Ln8ehnMhJa
CdLbwvX7BehqAjtPIVZy8bFmHpm1m1CjdYNbuivFsHmNpk4l+DXlhI6aFdUh0iKY8a9fzwqoNMXc
/nCqtyosFL66f21L9dTSzDl6f7HD5RaVA06b5k2C3kkp4y7XBVjkq9PuPpftv31d+A4QdeF6eBWZ
yQf6zHcDVGMejaqAIfBiiAhgXrnCgGREqpPSBbmB8BGzjRdAMGeaL5fOn7y5fsjKEIWj1dVNRIei
TidaLrxC9UV0FLt/QVtyfZfrp29KBSXRMMYmhVrOB3QKc8MrH6iFRReHVi1MoKCmOl3lN1xKrd2J
AlRhTX062AOzBYjnagsi6wNLHVBV+Qy1q/tyhbM7doGPlXukZgCJlPg/GfOJWEIl2VQO/bt/8eSU
r7WKVX/9k0Tkyp9A6Lhprwe6XKje03v0VskUFn/Fn9mINH3f43RM83jrdcRSZPkaaY4tDbgb9x5F
/zj4wt6IZrbKlge6g26XJAELLzGcfb7WhrBtlzPgG1y4j9exjs6SEQPpOuqsgUvn3K9SH74EaRIg
4ajZv7sy6oBQVOwnXoehEDxpUfpH5ZSOVDbSMFvr2M0akgBBq9iyJODp16evdyDeLPXczJgxUHpW
8UTufTbqkn+6xpihpivmJSz9bOAuUkWc2Wx1xAfGxBMCyyzcOpgA0wBtoymcZ9fyYhOzuvG83QeW
TKh3CjLi1UCrFA/wuEcpd8Oqm6pnyvtCbJ4xlptmPOSB1bcHNr8vtFdGGN05ga66RfcAWCc2+amT
XTdQ4XXIoDmZjpLNg839/NFWXGQDALTC/ox+uT0P/sv04AOjJ3j8yjQxq8vOrVyzXpbm2Lw+JP3p
zqAAYm3TyT9D/norvNFs+To3m25tVCaMBdIgR7VevzpQOhVgH7fbMo6thDWUo2vsq59k5AatNN85
iBxjCogrtOnWvYbeKCNFjS1Tt10mN6HkoJUD66CjSVq351/FF2Y+gFjBXv4r+QZrKLcIK1sKDwcM
N3560Jxo8ee6eIDN7D4YhcRaXpl2Hz0MxWVBsBtNv3Gd/2UziD59Rp1ZxIe/PRVU3Aq0UpaoPZ6J
c346UdWq+oqbIABYIJ95kAy6FbMNDFHP+QSsXqkVwKyDixH5FiCH8vJlyj7f62zeYg4hGwxTkg/o
Q9unCDtI0kfmtFI1smkmGLuVP8Vn9hhoF2hbBuMX6iZe7cNX/s/w/qSZFSzO2msHgYEmbaCe7UI2
irEfziLYBc6TQ1k9C9rV5iI3K2Fbf+isGKZG08TB7HdgUghtDGF209qlsX+lVn6p4EbBEbV3gGVe
p9miWbUdVnOyLGIvhjGsCR7j2pQHSoNE2gpSqnoa2wgw62VQ5sfNB6vH9VjW5pG1lNlxtpVV6nhK
ImuKS+nQviQKMuI6ztwV4YGSy52vmP6jFYQo99tc9i4HWM9EJO3HYK2SR12N8r5Ji5FGDobnINah
H0xhuRV/1E2JrWpjnBvy1wIGWoZZcuVgp7+lWaJG99kR4VBvhPyHQqzogmO2Gv5ogUWtte4j/kf0
C81vXd2gkWwr9cFIQXXKXrgGJJkYbsBDvzB5MDiYIEjc7d1id8/mA3drF1OIfQoveWS5OjV5/sKU
BVNLTy1ofTdoWVrHSA1znE9z29kOMmwquSIQn2Eg/D/n0NTdhQYLlvQMj9N8sy8aDKIpKEJQdNue
hjTSfXa/5kXXJM0ImYgwKZWlmyUH40IPyabeXl5Tn9tRwHa1mJngN+VHBJpN9T/KPxs1jQFaSrA2
KPImOez0yTmV2dqVj3IMo9ARL0rG+CEcYkWr5URNbaGr9LRtZMyssvZ7g2g7DyUSJF0LOuXnCxD3
UPmf91N/O3SzYbwV+SyXDJgUQ5FheNShv6uZtKeatnFNmV1Rg5DOkjwd41pQCcFpyazWMFROSGrr
EwvcJZeN5HlC7GlZUOEC3v+OdFwoiJ3qepUn91KsledA9GvALS/vmKrTicd3GP1W780OIe1f4pWx
4J2JIA2iZny8+WXkqNWuTpCJYBSCErA3Ksyk9NR58S+FE2vk6DrayigwEyUsdLOP4IHpvC1Iki4p
IDusfJswM6gOGqupdm8+4CQZSb/2TjuQF7rh2lxJ92WEdDRULPTDXujQ/Q4z6Cw9ruoHfeC4OzI+
N1u5m4tSSrVThzi+GCmc4rWrLunshyBzxRuVriei9mnOutAOImfBJYAtS+Sf8wZsYoQ2DDiy3P9w
Ji/AXugzAFx4myj0RR0bn6C/GPRPAClY9jYIE68jIYJNfLpqmBPU4FB+ElCgHv4BhY/edUuLmdnJ
XzGrthwJLX+CVdl+Jwo/VfeKZmphDNo9nou6fwQO50G4U7kA27GziSJwMM32jh0eHNL909uyWZSH
ZO9+fBCtQNXxAIqb46wVlYtuTpfDmZKOj3y9peHVV08H413RZvg/GByViWQUEA37dyT+5sS5Wqhv
NI4F6wxs5O4yLKJP1fth+YrhYvPBzdHfJAcQQUrHoq6vnyNZcNb7A6Ak3EAOJzVharfniy7lmVHX
boPAPQr4WdLBNF4DZBrqldE7wqHXRSTpgvfdUdO3mNuJObyOJ8PaPC8qbWCunkvUn8d7+/sDm18i
ltfyldJ0OS7PC84hUNj52NnH1ZGpraTRmVkoHetkae48S6/QAXqu5Ypnvxvb0RuTFuKmz41Wh0jA
ol/5FUtqnLYPoYKPyhhh6H5Ur+lngEg5KnGHONafjwrhE3tpFz6exofo/4AOSMBRqHwbqkEWjwxS
/l/MnVUon/Ad1mwDiTQec2sPJr4gLLEfMLgF4+OyiSnnddPrztHTjENW0Up6OiJQullCNcowlsnA
q+m7rdh25+tXYMZ65J/+i4TuWAYPp7YpfdehPWgzagfJ1kzmj/ghBhMoftMpOpbOkUHAfyyDXf/+
xdBqgMbcT4LuyzqSOOw+SEpL1LcOxwCt5Ikd2LtCnKetxbf+QwGzs+642bU77z1IzP2z26fw9ao/
2B4yfGSeUgbA8tSYnkQdiIxtLVDBqCZBPUg0re61k2Uhcz7Z5iD342VIMp6majOwJiNCZp/lhu9N
/L/Lb9UZRbUtABIyf9k08c0CBG0f1a9m2OhVdiHhlh6o3YwTlv2dGqZe0mBnj/Mcr/oHHxPZTzif
AcaT8so4Qw76K5yBJIigWDgiYAEec0tw4amgCYqH6pNUS5jL7JPK69E66MH8cKm95JO45s/XL2NX
/DDlOrcK5Z1b4o6RIBlnB6jSQ2mzFc7+YycgJ1KkkXyDtOx7oVt9NluUVJja6wxbFjsRAv3RGbw+
F4cUUoelTPFzg8vtiU2KJSfc9PqShuZyC+zcw39VZZifvDLffTsbXbPiuxeVx3kR8sn4PnfFzJQj
xJmJd3V/EgPB0tlxWVyDYDn5jgTMYMA84WHnq72GPE/1OCrfM9sdTknp6rKb9/9QWvNQ5A52F/mL
BMuu1f0bTcwYzoyPB7Vqu+7ojk/teKCC9PSqFRj1rkpKMmDWaMN6K4UaEi5zXOhRVo0P63LK0qyN
M2HvaKKkfnVXOoWsz3b7nZILIPuto+pGHM9Ddwfn/TvMMDLhdQvnR/l1AQy/zYAZEA4mfVSROiLh
Jdu6ESvY1Mh398oOiDhZgvxiPs6YWoNTDfmipY5PwsJ4LYuKhvz6v2sC58y5H5c1VWp2xhyTddEn
N/6EU2l6VcRrrqaTtOwKUUz8hHDZERZdv2N/6aLWziOEvNWLiKRHKrH84Payqc8lBiJFmBdSdvCE
Knv5GArofpe4gTaM1Drw/uEdCiHWDKbfswSwcPlzXkOn9M0qdonKecJwzZq8yqSNxGOz4RCgVs4X
B9AZB26B5OUeSmLuCKwip0xlsyaOQ6eJYogZBMaEFsaYjCHh2jy7qebW15c0zEmAaksebS9Ut55h
wdI6G33po7HgKAxWzEcY2eIHZC4NI0cKipEch6TdCjKd5+T8DWQu5YRE4xnjL97RBKMxeGnJqc/P
sgwUm1d1QvTHEy+88Jiegzi2OTKIh5QsKjE9D3LLww3XIoDm5S99bGOtXtk/eisOS0onXPkYOFmN
RDzkOTseiGvEzLfwOP2XSybPb8jBApOtwPMi9c/Pkc4njKFCJ+wkmShX2YgwdwxCDU87ygYcrzLX
fDyFr4obv2KCMg7hEYfsM8O2ONoZLb3FpgIDvL2cMg32tfJ5iaCiLvQfIWG8yYxbluwWIWbZkORB
BL14j+7a2nr/O7B58Mvhm9hh5T3ze0uBtJX/Hw5LVh4iImgBFODwe8lbGeKIcDKjbLN91Rr3+Qju
s4dZNb/ZbouGRDWybZkm07QoiiqB4mPcULcAzkS3WhzfMkEfB0R1kDJp3XEXWFKcRNBc69Z13dpi
AbB4eXEyOX7c+T0JQPd/6CcT7ERPRlmV/c2mkwgdQlld5p1XDpuUXwMJnQM3S605T2Gqri65Ep2N
3VsfHhvm9hbvKXO0o7CSZKQsNCVRMMMrSnonbORMl6oKfo3lYiC3oOQCJXVxx3moWtH7NChUHD8c
EgyckMI/Tkvx3Q+dDIKpBjmOgyWOZuhAY5pAVWMgrSNLB46Dz6Lh5cnp8T5DMlwQV049wc4wCbB+
psAcGkN56rOjAa2avShUnGI6F4xpmxb4iLfL+08eMrvTiOMazOD77QaOo6GB5bU+euAIjK1TAdHa
VKsu+EY7dVwlcXvtB04Br/uAPzAYGPY8vNT1vMuxcwcuJ79cR1wv0F3lbSCUqxoc2wslvvIX+vP3
2SQVm7GZXlna6rvG62ga5AGNcRBrZZ6Tv47RY12nAY64eJvcRhFxjQ15fDdX4GYD7UG2RpbiUwGx
4i3RTl6k9bZ8cCBVKh9EpreWwHQ68P/TvepWZuGxcfgsS5SOCXbuxQ0/d5wiIyltwevgjpvk2MGY
SvGd7NtEuDUDa3vP/oj0dITb9uG287bQguFyd97hEgHAWwhQlqrEFnS0H+S6aFzuFrj9GtBppubH
3xeVxn9ReS0QnwyDmPVKSIh4qATcGg05aCG8eUrcp6vm1kNUydsA3k5/6fBcUDpTLhs1nx00d8XJ
QB+/8EQLu31pObIcJd/PF9rd5haDza1BAw+TYpbEMU4bBcoBZWvEwvG2kcANpGptXfQX/2cXwQYo
NE0PTc8krDepzu2VSaSztZPYEOkOvOM4IMP3Hq/iu0XQ0dlH84Y0Rx4p5iip+dT/p0iwpPhvqQ1L
xkvWlFgAvkBFYoi9w+x+dV64GZB1+1spAJ6Q/FlJfowHNf2VM4HxonjoFZ9dCv4dk6Wj5ZfTAlji
1ZEscZLblr7i971she1IBBGWDI+e814EiEWrREb/j2fGIpqWnkvINQQGwfwitPP5dvLWTVTaKm8H
/w7E2U0R7c5VYhMVIdGSw0uXzDXJMbZL/S1+iD1RIU5yk6/zbbHE+4+2pBc1Xwpc0gz3Zx+FPqlu
6YNabtCjsFaVkmLKwu/tYSJ0UnEiw6HzD9FZ+CPo7gF13GjVwZoEWViLneAS4lxR/xSdH9QR02C6
MMjRS72O6IDVY7MVXUayMU38GINGsgJkXIu9AFGgD4Kxxs7edwr5ZQjxEdHxOpmgDUfURXUZxXUb
WXatb/ADvDJjvdTFWhpQFPmEPYc6Ix7Pya/67Mj5UEW5itMHFhDa5e9kvkFfBbwUGayD1ROS1RW2
EWKrT3P3+iCejP7esAAvCMLyqlOpXsd+kwz/u0VsOWS1Miw1ANq1qp0qyZrrhOHK1nHGFmn2o4MQ
BUw6KPGk4+PbEtuRcp+zg0Bmbn8yJav3fWtUKsjxgDt6PF5dEGQYoNUSFUkV36xdGANHGYakkfGz
ek/+KQvc7ucDO7l/35v+43yERfxzjkvSHV61sTMg9c7mpct9AYHOi8ztSbJ1PHOnjxaKOvHcWwRc
ssFYzroJO9L0mvJfK4FWpwyrjuoDRJqPbeImPCB4vcwNN4dCbbFFhuV77XtLrJ6LCuueut+rgUB4
mrotMY7vPEX4cxMC3TEdGVZh8NoSiyh2pmXYez9Ch9oA2pCB/wYzo+4IhIn8C2mGWmCBc1SqrN4b
3SrmgoUmZswC3olOSAhiqhtgBgrnVTk8e6vSvw8vgeCiIvJ7jxopXFxvIT7QcWD6GLCd+LO6tKsk
EkFWnOb8HpCQ78/gqubl+iuEYQC0HSy+eJF8qhdaE0f0NrLd9Y2x3q13Ppu500jABXIzzoEg/cIK
Z/IFVpI3duuKzITtLQGwR6/DkkRa8KAZYlNNLw5aIYYfTdT0XsM7vJ98st6r+BPAUHGRUcdbjf18
iNMWkHUywUy2yB5uBO2us+k87FpXvMTPHRUF5HBOAQ+cQHTDQWUoPq64++MWWhlq8DniVRG5eHac
L5dyN6l2P2bWEdJrkIIh+9q9DnPKzIG9TcH6ql2z3rn2tBgByozhkb/FnZ6k+0RDvRCVIx8/T/g7
MWkIZHIA+Od/SW9Lzk6MfCkJ4rbCRzbfha+jFMM4xa0GdXPr8px2q9n7rQQBDLvTBrrQvmK9H1xn
diQ9EOg8ZtOhMwCm/6H+ix88zo4FVKxqRUCNy0ydw9lotwot6nJl9fax/ZSmuAAkRIqBMP7zrarN
IjvsOngrC3zYVnW1QK6zHR4PVgH7LQmQ6cXY4OTq3Dmu9KDTr/SPm9Dsvyoe6uE7gEz/JgOIkVwS
EEqomiR83lwhJ3r1MFPcvlRRWmqzkQhLorvIBQIq5ox13cUEiStYdYGi8DBjYkyPiMjTuuNtE/mG
4nk2trYJ7xbJE1VWfJNbUJcrFCNw28HzD6WWc2EJbsBijtuKcCJwSza/LmuX8XeQg9hg7Kxv3KRp
VeQ3dHRoX7VI8smz1gX3MPgPeQeX8UUNPVgieuRawgteseJqiEis2bMxIRlBkZRZxImZFcaBLfDb
j375U+JAJVqbocXdzjuLYAc7txoUWigGwi1upabqL54U+CyjQb7HTTlwj5C2UkL+Bjw5ppmQbIWQ
nPLPxLCCCkCi2fec9qF5MxuxqS8JygFEEpoXr0hy9eYBs0EWLil35JnKmGmdIeYjhABFcL3f3CIP
9Iu5YRtNDlo+eEN/1ljFp05Y4L0I/Z9NIlmKdTz7OF1XQ+Y3Z6FgbDjPos+pHu8W0zWKRKlBmMKt
UVtGqh+MvHnXBXLgFVqwHg0xm3Z72ID6iiEyWTe8K+LprzCLYVwllCJSs0KiqIYeICg2bgwqP5Yy
R9+XeHmhMndaplU6mCLql+Q+NKwaHtN+bsDk6WWD6JTS8frQIlXGvAZSBAktkWW9z96z44FmTatE
l35b8iK69ljyfox8AY54jNhb/bzZW0lFTRtxXNCgyYT96BJfcIwVmJ6hJEM1YTkpPejnUAbL6unb
HBurV8QuVlYW6VdUQHYrhVi0N1Gf448EyDH1X1uqLRkhPIoID9zjCP9h+3qXWDrk9cpzONyVNBak
HeqEic4zfCihwXtJH/PvVh6prXpT8qnEq7eAQvgpEg27MRSkUbAQk/pD/ASpCEFwpoDsbXbM0N16
6nGrxNIYKafX+1BVozFyg3CNKqCEElEmRcDx7bz3U+Glg3447HErlMi7ea3mFdB1HhpsOljUPd1t
pt1qHN2e5zSH88lTvc6RjqAwz29O3VUvZ095fs15dW8LjuBDIW4WcsH0Hd0VIoBRMXbjP0hp/sBG
Asu68gjaxcrMGWhhzXt9X6AGeDXRbu5VwbAo+57DtfvZW7GhITA0CO/R1TyHMZRVbOHPJ+eQWEig
4fv/lN22ZVCrh/HVSHbCtDIEmkaIVXb/fX+AJ6IT8UnAV6kFjMCT0uuxsLIOJaR8Sd7ugMGJgmDL
24urO03d6HQ2LclhKJBflBQZQZwDKvFZb1fGkb2LHgdfwKAycRtWaCN9oWxHzs02mTa/cyHfJBZG
NJRIRUzJjgjLAACuZB7ya7suUkuSYHNFHb7yqLvZ89ZQUvLRt9f9DRTKpYoyqVkDBdWCkVs2zSVv
0OqM2IK9BeSuV5m04a5WUpnOfyDG0FcQHdLuY8LPbRHfb/EK56B7dY76ZZr4ALnKnJwy/fGjRsE9
AapXrsilnew06vAC6r2tRLMfMq6B2+n2kUckSPS3CMnjDgsFg9DX2xrY3P81UDx8FTSRzwc4ARgs
B3Hu39XxtzG4RA0wOYWiDgwUqaM2Eh38SdJEjR8e/AQdLflrWPQe9ruIXCL8B18gJK3jQkJ+t+sG
cvIXM9UtGGnAxfrKIjdO30Vm0GhQLoe4I0jVfIIjl4bS27ukcQ5sDJTnldtCvfTXbIUSlr3zOmrm
kPVSuAIY7B70WkoYGDvD3DuaWsbypnh+uENsE1u38X+ID44oftKJqtuRtZcZJ14dK75RTQNA1RrR
UVk5ryru0NKf4z8iemFhnWQaA5TDu6vXIacBksZ7O4+vkouacm7+vPe5VvkHkMeVEptCoZFxOHvC
JWx8nfNqygW2lMNMFjqyShRijlorip6wXuZvatD2RzVVbw3vtbrl3feo5UuiJLgwlrQKU1ILE5+T
0mDn5+/0fbQEjE8x4faBAZ409/EKj5CzpupKMjMTSfqJjkBw3GOrTBhO3n1NoAOotiazliiHshZs
DH5AyqVx2HUDKpBVYqhWIhBM2tWn5Etp8oVdlrIjRYxoKCVWs9esz70FFp6G+NOKzltVnPkgj3DW
k+PcPZuP8dheTG/aWmmRF+wzTO0tzxQ00Gl+XFDQpPJVrCYwx+YSlt7RBM3edzQWGOirCK1HRdFL
lL6QbZcutgui/D9u5tKGbR7v5wH06ppE1TRuvfs6qPPrTK5fCrGnRF1hpbIbME+Lq3RBZvzohgZd
nQavPobNDS2QXviSGEqkDY2UMvpPmXniTFdVuf3m9BRrVuvE94zl0w6R19KDBv7yLGO+u4wybkYg
yzlm+5+FvV4T222u8IaB7UYXuluIjglJjHsarNGYfDf1eR3PoIQ+6a4e9ru/aqsof5PJGauAlbo7
RJ6P054UEzIcURB7p6s1OgEVegyFYUbl2T9cAonlhca/LfLeMfskId9Z4i77tJedeDrfkH4tU+Em
mhz9HUglUIyb95FpV8ECJ/n8Z5wQkkAVx2e8B1vAZMIYBVZZ/boaUsv6ctsEM/U9QErpy09KAQ+a
hFJ4u2xxWJv5X8a4nJzre350EWGpWWXbnOUZID6IqkiFGPxuJ+qjXNvtBdcl3ZcCCQZtYs5C5iJH
HypbaeihRIxwC84nSQTBiILv+UrRzUGKn18ybxhQ+RNijLg6+zBy9faK8dcr7TSKajfsSG3552nq
3cJPj16glQIDe8NfRsQUPTpT0Lf6ixqXsbcFnH2+S1f42NE+hHTlRac9eFlK4mPFfMwBv9yfVq3I
mhGqd+bou+GEjzRYpPigy7usZT7oKEkidEXRyqKNz0RIO9uWniZ7FXZiMy9zdGn4FYspTMIFRxb8
U9i0rwaAJduL6MDfQM0J9Va90zIkaV6BkM625/tdQG7eV4qVOtLysPnz7Kawi4Hm74+kNwEnrmRf
4+eVAWfNxfHTv1+uhOMBJg0yF72ONGDLaIMWlJeTcF1/jqSlggrV+msV1+0Al8ulg3qaHif9oFfV
S3s1qVnnd5NQmaXwHjVWZaK17yV35fyLFQwhaHsCvGf4oLbmMyv4vnrLXpC84gM7/6jcV/1zKUwZ
D9smhBFweoVQi2Zv0rNNebySwm4xjR3IEMXUbtznSpreaULK1QUN70PEC1WfrKI+TBjBLeJdYq6d
oAABV2wm1mzsPzKcIHbF3Ph3rcV5eUb4fJ1ytkPLjRTLrg5CtE8m11KPIp1zhBdbTiSOXHuXFgHl
cE39tuHqxrPjfyLzhPZmh7oJYgMhVfBrrzDIJHmNwoPKzT3j7xYimhafSvWwR7W0MAllLKBnERbz
v1NvuLw8P5wh5aU+w8S/8QGzHUn1tVRuHraNlLSRSItgXq0Q7LA1mJzqOgR1dKPNoiJnEz/Bj//8
7j6oKwN+fJsw17weHD32XbB99wubDbu1GyVn+3/e4XzMulBF2dAOonCjpqPtnKsbsRJkaw0uHg/m
GEd0lWiTHYUDMz5Us8b41jLcsZK5Sr5qU3oAwgMESmklwCiw/cv50BXoyf9DjFPujPWjN0OdwXu5
ewLRkkrw8/Qw+3/SP+cAdAtKgCaoMQQ9g9RNHeNa7UH12ZmeUPiF+sR//XL9Aw8CuLkMkFUquE5Y
5CMqjzDRzDawya8asI1mwf+sFfzFOxWK7LyGQDJj5l2l7mAzolJB1wM9QZKsDnJkEfHCaPp4S0kU
DQEqdmAjiNgOhMeFK6+WUUqshdBLQGHuIM3GEIu9d24TUecHDfDwVWUukpzW61ydc6h8e4NkZowM
z95K82RdxaYWLtiFupU+8KybTGcH/Lm45tedOELclNVEsNQ3Uvqxd8s0itt5dn/Ojo6AAzxqOqmn
X/mQxvR2tRrdiwMgjK8EPfk9LAfII2Am4aUIWC0iBW7BY6LT37li8mMv0WzGoBgVJgKopNc8trTo
zGFji+XhGynHC6RegjcSIoqHWF75BtZqnZnvnES/5h1dfdw8hSwpowV0hkKMd+i49UkHdMjAUr0a
9PSNtUqy4N2AwdzxD3G+mFwJNvcOTyT+ZdDCC7yg8lC3T3wp27oAHrkOBsfY/GJCK15b/s4mQVhg
e/TUaczy5pAZVC760EXgXYZJ6ECKCih32LTIg687p+cnstwOXz8/NNCfYVlC27l0QR60EkcI/HhG
gJNPkvH/eEUeqtqMj0reuZFsum7HjgUgKmTnyiTEVo8boh/utukeKNfYh3wsBnvg61kW/fVYIQiJ
rgaKrie0EsiU+hbwqjp3C0j8dnsIk1KPjHSLc6wvSEj5gGnkFjVBoOFJuvxcNFtcnQCISku5tqR2
dO80YlA2PWI+B05rjSHNmHJqJRgqnJHGQT1akyaLSqEu4OpsViVDmRdp/iqr2SLeTZ78X0lgfLqT
Jk/qjePEWWD3vAuVjkpuSBRh/4ZBfXjIDAwgDHrduN9CaLKQIdCrKUgXgq206vVvn1YwxxZDw5z6
brBYI7Kcl0EUUvcS6RNMwDqSWKSS9GiGBMjnKQ2f64kQtZe1vdW1EL1vMDVRMRwK2r5aoVpkXK9B
K1NLu7A+6okwkf5tk9JYytXmA6jV8KICEQPeFFAS38lSpy3c5vh9GdO7ZL7hWPAUdKBs3XeCdX9s
nstvHAa7gruLa1T0KErQlYOs1CrcHBsf9kfxTwW0DQQOKCJbbOPzvHox63rrM/0wht9mI0yx180o
+cnsrjjoZF5ML4jd1VuCX/ZH4auk26TOh3Aqy9hPd7ek7r6J/PRBAuufiBfAQBWv9SgUe0VEz/fM
UvXVrXYaZ1Q3Pb7Gly2dq2afrLX9qd9QqeruLc+lBVjl6fJjzSFxAb89A4oT/p8696xlZeet20ne
29UT/S+FbTEXL8/TUp2iCHIvtRtDt5IV8oAS5GRjf0ZAx7tYpn/fTf0FUYp5lWk513CAWCkJuTnT
ckIJKk1s5O/bkpb8U1FXhJiyJLvdGiS4FSvUaFtgi1wiEalfPsapKAI0b7tPmX7YhUmaQtm51O0H
Rc6IU2m5EvG95OTBdekbv5cDN9CwIyTWcEgD+9NHyxOpY9W+2vWCQ5Qtn04L9b0+//7ovN/wQrkt
AV19K52ZXCnrYFUlGFzKJpKfhjdY8isLTI/8EB5idLjXeGQs/iH97ZiuRN9F99huD4VNCpnUnu6C
MEqiDkXn2epWXd7nUt1ECry5pMIETxHrc/dac4SdSoZLA4jd+jmyD0I4mA9b4ACVWqMa3D3ADM9V
UMSkkLlLkrcIwKuZoLPL7yu6ja/sqV2aoAvzUElZiSoJD99zhdscmHiXw985vID7ycspWZ610yc4
CUwalhrfc5raK/z7H3+w6JiPtblHwgJWf0rK19e/csJ1MuBpsTFjP47c9kn9wKf9YtMIToa9dYZa
2BQjg9kD24cMl1Um/17k/vlwzpoKxCftDYmJaTG9894Rs3IjK4bg8pAD0n/uMgwBoZAh9ixyfg9J
RnNiFQvKoZestqLNIBD/vYgN19YRG3I/dRxwkfCMl3AMKvEHlB7wFLDLtRd4yA7InmV9mF8nEm7V
T0k/FWQTePa9G0HtN9CswBUTYqIvqUWXVrqXhTFuOHSXlN0o3ymsvfR4R55crSRuq/Nmiz2p8LWe
jKMLCs99pJRNezU1or/oKbof1gwEdx0wqmnP8wLFByNQ72y4iwsVbD9A+JW7Ca7VN9OWzSnkgxht
yijtGDcQSqT7rqqjXVMub/blU3J/IHvLyFZgMigyFuhB4ATwzIy7h1f0oSrs6KR7OlaSvJ1Woxoj
OlhqRLojEFaW5Ez++qion3FR5HnkC75x65xUH1Hao/btrgEnzJX1z368ulHEmSXjxZoVgQTjKm/1
mXLMo3fRyv0+7JhxiUUv1yeT/fiG7LszIKT8quRgoGV/W6VLUfubA1eSW4sxE/WMCqdBzP63LwZr
QbX5fUOvhywJa7jc4EHWwmdScA970pi2xpPBrQ3XNmVVFYnAjKDhdHuqWbmx9Qphk/ZoyznYA+Tu
IOsqr/p3kVY3tb4uinxmA2mt6xEQz0prlPKDKlIZ8blD59FWoP/XBvHh2D/q88ymUoV1yi5JmNSi
AsXBQZ/l+/S/8XN6Yzv8SqbeZi034FobsW7yvMIorx44QWgndLXR7VCHDSQrq7UuzqIvjXGbrXh2
BViDs7WaL6Vx9DjWNnxd5TSr+MB29LCktuYCDkrsnuYGGUopKlwseWZj3oYcncoHJzh90gMlJyyn
iB4V9WH8BQhpKUbubMVPmXC6U6ywcmxCQhJM6t58bK9j2pKjk+8bGDwN0/ACu7jVNgrH10zqZbMX
QveczY51lzoaxQXtAXvDe8vme6ehj/vjTCFwV1+P308XvESPplzMMLWrySg1V2XSUpfNsygs1FoI
lwhrKRLLZlLeUtFWoEwJtHS3bG5IMIFW3XLnHYoJZflc0I90jFw5yCbZ9dIAMxlyOYcmzBKBC4uK
puBMrWnn0Lq0YSyiIJxEbCFKphQl3otUq6O/1E0DaIQlQLYmhe/YB5tm10qSdeb/hh+vxJ1Ic/KW
2Z+Ws9nv/IRlMtX1Z7G/TXrmRXINY69MvOMy0GY/BdqphviicTElXlTjVhctOkF9zpH1zzSn/RHV
pDk7vkrnUHB0fWzMTGBXVQSmE2H1XhcQCmvUDxhVxPB3cWIZgqqDSC1Ql4ZzLF1GnAClOTpcfncR
FsvrFey3gZLZhrIW5shMHEQme5crTmHFnI9Xlq5MT1CZCIpqOJFUAV/UBI5RMXxwqiqVCEvN/l2q
yVv5vVjwbsYSpGk64U05H8hyyiwkv/pYPthXf3KkKbZP32J2QOp8OjQUjdTLSFlfypaMZwR+5Cgi
Fr622stpLrzmZeyrR0Cvj/4CpgS+MOAoUS8o5dotkgj+W6Irl1AskAHsJyy9mPTMSblULjI6n3S9
wRoJ951dN7k28Af+RlcUBYblTLiMYhoGqX19lRgNVTMRImSgUdT0uR4fbZB6IiGIwLsZRw0nbjQ1
OAaZYWnfU5F/XPicDIX+xVUHpeqvGEhKuF1xFm8kaIuSXoWDD7OfTOlzCSbwZoTiZ82geyYGM74v
GmcYAX4y3LKvjZfixhWT6rMhv5xT2S8WB+y3F6M0ou9AM+RiDn4Za+hW/uv9H7fBkUujBvAHbpxJ
cH+xJMq8r9Ms6UNzhSahp6EfEzDxNpeZdHlL3QzPHrJZz5XLYc5HRIu/BOvR+dxjMRkcFliXE3rh
V2NSnSniw5zDQWvtIsmYzwU9E/T+RH+HFnzWQLB69rLd/P5nqgCr9pRhG3c2IPA+2k8fm7cwsYGA
Tvwa8vncLQf8jiofM/AmeCzc3juVJGJu+D9AE2EHnfJkoVMuRBNB9s8HAIK2nwJN0fu3kCczcAIV
Lzzd3byFUfejeTbd1O7R+3TJ0S2/8SLtLExE6nMyTp03cG6p7HH2jgGybApaIzbY1FHruiFjV8qG
e6P/YJN/yTjSTLseYdETZQmMqZXWkW7NZSLsIGaajIRWT4xnJYC3VQcmna1oM8T18+2+FKdoAGso
KX4KGi38AGOJ5DxJ6JnoUFsZ+KuAXTOY+yo00MY7RhQJ8stF4ReExXQViVg5C+ljJuZ5tc9Z8lPL
ANG0mkO+he4ecPKYq6La2h3n996Xf1QRej9taBHKlyDIce0aLziGDvTeRFNAa/r+LdTXqQeJi8OQ
oter7Wb8z8wCVsLjcCgfK5McUPm/VeHYhdHEVq7tw+0cuV1C4aY9nBUqzTHeOtRkR2DlO+zIUWzt
F10Nm9Q4ccXQIUh6OLiK6Sd3+GhZBxiLnCIsZmqX1z0N9HhQO1gZ/XfbALtkuQEvfmIpqSOZMwFV
RBZ5seMbK+B8VwwXivLZRqf2xHAg8ENXsy+IZQE+Z7ISrfR1ltcL99hri+HCFvX4paOsFg4x51hp
rKDxvgBS33UQSDsLQQAvnc0Uhtn4ZdN6bFhoftgCQS3Hc1oZTrGaKa3/ANbg41tf23dCs90umFyh
E38uoPS3PYQ1iUoGUSxXRg7L/qI81LHTbMx4qGKxT13c40u0cgcC2c4273KmHWhZloETQeIEKGfe
1hyWc4Xy4Lqr3RCp5AV8028+ycnoHpjU8OA3SqMYTR4xTe+SeTDHvHyqsldsy2qxigNqM6H6lq7L
JC1kw16EJP//P+pZ4T2ojTUVwiR+j3PCG9DDwzljYystkKuEdpYsovCTaN+7QI6RmGf/haBv1yOk
eHQfheglzpgILeNM8iMqf5KkctQtnEo5tRpHeJ7E/zmF2SOiL2x8UmAJBTH3N/BB/4bq1pDHR8oo
lVUT+7qSdYDq3g1asvtcoFc79qfmxDO3ZLU450yXdFDAobthYOScOHf7YI1bb7JCHyI4v6Uz4NOg
onHhOuO/kv/AAYy9o+fyugtd0X4XInR6x1BbMWLjvUBGkJfCLbSFdVlcXDf00XyvrCDbRH92yAGb
7NRDaCGztjX8UCIqcXhCaFkTGiTqQ63Ne2InpvejHNaIR3YfQSGdGRjHY7z0Tu2Hw3roNUpB2KFH
IVqwq3VnnTRxR/ZSxk6EsWA/9jIYUnyQP9r6WzS51cJV+s9Md4+i1L6RSbSo1Lvme+80I6Thgi4a
BQigKMEZ4IYhBnh8xnAC3OzQuqREZI4dgqxA5mXh6cPfIeQCJ0yh6inAT+tlWBC9ovkCRl3WOnRy
omWH0pcX3wpC9x6byy/TxeFqPnQflolp2tePUPWGxuZ7S4Wc+mSoO1NQRDiHJYjgwmfUz/dY46Lo
0i4rvkRNDVGYuQ6Xg4p8J+VSKRu/n8RqV7r1sLNKaekuUDSJGPCS7n/RQErpEW/yev7tYYFdGvDN
pRbcmQQKA0d7DUEjznYnTk4e2pKaqJhYAw7Lc/Ue0c/fbr5gdu34TTqz5Jjep/H/hP456K/hBd4D
DTjsJ926cGO41tKQi6lL0KnoZcXyBLH6gq5nz228aR6E2moRT+CcO260F7//rSQnfqSAbR4z6+YH
EgVz6M7imZtvuFw7T+MsJxfD16TW1NQHdiO9Mr5TpuUFUUhmiC+Ytu4aXl0Wn4hKA/zXHMgQUumR
EMrnM6wfouRBIhoelUbVfH5De5pSnKRjXOmCedSCNfqmejkmPVCxFuB5QGFXACW9WeYn8nNcLvFM
iD4uKkJqAw8DNkb89zYB91Kfpbr9xB4dnrDyCt9Rk2dQuv+f+abbbBfo2bj0Fp0tlI5f/4/fzbIf
AxG5M3WfgWvmMDPXlc+edajY7Q8Muv2522NkLVSv0qnt40qad4UAWgaYqalRTW7cJb+6bwKcG6jA
EuzDBfQJTc97InCcuPixUotv4PK3xeaINbyVNBkOoahPdybkSt1vt5/F17gXm+fJBl7oa29TxEy9
e7nIqxXgFngsg3YE7dSuRVcrDqIx8J/Ky61mi6Rly5usbd7E1jRM26KVJYgMfp5S2WnGN4KkN/WW
xyTpE2ES7HMF5oUaNmYnFHf7T+ueA75SPjP6C/tQr2WbWZPdqmUsMIuYCezCM1MJ6WdLZC8nP8CB
5LF1YweknkMoCgV6SkXdl+Cqb/90Scmg9yzYxFDhZPjKz27Nyrn2xFYqR7LtfPSCqLY6xq7XSCo9
27vgoZBCwUnpO3nBqW3YJHmPQyUvM+sH7BGALzM+NgBuaUG8oxaOtWukw/0qe6JKzx69xONg6dB5
zYt44X0VC4pKNZoB1nNMgKRJDHO1mA2T/BtqCAnRi2R7P0P3GQ95Hct749RhM3rc6UFhPOtVzSAc
lBSeMRxizNY/6ResRt2mlzAqS8l0NOs5vQUKLXdsuZwCZc4CYe1/NawGbPlIm0P5RFwf0/n9vdJ6
05KkCXJaIR0oS8pV6w8UYGsiL8TGMwDx6fuQJnXTDT6wp4kFaQc2AdG0OloCR9n1f6ql2mR9PaAL
81YotchgpreeEQ8KbxG2yg8L3svoep7KX8lUuofPUJX6ZS7oRpgqRQO5t/c1HM+rpocFxESvRqp2
VT8YUqvQWYxZbFL8PY0fB+xYLKJLp/vPs6wtYUPD6+NUze3dC483JDAQT8ZktgX+g++DWTd9ZjMg
l5E8CI5/BJo/YiUiwW/sITHiz7flrkWsDxwcNgs26z7RUpCaEZ58dpC088ewNOUNMI2CmKaady7g
MD8udtDX1qMC+ST2eeIMV4Sg6oAw5hiLYtGITvRm+0h/bDwbS10aeN0L5ZQ1lquL4DroWmZQxTo5
c38oGmcxtZMV6sM4+ZKLOqR4VjwfK9JdPKx+FRxfFB0Y1nqgayZMkHcg0clKJ4a4i8y8RFm0Dg1M
5Qn3QVMn8nZYPUj2VmRDiTXo8fMDR8FPfYh+6OyPwH/1+nefOGb7oyWpkL/SCdwDg2kXiQKXki6U
ezxtepNPXvzscLQUXc9j2F7VgHrySts83dQZqBWpR6xmDQb3li8O15/uslNkPJzqcw6ju40JSM3r
wCtsvtmlSktshalL3H0CK+saiOpkZaukvLY9YZ4XwnNCB4tZBNbV9TnLCfUqMMufg3pyyRLA2VAB
UsNSYD+S7SO4VHWWtX3T9k8FK1VeSsQCFdXD2+PMrp9iDE+xvfYLaiqLdu6uWeqLyJ6j/ADXGKYn
KUPeZur/Oprtmzcz0GacJyP+QqJCukoctsAqmKqmVjvqvXLnlWWXMN/WqMMgzeDC90jtn74c0Ahn
diPBT2Fcykxoo9E81lTfFKWNd+/lWXae/qMLGz3XWMSNRkfWNYVv8pCxWMgUEWbqscwcq/erADpf
RuSlINf6neCz5iVBZrM27Y/Ch5W6tpYeOO2cwCGsEkhs5BHynmDP1TbMzSOoB+6Gf/KKpl+c8J1Y
GFIy6wDJRXx2uMtA/wtCNh/bD34Blq3L6rf9Z6B7XTNSozEbRlYJFQSQPwOaAF1ij2dfbBotW1Zn
Ri8plgkuidS9mjHM+96zjeh0/cTBObO6aPcfOu6/pCHKKdFlilI2kBFGDUFx9lKNiN7S340KN0wF
xQULV61WqZQKmb3CfbUd2HDyZzKSdjHqMPF6lJ46DR6dCzi7MqrphY+qaVjbldlASDrkfw1nSvxC
MavjRpCWUWsXG2zjiLFcc5kaCpu5vuqDj7IaYP6lLT2wWOYXIIhY5fsoYm3zfpx2lzYnQ52g2LCW
k7RwbhjCnlWvmBb4utCvagVLUCycRJ+o72UqEkgFKZqInJo+Wdj0D+WCVsC8qV2MZy4w7Z8lQiPC
NyUmHTZ/Pvni85iLjMtbcx4rXEkG90JCAOjCLx5qn55zoiKwoQSeuMDob8RiF2Uqlrg/f6OE9QOm
uKsMN5NDucOlJMI5Gr6QEJvLP8WFJXbSzFMgpAMdg8OE/mnIy7GbvvX58VQjrqngmCnQNoEJMc98
LPFb2XYpL3B1tRG3QMnswo5tt/zQLHLeSbvVRktppp/FtS4RbBEuqISWGUPNo1AZpk9OZ8ZEwy7g
cihucjdZDv3D33L6eVhXlh8dJhRYcWcVtdtaxzfjj1cYkzG8bOL+fiYmmpBUdB7AV68LnSXptthQ
tmgYFZtPhULtdV7vPeqHjZLIUhGrfhrvPzU7hsy2oxt5Un9AfaqOEWPW+ZXd11gs5oCZ6ayt7kL1
z91LHL/ATIyby9K1CVzL8Yjv08r00vrwCbv+I24dusKQd/r2mg819WOh/3ApnD6g5gr1G85UaQvr
eVKNXAEfBeOzwlL6MtXpbcDXyC38W0qcjp642DSJBFnD43ncb3kH0Whx3k5LSlBubSb2cKWsV36V
WQsFBJFlYem6RZO088D0DNYFnz33g/qBtM2lZQIeco6UX72uvGeNpwE41kGZzqGW/zmoYpL1Ze+w
gfsrBJokgGc2vcggmEnA2IuNdAgZ4VZN9O2dSEEkR8MbhILKjFwAailk6v+xU566D1nDOSUc6DjQ
bhZcinqlWR/o2kokfKkvr+XuXtwEs035Nk5WFNFFZ7o/CNvatUOw9yKlGVXep8igCzI1SIQJQFw0
Z3XuI0noCHU9RotdhkIXp0Zo/qMR30NE1Ni6YxoT/JOkqHjNZeeXuVHGfk7KKNLZI/La3uV78Zwg
ZS6LJL9V1JQ7Q3TN3ROGJlHDBx8TqjS+fDp3Klrfw08mFtNRpa++XVDXOGJWU3MFLj5FU/geqUru
wO2P/+9lIRMYDPHSJN9MMUYWfOz3NQQZR3lkvkOiWeIpTCAWHUxK7GZIZ7bacEWKV+pU/0gYHpf4
CbOQtaKzKb3s8zSUiXbtUFxr+1hYnIXXkCDSdHARcMBJvWK8P3smdnC0+3I5SSauVzAIy3u5otzk
JlsMfXSeiE+/FTL2lamPovLztJ0chY+k3mYTF7gOWWcI81l63YlJhPLNmvLHbApXQZsAnKizELU9
jLv3F2P6uzht8xF/KyQlPiStBWvu+vek/rzTKlzZYS0KALeNeHObEce3g2Y67Da8Ycj2r4TAq3VT
dsovgkA8sXeqdKU74SjII0t7//JiT3sQD/vZCQbKcjYQPURRogEFidY2qK8pUemhzZ7WqOyxuQxf
PeH7TUeK35GyqhKh2LPS2/nIwfreJSsv5wvtugRDP3Px20oapuqRyIVyl+H2asSWDv6wfVu+CuxN
ZMzSOeMfqASQ8IYcZ4b0/ozzfdI3j8owerRON+feb1NDzyGaqn9UkY+D05Y9m5hzD+6jmNXbVqby
G+jt8bxkTWp/+84UMpqDGliGkJfvgcEySHJ5t27Wx/QaNe2sJZMlGYbqfnobAUDjMw71v9M4SVfI
IedSkmFAYgEEExN6YQ0QDxurSGL4WANqsEUMAMwUicfEe3yK4P74cp8QuDx4E4Gi1b8lREcdaHOA
RqZBXRxPaogHfoBA6eMaJjzzP+P0kRLu0EU90ME60xPdH32ng6hYSiomjn1knFq4P0z1dFR7wfkJ
KiCGY7oebljks9FVKCFbSfH1Q4tW1sg+H+nD37rNz36mYFUYA4O34N5zqOvSf6tquXIE35Q1VtEO
Y438Ry1Q2q0ZpU8MrhCnRo3GLMXhmnmjhkmGk80K2DEhwxJ3F3P5iAIjMZYfuRoR7m98C+jVHowb
eBILMv5Ng950KyIKFPJaAbhYosmBDjOFrdWQgbJ+fMFVPKZRxAnFq2PD8GSvQwd3rYRyVuzheQ0c
m7vTPuartTlCtI4th7PiscLkm58wi4klE7VuljreVQgNsvmaLq9CpXX3Ik13qL11+jpQIqO6gR3C
aE+Kaql4CR4rK/FvPZyKWtTFNPmpQXinnbAHvKH1kRCCCSMCF9ZUlHgnbnLjsWPkWcQDc8MqjoZS
IGFcZ5AjB3p0U7xwPJ+9lgMTITazfybpXCij766Y1k+etswJCZ2khLXvgk/dnlh0zy5mTTbl5qCk
Add0VfzI1e/UFrv2A6oNtemrwOqwSt9UTXUBYQSuQaK9upPiY8HJt9yAuj8e3LEsRCr2X3hVV14w
Wp3Ms28v8vQe0rGgob1sBGAhszAKaIs4DiTqBU+/RmhWX/emIzpSs7EtDRqyEo8IzCotlNMFUo0+
qhnaNccJ0i0Q/lDt/zMNR703UQ1ONldSw/WP2Y+8YsRo2qR1F1zoDOO0HHkLTd62QbGyYNS0JrVR
Ll/Sokjj026lFOAqYc9zIAqgGbezOlTj2fYmgUyTf5Ufkd8gnaFT0q+R1mrjgsEeZGNmuXc4xgT6
Z5TR7BE0FmhtBN3heeS1GAddvuTXICitXWVIFM+qBkG7xo/TGJKex19tWazOpme86aTcjEq+q9JH
99D2GZUmm19OJoH1qZNH49eZUJVnnIjPQEHTQ47actxrdvkGoR9I0fRWwifWOwE14dfPMLuHilTs
l+P1DoyfZMdWtrI0A/PmaKbcbhwJ/YjK0IBbs29NH4+snCfLIy7cn4Q4zrdCrSVAhF42qQpxzvNi
0jJkIR2WLfB+01SwJwoA3AHKXs1bsCJZZmtYMCPS/gEC4LF9uJDjHCpvTJFpp3/D9ri+cdAvlsx2
DtAlk9gZdk4S5UnAhcIqfRMaP/OBbqw0QBy2xU0kmxwn6V3xeGpO8Kp+yof3HotnhIs+lSktAh1R
+AHg9+pf8+mFHx3J4tCJUxlUX+6y1JrkWuRK4PvT0gO4CT4ulFrFYBUtf10QSkcHLXAFiSwv6IBj
0jpNHVLX7Mv0htaMR+Vg0R2lxWIeqP3Y5mT21SiMpTYQUbVdVqrk6gcVKto0crZnsLr2KY9Qo1uA
QJ9oSJ/PaAkXiJHSYjoLPK7MPJyecHpr/P0cD6S/OcIX3v/g4spula6J49Kh73SrqLqA2b/kB9RQ
uUxHmVaMvIJbArC46n2ruHIkGgajGMYoEyzqA6ut331wQjWEOb7LMRXfGusy8ayqfolL8+sCTohx
QRb9Pz5vV7lDpY38SvW8Pu6szoA7rlnZeu7fO+ILDj/xEGfG/CSGUlwf7yZ1i6bwIDczbiQE9lEO
4oX5AME76ciHECXYARm2AsUVrG65a8wTC1/+TKUidCi0JMapwrOtJmt564ueoXAuDqnV58TCPVEf
/Y8Lzy/OvezX/szwY/xkuKKPKfNviBe8j6uWYQwgRzfPI4of0NRniqjXRK6TVFMdq6+AoUfHVzIz
gOOn0VQv5/4AgYWKRosd7cuwK3TgtWBgqxG08VgOoQzlelCwHA2Y2iIxGO5mSrfyIJtHwLGjMUzW
STCsJ8jy9zjDoWgP1bEV/TbviySloP7/TNVtIjf9tE/n0FD1YKe87WbXzBnJyhUnC50GibWtofMD
eAfq9eZ+uJ6L3A7ityD/MjumbWWMyQ4tYJqehcWMRkJ98aFQxaOhdruE9T/1RqHyFajsLX5kQLsh
R6xdz/h9uyfstjZTQ1Y7VT5BsC5eeBuu+BrTxXlKqfQETTpfbIt/nsveJbB/AChN3nnR7TIxHrGH
7CGv4p2vyTGWIEg7VFnUax68ssWyZqgDPqIrCFen9axwj0wknJNXl0il6aBy1njhncmYgMsUAIw5
XscklE3VVSZqUEfSckZfJFXR7ZhWYrytOhU13gYYv91dWA67cA0Fhk86Ez7dw0vNBYsOaWjG0KU/
QM45NnWxGM/Tfy4diOnZzS5ras41MZIKFDD1YqJ4q1hefQ5lTUHtpKxysP6DcoSnhPP/6pjgeltg
aelIeLEZNy/cT+Z2OVYivyU7VBDovNZmehNcYQsXXM+60zHeGT7vnhz67GhEQ1h65HFUuJDVCZga
9Wx1DWYXNLLKpHv6lwfzbvwXiBToDZueK9+Wpnqa/ENt8Gp9K0oCb8qr/oQ9boMV83UXM2u2aPYI
/OowaeJbAyE3M7J3Ngrng8Z4fTb0a2kKcqRftIF1JKE5UGjvVR2mZTdUFn0eT14TOCNGWro5V4or
jYnvQuiNx70+j9AOypOd3Hr/7pIGTKOqNKSl+mYEdWkbDDpwS5HtRtwdl6DQuxDMzJTd2tzulbx0
J0nkkv2fAAjPVoQJtAGrO42ariWXVyYHdFX1DOlSPqpl8PjodNBwWc5XMO8jG6LF0w+zZumx8as4
fVte79T0JKQRRS9yf50XCckLXHDWdTm+bRK5G/IIxS+3mGETmNhu1S8v7Y+PqlO3G83BF3g47m/U
+zgRY01d4RKf6O16yjG/ZLg+QHgmF/ewl0+IyLEV3YAKPHJoG/D2qXLS2/b5BddgqorNsRAMWceK
j5mExhT2ctKwSI9rCstpQiRuVNcvo53DpXe3QEBVjCLapEWxeM/cLbnGbhHuRibXtmB9czVDU140
rjkOGax1V2LfaL6cL2jhmWR7jTTtGCnGsUHMm2OUfOy5kSs9D8N/VeGnxFi4BXW7BjelFrBe2tMF
h/kwUtlpHeGnXP5UNWcUGailBt7Lnq4bNq7N8CUah4XMoO6fWx+wSqT9D3nuOFqnGwY7G22elCTT
55YRqXMaEZy6395sBidoc5S9jIK4Y1ka08vu3dCOpuE4Ku/y4f3Z2ijI6wiNCsibSvPtntG4L8GF
usdWy+6SA0Pu/+Y9L6yuatWkwbfnOnqGb1vx6LvvubkpoknnLDsQFR9ElzVwwK+yJRxi2r+eVIDG
Myi+VvkNDTefpN0LoDRXwToIKNKqbs+hxBMnJWwrWsVqTg4/NOtj5hUF/rYmOqGnFeSdxCbXNZTV
pXq9Ts91KxV9KpUf0Dp9usGi1p4YODoXM9LO+HkJCsajul2PHi06XRidCU4qCoT7qL9di2nDO0yQ
bAshtp2taXCAMQELXPOl1nxoglFUfJ4NFb+0yxfbGikPIPFjFr9eb6ad2ARL/kkMzJy5z+Jeb4++
gghXbSAWDXluFqKNyZ+WugqXMVULLX6BEpjI5r806hUIjuXUuDAUjMZRZEPQmCVM/C8Jt1COHzg3
NJQgdpvzo1sxoG4xez1uPsLBJ0Dsktx+Hmyw6ddPXiiWKBN/nINkhSaJRHnuudC0+bBtI3tj2UdC
+4Nhie7yL6iW9jtBQPpZD0bVNsVThw5qHiSSBb7NFZHDrUT2lo8TlZB8l4CCVASu/JFaVRoG90zO
4UsI6DW1wJDmfoyubGFgijWN1pBxBv5/lJZUCqxQoaTDjOeS2X0tiu1V5yPWSthKb2LlUuETlVOu
i0lzmC79JALjKhxMIkUVs+jCQHW8NjXbYUR2HqOdCSLk59YAo8qEiontLJxGPFKrWj6wXXF60Tgq
LDN2LJ9UBrK0NhWkuiLrYoTPgLCeAWa2Z0+SyefX+fLxb2mNkT8xf1Zn59d/hD7v5r1VlQvuXvDG
QYmwLUVfEJT30dq0wPComa6oqW/O+2G9Od2ItbV4RsiIvRaondVjP0w6SKXvHh5ACq5t5B5M2HMQ
Vrog8RUZ8D6H4IWuJsJpSJybAj3scUciMXzJYeumJPEsRUJeaIej2QNjC9aDV1oD+g1sv+5Sx3S8
GM9SS+Hyc+1sLiTmam05upOsalFTdkSk8wcTLpG5AepcSljjwMpLHfKOC31TzyA69xNwf+sbzD2E
3GcconRU2ofq461l2IbWVuNhT2OnQ32cO7s1un5GP8dumg60tdp0lA7lKExug7WH1dGiX182h/SQ
3JUw3lkle2qY2egY2NNfWMf6C5Dhz7+Ue8PZMBKVYQH6JCDYt2Usp3cLD24q66no1OoAU+DPbdpw
cA5mQoXdKWnhT2Bd7JodVU+7td5HmeXdrQx2VHXANbi8XbSVm3yu8+GyGXp8g0A1zJKmHP5Y2sQQ
ll7aSo/0s/rLuax2n5PznPpOkaDvaRzuSp63ca5VIZBHoWwxlaVmcVFA4Oya58L9tMY8jka7/+43
Sg4vdIQ8mYyw1dFAQhOzNl0RZXmd3ReX3H8a4Uar2MGzdeKIL7WGTO1Yl89t5TqKCtKgVdv4k9rL
AEHOMBtq93wbJTcv8RQ9kJdpQ+TotBVlOY07PUjx8TZHgJUy59KtteuRqGK/ZQI/FbJ6X7GcuK3G
iuLEE51HWJsOyzKWxHD5s37JoDPmLsA3uJtLdK0NOtG5lzdviytvlCjtxcY1a7sA2hmQtpbzZS5b
nlMRy/C/+JKhYEVVGViMIzyn0gg2Um8Vt8qyABcIGBQedS2UjvLqD7JS82Ha1nC4FSb+EKBRKx13
7JBO5MXATZbIfLgFl91RHLbSFpa2Z/wWnw5MWOwkU8kWBwu1usf7tJ9Ju5feAbpZrDzqww69NFnh
VeJHhpOwsfM/u7SA5ioXegXFyJnfxzSqAIGQ2Y+yYaRCgAAFTJ9F3mwrygKLnQXJSggqVeNSVJiJ
c/vO6cgJr14w7WBYcGJp+JrZ6Uw1n8Qc1LS0bAq0oUBA3Vj/0NFx6mIusbSWQbScB/r0HSwuCIpC
WZ8WBN8qq2j/BkF0b0iglp556QLSB2eTj0UP/IXSpmwygcIXmyJ3MQJ9fFMLCd1H5nW3h8LZMri0
8ROw9qrqdwPLvQDTDSUnyD6nEV9a8Ym6NwIUJsGCfkyspO6Muy0nFUf8frvI8HGrjg3JHL1uwq45
a/Mqku5i/tlMUHoj4VaK/pW8vC7iNvv5BrlpkPOnghcnezB284pCr4bzAeXF3a8W+Gucw1oA0Dcp
zVKErp4mk0jE2O1n2HTt6TG7lxI2ZBqNI01VoWX9U20N6bR50MYnUpPPNQicEhKcMw0MYq6yayI6
TCj5vR3V9ypWTLTrLxoRNwCO0/64MGm1kYKituFQkWWZHEX/PljnoMLUE5C9G+PgSJGnTpvsCAwc
wBm1Ls6J+aCg3OXTOQAx+OZKcGmw9ZXj/+2fNU3L5+jV58d+8pMcf6qzdT3nlYKBJyaPR1re1FAx
TW3BIHG0XIbiThvn/rY9tpgfiT2rFl26Aw9h3iWyesnsC1VCTxHYKq23SHQfnEbdgGrcWIc0MMuD
kAsCiNBxZYDD/jXVDBVhW55/j4N6NWDcYQMDExduwQaYaXdCIV16KNVSgIjSNuuJJWRA5cB4m154
338UeyGypkpvkuJaSnBbWeJrwOqJJYFeCxIJVf0XruGAeGfwMl9B7ld2X7AlWyWJwZnESt2j0v7o
OoBahZkxqReXDudwlJWejGEy+I0qlK5+ACwBxD/EyEcdJAQ4ViOfycUoHcVanzVE/3bgMbC/HckQ
4lY2xm6TFn7QCIy47jDb/nStj+P470HTqexzu0vqny/pKs/QSz6gXVwyFWJEqm/A4cT0N35zhLd6
Zup3g2HSjh5llG24LBS4ZowqoUlkg4JNvmKidrKf6sy4XK+Pa1Ij9aojpVkackfgoUeBWAKJ+cy/
bfruZSsOnVyHyv8GjmfP/lWlZbRStAGYhV+v3MCGFUqEpgmoAcfhT/Xo3TBE+vDC1mKKsH4BRwt3
BgiGpBFW1onj3GoJqytiTtmMVH0PPRTKQnpdjsj4wPzndngCTnYCSlyAa18SEaNf/66+n5QGTibV
4BO/6G5Lu0FSz2wWK/Lu8+/qO3SSpRC8Lm37otcRueWrMbGUaCE5euo4YaPjul2YsrA9PdGyZn41
Nz0JriyEQI8dNYXK3jkaAzCgPPbNZqpkcehd9Puvwe437bFGjBYcaxKOIcBERRqUQqQLn5Qzk2Yn
m9OEH9ChVJy7D2JbpFJNMqOWGpMg/XQQRvTPFhUhfPioamNcYESFcuQLoyRkSB8XOmaxb3qKAMb0
0GrUfFh0VxJRAO637I5ACBipkMhH/S5BVPY/zLzRIg9La99hMb8vMs65krVPK4ii7gesbuUSP/Rv
R1paFI44ddOZvYYZ9swuEk6b1iFD8Sxighgx8pf1kPuGaMwrAS2SxowDuuNFJM664riP/RSV5lF5
NXu+AWrvJ2eivd7vJWtbLdmV/bt4fROF2oNlxXLh6KqPMVluu+185Gci3PD8Oz/TaFev+mPR+h13
ll80qM26bUNV3CG02kRC2ZCvw/c71oveAj6ZC1tHVAdgPxesCpXJq36/Ii94LNAukThuW4hsED9q
YfVDg7Zc9m90+zzn1Nq9adwA6Hr9zb8nTljl9hBtM7qLX05Mea4clPlXnOYv6iARbhBPjkFp6Y8n
hfWhToXRKpKrJy4edvhmIAGhk357BqxyD7R04jdaNgJP7aI5sBIr9xIAFwpF6Jwtch1wQJS8Vjkt
7O/drZZ5sTZAE9osA5QKCDJAyTr+ox0z+MR32bn5o6t6qY0AC+R+7O+v59eluAiRzTZ2m2iN0T44
OiMsnMzDh8jAmzdHWsz0v7wHJkTEKY694loqaVc2IrjZADOPTjyhzyK0jgbMASMZ2bLyGNm7iX9Y
9OFTfAQwSlxswdJeXX56xVS5g613bQKDsqrJtIr2C05It+JdlzI8F6F1omX0c7L4EvnFdAuIoSUh
T5Y289cufZ9yigCeHiC6MzaEKpCHrYkJrGA8sLxsy7rmRy3UyXT30BViRZmmSnmWZeVeLlT8FnsS
I9rXKMvnrGQ16sCJMevmiGXVf8kR2kYlBnnIaL46ON8y4AW67b/3kicnzsMQgsZh+CP9PnkiWkhF
/8ZjGEJo6Z2x/nS4f4zipVmpjAXMjwiWHL3vVB0DxG6uSjJ1kzLFsBJ7l9L7GD0T+VrL1dhElZEQ
Ukii0lQsD1uMMb41Fn8iIjYceqZUyg1Zp758YljujVl+y7Ost9MOzRp3HM7dMNC9p7/Fxt5TGl9t
ybyV1l/78S3JzekH4RqcoyxqFc8s5TjXTVH+B5M1cfUG0m4cmv16US0WY0EK2F+BPPNATi3KoH7J
YHWSyQACcj2PwUPw+xVloTBILLXC5/3C/uND4fFuhOdGu+sCINeuaOBkZICY3Oq5pNrH4C3ngeql
Ot88bWbMHSuCppil62KULR3hoMX8PWF/C89ix2m1M3pQouwrgEjAWuMhcoZmHVBkzrlmfXlgcmk6
qliVkFmNLBEzSWmEVv2CV8J2wp26TrnzHW4pcTYmAU6HSnML2lkttT7aeiSmzKF2R1npSuEaqzm/
J3gy66iTtBjo6zoRyg36edVwx3azLkhe6DnGq8JN/OP2Towql6KLdW58tXMpY8f7VSDmr2ggMmDk
eduo8FP++dPZoF6K4gjCkxgrKzJJEXi//WvZMXDFunF/yCkRbRG49AojAvkNo7gRmCrSBLo0JJMn
Ug7pRNk1J7entUYpbImOn0iBYrNmya3X5pRPct//PUz6wXQrW0i8MRycvZpAK3ypEMZXRxqB2Aog
AHpbK9/yIULEB7E6slTtPlI/oUlfkufo4U89lgLAavqKNJVrlilcBl6to6MjlOlhh3Ju2HC9Vx0j
hP+2xrpi9+MFdQ5XtzyDlCNvFCKS9lalTh7gBsRYPgL5sdNbBGfKIFiN5hSWPWtaTLh5eVWmnzno
ZLUz2mYtVWAqnUypGL8ZPBo2NXzaXiJPMEc7wrF8S5ugmoWRD72NaEk5kBrDsk3w8DlArJr6ykuF
Qp84LRqckbx0yAp/fhDNudxdOqky8W08tMtiXoWxLwB9RqT+SWy4ucNAm7w1PKvS3TW3yZrWJs25
A5fWMGK1EKXf+goqO+JSAoNkc9qUQaxLldP+d2UWJHI/l+czJ74cJPkIC2Cpa2MPw/RuWbB62XyB
I6cTlxa426+w1Ohwyjfc2dfLz8axvRrrWgR6OMTObDu8PrPzkP7ktsR1/dzFF7CiNcgZ+UCeE1VT
/OYM0ATEY/4XA8Qc0u5wh5HFSB1kajZ8dDf8GDQSKfzlw2J25shhlyuZrJaeUkZXTGIIauH2dGHF
Ohm34bGjZ+ztfesktaqkivCJp6rP8LwbY82NSd0xOXJDi3jAIPO+mEIN9rYbooNDC78Dw1DJzIRv
4nIuUilHye51vOb8Epgj2wgXWC/0wQiUlEuz27vtpu5foIF2NEanD8ipzhQY3nQiePUjDXBnjnBe
NnEt01GfIc9evVjB2Nv+RQ8Fbwv/A0heYy8SQpA4fc+NNIYsi8pOJxyLsT2m3WI3egB4uUmUIq6j
In8ohTco6NBrKlgSmUC0ey3v5LVmzzJg+9W9vc6QoCKr5GFuBK04AIqfH/t0rK7t1nMhNB1znOyA
RRC+jhr2V9h+XvCYEfieJoPcHZtEPQFwf5tKIRUCznj7q6FjWDQws+c64h5N74ESc6iDff9NKwmW
gCgE0qSmX/OvQ5Hp5/R71KJDLEC3C7AISfMzH4CQk6qr3p8iejU34HixdPYWmK/nnvOEk4QPXbdp
a2LgwpexfskMjwKUPwRbVf042+FZoGoWcIaOdWllDDJLHC5R+f+R8eQCCfsOZ1pFiPd4Hd59JWBW
k6N4J5V5Se9sNMUaA53L4rEWelJ/XzhoaCFGJYUUe/dpXLR81TlPVQQp2i9P9oWKwWPZ8iqxYDr+
eOThGAD4lQ6nFp+QKI41Xx/wmmWxTNqiorrNEXQenAzXxpzPlP4CFLFV8EbN8bk5X+vaoPkUjjwh
x5weAhHtsCY21Uoy2ARKuDjgm+QfR6u+Xsr0HsNp+UPnqNRQwWOtudU+kGCK8dNtu7XGTgaIO2cH
fEfF9kTevbYoiSE1wRTHXITaFwn/EWcV8zc3GrYc7cVSRvPtB9TupChn8t+BN0DwB11fV64Uwccq
KRjNe11jvzwUn1swckbXx/3rJUQghBF8I5P3MphhlXcwmcNeHBSOrEEoR5Gjfqh0fF24RJemgXX4
eeBjndptMIMSuU+BP++/0XjSDN2LP/ul09ENUyq4Mzaq/cfw1Jx17OL0n5a365R6V4abgv+iYFLO
eDiKqIqa43fgGlBEB8k7Z8ag/ytic703bGb3NyU7vjPjsSUUctxlcNPZnO/aUxj3VHfbhpNdieeq
o/I2oPiQIQtVPfxzIb/Rk5mhG74xkgCHn6jIaZOjGB5QDku/wjcLcbEKiwrto/c0VXIcIH6BpxxZ
Ijy44wZ6LNiOKA9DcR3A8p72Z6u//LBhzdHIDX2vH4SCDRSLZmnRwa3GGKCpDlgdKjY0ebeJCviI
DAufEqCe0kaxDbEZFMrRPpokupZ5Cp+fe9LHoCIZ9fV2JE4OfTw2FSJ3SOlaEwCDAG8gSkjWRcYg
tAaJGTJCkIeTTWjXEuwgH7h/njXVFBM5vfHyftjei/X1/h6w8W2dDuefbmyxgWonD/5do8jJjPHd
mJRtnQfV3ejpaRsttyBF7MbFs+wQ0FAjKootev2tfgHaEB7E0OeRFzEtsxaIvdrP5DTS3QCLpioS
x2ZeJUeUhfS+cEhDJCNbdPXFlyviiH1JvnVaMqWQK/+sW0Nsrf4dGGPvo7JerKlQjvL8pW/IlLfu
WHrqs8mWPTxD80F5RzmZkak6vg7GPetYD0h3LykOs7/ekvuZZUG5EPFss8gyx0dRMrFEoJuRKbnA
xlv6NuqSPugK+m4+rywPf/dkE5LQbB8P9/gsKMpDrDlroimO6s6QoKvhiyZrpUQ8xAERnz/FjhCs
I/xbswwLcwuTe8C1NC2t/BXaUTotvRzcbEWRx455iry/ThRx2nW2F5WZzBfLB8ppM7r8LT4fbjYd
kRXsp1sLvkeYtmlAxWT8RFp5BBYD3/4IihfK76LqPhE8WGuml4Zr+WeTKo8Nosd0F5Urwzd1wM5Q
RzjVLlgAeK893viyQRGz2uKScAPfCX3SUQb+h+wwa8sjYUf0JuWy9kSHh081tjFbI9RAXPLFvUvM
hGMafjBvggaBGwTrUDWSTFVHBO/vd7jDlc10AnUXbYTPko/6pspaTw+JyBFlzNFtLsTkFCbMgedJ
b6CdmXxm1ywrmBywiZItTqB6fKLOLxErNYFd/0CQ4t2Q5GHnfD2DfvJnQfj3FbxDW18Nq4BL+/zL
PoVXiS278Z79eXqyqc019gFIrko2CjUJvzm+UzdeELxwAHbQ/NK1YOiAT2HtBfd9upXNfrw96UOd
oqqWr/fdu6gJVq7y25Nq0NrogcvCHn/XmNkGqlbM2laBmcO6NXJNTcLOi4a6V4li0ieUNgYO9N9I
ntj5lBnb+rcTdQR0tNx5HIQalKGJx7l+5oz6M6Zie2Pz/EI5/fsqvjx6p3kk0PoeF3hDpNwYytyf
oiqo0HfMt4r7GieaFuUkOfAjgBKfVKHCGvuibFnPTAdkMRQVCV2/fej26/XazDtODlA0O8GLH+Kz
7ArLUxryhIDutxY9g2EnrQZr0bOVE3fqSjJhO9bL8v3V48OEaVsLFsuoEHsr7YslmD2tHmObEtPs
GhmUM/M4bOAOPFLdnwxg8VUR175df5zhJikBqVjfgKiA43CGJGsw6JDX6mB0+FOKaUCFQyW0EGCx
1IvuLycRm4rRPoB8KBjMaNWwBrVUlMTbq6NNg+x7GN52NO4JREh1EQNJtJpcdJpmegEqQJYHLCcX
tmSL4lM2lFVQtetWTEOC+hD0gz/T/cBYr0UekQifJBPbSMAFGpZ7XqqFTYjjg5XaF5Gik8CoXCot
9kDfEzpJ9zuPm0qVBV9GbElrESpWnCs6+O6Hh9kG1Yr5HbD9dnYQ9uJaEbMi3AY79oizetB1wwuC
sUOD94wEneMY5qwTongu+DCok6loH4xTMOkeH2ZeUorDz/+1ms9jKcZgLdf2pzbaQ74Jrg3AkPqo
DDoFT8U1RXVjLcaNJuiA60sM4CqMOCXotCIXdP7yQocho6xG+cDOz7gM9UYuSMxu4fQiAZNeFIoU
5xWGjnYnWWU0q/qhueivKHn2lJ8r8SlIiNvmt+2sCa/SUi5qLiqGJWeFPDY1tOhkC4V7t7XA7fbl
rDfeiZc18B7C7m+qFM4T09itCh67kG+o8i4zDMSwx4lrxRtegg+/49k6MpFkxOIXJ4HDzrjwl8PG
djGXpCZZBTGycHX5MJHC1Br6l5IkM6CP4eh2an7RBtHu/24bbISLBbOYgHlxPIHVsFlwiR7RItB+
7qsz3EO4DUZBBuLCgSM/ouMC+Z6CTzZB/7d5UcbAnnsco/VAOdcg6NOlx/xJC4+jsxGb4QMEqzY3
xuSGRIpa61atIIryREgggbWdIGpsdPaxZZEJ9u0ZabDaSxUTW7tJl8zhfOcy4yZrNi4QU+/sufhI
olWTvgFfUgLvwpo3Spglp0p/5AHNBtnB91EEMOyHkXC+zGseajXnjjfUwn8wKNGFp/mI4pANL147
9FKgrZwFlzy6mcvEvMH2MsO18EAQhuL9A+XKFmLX07btvtt62vvVWKZgxdXeIAPZGVm+mp8Xwnop
E5ZkrVddwgwc304zFAWmn6p9vSwtxdL5DYN+XRH9+G2X+3CXiEjnoxpQBHXCoFvUcuMPICfEcw1C
8cKuhYiQewa4mqD+a5eilDyU8C57QlOG5xuPf6eKzQVETAe5jZBAPFh9ZaUGBcnOBYEHXNg9QJdP
GUsREZzNpXZJZltSHYagVjyo56dCKLBHM3E03gZ1CS4om9Vt4Y4gGwaXmJ9KB57hoWKEeOvsuBFR
LZuwHlmFMATgdacc9Hv7vG9R6X5aOrHdPe5FZs4JNx6ulzzgdIENyT8IZeh6/jNTLnzl9BTAeCnL
B+YF9esXsSiJL5LUwx57t5sgBpl4q40vZ6xrgRfX/7hRKLo0g9KwxEkaEsbujiIH7qACPEteWywd
LxPjLwEfwcQXnk6o3KRx6IWV+NYFiYDzXmoDsi+9T7jjLsrS+NxzjvRPnY/1c6s0mp0ScK/+40Bm
IuAZWKDV1dtmmarjn/BOLyhw6nsE5WzKbDPmM2l1mF5n8w2bMaiwdWTv+aSsZsOx7Ysx4t3cT8cA
Ivx4PLH3SsnXWj5/+a+SnPVMCoVVHV7x0TrMmD+Dtb/KdCKQFStO/XmVA0ipu/2GsdNRK/EJHr3s
7avAYdYB29Gwv35vhnuCI7pq0YYaYactpfszbOjqOf0IWuK0L8xaDmE8xuEKF3TV8Rlj//h6/Loc
bDDDNcYCEAHvxYPf7P4msKUQbABNqLao2Ej7TfrSuRoJgrOFTibEwUL2giEqb3RiPLegFmHOrrck
cCePrrtWN6OAGewjp6f2VSY5Vx+yy41GYdnvjE0Z0o0d3/c3LbdF4E7pZkgSJ1BFMFeE83LwOzWz
oVCmJRRPhKQJ2KPs9RnApcg5LCokJEVTyu7jwrTxA+Ynr6P8MWiJpyO19LNdISKkP0EWbNXf80vl
dRVW38LNRM6l+On6cCUsJiOvP7N0gYtXdoAcZt4lVEOU55yQ0MgF3wq8aw41+EZyiyt1bTlL8WqF
EZ6XbIYn4x8lEcXn+EWPZOWs+Qp6CTJVzPjPuRMWoTXJ1bWYYpPxVNRP9jRk3r3oaDmtywxQ5bjY
CF+4pQ/hDrr9Q5UVFaiKI9kkhSVQKqAvm5/Jd5EfUCkKjCYD33n+XtB1c69k6wlqrD3ehxwPeaby
v5n+yUSW/pgDhV4C/M0F0Qc2z8w7nJlWkssjm1uQ1b04RjTh8nDQIpm6JQCd1+1lMLTW3fKsZzoO
EJvVEI9Q76bwPJtwaZLBYBXPjdHd3NbhiYQgm2tMbUhJZX7EuH7u0zd81danyVUrZdbjnoi/bSE8
dSMemAJqrHQgpW2tMtEMYHVPefabnSfiFj0LUZrk8IdVHw5VOVSwiAMjLKxZ005/bpXNyVC00ulG
tp7ksVIFyuGY0piYw2BmuV+BWpq65ytJytmtNA1YMRzcHzvueQducTdTM+c3ulwTS/drVZcrnV2s
Rzsy97uj9yaxow4EsS92f5IJSkyfR2ooxdmlBfgkeMuQ/YndTT8l3lBOH58LHtghZmXiexKxDvak
b5DiGObK0yHfhu8PEX5eF5uG0uR/Ck4iHSikBcf+JdJyQP0X7ELsubP6vO6QSny3vWBInutLSBGv
K0S6HAyEwNIlfEwVO1HPbiC3yv92g75K0r2g59HGPY4Eur5bhmQ99rkYK9nd3EJr21+0LfP3a+bg
nHcIfppKdae7O5FQYH0rokbodd55AZxrIoLULGvpMYqJmmxwzkKBUkZUgew5aP3RYOnFhrcU+Hgk
V/kMO7EuW5qMX4IqWFCNJXctr4cHX9UHoU9YxFWBGHYFcRAIBqwjn643oGUui/0I/pS5Ou7EyMX0
zJo1k964VyGDM6VvMz0FjDqw+J58VY+X4GYqbVL0nr6ZcIT23Fdn/70I8kecHYP0FxNlTuwZWGoI
ihz0njkRJPpjo+O9BY0TP4KQE21bLdQ+G8edKQPzlmYjlO3tUUN2IlK6QB2hLYq5Z7j1/DCvwuxu
HLDDNWEDKvD/PPhS2cYWpvu4h+QjHJpEb0Op0KxKRMg6g1BvkR+/fS2eMebDZgyZcGqoPyGnLqBQ
k6iHh6YeMkbOpjfzp8Iq+XRTgYOZQwCtqmezDMlEJsGwWCDMSbokVN3NuhtDNMJN0BARW67ca7pK
tEgwSJDdFM5iioyXNuvxab22PcwV2IgshP5uVIwa+e1mI/zmyDS7NJO7ojrf+N6HxrC9kyW2D5pS
17uAgpzYqQoq0F7He9Kp9rxvx3uB8374o+VGrleB1r298D8kTSJtJoAGUdkeD10ysz5e027rMCyU
tTKC/KElbdUyWjvOKc8RKksglvZqopS/C+xZJe1T0l3IbdoQd1SiYgPZyh3u5qprkirKAzNZNxj3
SLl//HsguQeG6ZWJmKYMkNxP6vbrOyw9qCH8TtokTtXLCE3FnlDB81eu6Lx9bF+1YIb5Rdi6UEnk
SVb9eJUSY8Zg5F89bUmfVE82AnqelbxV8MnaKnWFIpXetgd3hSIGrYiZdNLR9Jd3Ocdlxm8SFUt1
fx2fGHWUsoCqdwYGmU0+cA5UoMs2BAqAU7TkJjYD4UaC9IN8iiMNysQQmaHnBRFu1JrfD6Vn6Y0D
J62ndizXTEITJWci9Zjv66WUVTh8WXCuUha9eU1XstDJmLcA236PxE/3hEA2ByeIQDisjm4jlT5n
wo8+q4OIFn5ZdPKDLNitwYmYmdTI3QMAWJ3rJ4qdgCaiU8inMbDS1spkNMtqdeEQT2ik/8HMpxtm
qxs0a6jc2TTj2tCGjRYZ046Cs1gsCFW3WDuLC7VwPDsKY5tn1paRFoRXDY6oU2AZ1q2W6wjiMFRo
nQg6Jv/Ok3jkyg5AZDsHFxVncYdcTK50AK9bjooZiocHL7AkcsfpANJVhzmLvcm5INXXHKgwy1Bp
gOdeniVgFez+3CdNYTD16x+n16dAyQTantMIBQ4ZXRFyhlP7o78G7qAXRBFdfBF3fCFDWziSX7/i
MJ4P4vFyPyIcLULTdfPYFOdU8WPwQ03f/mj2k+vvLYwfNAiRQt5ufJDiTuhnUNCCOTCeOfJznmNT
DubLZwBi+3ABYBeL3Y6KpRvxfURKmygTn/+ykZCXU0SNbCfrshndFG+sxBpyDg25ikWAUGkrmEDU
Gk2GJHCrTZzg9NCMtP6DMLzBr6WsIq1PKt8VzPDW7ZyJXXh7SGOOrnq4XmgEjcCB+tTMAOwGmLMV
53ebwgg8T4dgyNtVut3lbQ8Xg6Ky4fOOfP6hF3Yl14f37cedniOIOQc3J8Anv6HDnVyhYEGApTP0
7a653zcWujzSOH86HdNnuSNo/h9BtE+s43UC7EjMZZVIJ+39jX6p/AqlC0dAunPy0EYnrp/0ZS70
ZtlxmWAfbqI7kJURIfMZSAr0smVEaTTCofoM/ikNfGQKQoFisNMxpErGBOcFtUc2Ct+T+pcL4QF4
6lqKKgt4iPrRT48/H00RGaITLKXhR2dH+cjetyF189Igv48/OsJDYSvcb+0Y7wIUxHlU9It+GjF6
ggt410kw27iCcJBjYYzMHrbsIFp5tB2dQ5FyPUrw7hIq3fcgl5s07OC0SUDd8E8d9IfUkL8VvpGJ
OoBuPFwLCoEdHfnml1ud7oNuDK2/qE9+i7tgeqSdv6fs+wURsG9UFKWfE1WQDvU181C9BzdtthmO
48DSqsZTyzlEVBpz78Wi+6B6wwoqBPfIZ3Nki0SanZif4YDXliYgfBs20ZOBREdfpde3QoR9odE/
iiWwPhWR4SvVTkIPjSNIteCV6JIAsJqVaAL+sEoQmemUzmz8FfPJTnvY5mxQFPOJeS6yG88Z2L2l
HpeCiu9wuC+JiuisJFVMOh0CfRL/4i5hceG0o28kPbu6iw7LqRN8SvN8M640m/h1/Y/MPePpbrRh
cZR6Jl1zbxktXb0YtYuNnlyU9W6DsU+h5bWF9xD7LWf7HjvmfLs96E9pcxXucasJu4mmBNaf1RFD
R9CQsi+k8YO+EabiqRVg+OiF2mOElrIYi/q1Gt6bVkFo0uAGwSiLH+K8hsC/NZ8tOLd7m1MP6sTU
m6SMUYv66+A9xq6mXgGx6Ffxx5V4v+HSGXj/yDP3G6o2II4bDoO4huh5/iaQRHi8lcUu1VmPl+/x
udiJpa7YpoydR+ff8QuoKt3uLXGhpbLNuZkKL272W2RhbReB5HjUP/9b0cga0+SugH8NCwE7cV97
Q2nIjPQqnalbX/j+kgeCmJzGCaGLIysds1twlPcWHJQR8YgiTp1pSriMlHvj6ox05JsNu5KijPnm
StjQTEAPUZX4GsYfBA9isoVKgIKnSX/bByUoAYbnI3q/vfKgNrSIdWKGozZJ4AS1LEdej0UueMK2
OqE/N2ycXxgAPSfZGa9Xd/EgLYLCnBGFduPsNdu3rWCgcgsTjvOj39khJ9kSM1uQJhmwql/QfMGe
neZpFSyHlgO4kMAMQECKfJyVyD8DWnpOBSBTv1AAjqzn1WXSu8LvbBCTYkKNzFrZQpsLm4qhKNwq
ZN0oJoMH4mE2vDaN1A5EGhs5Zz7I50xJiIGi4wOw1V4+wBBCalySjdfZ7bln/ZrcWyT7k31NEUuM
ZI3Ds17ps+7Zs2oV9QGo+sN1SS4btNMnZAfKqXHYCuqKlHxyLvrbUjU5JGPdd44a0ek7XQgy46fw
jNDRScn9Hf0lWJzl0rk40Ghapz5Jj9+EuiZCI45Mk+4VFs4AsQkeSuU7Yr9cXTiQxqqPBvEdY8JC
Uce6jVI7H8F43vBpMDAluEXCoBpy7BJNxpFl3xVoDleFl9t/BOwWPRLnYE35FTTluwMbTsnY3N4l
3MMwhDgyhMLJ/NjgqooMX4qNTKD5nIZenvzvl7jozlaSRTOhlI97nN0nUKYQcn0AzQcDq0F3UTdF
RyEYh0vtbSNlkNl765mWoxZrj1THRLwOfNQjwlbZ70MOB/fGaX+wviWrYQvhU2iqbkzSUxdaNDNt
RUyMN+sM8179y0Bx+2/G90nhJq984Jz2uX4xSWs7GgSlG2Kx+ZAChja2ouYhv0VlFSuL67/iTw2Q
cj2nqBYS5RgxebudJ8Dz4RBI7mqRVs4Dd/xsXgn6UcxwdvB5eut7SYcpOSq7aNzFI5L87aSYAb87
K/hgBieNrJdsFuv/4WLOP73SCxQEGYjZR2lcoecGFoEDiPW1PmIOXA5S7UbLxNPS/1bA8nSyr2Bj
6fG8JWWwAhVChtAYObmx6StdSOzASOdVEtgvGyo+1WCHU6jcMi82NbQa2pA+JGB0LrxcXOoGb3oI
ziPVLyuZLOU7GHUeDwj5jqXirLhhgNajudza6aLYij5sqJcosSHSNjBHqVdIFzrMum5HH0clMwob
osQsTNmaK4bgYqRk5x85bS4466IrDmMTSkoY11Mw+lqTXhxlbs0O01mlmUzplocFi4FJVWWk98tc
CbiIk0skzNHpv7+A0L/ITkCE1e0keJDTaqr1qyMYGKpdoD5GT7oIBzn8wgTukLrB5GBX1YjuD8F8
kUt8zxsxQ7v/WRlFZaFN1WXWn/0X4SUD6ImaNyrXw+clUUHIxKJb2PjBhPmsZg5TIsTDGuHuPb0L
5CZ2wbdylBv4dUCy2v9t+iD0Lsi9ENGnGGJwDMVut6epWWBGpPEX48/ZPh2IM9jP7ct0evrQHNro
i0jVfHLopLr6YFBo0XfzjR0Al+01aFrNkLp/n/FxH907NA7LBu8f9tkbpComruOVgU0jw5bQjxd1
Kjtz1lnX+XhpER9szT7iyzBzS/KhIZLac4fjZ7ckSLukTYrYklR9pHhRwVi2mOWDvL/KvBmL/mN+
szLI/zq3wP9iw9vGhkbPXgY8NQ5slIa2KQbcLXtY/ojosrZke1YuohhwgDELZyu37PON0RQiGaL9
+Q3dr3A+Gm+IL0bNsTjJKojh7OEFWlaZRR02M+oDFqqGiS0hOlm4MQ5AXNh/awXsh+EoS2D+9wZN
JQK+y8a9nUqcQRRXGBm7BhBIkv+R1aAkr/boAPXyduMQVuCChpoefIR4HApvkR8mMTPpv1c9DGQr
JI6uwW1UbrBeIYVnfRFbHEyrqiD7ht3y5lmBSMt/SRU0JU0no9qtNe1P6CiGCznxm0C+MT0EarCk
VtvagjGschIllL4e3UZTKLcjoDCZPcUp9r90LRehTNVw0F02+RkY1mE+S+TBOyGK73YpOgAcZ6lm
ovc7v0ZFHrhLpBhC/R2OcNDpw2Zkr5OiZCozXS8SEDiH1KvgHQobP/O7vgAb5BigP9mVnkrov5KB
LxVLxiju0Y1sMAKvsYHDQkR4Rq9jkB4aFPrVCUY0g6bA2Xp7pNecn1kfPxTbNAEpa04qM7VAiSho
ZkQVMbx5BvD8AFlZvsAvJfulvcWVdR54R/ysva7D1dJb3qm+PWg1F7d60HgeYejOL18m21+yDiel
O5a0YkyFsmxb28+Ki+xDloSfzi9ux1nNc2LOaCM9Jg3TohsicmMjkrz9ATQhrNAwEHxhZBzcdz6/
Gh6LLDXbGHE/RMKQPEowxJK1CAx20MQh1kogQkqN5kog72maAQfYuswtajZfD2dUppkS97NSoA3s
UKjrt/OW8Xij2vtWaF8mLpOeSE/zUVFXo/nFMgbN+5U/4+iiVZJoRdi+MqU1qDMtGQ3TLTolJPZ9
/t4OCYqdVZY6UoIWMQJ/+C2TFCkglR/EPO6ItUunIx4BC4eInbEJ7mn1ZY4XxKn9u5YpZ/cXAgk3
vJz3CdadBIHHptSLo81KzA47sqfZsz7cq6MdYvONFvFTGyiZkkgrjIgPytw78dwAmcJRTjFHTQ/3
wwiXmpCe6CBhLYjAh/uQTui/nPMD75BDLJLsq7e6NdnrObO+jiQwFPkSgm1cOgkTkWuIv0A97bBf
dUotskzlKJyqdczKLJZnq+cFpPtEhY8i7T3qVqXuWV2TReAPpZgypdGh7HYn0L9zr33v6WTsiGgJ
mcydZbigzLGc0GZO2f4qKGh5TltbwPXXfI5d9UCXL4wfLW6lug/2X5Pvuss2j4Us3j/yJUI0PhHp
3/IdHjRRl/NatVt7RuA9pnRxGFH6+YWs4qGRrycTXovNn4oIJJPZ5ujJNXAA6AR/sU8CcVYLT8AZ
+WJPg1ATdO90jlTGfdt7suAlegSmsbW0uDIiYSHoPBJPj5I7v6tJbnwKj2LfiC7Asi0507SHUxZ3
u+8g7BmzgJyB+8efbn9ZOjf+sifChMXKLGKTQUzWHOP29P9/QQRPUuiscmVCYb7NLfCPuh1ElzuP
epMVFj3PsEnhkW5O0HOn7OdkLEMZjaAWT96hCVt+T2fZiMrUMopjEWUzNP7hmmA64W82iOvO4DyF
9rmuPPRFHClCiyvBS9NKi0euQhSgWkCWunkXDPC5wXfOq5llrzibzD2bT+qElb1KrSA4M6RTFQof
/KtX8/09juXcwwSm6OfNofg13niWHwVAIweKUys0Nxu4+yBBXHGEuxxiv4kvjKiLES1fD2Sn+Pc/
YJSw8f3lxVqOc/EsXDOViuSRrJUa+hJKtagSc32Qk9hkHViElVVFiqVl9quwHiMDfUCtSFRT4Eew
Ktc6DDKOW+Npor3uBSZ1qc/F9a5jacWPXRhUuIXdY1V3EtqSQaA2aIW6WVLP5AymxrKFkc1zw3hn
smkR/95jQsRwTrbKcXl3kGGguQN1T+r65l3YaFbne1JtK3KEGN72k9MelzR4yrwO38TzbMBADCJX
roj068u/3Zu6Wj9APyZr/31ZgCrzL8IBGYf7fnOb5OIkfgaj+Wg3YecDcfojm4SeshEaxpRSVoyv
2pFO52X8U8y67K9wTbx3PDXL3EDbkZTdXKsVGWIpESYCmXUwDPgAjTwQcMLXGH8xsietKkAsOZgK
xBR7E7RSK50IBPZy8WW7BHWaleObtOAgCNzce64X1R079CVGvFypmJEhGYj1PvYXG9MYxEEJzqDh
OdNmq9PFYyoe0VssvgoXMiCf9Nyu1EyxSAhY/fq19OFJ8w74kloiOvnpC4DZE+xw4dRUeVIUiE/7
lS17sQ3FBXfAAgFozYyJ4FUjVqWz5IcyOD9AXnRkZGCZ4V2bM7ntR70HCaAQgcW2oK9aAzbksykX
Q3owdgwTOwo7ME0LmVAZFWbeej0sG14RZk4BwQsUtzi1lTNf2gvW3jDYY+7ppW8EkX21EEPbAPSs
/2++OoOw28Exgm3AnbNQ4/khzZJPqDp+N4jthArg1RHjqf9ndZ+k+1d29mxCF6mdV7kTQa2Omaaj
+gJdKG/UfjSnJLlsWbtagfUKBVN8ASbOd9AEcghPHyqrsIc867kyowX2JL+H2Vwr5/r0QpRc2bb9
SY7OBW7PpOrACVlhy558Y0bjNLJNQegYwcfsZ7UZpsS55JA4be/YPhbyv+GPE4ysKLyeaVc8hdD2
vr8nYOWOIgY8kV3AzdwPowCxdPzCTRqpGx3y0JSd9UizxnptwjC/X69MLOOgsl1nu/aGnnLJ7rtI
IQ8ZTb6RPIaCX3tIw2fgrF/e5k9hEWp6bPV9c0vKNRFF4RSmKWc4BbfW9W1Tr2hfRNfL4ZQtghrA
bo6mEAG6GxuidYkwLIQGExMRD6dXUnN3LeDJFRhvX5hbhGW+dZQOounVRMfgW8Y+wgkSXW6pn8hy
xvUXxon+x/xDq+nvLvs+1WOm7RkLtMaL5wOsRBcdoicYiKHeAch6+0WZnZO+jlqt2JNCJo2HwSD+
QGxY7ewcumNaOBkCOLnxNkA7s59VmtiFnQiRjD7iBg52k4ln6g9Nea6O5qjQTImek/upMNLBQzBt
1nxSRHZzuzq5P5xkTKHXGcWX6KbNobY/jyQ+Vrt5GxpSaYm0nWqY61NPYD6SCEYmOCph5RrZZ5Zo
fHV7eaHKevnFgVP6f9AL+DEWcxchUcudqXL1c2rtAkLebhodVvPxVJ/MMCATltFMhuKEifutFclc
HDrQlk3jOzRWELQ0cdzi7c/jywwZfrH0SjPhLuOukIV9ou82MVOREf46f2Yz50qa9x+uNYsnSu9X
ijWUn+qhIXFrDSEZ1gCzdID+P5SuvAO+tDHeLJh6dK8SE0HEqo7coOkUITNcIlGQl8vcB9Fo5x3C
NhRPVVt+HAmf7z8BLL+XsZU5ERnvIKk9mqS9Gz86XlfSnLRbfpWRepjhIE4ZTYJXAevbjwO4A1Ym
YOjdvY0lGCaz2X2dKWX52y/qIhf5P/u8F1nyub7/GdDzkI/0XRwJbt0owSdirEcbyncvkopJA71V
3zFOu5nJUhqIZpoLvdIEOhzY/6bKQo7H1UR0bCzIvuRl/kZE+6G6hSXmD9enFeY0/0+3IW9DuK7S
wsffRstzqSAIUsMv2Rr1oSbBl/CGykFBI7/PtobtOIQbcqHALtXXvzH4iIKRDMTAojxh4W6HRBUM
65bDKOfJTTa+d76X2drHW5DFW2tSaEv4RsLZ2lX5QR5xlXxLgv9AjAXx+JfCLfb6yxkhHRL1jl0g
kHddUw7l6yKGpbBZ24qB1KLtyhDv6x/LT5BuQgzjQ9JlVAIyCWWD1I1oqRRSkSj+mKWX8F0B2Pps
b1X2/p8UkVFLQBJHg9qoh0Pp2LknY+vQCqNuJx3X2OPTypHv6pL+CmA0x000N5tLZvpFDUlY9DCa
hFz5Iw1nhg4IwDUtpUoyCKhhQBfhJdqM0b9SWkaQMvxnorg5xDWAKkR3zxui4I72e3CMvzhIOVrE
LOCCoRmDS5S/6ByxYCBMBQdLzOCD0kn6A75QcXQz+7eQwh8ia9BiXBwgvU4lAwahz592MhmVd/Ad
3ljjDcw7QYi/0zXRIGfvaWAJDKTbVU7djazr+yBoO+uZjNFc/vVX0HhVD0YbVM+NNKQrN2kIDzQE
H2YitmrNY5yhaw9ND0SLs6ibdXq56HfZ6JlOQU9q5XOkVFuDVj53wPGRqOQyBA2zyUMhPaXNydca
isxaqSf0Jeopbo9CWm2CIraGqefvuP2CbQ5v9sb0Jopnr+ndD04WWUI3pyS94QCSerEFQveERF12
5BVuWu0HaChqK1YYd/AJG+8DN3qWt6G/rCl7nkudJri9oMIp9g4TUr9yo9xdUGM/tyqtH93yd0lU
0z4eptSUpLUxTbt0ZRjYFrmIxBUzPXvSBxlgo0ZNNJsG/fo0r/TQEFUnSV6ob5qNDNpuIVaq/blU
uqtvuN0ioyFpV0wCEYgM6gJCyTaS8HhH9bJA6MOPHa7Y69LXzLWUQdgRL8Ei1UpNni6wLiN/ll6W
Unc6n24sfzCIcW04UWD5zzCKIZblHjpCCZ59/3/9QNbB6yP1CgwcT45cpILtOgAuOxyBDQENDWxA
gfCrqwthZ63ol+9f3u3Tapv7SK1vnbPQ722ReLxHETwpN2ajSwAhSqdx4O//n9Qxs3GcI/cKXsZw
h5nHY4vAlm9z2U+KpL5aLGyM3c+XsMYvAGPKjHpmSH2soGw59tdnu81tdOioFplzwA5sDSUPMSIR
hdufbSoOvGSrqPtxopxaFfa/WnuCBOQDhGgi3ShMYG51IE2Qq3eEnPFJTPdx7GuRgBXFov/R6E4/
+YvWRlGDfthfGAsTBpoiYDkHkmd3R6P28Kh+wNN2Jyvmoiqoykw7JEMwr45dvSnobu6tsKmLvPag
OSed8Q8uB8ntxtPQ8oAkrKe/3/krhu5rNGp0QRD/VojnAxgQXmAs3XiaBotyyVU6GyZ0uzdzmdn/
S8QwElTSNITo5kEN+zQ3UJoIK/GviBccIBI7g1KURekZwvPOKU6pBONdGSjTQywSXMpTxbqhVDqz
YPiYXdLQ8UKHJSmW3MSQJtbSO3FuJ+smxMXm28KCXWAt9ds6s4J92qJ3YIz8iqLUDFKUSgn478vG
dqkhma2+3fW948X3nJfigbeGXd8pATuUDmDuB3Iz5zfmMjcJ7xB1SFspteJvZ8ZM71ZBKLAQKlse
6SE8Or25iEe5TacLEz1Y/eW+/Ja7yO+VMBjm6w1qMe3WHkVXu5cEPo0dIDb7A+XdOLGB1hrHd/XD
aUDk2Oukkb7Iqn3PBYrPAYwVrXxTGJQ0eMaoKEwrwZtq8nKY2YoCc2lICvgO43Y3lecuCBNNHyMY
lwzt0QglGqdBgPwscr3JITj5n4fLob3IppOvePADNQShSqOkKB9FAY7CXJoKoWxgMhv5e327WTJP
Bb25dkhDSnCk7/Hwg8WkYb5fYHC4vY6bHXeE+1F5TDoF1Dfwkd4TpEuZhJqmcVGMG6sZGK1ZJ5m5
6EVAHMgUgdXMcKfhFRrrhiQP338UjoMrIjo4tywlq98hOwP5mMtAWapYG8YtG2YS2uFHBLant/dc
xjfGymaHz7QDGAhp7dhZ1WsHjvsdCoif1mEwif/2XQ3/ZwSsUTgq7oQmRN3qHKi9oqbwyzEMziQr
8IsJ+Na/7LpMMoanFYC0E6QW7ClmBTeUu9jNeyphLDKYYmSrdW+6nN8gbXgN3v+/kXxJvzZUIF+a
9JdRxC5f5uOHB2ZZMT6F8co5i2uiND4cE1JAvHMQzbEHItqBgtg/42yyE/wPBx/6B/FQbbJHOO7f
iJ8U5d3z4qWqMRCHZ2zg7PZZ32y94O1V6oNWvWxbMulbaKDPvUm1aTBXhiGBKn/WVRdP3dAKIGty
Cv6ehQlJbIPtcSpWE8Nl03eFlQPYuf/tvcIEnmJLx6mbAHsOAri7pm3d0VNTahtGwZBlqVNkrWew
XjKfsptVf50hEYNuBePZP2JNvAJfoZ3mwmZMZ+sCf70Ok2H62QDEU6d9pE1ir+fzhVAuz3duZvDp
T2FUR9y09fJtdnSvbV0y3YlkpuBa2PZtIA/yYyD7GcEUCk9do6EsdaB9cjwI38f4tid5vqFSn4x4
rUvN3oRLKXOhU1F27FFEPLDxIoUbHfyhzWsb/3ehjNuczhkqiPKHyf09bzuRXUm55gh2yyB4T+rh
kZAYgc63wIiKGYOVlp48rktjrQ44W3KOeqeOHdxoSeRDX0vGHeU8VNDRepfB0+rBJVrDJydXSFtf
UR7QmGWQiGTJyKnOACut0kUwOqpt5lVHwpYn6TbYTc0RTjm02FsqKUT8t0oLXTCm37FU81ubUd9j
6Yi7Z5dlASyBAJNNCz8Ujm/UrIW+7r+NklLAo9Xg8YPeKpzWTKuRD2vX+tGgfcrahSMVs8zY2/Ci
T4fAJWWkhiawsY+reAdEaJ5RoIqo3nzSTIIhG1bGf4GGeYYys3TxPBQ/Q6LKio7oSRurtc0M3DDu
YXyJjsyFqiwLCYuqhcWMJFGSpk6+UUEFjKbSOpnh/+NhiUrbZPebTEx2lYWm3Obb7QEG9QJBuIWm
/VH9NofiBG0nLB+d9HGmFzvaPRPLfE3kiEr84LLhuOfyEDbVc4lFKS2DgaaDq9NvxUNQS7e/KmYC
LpiaHxYLruqSr9zJLbTqeSY+FWiFxmA7OkuC2RCOySqL/E6FUNuEI9efCEW5gg2rcbB8ZtKmIqGS
Diouc+m64oc/dWA8s2bJYTTewTCSF1o/P4tKvenQhkrZcBwnoFU7JvK6My/+XYbL/+AC4TS0ntls
xpGBkagZoa4KnXirGy9PgiBaQ2uabMSAN8j8e4z6MZQTmlGadHT/a9d8SNnTj37sAqdC24QnSd5O
NhBUM8O/yjgafgLlQKstm4mK6a5CQQMTty/Ah739uHkV/sHPiddlxDVHZftuEpDwh0rZjJ/OpQcq
XfcRXYLHjLbYNGiFWBGgk0+W+NcGK/wlxO4kK9ETNemdVGYKRMt+5Zh9/kAj9bcOGheWhV1NYctY
eNH14SIh3A6ygmMA5EG6krNlzNemJ0FMZDgM45o3symfpnNrVJ8SHRYAcgSFUIwL9u/1xhIFnBU3
mSvXYLHdJQN5i4m6/8lqoHK+UILhRIfg2h7WpcfZpn0COeEJ71H/Tu3ZiGlylkrNIFmezp8Ksq4t
Crzkvkmlvd9sep8NhgU7fK+XzupqPX4s98QOppYCtywbKXKmzllVt2K32OzQslQxJ/9cs8rU68FC
O104X3D6u3nDre295Uqdb0nnsMlXUCOrIeumXVp4Fe3po/yk9Ckcj2lSfHVL2MjjAOvmG04sbSC9
uUb216Ca6CorN4Z6wzqXCYaNZ8UpsYUpoNULO1kuHNlfDKr83kIkNFTVBCNPlWxw9utv7947ryWX
tz/Ok3lABf6yuzBtsqoucMV8n284T/fNcx/Jt86XWM24yTAG7fPteRB7IDrxxxJRKkaPdPB57tua
cSf/Q4G65R/W/X1r18y6v57w88TN1S9iE6//LrOw849oI2hETerzV7eb16/DWlNS50+oMQ8LwMIF
V+KOGuyVbKYWRz0teiP9GKsxB0tmqXzTtwWI1a0haVxiNdjCxNHv4VwuOx1uXhrBBolloSD8vqoO
WuefLbpsL4a0VSlSU8s9ClNEtAPxj3v1hNQ1mMReioFn8ixIARvcPyTiE5+5oTBea/pRBrL8Aqcc
UOC5ySFcfll+XT1Z2IRzastpBMdamIHka+r5RmT8EvJ+HgJ3iO4oj4gTz7oczg/Pf7tqqVPuGpRn
3DE1StVvhyNc2GLa0YqWFBzSfzLlgMicc8bAKIbCYOXALaV9JDU8ZN/D2oxG0Rfs/lviN8dXuba+
Pu3CAegXVJlyd7huDksGtGF+ev2wX5nxaS3Eaofy2/Nw8f7hdVlefuu5GCbhHaU1nnmhI88RYi7f
yUaZfocNCGICx81Ea/JEqWozHYlokC7YAzGWCfNf+UAAqkBWZyBYFUb5pmdZYFcHk8nFTu7bmyOk
YIm3WSieLhTO3rWmGXJVoasZZPc9B0v6+JZ+wTpWkX2ClMgS+zGlTHOxgaIYUzJVXGtQSimDZ/eV
X9tp9/emyQj+ImQh/SPu3R/M1zYZ2XGBZwjQNkU/yjVNPXeMWNZKCtl/chtGzETAfqM/Kx+nB7t3
iacQDUUkpOJICA0SY1t9Dz3P4p4UXDZlFGcXvFr66AoTJxHdHq2Brhj8b1Ifc7wGyK9PQACF+PMR
EYPvhqPXc4ZAyFaBqnqIL2pYbUdjFEj8UIjoK7enq8f1skBbG4Os135sfZ59+KgYa32R5Y2G+Ini
/XFUzEEYolSU3dErn9R2Y5CgRQlxADK9Yue3KEsxQmMtgfzNw1zv077IFmwmY4rq6NA+gEFV1KjJ
RQCoQNAWNObZ2ayv/RbRdQ92Q7EuUN27tiYUhyp1mMgG5to9D4Uk5rWPGnhzM1YtJNYmpymdeMcm
yQgrnNF5M/lxnhBbH+PCLirqp0WYohUCfZHZVJ3Jke0ijt6ObkMgOdwW+bUgN8Niu/7HrWYU7oCU
ZJHx2PpEQzstoKsQ+wCRrFb3LgegLmgrheqZm3npLLejGQLQQMXmZeo5w+jzNNYEN55hBjdNFVYq
GcRDAVwr7sDEl/QmU/PeagyBPe3kSm9vtnQ5B7emlKWbYNj06eJxCsDmFx62tm2wfgWzOFisH4eb
kXq+5235d6XXQUfXmk9PrSK6UEmXZp7QNcbfNDTbyIaN271zCcLjkRZhCcLFlUNSjTh7B5roOPLS
fzMzUcZ4J1QYQJ3Mu2AKPBcdnAkj/oFK7Ztemp4m6EXERLGU8KKf/g9xzzGhUZE8EXEBMopCCh1J
2NjT4txBdxruxfc8WFlu/uQpS1xazIF6JTkdQmO346FUhv34OpCqhD+lIau08+zl++/wABBHXlwd
BA2AsQROLrphDKJeEy8c4sp3R8j98a1a7EBOVUYXxV+/K1o75jvsbUxOVR+yBhwnyzUZbauIHmgD
8MPmZHnDgu/g3SNqcPiXv0tDwlnM0wE1DHf/tN3JnAspNRztkQJLP/wcxzr7SZMm5rHD8hwxdA+Y
lYOjaOWIfU0ZvtzGhbfnFwQx6EMqt8aBC12zO0aABK06sQlQRb4qmMHymcIS9pITwwdiBclWer11
0ReUttzNEj0Gh6RZXNhQtYEr8x+GuwuaWYeQx0px1zWuybHe4fuNgP+MWlfcNyCDwFJ1NrF0t7l4
dHithwheXzm13MSkj1NJB85sXUDteCEdC2Vvew3Q8N3Xj+FAKoUKohePig7FGxbR0gF4IujWjlZZ
OIFuFt8esdrco8ECOc0SM5wiiswPwAhnbYPTOl+EENVBwaYGqnvdRRb1yT4cV9muOtBoDj1zKwFV
PQMMknmvzNjYLRcCe8dR1dAydb0V5o1LAU4uXg4bwHvDkmc96FuvTFBNXD5Fc2pBTtm8hgCFAGMm
vbZRF+i0VZh+7aKySLELepQ4w3UBblTkufiYUeGyW3r/xCkV20Wa/5mKlO2RUEWt490ahfctKTyV
rnOsq3nw3f2N62X2Ew6EpB7FDcl4Sh0r0+xmXWzRnWFBXDBbeTLnRSgylACnIfZ7imXG32qQuKAl
++gkrz3sGc/NglKfAFII9gTvQLwd5tMhlh1uX5Q3YfqetBqMx1kYSzDc8GMbtCBbMoDJ4dQA0sM2
DrOc3YSQ3zMxxi4uoSlHeizkwWl4ECLU76LtIqqPaJrQ+CREUoPQ8RmYDBjKwHgS9v1JfkFwjJKv
DvTBsNVUAQpoiWMnd3/351iwWP95DYi0WN7JwIMfW7WV3A5sVBah1II7J/MeNwKwwvh6Q2H8iz//
m0xh42xdVqD/7gcQDUOHKJYVXABD6/Sl7O00kAYHZQhYGgWBb2RyuxAFEr2NSoUjxzWWFicD62TS
a5GHB+1VHg6Vm9sOsIwaSuiLCgcvq5OllmfJNhBo0f7TznDLxYnH+k1by7SmeFovYpvRcc19WIoP
lNh1XESKolRPIlZ5Cy4lM11MPxYdmRw4y9b94pPgaljV08jD/R/l+zg8cbyXdtC0hBC+cUxQnbNv
b806vl80xHjWNcT4sAINTIpx+mXobS0CnWulnct69pkY1BUfCVVw3BvDfnLpihidRLc5V5AdZnPI
GFhIBgz3/qIjb2z/Nf67iawrBoYplm2YZA1oRPyrA5GvReFOARbDVs6JyTmNvb9Bcnro5dgMDTFV
biUgvJn2yyJCFj7kc+dB+kA+JO566UWV7kWPRygPZ2egKvPnmpc7PFFNaYtb+KS4kyC9+sKLoIKL
GXJJiHhsz48LnhzjoNPkaFyEj7aFfFyZLv11qbGQIlufly2+Km6ZnZTzYS6ximGc0hkNUp+z5/ik
ujqvTp7PKUay6pROu7bhm1oLoxFIEYYHmt9LT8jVWYWGum0QRrjtJ3EK/zoYRA6OPCks651ms3am
sr1Xzqzsy1+mgPPjUvNuZIuNWrCtrrnL8x6hFqZKb/SW2HF73g7ytt7F2qzHUbD7GReyd+AmpTdL
WQWUwiB3yoRRToYtoOw7BNchkd7jb83D6Nc76oEoPfc3uH4wDsYR7+CWf1wwWMiJc3GaRnU1gAwz
yLI/Wxu56eLQb347/EZKBI67QRdDDO3O3iTIZqs361H4Jy4XY8pblL9Wa2opB8UBmKhUTmnvKlQn
np7CEZxdy0a0iWoo906+smJiZi6QjrLa/igH58Lc0tPRor/y0H2u9xHsUious6a14QD7WkYl+8cd
E0miQsSQqbPhDOctGtk8LdaADqvkR808790h0lup5CUyHzZ3Xb5yMtKQsLZRn7Ml99F0uzbc04NW
z29AfQj4r1qdKhh4bVJQ92ns2RAQXNVQFfrrzvgi5mVd2xYpSBhvbu7Zc6pwGs2m7VgiSFFhWECv
S1Ya4AKOPGEPqKywam5D/kfoLIXG284EsEu+xEIhslOIC46AjPiP+fyebvQx9omf+ZWRmgCk+Obw
haSUC/pPsHswDBan6zyoyvz+Zu+DQNymHdZiZEwjMelG1+6LJCCHygVZXRd3iTMgD77nX1aFvmfj
9MS1xdhPu+5NbF7SLKRhF2bVZf1uK+iwMQhX+d3XujvgqeYUQ7h+Fd9j52uTOqXtKfUFLLdnk4yD
jk3rbLWgXU/XlHznOcvM+BIF3x6aNnlrUWfX3xIzO9R9D4oX4HOoWdnGsDNxIrwmEMGImk3dHZYY
QLqyztzbUZ17qhf2tuttXMe+rqP8Mzrl4HAHB8XY68m0SlXghiA94WPhd0WVP71wk7DrJ5IX9fGO
VLdNjupxgI/jrU7r5nhmclRTlnHeIAhL8yxKs8NYp5vzMk+RXVyC9xtDeIjkQ6FNuusZt+omEA0a
8+p8Bnh6mC8f9CUNSYDr3hvxtZ11rvWyqtofGtNCgLpeYMbRdmClZ03Kj2K7OyRIpZW7eeFy9ws3
wXFhviOKmQeHdCB75hJW3XHwq0UZHldQGJkybpK1pD3KthSFUbhysl91ZwMc8nFmov+3+7qsUsM5
b7lIqcCFuxlb6A0flT+ypo4B5/0MmLYK6Cw7zVIgepASwO78VswFAQ3VvGTq8kEhOmFeQA4sViBN
c5UzG0NzQbFH+f9pEeQ1ZERTyyb9d3rwzVx/x7Etb59L3+E1oJCx2bNJKRH49P913J095T9R+OCS
Ry1kRIdIUCrEdjkbbyt+VdD9uznD11ZA/bHxRvdEhXtH+DfYllu2JmQysehQCWJFnPAbr72gRPhw
MAvXj701rVOXJVs8Ll5aMsQtmzm6LRsj+DV0kgNv94mXmSaXZJqqJYyZ6oGXIQqK8YoHBhjSGZpv
uADnhlwD7dXV3/rn5aybv6BIKTOYtD4kqPZqT8j0bnnvM34mmGzYFwt95yNaR/5/EDLIUGFrHR47
YmB+5Lx1aqnkVWif3hNH91BCvJOv8J3Ut1Ll5LuoTMEdRVR298zGBsyCC4kerxTSzw4GtmFF7uHf
EipInYHUTugdJJC1tgR1Ennl4N0lQAVPE2Lr70nXVS9h0lrwxi2Q7H2i3ahezkqmPhgprcZnblMz
lDF/JSxr52ahott2C/FuMa4TB46xbra39yZWFVcOkcmYnuP18J5vqLhP3N+HjIXXNF9CnYaMdFTP
AlxmA1lZBYQRAeKy7kpADQD/JK2rSgs6OiXhjA1pE1711y+T6QM0iD01nnUXP22dOgjqZVQXAr1V
2w12DyaL1fK284sJ+W3BMBGhW+3hzwU5ZMrPPaZnDYmJTmzzdIQ8BCSIdoPmgVL/F2snI2JO4Ghs
PaNBhkfqB8XggXkVEs0Sucfou0gEED+ZgXbK13LK2lKWgLKJ1xG1h9tPFuWteC9nPkkuBSyzUIbq
Le9FcjNq9LJCsoqyQLuLycZiqanJApaBIw9tPk3yEkaX3+w3NepdA1NpZ1l1rU0mTulNeoKVyGrj
I1nZJcZ1YvMtMrGd15cTJnAOc0OZJef2okYRhKnDwS1CpgfvW6wOk+uxR28ERygM1Kt0Nk9rJS/c
+BSSe4mWEb64XSpiTPoOVxwgJU1L+/C0D5N4MaucuZKUFhX8gQY5v4zSGoOUbaXkyFrgz8tQjuCb
cseEHHWnvGnJu8p8/L4tSJKCet6/SNhvB8HJAo4j9tbAw9Dadp9MtYaQqeahlzy5TSWL2AH/Y+0A
mKM1zGLNGsPZLHgd+P8Bp4/joQImcUwB+TI4lE54AVTHMpYkuUnYNehUxjxrsOKd1w9Hd5XZ+/mG
4X/e8mQZFTk0TcggwhA9l4wZPZiLyuApY4RFHocyZN84jAnV/L1Qvo4fUD4edq08HGvA9PM0Maav
eUAtZQcRH8b/lBKyUlwOLaO2rMBxCuRomMmWYRZ3is7GdSHNNnE+e/lSGM2+DpUcktZjOOEP2rsb
tXbrKEOoZG8wxnTHrgt8DROgD1sba7edU8P/NAIpJqCqRn0fgGGSvNfGZCzlGfCSLu3viibhZwC1
akTHwHz4BKoOXywKgQy8z+KiBcjxcYLIK7AxlugduyBt/mJYmgWSj/6u/ZpQWDf+3ktYjvl6SjKb
CInZkuAjNqGBENHZwLMIMeq7x/eNUtqnKkLmFsHt7mgAxAfiB4WX+1eulX80Kq+3z+XxMH/SeJ0h
oJaJGQqQY+T1a+IbUtBLxb6caG3kBc3WZHpntAxDHr1BRpkti2E0Q9RDuPAuRhpatrP1iYKqWSU5
36+unbRrKXk29GaxrTFNutn/DOjysNjyR+GcYA2h7kDeRmvcDPc3vh/vXLl9TJzEKPZGxf+Ew11b
OHdsixUxUW09DBnPTA6cwiGyigxrMJOi2U94FFw89YIf3CfgbJxi66m9IX716sYKLnqNztG4XNeL
LXvWBjMzRO7VxZ0sQLam5X/GLjkrve2cdDse2k+3lTvq+rG/AA7WIbJeY4eHuPgV24+z7kiZcdUS
8QGtVpc8QfTh8Vb5IIpndE1ExA7WG0VUDINW7mAYX+d6jfth5DWWc5nI18B0+XBRl0BqXqLEF1B1
0qOjzfOXctFho9Jbb5gvwg9zj9jIOv7yGSxE7TNPT/SoLMAiiGuml+d21E/rAQ9CsCm228y6rUM6
8lWFejEQXwVyrYmVCcNomYVqzfTGsLvKFoPm6GS8PJNgTAHaabdoxDbLvFnqfqw5EB/LQp0PSWsk
dnK7g7tTcTV6EFkpX83ijKKbNTkJMAjoxNHMz509o6OwImr4bY+Eo0Q7OneFSYt9L1A8s1ETcrTs
q2R/tJDHzFbuzZ85Rq0GW8Rj0OVy/0JMihBDWTGQW98HjbLhoXhl3UU1klOhaB50/qJBHpFclx84
ApUAdPGhCwf7Hq8kTTfotApSBKWzt8gJODR1JgLmWFCHXZESz/aE3zJ8FYmVxR25mcrGlI34J9Tl
laAM0abQO+kRMhUXwl17kAaN0iS2Q9CtZhh68dy7rW+fkYRuAXi+8YYI+yTdfOz665sRY8+PjSgO
qXPJlXwIllNI+6o/FfJkFg25XbYQt/UYTSPjbW/oE/jzC+FM2yaX91XxYK71zcL8HCQZlAM5i6j2
RzRP87tlvCCp9mglZnQN5KwUw/AO77bpl2iNhiJl4ha2n5ItoMitWYQiCV8osydshB+6ru3m6ITI
jNYLPnVqN2HOWJ3bJnwPXVdHJztV9U1BXs2jIaMsppt9j0/FBJP8Ts4CAfEPTXRuzoL/WWmYT0Qc
MmCI/U2s8ILkhSSaeMQn/MC96rNnIcE82RNZ5L31z0ssgxef2xpemdf3/PkOiAO8jZNH4WrsQs2r
GOliG/Tm4ANTS/IKlnhNywSS050Zz04JM0V9uBOwdi9uHEJNqWR49cDnOi4tLtZ0HaM9yR0YLtai
DVXqgdNcz7t50ZWTQkJD3FO0wtfuU4gX1HhlLJHoRp08jUQxfeG6AqDHYXJHT3EnGZxG/Qt9iw3k
/DIvb+OyLL8ORgGn/BGVVe7A6KXf1VzpgWo2NmS2Wtz1K8YZkB6yxqOQ2tKIlFYxWKV1AalGupwg
eZR2PUDQgJBnLCK43ztsPn6lclxqBnKcHcQxsDydkITzUB+Ez3+hOmxqZvMNaVmtyLclWj1szSQI
Q9jh+GEHjOGY24merxV7G7lptxoXYkWK1Sa47YL6FqfczGhSr4wgm8ODT2HRlnJ7mdxvDaZmkRUa
cUP8EsT8Vvty047cY7GcEWzeoeQTzztRIUz7peggtummwIjcougM3yZxB9BPs8ehPAIkFN/2WStZ
6AywhK2t9JsJ2qXdXUDD2lybKRxe5pGChaZYXFlfYkyUxiiiVvVUKp+M26wMyJmUzMACG/OQEvPH
zRxkWv8gbadlzXT/oP1O9D/JBN4LCKmWz5OxellgkgO4yClissWh2KxF5iJFjj8b3/pw64vLchXi
ik5eHm3DNW6adApu8luRSAEEarVTwHjRNmd8Y6/LtGFMXWs0e5ABxIQzkUpDcDOah2rXb9EPNzUb
8YIlmhrlSPxC/8VkTA9Y78livTyNQOZExV/9YYYcHpei6xPzTqD10A3teVmv1lNDRNCV+FnKOH9M
yltGVChj2/GlzGDln1oUB2lvNkJWVsQM8+ft2+OEOwb43okPuoWp9UQmsAinJN9OOCMPfLR+8mgo
ErJ/rYcLMakgPjq4GfCesAIZ8izYOqQ8rc2Si8jLUl+0DKsylx6U8bMRhm1z5eTer6tny0wmIXA3
fLxv2cLzLXsCgVqMKA88MXbSNS6H2hk/lCWP/qFLNuQ6jvWLD06B6oJ5NkpKYuK/E92po76s0kMn
2V2Kkh6BJss4wwPSUmXNwK1DweXnFf7BC+psFeP7hQJj2ktQUNxqWcOi4ECMtYJMr/nRDFVMhj4f
nrDDVLvQp0k48gbhajSlM1H1QeUk1leoQo/UmqBiKC4V5m94PVychhYW7jnUdV+RgMT1Ax017xAX
s1bdgc08mzTgTD1izFsW+G+7yCi6nATB9jcna7Hqbn/T7vD1UaJ7KMGsAnWb+ibmXM+H6ToUiKMs
2uQwNG9VVU+r/APl/6ha8ourNLCKqVO0TnHftuY9ifkvr2TdpqnvYACLpO3y/XFTesukHg//UA79
WvTYvIsAascUKQGVZpdjcJfW+itGBYD/zfrEDIS0Vu5Y8zI5Vqqq9BEgEGNxbgVjQ2AWxL9YYXmI
N204hFyW+TUIXBdhdoxQ1m13RGlBvDLEzVJ9O6olA6BJxAE5ERnTA+6rZK5S85ZABFlAkx52s25K
FHS1jbT/kC4+7phfInRI3x1QKkDCgphFVuR+UDwg0ch9XiYyFkURn40t8DYjl2L5n1vdpJSK1b6a
tba/VsfLpaha4q1cN5EX/XZUZtrkgHG6aSNA/MgG0RpEFt3KAXMWMdtyaQd42eYYOrkxH569sbhq
mbJbT4Tjbu9r8O5ADmpzN13ySZYZO8nVar0iUEgdss/VToLEwhXFSYzAAaR1nlVdFzdcDehv7lrZ
hSotxUU7fuTGsDweH0DSYqSv7DyBQahEIem4vrdEVMUt3HFlvQUAUyw5tRfNj5Ve0U9bNNN4n/G9
NgdSBx3PDzN0UV7GXAiIJ2LTRxTaXcHHCtEgcgGRak3E53K1+7rJJyPEQh7MbV/h1TBZZuuhI4a8
GhsCwVDIQhUSF4b8A5f2JPv5GXjo87MyNuXug/z8Xfa/5LpnCIaX3uKz3aBXsQjdnSg+5gdttUX1
yRfGXKD1mAsfn+V1Q2TklFUepRFzmHfAs7LXdeNNAskem10xw/I1AIw6k9V9Gbvu4YFwuyWRnOzy
O7kzOjUGodT3uFd5/sfaySZXFLwGuE3UH0i71Bo3Yg9p7uceYUNI9tgPdkAjFxzic3va8boA/Vdm
OJn6I56HW6gMlBLXtYfKov0Nf8HlXXdS+ahFI9RS56VfcFRokTdnmIRMavz+UFR3ObbC3AMv3zQJ
/js7gALrjkwugQfaD8in20OqRRx1iTd3plTX0jbu0B9ycaA5UUQ8sWrn60tXW7r1AopSuPzpDRi/
u5NcCqh487aS1dbUnJLUbjDJ6tBetdrxEq8h+gJ++ygDKX5WMOsdLub4ue/xpG2pWVVO5AW2iSQm
m2kxaU4HsPnEQH+Neos+W4qG6jVOhWFXbkdic76FFRWTHzseWL/KrSs4tbf/jf/PU1B6g5AG4hyv
rDRZY4hRJ7RN0WaDH0ZaPbRD0wXPKHWIS/dkT56JwDGbhyGmpzf5u9Wv0PVkbKyt39VfsD0NvQrr
Kz2I8uS+LLaZ5tUC9S3na+6R63Yv9s4cDUgMyTp37AoxNPBrcBNYhfbnD83BygeD0qN99Cy0J0Lg
VHit+AaDMtzNP2bDo5bbyBq3AWiaUZFuxdvHjx9XTv8DZrqoNFBToMeHrHJ7bSlFgsTWJ26/F8y4
MQrIw41uyU4t1xH3UeOqpc5mjgV5yuP9w+qyEc3guexmAVbLafQzwCHQbaRoxWMgkdROEKMzEVJk
+53Q4U5qUzUKIcxLpy7UGPTVDbTzSo5u+OotviWDGYGU/asT5jZb2rdwoY1ggw/gw9KpJ9tDAKtg
1wzxaJTgV20CgsBePQnBhsxN/XnyxymUy6bZzOe5R31JZbfUVQnZzMXzyZdOakK4IryB2PIHCBpo
NGnnau8loja58eb5ZUUMKDcwdWbtXeOMAzqs/z5U9Iq65Y4ZxOcMtsNTCe8+jNDxqdksV5qK8aSN
/GDEo/eH0Zr4eqSt6ZmUgbiG/jza7XqInl931K/JQTiloiItRkf1POm+3CQbVe+twEfzrTAG1e/X
YlMR8eGiLsLi3Q5ZtC0DHhGni/BLjRDT5pMCh1U2qhwffozIr1VKyIMFImxTf5GVeVE7IYaTwJhU
UDC944c8Ao9V9SHeoTGjxFiBnrlbu9Cp9RDv8sIK0UIL+5mr/B2iytapjyNnh8jY38aNnLqfcGEl
G54rlqc+Zb+ao283GX2Y6lONFCDFO1ZwsQG9BVIUE+gnrS3UovkpEMgQ6I45SKJzSCCXiQ1xGaMN
r6sExHQ7T0YVjSnJZvgS4/RcfCNe9vIaei4s8gaeRYZSWIkbN8MTW9geo0rfIweTygRUAhOaZGFr
f3T0m7lLqy8iaqZWFF3d5ZyIiz71ctorisyHUSoyypVy/5eagNvzoktEFrrP/Vt84DK3JwK+6Zt8
8/YK2J6hEgEktc5dHZhmA6IEaSiit6X/IEHCD8E5TV/m36Pm/3SxYVQ9bkWj3uL6CM1Olkol+Ge+
Jl83nlDOL9VJ+in2q76WbuWX58KuJtMq78ETZwp1duwdZEA+t+P0kUoE0LTXtnzVL3t5/HpmH8kW
Aijw06MrEIPsKGakUJjw4k6C9cHjd3o7D2XX6nP1HeNgnNl+lO23dtZLQLjz0Jw2A/OekeKpN6fi
9W8GIP0uWGj5faeXoaeF8QCnyq8fqPkbQ2TNvwvt0wRTjgKswFXlaV/LTsVXEBIJwoesQFnIOFD8
t+wMaUkKsX15qhw0XzNgD7wFRKsd+LwpTmrijRYnzeNdcFqqyH1TOO3PimIlFiuLybKX6ACS9ByQ
fB4i5N7NAEAGMpV/SQv5X5qv/bOm/8ts3BtSYHU8buCgwcgfYFIeXTxFmqgoFJoalW359m7Xb0Ww
/8257bTdAvuf8N51s3mWJfQ9Y/sWqGPSOIzIQggIjTC+/S1iuM2dgVq9n8+UwqRLZYCt6rfUtw2Q
VV/cjdwI9AWRqMoEKwH/f44A+9IwZfhx/PtsaMVeiHxzbvVwwdCj+TNwDRX/g1Pa4+wC+z8BzM7P
ND2MAUgRbTCzspS8DH1K1KyJR4UImuLBmyLts3t01UoPne7ZuHsbAuV+d5j4rUHTImtexMe/fSsd
RoNYeTf7TPLSfmqbjin3cfVXC9JTvGeT0at0YOqR+mKX3jBK0hNelQIesUb4//KqPkx8RpRFsjmw
v4R1RUKwHs/mTC+Glh6yFnNtB9YGjOUrZlhy9QNt4prZsPmvcULwxi1Whl70ZcUgdrPe5zORFPE2
F3Q+iEJGkWePEZScF+0BBS1qtwclCBpV9YM7VuE7qHaeUHH1Q1hw2ivIR+Nc+fyrUn7K0MfBXGIU
hhqiIQ48zeCJdRKT21SQFBvdoIUpKjUabCUWc8Ui5t8eIbgcgNg9RAT5a/nehkACEPukIv0V1hUH
9LM5bQyXmydkD/gqpC4kbrXbJvD9BZJkdEjOX2d6IVaYDhhITtzKg0V++RnPBx8v+9GJ09O4ptgN
kyN809H/TDPAoMZGkIrAbEf5I8ZpgdC/Hahc4/hqlEuEcL+8EH4ajVC+gCplieVkwnErvAcVOr62
VlVSdoBvJZqlz2S7sZgeAXqcFQBSust0+c8Z61sxod5tJx4Xy1VOi7tMmSpgmPw1IyBzAY3O88Aa
Pn/7gnKGh8RaVNR8IJUrPNnG3Nv21YhnmmMKKA6K6YcmmAC2r4Upu95tCdmRUEJPVJVO2qawASCB
u+Vz0/Ut4GcqbQeJmP43mU+A1q6+3o3f8kd7QE16q5JMd6ptDHaCCUusoVY4JncjvnwpivPn/19Z
+c5q43RX6DQrAXqCV47pcH4p5U4vQu5TkgsW9KHrBmHRJiwe+la7Sz98S41/Y/xMwj37CK6+myUh
ocKEeKqL0LC+ZXxzEq8evVvF8Xzea+bLWkkcF6tRvq9vSTXbijtXvy1xlmKEuB6gF56mbchg8h4e
8cLmikkQSgfQwYGthuON4hA7dkxdvoHZoTtPSXkQL0KSqv9AP3V/B+ls56CpsOb6gmIjND/94Ioe
kIVVOTE8ziH1BW5MzcAFlJlltaozNoZkbLZriq3bPT/FOdv/E1gfcISlgYN8ZqgGloVUqrgQ3RbE
Pcrv9JQ3Dwt38XsUL2rmjgjo4rxBAW46QjDgNrj1vCLdvGAiKHnq163XeJ80VHOCvWO6bTUGUdKh
i+FynLUZL1Kb7F1UqrDKDpIKLxyvRpdXH797jLsOtwUmO7UmpA2ep2UnA4/MaBofQv3pBg2wwryS
1N35mRqA/Zk4/8kvvnT4qlwVJv2Q7sknx2StcHf/slHZYzXqlyaRBtFwyRD0yaTXrhh50NsUzjUu
Xxvm1GQqlBJlQaPji11RB3yeB2j2bK2pFz9w45w+GejZm/1NqCUVudBT6VlA+DLXq9IGE+l2WTY0
PztVSUbEX+NtT8yGN/PgOtFBxpB9WJ2XWXd01GWdnXqcYPsuttEpkXvNck9gmf646G8vESv6unnw
oKlDD+Hu4hdLiiFqruLzNkRnQGEgUKj9CmwsDtF1x8DpotHbtSm4WFg/sUE3N4QTe2KKuV2T2Yvu
orB2UcE3jku0w3dZ+P+2iutus7HtQ9ord9s7GPdpNjb8LNg5nxUmzkOcxUHVnb3ui3xFoELxMdnd
/8wY9VpsDqKvxr7JsJ6u1heybwLjhcLQdsKHeicTBYiNCvi1IxQteoDxufUD9hTHPsKBTi9MU7Km
mjGNd4w4+sML+Gx2Kbd7+5yPFR3FBFrbrU4wT/UMXoORFBhUvePqIl33izEO3ZvN/Ywb5ZlG+pLe
ulNDqzDXRBYQ+ZiO6SoPOGdkj/1l68GdbSTmYr1oqgeB4atCyNgoiT3uOboGKhd0Ke74iYCly5Es
b4v/xu2iIgMBwfOprsL2RjXNmzADBrSa7M9N1tdaBDX3r3PQlwmwsz9HoVJglBAhkFYb7cwVLRLa
0VzxTp4C4+SShXsRbc/6S3Kof6NV6nE98EJ+wh5D3tkUq0UOdVjGAIEuTpqz71f/CkrnrOO0uSMW
lkr8HgKeq3NwpAtJDSyEiXIBWIace7CfvXY49l3x/vkLXa+/TjVnT8rAJ8dbNcA2YiKszN2iwM2B
TRZwyvKSoz5rwaJPMs8fKP03QgcX8b3WGuYiDvofabg4c/clnAErXOHOSRF/mE2h2g8GRwlY67rH
P9XbOhGdKYDeYA7v4gFJ4G3cWL/LRjC/b3Cw4oaEvBskvgQTYE3O4rEMuYvy1WRYmpoYYuTQ6Lyp
6jZV6rvSTAYXHrLRF/rIxbKqOKvCxAdOtG+OQxf5t1NqQnlt7d3FI3uFnlxIdhunAqwi7N3kJITF
3XbwdYcptcGg4rIhRS/72j4ZcHt/tg3lwLUXK4ks/pjkifMr3akCc626s/7ZxWk6vpv3sqwiUqcw
WYrxhEaCmF+HPfoVV73YGnmTVBL98T6+mMSqEMpzMdXZAKYrsMsX1D+4AaLRhk/INmbbgiixzeQI
Qq0mmB0Of1N0LetvWpPSL8XTHI/LDpVugbMzHs6OnfqumIHhrtndIvM4bIFYR9F/44Ja4qySANf3
pT3GMcOENRNDPW7O3qBttEUXZJ6NXyKombxDmuCtYsaS2e6oUcOZmiZi7TeSXG/ITm5r1poe1I66
MtcxxMkTjB3YxPlWiE0lGWvqIvzElC3R2AZAOu053HeCBO8G/mRx8R3hCAWgS9eT1kuv7I3pKdbT
GEelscvgYKCsM3+NfSNkWl4kK+eNxFTKH5Z/5WJwKNcw4FKB+j+y8eR3bOHQoeKo/+iytND8Wa2W
ap8/BUSPtOktGRi3hJEbKxx+fSf/LZRl9Yu5b2J5Mv9xJysYszjIdStsGvZy1Km7oUIQfxOb4DUw
LUkwThK+zQszob3Hwglp5ryqJE1B2Ju7pXeUoEGbaNKyFgU8P/kXFXEBShYnGnOXNNeC3SNAtQTU
YR8u420foczARSfARFes1pamBbfuqWm2TWy906P1xA7PNUAFu5m9aHiVYWxdpegBdG2DL9JcdnqD
p2ohsWYwXRTud/KbpULAJW+5JVWdxfwqDkZlI/j2smCcmsllCBNvyaTlLpo6qNxG9DzCuMph625k
8ogOn4suWn1f3mde5JT8DbVvV7MDH1TPzN9OMior2tvhfm5kdLaOmXMY7jemJnnyS6DKTSJU8a7f
PATaVvm09sYQ/kfbV8Onblo3a+e5GW4/TaDBN0hFIFII9P69DXd3vdF4bCOAaLIGP7g/5K8Wxbnv
lFXOKd7UMBkZt2FH77JggoVNJOwwxOJeTLVLoGxuxHEtJgO5HBXV2884xYDA/Z/AGW1ppsaG0nV3
Z7OKi1/wIAPKpi8IhQvMJAkx5iLTMo/I5bVQTDAPMT+JPQSru29/dOisANzTaxl+DtbGGGqdjQTi
oExjaUG3Kxp0RtLAMLz/mYqW5bllNrzfxcGcf7r5LobrX/JTfGs3STnq15xh/iZrawR24m+5DSe4
+NrJ3TdZzKei//h2ia/vMo7sLOhTG6Hxe36Mrp1Wx+uotGsQ11w9rbKEfhO7jphqz/eu03tkmdYz
zmxJXpLUSSNISx32FeIJpeXB9z6UG2NOlVG8MsHxy3O2U61qmQ0a5Dewt3K5p+jPNDn17bvu/Wbp
DMkiYY7PLHan7BmcsDSXpSXDyB9xM0rj3yBZ054VBBs5sa61ZORPR4vgqTPAILZ9LdzZiuD2lLBs
nN4VmPesAqh4HZzK6XwiY0mLox4cMuiMpJVs58K0IxK1NPTWUIEQwfOAcW4OJJnmTrfNOI/RBDDD
a8pNBvH7pMzXbz8QDql8iZS4J4JzKG3WLyK00xRdF4Wq5JWEVxGCptZPAJjrpXw2Z1WluALoAX/K
7uPVaamXYbJhb7/VsSUGF830THUnGJYTUmEoeIMAn/AicTSPsk9YKrv4Q25jqpvk1KP+L1nj4c57
Qu4Bj1biXRM/A5o8e7voNygjx8Edfg/UHtF11sVujGSteR02V1HbuEanxoTWgyptvMa1F7e4HuXI
4wJrD92fh7nkRWIj1AZabiSJH5AxX4qPJXjBMIWDqugp08NIQuuYzOIedcKOUF65Kz3ewiasprzY
s0iSVnIrKYW9U94Bp3owOdTFODJSLEYqKz6o9dwttQkUDjgqoDRb3PgzTb4JPU67vF31VyZKwSfo
tNnNrCOcDAqI9EKBAZRU0fEXGVbP6PlziimraPChuaKEk4ewSATEtZMd3f2f4b+nHZmMWtezEluZ
UZGmpOMsslWNoWpBtBx+4au0hOm/6A68WLB7BD4Xq2yqZIHZpNAMJbecqzt/oUDwTPO03pKg1O/u
zcxfuf1gsBhbVTQ9TR0aqubnjJEX6AoGxwtAtTfQPLf5108QG8nwoidXBt8D4ZiOxBBCwbpnM2NU
Msu2GwsQC8Rdws0pyK6pp8jjZHrH45dZqFPDuiU8+q20+vJPrn4k9YeEmyEycb5oyJm12cSwtNj3
Bxo/uIfhrxvRtXQeccLOuM9bTU/w4UBPlEeFogwhM3tXD26badFLJyS1Bw3sFKuVB6I3FVqgta8i
e0eioe22VW+5rd7Dm7yjDffn1uzVUUuhn92ghzpPhn2UYlBxaNBCcx6VLUDxNobH1cjfr6PySSka
vQUFKjHensT3buZKJO9N8yXbKcTyLY+zV+ACWUL+JxIpQZjtEJt4HuhvJqBvXnaPfuzdCwAl9M/L
Spl9kCN9Wt+DGRNSg5wZrizxi3fUgan7LPttQ7uIe5+NL4bwLmvUbeTtiUCX5fOVWuwNSlxmpG1u
ILJiI3behi2pR5a02uF7iaN2PWUzJnbNsMNGaIAdz1CFyXRzKrRNPrHxI/N6lVkTN4K6iYaLpNY/
aR25mo8ksfWsYLZ6ge1BMze28fgjCb4Qz6veRYLbeDKDiyYJ7/ZnCRcrrG9+t7bp6ntAw+TQFQ5P
fau/LQesvi5wARZIR8mKkLbstUAP7TW1XToV5OmumynWiPDK/WFNXOuqBHzHh5ulHmC81289xXJ5
mHy8AZo0ZzRmloaTruDWb+dZf8md9p1A8vMxvdhvxJA9NOvYubGHYWa2DBdTICV3fgN14LLAiliv
yyA7Uq3WaJN0HN2D/VqSAiu1tXGFqmKmMA+PFlBjYua7h2glBf63Xb0iHn66Tkciuc/pYtzWH/VK
7IVOJXikmfunwmnQbKDXSobPdf3mHfCc2H2shL0vSxPPQ2aELCku7fIWMmegu+cZpzz0NOmAKU32
Zp1wHaNsHeeNiJvjvQpZrCUKTDqT3OCwBiKL5GborrVeuGmlLO/4IlsqqEWwittL8K0/ASQaPvsO
aUO7hmkEvPDrLF4pHPhoZNsyQksdwL3Qh+9NuRDSH1zthrQiKntwRruzen7xYoxpRoWOfyWHAKUN
b/e/eIja8DbH6Baa3yr+DCmT8qgLxqmse2NE7tvb557OjD1QDVmVhhhE2DhHxxWUioZUIYyhfV0H
C4WQO146fihcIxyAnvi0kCPSKJ6/bM3h+eVUK0kvIhAsBGHvqX27l3JoaHgEh/J3AbDwIZdeMJ+5
7T1tnGWA2YAA/BFc/SwHy6aT++NM2s7LbjVtAG0KiEaADoGERhm6E8q8AOF9rmToJTwhAvn+Z2+h
LPIm1qv/5jXsrt4W3fHOOptAD703olzDvYfyL154f5kWq+68jrqVetA84KpeDxtINjqeFTIj5NDg
rQeGZqNMWLzQVoBdsy1DICPQqiyuZug4zcGLa1AtJP2X67gZp0dans/g9FKKgdGCVD8lu9Bc3lAM
6Lid3lvGPy2zN7vOTynnhrtbb4j8vupnvH/sQFq3y9Cde0MMGBK1Y4GJyHHxSWepq5ntP4Z+lxpp
RtsGMfBkIc5+13LG/oFdzYiIYZ/NXSPEjS1sAv/iQ3fjnt7lQnhyFUMJIybjj8YOWcvbdNuhuvph
IDBJ3GeQKl5WyvpM0JM6w1kTfRihHu9J5LQ0Pgzm5jAZILlN8GIyxxtAoQqrOWITIAzKy3+BLIu5
bLqJhCDH05KuNEq9Kl5tAh5Gy31PQVG/xxsE7TAndb7RxGP8wfIlJ8O5JdCOeQfho8e67LU+dlpO
IqL8aMReIOPQb+UrjygCbJs6AV+wMM7ZrJi9tKTXMnsnOB9YueJuIWNPoKWDrQ1LxPxE3yNuWVjF
168iWqvIi0/20GUZ1AKVasm4kX4nd8QsCCPMCq5A9GQ0evlYj/Idm+GJNSn8TBMeulFB0fNf0VKS
jMdafjKxzukXGRwK0YVD4D9VRVd6gJuHF6AavsF425Ol2n7YYEccB+/GG/UvblnjR9qKxKjnaLzp
hn+1Sj9b50n4Ic1IucEc8eL4XG80tEKnJ+e6jYBprVlsQLEGZXC5vZlFD2c/96d6jnnwtRwp/Lj+
puqEk4ZZFcNmNXsrPpBVlThELSEtbXNgyYvMb3dTYE8Mvvq9To/Bn3pD2alhgamg7G1DgDssY7r0
eN9hW8sESpN6/gq9iOZvrePMF5mArUtzcvoZHY2pf6sejcW3GR6+jz1Wd8ixeOJ2iycsuZQcvUOv
ljP3E6bOFd1C31No6X+Jx3ewataDr6JkadUgDMksOr/TdIDyZkhnbQKXPj8JGyAl4le35F+AmGc0
ZnRTjuXtaXQPmGZNkKiyHMouSKqSSSDUpKOIAJwVoSLXKSUe13UP0w4959ynB4QZuVtHrjjg6GkA
IRpmjwJZLPlN7wy9cuvv2ofG1xiLWYyQDx3LY/jFvNKkTatdxj+OilZqjlftH+tBJeE/PVUsFwOM
oF9FIbCKP4kYLK8ECir6OfT5W7aakThcF1UKne94guFeQXqC267RIWtUcJCTscmUdP3XZz9UuU4z
dHI4Qut4liI9ZCGP9xMEmkS0X21IqNSuFJg0E3lhaj90pPVTfTTdeHb4spNpikMHZ8Z7w9Jl8ODH
8bUA3Rvqt3rrChMeH6Ro0ExLR5bHscOUsN2O3hHU4U3jGjG8YXGo1O7DRKaZD1cgQ7lvt0Hv6aHt
Sv1ciceXRI2qP5gsfuiu6DuOQVgMEVSU+0TTGXZ6FGtq7d71aNn7GsDobUctoJPJb1y7iG32VqtZ
pHMveowIFzzXpfsWBbn3lKKXX3HoqUnyIxdUnmz/sv7+O/R8N9b4FYRKYuVoNRI1qbWrbfUyO2zB
3Sbru6RIGpHKMawPMvs6dG6lu/8G3GGF0qOcH5fLpuaGmeLyN7JmffioxA8oE7IJKIUnwoyGXVmg
CUCVQXpBE6cdE/rp2KUmdAeMWnqHxAAqCOd68WOEYjBV+qF/Y3N8rq4bAktb77ZXV9Fp/E7A25Li
Ng4wC6aY/o2rwUQ3bWxXr8n0ox/aAwxXeWvxM3LPas2MOhI+6+jw5SN8fqv23bo3LUSvvuOrfQ2n
9rH1Tk+DwHCh3x5VjibkMSROcrKVqHpaAR36r+Ghvl4w2d3zi050wB6JY3QjloWczizLMtZ5/rWz
3xJ14303fjYAb5lyKF0+o/t5CqBp83eRoqy8RhlE++jNO3ioYxmqObJRYoWZa6kp8wJPaNhIHcJC
yIObURL1VLPfd+Pc0mNRmildd3ks/b2h2htR8W6BcqMyZV/hlhbwL03NVr/XrmrXKI2giqX55pbS
ylIASvHbnFsCa78CA6U3SfeIoo6HrS0//Z/w+k5iIOlIcertlHODzGQ8xRo9azAT0SUl5s7Tkn7B
yiwIjZbDtY8q5sHceXXuN3ikbhWb0q7t1L7GkToDZq79pm5NULt5a64CMdG97ox7VAiafifMVEq7
cawS0c6FSJefqTeZvfN6J56BVMYso2uaryHu0cnODp0+eA+ZZ++hYFJa1Bm7HMwe8wRTJQwxxP2t
eOZznWIayqK7ymTzWXXKTgV5byE9rJj1p8I/4yRJsj7Q+DtUBwnHlUHs2ni9NfY/5Dlo96bdoHii
/UaSwwQbQzOprZWEa6ET+TJmBzu72Mcg/hf77fyuBTiom7vWm1SKcg65iKbFVI4dSCkOHrwuekBY
VQ9PmqnjSN/o3aEwDa5VDI5f3NDui+nicDZL2Xhwzxzffojb1EI2Nr2g8944JYSzvBb6BRdfcZER
dgjLC/bJ+TTpqDpz7F3EooI/Cdm77pLSgKWHQhXo/SjvoRpdP1JLs7JeI7o9PWyfRXBJbkM5dA1I
9YfkP8Ss/z2hiCMtS2+u+42//mauFJR/oqx8WTeZT0aiQfzE9+eizaR17E0pWJEWjSsxJCl747ni
4XXz1Xa5uoZ3oRLMD/c16rBD/8HGFeDAc53OaMTyYH9pmobnQ9B0MP31Y7ZsdV8olIqZ3u+ylcD0
3RXRo9dfEXwqyYgv+qINHiW1k2O/VweFcQk6VFAivWK+wRwxNSu98IXJsmsxIz4KEQD3cxF6SQNq
qbnOpP7cLfRZMnR6t1Egt6wFazirojkx2RiR/prAuPN0RZJPqWri8FHIfgGlTHlo1pJCEyh8G0o+
EL933TWuEPLC4/zqw46Kd1kN31FDEy5pvQonF2n4Dy7KlH4tHb6DWJFPJSQDpBQ086JvHCc8+hRg
3Un8CmemFELnjCxP2TmkNBkeYB76NlwyQvyiFjEfO4HVywwwnUFKDBfuEmR+rzyqKImsXTkUBQBg
mYDCbtFsySoDuiKh3ZXPUWr6+g/7WTHTnyrx/pwCo/Vj/I/334sZrJZJcJHHijZQAXQ/IhO4WhaU
QxwDoIK5dCulMiQFBb2K/VkQQHb+55HOMM5pIMdLK5u1v1eT3FFgZx4QaLWkGac7tHv8SU95lt/u
z6FwO+ph7i6uGG1o+OG6POgcp8XhYmQY7D9teSxK2Spo/ysr8HpIIoiTc4/KYK5iM/Jx+syc++lp
u6wPSP+X6gxTRfbBLTiIR02QvAAeiDuBlvX9Z7snXSOEkx+lp95QamLh5kNo5hNBmGXu8GFAjzUD
g4UIRJO1On86PYWLu5HNMRvuSbO0qU2j5by0xXWOWfnGbDZVDCWB3s7kqRkK05k2O6RwD+EJ3Mm0
6dg/A746IaGeX6+JvyATRj09+ceBi2kxx+DmJYhpFw1wtKV93HffC7BPRAhJOcdyzy8JiAdJJxgv
XTlDWGlARaUcpv8SMflNHvOyl8OsbcO+msnis5to6qy8XzcXmBwMLsCuDXrKd/T3cVOUDeiVkE1r
t9Fp8kP05hpgah7djjIfKa6wL4sZkxcblH2zyMqp4sGxrjd9dB/OvVDSHSpP0zRrp3GwyoxpHy3H
3d9VaM5W7fiRS1cE6Z2q9retYa7jfRgOtnhhRGKBUS6bPomGVnMJsTLapes4LiD6IPQdXs00aHhj
tpaafhluzZFdkrk0SQ34/oag3Py5DirW36LipSDdtCWIyKsnk7jxOUwc6v362D2Xhio86ryjp7gU
T8JEqJDDHMgt+B8FqApEh8P9aOVx9ndgEqV4eYcL615yxVSmxG9VGkcZzjvnyCHPN1Os6QvMW/fz
0QGbDxHQQTy39D5T9tRd7zFvPi+u5W5ZbrCDbIlCnQDM5R8noxyxoev/mPvi3+Ew0Tp9H1or6Xaq
c14O/AhVpkpLhoTRmZRxwUVubq/BnKhocX6jkbyZCbvZ7XghH+CX/XcenFK24Wp3n5N+Rxumf8uu
39aoBtH6FVh5DFKVxJP30gmuMO3aVSPuNaZguCU3OabhJ28ZH/xEszaRcSau7ELUgoGwQU6IDK68
Ijo83SFfAfczQRnn65dyYlxk12p83duVo0J/dAbDRiXRR7pPCSRIoCKuztWrXlDeMjcv37j7IokE
wF8POPohE0pZsAxIsxHlstThyH19+GmkcQ4s1UOVnjMBXm+bZP94XhpTh1hAfslVV/aIRZBj3Bsv
L5cntwT3h/BLRR95zxlk/3OTTuEmgm8r4xTMXZrEBl0GhdP+5KRC33TEeNaumzSrmhxmhJ5fr6Qa
ZA/4XMqIA47waoOon688x9KLGf2v2B3BobXgGR0Hk2CXioROhzmnkAkjVcjAUwbfMJ9QC1vxPXoq
f1J6VW0gL/4xWcoSUdGkDnNNEIG874JaAAV1V0/HJ6sBkqFzyT0GKUSEtWz2EKxKFpPeueBGoCVK
JH7bkQ170oLrQG7aX5OBgU/ODnAtyKeqg1eWv57Osu+5KAL1zJjHcCL2QlUk4zA+55zHOOCxfxWA
8fHI68Z1xMEQeUWhrZUizCyGB2pilHXNhpfjS3ihgSMYKtSLQ3SKVFi3TMPc3+FhaavtX2WWJkzN
n2BNkFlpeRGHnguRbxnBSZimKFuRS9XbYHWutrU17shbdi5Qa4LDWyCrqPc/8tj94QgpPtapxrCE
i98keEfbIjpVRa6aUHDu6jI7RyXtPG+3fxu5hSW60Lzky8jIM8p7OaeskmIdarA9oxkZiO5cMR9N
5kf+xVg0xm3HXcEvDN8gFYu4Fs8uogBqLsxEFraQrvXVgr0s1LNS1PqVAFLWtFzJEJZWGvJo08qU
vMBUFGPAWKHUZFXhyZxjzoInef6v2rTj/L//bY2AM0hODA2I1lujg2PyMfmuGd4sBgGCCAlG1t+M
vjJgpeWJEm7wbBsdzVu0Bf77HBWAHSDKg2vcycoB/g3drW/oJwBXdUjzEFctPIybnhMbInWzNz8O
EBMWKsFdfP2WHII8K1GaeD59JM0pq6jeANiVmdEisKjPBYgEM+wmOwQX39aDMkFJo8Ih9tpDT86m
70ojRsMBfH+7DVFJprrE3Kn8rT/nQvEr9G486NRZ9NnnuErVI0AE7qewPcC2Mnwmr0CUnsQp5Z2h
shGoKePje9R5xV4AnPUiYFDm2Dj8r2Q4nPjnjZLSxJiMKPyA44zDtOfbBhvanzKEzS308Oyg2i49
aYMtgFy3AqqM7gb9uz4++vXBQoXAvoI8kD5qWKaBKSeOfCsb+1Eh9jNLbntQ7dREFFllBwfv2l1D
GQ0ANomEBt+wPDhSPQTcqxZ1kvZX25c3DozxOp8p6wzspdtaW5/is+BvzQeSNvl1NatfN36vP3uR
2JMX2Ufwr+6Rgs0WS2mOz2o8cot1F+22aXKTJFGjsf2voS59lbdGuh0OXX6F+AfZlAzm3iXe88zw
LDmK8JFth3H4uwVixDj45lOGWMeXe+dOkL8F8BgdaqSG9C1tW0qksEcrCQi68ajSYX/071dxKiY8
gBRlc7J9SpgkDmSUIBeJ98nxHj+FbS829dr1ySzn5jqVklWb5W78qq5S8NxaWM3gChghNOPiSFvN
j2zXTJ3PmPyIwxpnTd/Xn4xJC6gKM+ViBFGu7pxMYu39l+iYeyDQMfb2nhdLcMJQ+G418JJ5Ft5B
u7+aVPw7+sm9rSgxfEETm5bJYU4kVjcgld89aOFNONsfFziyNh3ViLK81FNu/jtGDuqhQ48fXKoL
Gko/7TvH1bO9vtoVf5MlcqKCVZnzwXTADHji0c08pYMY/bcL8cJCOntWJHB2cRliv1R5nwIKfWco
MEedaU2JD9WAJVXVo0wmNQGKlzSTPX4iujmzFQbznAw3nnph6avflB4Kik5UC4EBy+kHRK+nHFtd
ejE0aE1goLzSm6VEFSTgVnLGJUwGxybSxAJUbpuuL7NazuBWzpfPF07EqFMLWqAu1jhYkWqVJJo0
QqndGv0VPkbAa8yfxAOM4PPmIOtJd9/bx8Wrbsei+3xJMuHtNGW7PlfiqVKy04YIebpUdHO2MIQ6
suohcJ7KAlVRsuAtOjfe0SnDkohoRcPuK0lizRGH99OOx9W1xWnS4dN5ahA4dS+042BCc7XjoPcD
qLhSrl1qwyp8Ej5lqSSvmNeeA0ZnU3n4YCJcM80cbwGj9CHLMij3jVeJv03AuQxUWDS/NxjdKw3C
8zXVEELQEsiW7kB1eAsnu3KzeYMY3V5TI4GqJvjTodA5Yg013EcjcecII2v70pwYL7+TvYME/fw2
AIE76zUdQtwALSHngkxj6aGtx0YuDw5TRwG5ZfMS2gE/gASlk4mF5PMlhJyvEXWmFNP+IidiKQBG
74dSWUN8/Sx9GazwXxoLAM9ZgInBuAh5blsSghIzdTSGYuzMFeU6+hfoZIXydkRv7CwEivs7QZJw
Aic0kaG1fXsx0SiHwfjfr76LxSVnD/Jt33GlWjGxgDNo5LG899muzv8GeAEdNBY9DFtXqG+IkbFz
zz4RbmQQHTtRu4kfGOp9DpncisoFKCDLpy4iulFpsJc97bzrWPd3MdHAJv+f8+SINc8UDVL+RIQJ
7N/A7L6NrNxpALSW/Iq/+ZY9FURR+Qx0dauSv7fCfm6SMIBPp9zmM7Lklzs0R34IWS+Z41gPc80a
q4+Tox1fsPphl03OK682Vsy6ZkfpskZ0sPBzqB+Cq3M0LLXYi2LzrdjK5RB11TZGuIxjz+AR4DLg
sO1Fvkf187cwNRp70hZpIK2TjlaDzy/gzu/vr4DF5+laeukx+leDhgSHIJVslbvYsWCR+NfbWGwq
28kkyRtqZNb1mtqDTPCOMumUB5ypeX9DZnUYaxRRWFyKqbLRNKITZXuD+5zcD1ZnBb3RFAPZkjnF
iyI+IctKmVn2cqc+NDI6J45EsuVzBkeOewAAOxK+RFYBMOBID5+rO/zRFtg+eI2G977i9Lq7/NE6
E3J10pnGHhw0xnjicHM4awmt6EjpsednIKUPXJsLeUExhaxwSVskyUptIi53vJOw2WjM/pLDQ6GJ
UBWBdZ8acEOSs29YQG2n1JB8lQbelCdr1B02POdFYQY0PZl+piypmlxVMh/2UunB/5zslfW3/Iw0
dQEd+DMzAv0u7XmlqZEq1rfuwlEVvJkfE2Pe3dIgmu8Mlrw1CeG97czoiL8uBq7rP69B8DoGibtL
6ZRcLbUXxDd1AvEpnOt/vKxOrilwqZZcXh1VF/Oo2st72QL/NN5GijfvKClSszv0OCjN3HK1oUNo
dDb5cSJ0VU9xpdJrz/V7KDVXSmwHITJj/yQR9X4CuLVFfbbSGEkruqPfLP4jQIgnn2IJxzK4kin/
6dgHfVOC8v7kg0aaJsqrhp9wDY0zXfiL7aZ5ZNZzV+xvW+244bl7JEA50UZgtSQ1EJbXO3JVhKNe
YcXfA4LzSU1sP6Win93+T3Q7RJNRTsqXPdJ6uhuPnRNJPp081FsnfQbRhzyOqt+HrAHNNFDLpCdk
OgcZATbDnZsJ7Q4xQqdFR32kxebjuzlNuBknO+uAiim6dYRl0CrYkXVQ5kwS6ES++dg3f/6nla9p
qKXAlUcZ67/OYepU/Id4JlfRXCkOE+ShbaLKILhLfWQbYqhf6hwzy7SE+7Ve8BHrUanwUxjrEWnJ
MEQ7G9bZIxio5/BmKoIny90/k5R75U/MPvJSFrGh3uggxS3LyQJXoitfZ+Ki0SoKQUO2PW/eal96
OrWVgYk8PDP4QWfEg6c6pFYHAkB5q9MsOEqFwR2aL4CaJqXaoG0FGT++X+yG+a2rDGpzigzUTbeZ
7A2jd/a01ifkOlZPjnlV/Oxi/4+meBQ12HF3Aob4aKjsLYanEjQwKavSJK+N5HFLGayv6SK7aVeI
afo2fZOytUxN0i2k6cOgP2xzQS8+wIcrXDOharXwblCsolkQ5FyHYUDP43l2UFPbOzrR4IrNg2zg
xVB8oUrqbhV3Wp5pNo0E9niO+DHvStj5G4OuPCCJJLDL/e52sqQbm4i2ZJ9CrPLSoPsU3nUildx6
k89ouzbnvNsmoOC8JAn9VnGFSvs+ERZ70JjwLCWSXaovhMc7VE0KMJ3uvXaJGIV89XJJhuZE19iE
cnKkwtRmK6DWx0mDF859v8CTjGVySKZPbwz6/Cfhp0EZz++d/CxpDQZbNjnCp/WNFZW4OLDsB3lR
lpcHXIVM3YseNmLw197mhiAo+Acdt/Cfmzc1Sa3HCQN+BI8LgaCpnfqHzI0XBX3DqByXFa+YapxS
wyK+lJ5ML0jsZ4QBeigI2ds3xSwQzdzAW5yXegBdoJ7ansQFxjmeakHh6sqnPHDvBpDHZjLHWFCy
VRzHMMGPZysL3sgp15Y5tSxkeUzc+tMQmbOcpdmdhFjeg1WU2MLZb5bHH8I4H5V4BS+X5/lCCAfn
SZe7t5+0gPzckNRQqT6Bq0bGnNBEbZeT7pxqud6/KIlLG2ixVR+LrmCjXpNmFy79S3L3Sz6aEtS4
eAZ5tOAw8tJhUjQHt7caRLipK37GsUwYYm/O03BqjNOfynBT8neLVFq24nrMdL9cpVZlynSKnKBo
bi/k5d7SLerJcES6wMg1YhGTspUAqfJOmrQMgH7zwBtcIa1n7DtBVb8xrTN6dKVn0XFnE00XDkyT
Edf2zqS/XC51oIjpWjR99OalTJJfCUwVbtQevP4f85qDk1A+NxKZ5SLpCiYIG4EYYtivNrimesOS
VAd0HaUe/GOWiCoko1VrkQXDY4QOwThvmb/wFvD/UKI7CUvJMkblLBQawNOeNMpOddnfABIPuDjf
Rx55VhUb38P+MCOqkQOwsrvDdpC/aHPNQFu01/S0qeTEID+cM+qQ11lqb/Knxcxt8FIOKRyiU1op
zSQtPsLcMWuLnRevKnMA3ollmP5TCZR2RYRZ3l3RPjqUV9rGZ+o0bk+KxvK65Yq8yrpnuo0hxgyV
Bx0Zito7NqqfxbHYe7Q+qFH8kMUpJKw2TH4YnYQG1sgpUWdyUPrUktj0ZQs54dSlGf356/VIaywe
BKTE3vNC43DY0lpRrVg4f7cVxbzf/4SvGMFafdKZdcqAZUa/Jjmd/uSP3NhAl7MwTg4/KuT53jP6
Y2RD26PNkZfqEIMO8Xg8nFiiJALQawZVJYYXboU2cLXan7YIoQCEuLZuHeSGOTQW1Es2Edk8UiWf
yE8EVTCGQOHDGV66nBHwHKYaGqMyV4dPVEYHyWVMIhZ+IoHyfIXAR2yYR860x8rCDKCbuLlzYVXu
ptmg2FMtFt7lLJej/wVWG3V6sEpN/Vd2XUayUO3kemQH3CFtcsPHcZAOsxpYfoq/+SjILhXk6LkN
qrnFn0BYC+T6D5zt90V3fTOmwPsqnWqvDcbC8VRDq7cjuWW4eEvWoxgpu/a0TsqO9FV+aAslioq9
5kOVvpL0Teyl+t0UIyWIf5UmMcoEAVJx1ac8k/dMukjtVOSxX2f6x+xuNH+1OdSF2suxPINGhlkl
4ezqSfwyR8ZpTyqxBHe0bU3QmugQMZWoL1XDz3xJHANAu4Sl8WPTILeq9dgqxoXa2bvITM1K68Ey
9qxRgEofMSjmXGptKO8ytp1t6lv4ohTGfAXQWNlbTHCy0+FU3qfxKZVG491nrJ7jGbgjhHWx2bA8
/Pjyb60Qj0RxGqu12bSG3WakDi3Se6N88l9NJiof84PLRwL+PKmuKXSNiI69Mi1KYht5xiDMcNmx
oVfG+SRD0DvhbKXucEkxut6HKHKrbNBLdpSseWxjnZMHb6KfA0ARbGtbyYy+vb349delLWMKoHgM
pX1uAItt9qzdybFDin328IK7/KbI4mmSMlr95sZ9r9CL8483vc1c4snBvJg+bUIifQc6JKxayk5u
dqUt3QAegpW5spZKgwvF4bMgkjivGyroIKKuxdn6dglbfLlBF2nMRJTFXwkSKK2HHfYXa0JWGnH7
BVIE92O8xuPVPCYq5hFbAjLI34EH4XCKEucmhnmqK6qMz3gGbseW6m+YiDh46piT2u1JXncNNFel
xwEd0oXcicSb3BdjquMKJdNiJkx3YJ32HOB4Vv+jk1CMI3OuZ95tGjK8gEjABUZ3+Psc8PItidXb
wGG7dixf5IDdMncxEJy1MgT6lpyv0Aox0Gp6oPBpwAG2UJFd/7nhp01B5s+gcGfQ1oNvS5OnoMvB
SVURBQoYvKeIQmVbhPuVhj1rXVF601vPdX6OYewYZt0hXkw3BrZ0MOzwVYPjVpXXmuVF0Et4XO7K
0Wmx3zVbFddFR+JrctX2t/o6JoT4A4t7t8mv4+W72o89iHNmu1Hc8smSbwrD8NidZ0asCniQNTcc
Q2ysc7m1i2RI/M8g0TCQx13HLxBtiOV6y0gTPMe+Fbh/+RyAERX7QsEx1BPVGg8A5TLTuysNnUh8
Yq7hKhL2tUNhVaoCP+EnTZf7rzfs7FqYmBEQwG/LdvIBAA21YV5f4cU4tP8RqYgFbRfA+YG7CC3C
dld7YIALGGbOot+/uSMwFJrfu6HAV8oNuF87iMeIkhx2BJrMNsKnJnHnhGF+cMqL5geFS29QIkBe
MAOvR8X127omEwnc6Nuxcp/w0vlSNhIVc8GjygMT/bCSZUzp7M3hhiK90fJOG52bMk24cgNHPJ3P
GVb1qbTypwJg1kdlSYF+hmRKOBZm1aOiaqpzdsKsZo9dRhH1U3PeJBDtxinC6pKk0F7Q0ylYLG4Z
eKuumtTMaxo2vZ+jh+sMSn5Iu1otyjUlcprQy0ObKC56YOafZiPGvwgfoTCZ/P6DdUQINdS1ygVu
I1qCAxBF1bhnhqIUJYUH4EyMdl+NRm9QmkmD5RS9IDQzEbFghuNuty82JUCpniecDElObZd0x+hL
yHdoH6mCa556Q7kT4H4z0jk/5Xo0Ar3vSDFsP0tSTySwLQTXDB1yP1vyAth6/GY07+omN7n+deTg
elZXhclafJDzYOJvgGdbL65lhqxCKA8gcCdsyKwVHmlMzSBWE4l9RtD3z66LnLcwmXD7nOfJKDXF
OQdzj9USzxmG4aunOe40SXB6g+QljIU56IQp6Lt/O4pHYCeiFovXofLs/B/s7Um0cIYW9jMJNiCo
/dPGGYgfaYjUjETbcazYrsz2n518dRpGAMGW0NsGofeODUTjmdawZx/EoEXVmNrXsBf5/fZ4COZi
j3st/2XCy4WmMc39Ce94uVeaKUmdqlmtTkw5nZMIruNz0RKFZkJK78cWZllJnXwA5TqzAXNGwI7l
+9paw3v3XEEshZAp7svVVZZ36VBq2OoQy1o3w78WtNLI/yl1VUgaWwafBfIyiaWePgjuQ8yYXOAt
ozTGYrVLKVH+H/cNMBhiLN1S67LxrT7n+78Ychn6G40OJFEDkhgVnkw0eueurcEv79pZqKnQiW0D
Zx64zhLrdbrwd5tmOQJuUuUZ3qtS79qxhBNGwihZtcXqSRPZuujl4r+MkhmO+8AoWDSe0QxQG67P
zfTP3K5Nq52c6wneW0iTHrlT6/BPU0Jzvxui0loq4nZCo4cBfhwdgNxWsxO1hcw1H8+aLqKvK5Zc
CI0UVFNhiLayX2haTF4qZ9A59QnCGOmVt35JdSMrAHS9o54BfJuYGWpeqR/LOd0F9J0NarxEuny8
uGVoWmdKNRrrezmIk4vi5ynZ3ZvCLICilpaUGnMUbISjZTgv0tKab0QJsyVEL6CcEXy/gfNUgWXW
tlPiTODLcHpww6OaEHOFw6JYzTvrEa46frzPDK/3WY/1j5E1PNGbLTHx3dCENWmaZuKliQaZUmMj
/tZdZwLfiLZt1WbXIbEOIBAN0H/brGlEgtXafpajgWZ3ACeAaxECXMPrPxvh9FxvM99UVsvmm87h
HJESJ5tuRLvh2J+AcGcV2QhJJKEFzqPZCM1Nq8b9qvJAN0ufaIDuzH85E3tA7tWbu/X+HctblenN
pd8M4OGfFatPS1rmymYzdZB2iijCiNP0UChkcAd2jxOfmKIyvoDbgO1jUayLiAR/IB2bVgeTyOdZ
KDKdIsegvYNI/IWOREyDW8jRA536wFmlQXb4zkUjQNoVedYtmicIgAfaf7Nlbefhxqbr0mch7epr
+FLX+S8DMCUk7oUOOswiWmJ19szPYF0vNEKrgPGczLdpwmSbOdWkBVZKpsDoXhGjMR10/UfSM9iQ
erygCaSRn2Ixm10RqdFLmdAaXXX46hXmqqpbhrYoYiWWZD1GJR7vmN86p5iA3OGWr16k17ffYvya
aPlXgrBsN2TErgfVuWbzRWfotlxUKGDlECGxVKI7iLakmEC9BL72fZMlBgvyjmN00a3qk75y4k9p
R2MjHpnBIdwGhD/6OzZlOGDpZbDImJJ1HM1xbxJJh102mXJQxjoqxQer89rWz5F6AQpM0zANW4c1
UZRXu0pdbXoFFukMh8GuNelopy7C+lQqy7QibGBpBygt8MuYNnt3tQibhBzEQkiVdFwpBPHGt1Kw
V9yoswcCM7QaRiQiYtGOm0NJQ56xcQyaTP3yDqPbpyvZPnoKY8EF11MXmhegzKyDlV4HiFaBrloY
WfhZVPFC8/Wi2ha5RlhxO6XZPw4rTPl1NXGNepoDwjxHh1edLhVR2yhLRtV40QigpAUyR06Q43tr
fQu2bitRxi+HhMC9mzPo+v6QdIct/3niWyepfhHhhBlbscXq16toyDzX/nhxuDUBSmWJ9e9/NWKX
CqE9a6FVh9pY9AxugKeuCSeqyNuz7q9O6NO+JrBYC3JC4TNU8lDTIAeG5QwI5LIT1IQwaTr8qTfg
Fv74TgCjjddfi/sNV4yhkztsnGSN0aLjRcyTjDuFmL+t3GALMTW6sueGDj+DsA2pTv1viUDTi3kF
wFs8iCh+8UuvBy/m8mfFJG+sHv/Ys2g2TY7vLNUOliwV/twDOvUrt+tprPb9UScbKF91/qv0Erqx
UnYzQoI5WvNe8wsgrP/gTImRaf/8LkFfhXrINBNoN0AwR0c/DGbADEVwfii36Apawtc38+95KOAs
Vl5o8vv5YkN4JEv/w8Pz8QFjnPvotf3XJjGTj9lsan29EsMmNlOcvuANSFhRVu1P6eU3j/Up1pxB
CK7E6USUoILrGxLMnUMHfifvq8Xzs4DYaMjHNpq97chh5UAnH3GvHRVKgkQDYL/Y3KiTI9gmwqV6
oAcps6LTAex2MwA8FR53b5FaFO97KS2iL+9nw/8PLTgPGpDm32RIJv4p5LSIw8T8gyZaDSgVEvvN
QZlmJWqeu6WDj+b0oE+0t29MyBpoyYw6JP5tquKBSh3QGw1PJOxSf8FwaYxyncVT4TjZ/sEDtlNN
PJ6hpXn9opEqctu84XPxRZwdQszTo2UGztb+iicYCTXF1Qp40VavvyZfIweu0ByIa4ue/Vi1yFlz
/8Ab0hJIirFK3w4cE2CtlJ6uPuf4cY6Vlstc0Trjpl9G3hHDDzselwB2YhWqzjgh7VKucFBhPrgx
NLFTPxryS/xbbLblWxzu+WeFgJcZt03LZGxyK/8iJ95FT/p91ZZzfPSY/2lL/QG/YuL2C8YwKzmF
nVkebSeqr5OVZynvRABV1Oac01WTvy9j2yC9KqeSyvJmoJmLRsCd5f9tTV+84uZ/UEtJ+7/Sc2bi
ScqQVFEqIkCC5mdn8OqzhH/y9GM/zdopneebzPbOFwW0KStBlLdd58DfkyUeOUfYVkwjmrYJ2lwp
JDycGqf7qih/RAcnZJUyGiuz/cNEnPXqxv59MHlnBVYOaXHK3ha+e54uUKsYnzkFK3MS9GXsSubr
LnUrEQQzHHIMm2M6SryFJFDtOqDDlg7fHv3e9bpF88irvTrx7cdO899X5GDHzY9SBF9U3MkQOWtO
7O5+Otu7ptbQdBowzgTGUUqV0nuHnx9iTHOElSHQx+CXWR7Xlm8d89BWkAkwADeupHN4y+W9+z7x
7Ka2fj8utPNpskECa31EHThF3/fGdS6RbrebTYx6YnUBnZpRpq3PE+lO9Rj3Lx59QJM2JrMVkdYx
QWxesqzWdRrAwaCy7cc+1QbFj++Si9gdtt9vChbW5YtD3vJwitWLhoC/CscHUEKbMZC8FrB7p95X
EyRajSMJWWIC7dOhQ381PR5J3cKr5vCtWtrHmh5jjwAIibNx1WnpgrFRW4tldcbJLB3hjXBm+36r
04dyUxkFtC+Zu6K4OmTPOZWWdf5cda4CPbcCRcfPm0d4ut+n2Yqv7zY0XHM1zUK7aT41MhHofM/u
6izak8ovHhUUkUFhNqLS+2ZR9geD16ytucNk49X+LcafSMgsZt2NV4bdL0u8Nixnb0r/abr1Yvyl
KU72wqhj7Vee/pDkBw7xDNti0BMl5oOK4OlVdZa8RDXr79rpiXva1sMGpXQ+p24/m0Sjsq5ouf/8
usw8opT5n+ns4xv+Mc7km9dRU1Tsw2u55VslTsVv5/FoTFmuUZP1cYv7kkCtUAnIApL8N9CDdX5Z
jWeBasnyGmUFuZg6tI5+1Ic2UXyI6fXaS6fz/gwrvDHdRf4pI+w28gqfxySVNGG58UvaUIQoBsmx
x8/B1YH8ir4djeiINzUrKvW/pXI6fBTLet3vgWIwSV9Lf/OWTiYH0n5aX8gFYGHbQJEo9BK15tjS
/6P/SRczny300L9mVg2L0AwgEBqMUaK0LotiYQqD94PTwrdbykw2FSPP2zwMvVCAihZPbb9UutjB
2RYcx2h04pYWDK8igBlfs4wvVwnIG6HSqqMP4S2CpJpQGGylJ57Qn+3UDBTTY0L/mDx2GRAnS16l
jt2c8TX9XgPM8SZI8Sv6A4W5t1ug+WvOm/8ThyvKANAK8FjNCjE/vK/7Ef1bhBctbZurXJn3Lk6a
m3Ghpz6GsW2VHkLPzm/tMhSXEFgzWRh3u3QqgeOIzQmDocm07nXZlIe7DUGrK+RZ4GgrZi820K+G
Yt4orr2RCvR2ZZiq2/sWEpEVd78lczgOpZ7gQvFyUGaLJAiSrOEI897tzcj6+hKA7cI8YlGeZ/1C
zCLt/CaHAwapbiBialGLNAmKneY3J83RpTFzUDFltaOoG4CV5vaVvZUePLhvq6zf1XkkJGE8iqvI
Z2SW21k905H+pl6pjfXg0yuKP1Jxams4k6neGI71MsEi+JYPkLP4qyr5gPhjti0HePetgX/fNIgL
9gevgAFG5VGl8Ab6a+NIDOAcFlECXLiAnrEyGp1EjuGoOMe6KKDZejIimcO3NnJuYv6uXNUK0MlW
htr/Fk/jTZUIokV5t4hbMSOESeBPLUoAFJmjkEjuU7iNWJC4JtCRwtblYH5KxQevh5HSP/y1kuNi
/e7fuf1be5rDbzdw2qf7ktiTcpcHUXrBvcw+nq4eOEuw69s+5PPd2LwYxh7dG9TGYnd9s4zNaNMo
sJx8dcfWMVZXGrtUnBdZciL++1f5BBYKq9riV+riVSB2+sbWRdAfWAHxKEMmGW37DjAJbkljEuG8
dfEW+kxkr0lk/Q4J7YF2b0gbRhxHERPgw4LEgxPsdaPxk3lPT7TuUQHqILyA/R7WFBLxhTaedM5m
3TcG4hq3+zt3AYSuSXAEUDvahU2k/8epyAeCqMhrOekF8BNKNQzy6SCToFOQWWQIPsJ2Z2THy9lp
7Vtfq2HwJDzkITVecssJqTM/6tDjcFsGiPL3MihEbZB3uJqqbiOgLyS3MXGdBki3ohQYmfmj2v4U
+5oKfOFAPGLR0NQMAZgnFAK+UTkfSJEGsvCLOdDy0RMYoUJwK8JjpJl2WB4iLeFrqVa+07+syTYJ
l/IKfNWuy6K/Kl7WSjNfIWWtUuPp6E4F97LFwTsxfVDJf8dVCF0obXv3eCfpL+boWhvxkbiY7//K
6H2Twb5XPu9onQsJHKVIBm68gIPiPolmc90X/Ea68cIhwMSUrTnF8EvGTrqAfafP8JavDvmEVWrv
z84hD7b9+Ax82fNs627tPBdOJyAb7EdJ10hu7Ax3WTzdgaLtGKWkO2NUEXx646Er+i9muxETzGa/
yLG1zzj9a1E8uEv3Zf9nsNupbVWTHpH3l2MGbqrJuAMR0L+LNiB4OeY2YkTd17x1zhkWB/ysiri+
pGaIlbor5v8kLhBLHozUzseE5d5cq9sNsQxvQ48Fdk05uiZHRYLnxp4euqiq94ZYN22MhVhdVhP4
QzqDJcRau4Y2xAiAyF5p3Z+rN5xuD8CKUgz0snaNqrHHAzpV2YbBXQRbaTdEyOpRkWUTOPuYNxwC
Ymnbm0JGUz1ux3+/BWSSsT+7JaMDZfZwQK2HdTII06/ITBfiXnuhSVc49AzWLJ5J7P7sBZfbjoUy
XIHug9Qpn6HR1mSLMkgAE7+/E/ZmLnfURxmHy294x6POtAzXFKrYT8NX0y6Epg10PHzPo5dumxOK
JtdA9vHpkE0ACapyz/ryQarMNjSpujzyfTmKlOV4RT06WMo+lN4BJrIFyOVaw67X3pao6L3vBAsN
gyyLmDc+/k9n2nPGTvvjrWJivtjQzNhqXPTflvmpmGnf4D96K2V1GXx3XDBESqfzH66j6VN4qh1F
SEIozIivpAhB7pBIPhlbS8vMp4PGBF022XHKG1lRurGNwxX2jwrbrxGi+lJ+9heFMwshXeYJ4GKq
FS0fIa6BLaHzZyAaQhCAnQVcRcs9DcSIQBXYGny4WSN/McsR662Ra2Zbp6r3rXFk0CQTIoK+4b3c
FHRwlXI2r5O3irGns1AXbb85e2P3xW1xAcPaJA1UXud/wlw5AkKe6z0bFcdsoSZJAhlF6NBzMHBI
DNGdLK16TL5e2f5InpuWI/OSENko747zpp47VuliqaLlXl8OKFnWdpC0kuDeJvx5fJhUXnf4Vdsc
wWeyxUIU9/8w7T1kikZRybuaqGdR3AXFdzU6l1STqC0GJLmaeLsC/y/l5D1ex2QGKIrTMRCldbVt
wjGFSd6wuItA1xLhZUOT4Yhqnh4uCojfyHlhMTjay6J0mD9HzlVic9Czu0nmVHwb+MqxFiyCNigu
12QShAgVOwbS0aIBSeANE7TB2VojM7WAKApIxp9OS7PqvfLQcZURu3c3ILvthf7IzSjvEATNBPbG
97oFHYnczo5vAh2NxZ8TcnJUxKkesILl8gYS/3iyAB2j1xnWQ7bYEoTlUwUOHbi5536mAMaM9NK+
JszUjyBALLtIXSZl+3IVbYTxMdmL8yFkRjNSqR3bAeCOSc6grvsEsp1PcncLhqexiCGfF6X0dUv0
mG0Z7ibgkcEjak5X7pVrCAaE/e/l/Vljd/mP229phL1iU7vblGFS8Ap417v1DvAK20epr7lzBW64
jYZJK+kf+1zCLUavczWp4VvzqeCNuQvQpdR06rvrjFn6aXakvZoKy8WMizzkv7nXdr5k37CGephj
aJcWLrX49IFqni49YNZ6/mgO9CSlLuw6XDKF9reUoFtpMmeArU/OJe0iWKq8HzMtlLWGftWqgJUz
tuDakIYqqeUFLn4dp/BM1R+FC1jsmPd1oKzJGtxxFUMc2GXfjghPw5Iufl7JLMbZInmczH7SVg04
yAm4NRQiO6BE8DZTCMcY26zFk9C/mptF+2PS0IOXqSpX6ou8krbtsAjaY9yoypioDC3/0l3a3Or1
6K4zRwAUoJ0wLIDPk+cV0j+Te9xTEslsfKmAySg0/SkBvTl1gVnIEMxSshQ6VVzDy7NFZVUAJtEL
WHcT+zdfN279xnplYrk8KVfw4gYe1sWeJJAmuejh6b5VnPVB4h7a+2/RvYYXT51Feswg0gT/4cxD
9RC6eIU9PtwKgaGTW0QKks7q5NEdn/r2vAIokJb6HHUdP7TTEEwAIw0V+6jzD9245efcHxJVYbcK
TwNuOoSrFMCMXjtVBTI40GQDNWJ7WcfU3zZtmIZuhx8AJRDZ6g7uSpU+9pfihlutZ4BhrgpKv3sb
oCqpPe3bI0QYYO1KF7NCcLukPo3O3sYVQiTCncZ+gH2CayB16JbwWpfoZMqi2gpvdh1rCR8TL3Bb
6Y++uqyZr4fVWCPMXSdDkN4GdZ0VMpY2Nuh+Qsri/wpo84pxyHGBjI7aRPMPHdyhTKyh7VHovDG/
hLPjayP8nm/CR53vUARrpKFA0kvSlQg16GGIXeEUelRlldgBrK3C10r+8Xm0boeEsWLw7GxodN5M
gczKKjccKcUMPhlaQ7Njmg+o7sbxb715SEYFBiyf8viRJO+ri9Y/E4RyrXSpTBb9ieAEfXzIQcNu
pGhpSFDgD6uZETOlvNjZ4i9aP8kl7/jK4S+x4qM6n/JsyaXB1v2NaPx82kfZAK6iTHfZ6laYvDIR
7SaRcJSiDsS1UXyrvhghRe80SBxhVOHTA20Ta4OfbhR98Np2iccrt47L4NER8ccN8WHeymVkD5Mu
DmkzjmzwFkDzpOSrvpaNDwzb+XdRCIX9zW2r8gtnm5NWLPkqcZ0YV9KeqCZa3k2Q7Txf6yP6C+6R
EtpV9B1cer6PpYxmwpytADO3KTm5tXf0uWxGKf2bpsY7MjloyRDISoTTsPez9CFsB+3eF9GQ9QWy
r2ehtvKqu2r4pAPO+sXKPpPGSorrMjSTONRBfditnV/AMM6CRMLWmwhBY+jd/V7V3pvYgeUF6GjO
5hB9XCN3Z/OCDWk+4wihmefUnnJKME3YHnin87tobsCffinCT1kwxROnbRUD2G9GuRsZEkMl75/5
CQoipjpD9rdECWW1Oq0yc9C/WOarXVZ5OnIcxlMGJ5Z4UDhuM/zneEGcL7PNZz/raP7cGWlzpg+W
3aEcEWHVPHsC6JuY4bxu/1GGfo+Xw232XNDiYikWc+vGiUtlGq4WCBLScH6MOvDCOfMsUbsFajVE
7X57diaGaKYMbMM9axeANAHL9b+PTPhC5ByFi4Iwv2MFmp4OxXkrWWm7TbymaRVL5cO5LbQAZWDV
vh5T31eIVSvY6G62ZH51QCMgmMVNKroOwwi1+X/TMo30p+xx92c6dIbYFPoQNmahK64cmzMztRIu
XLJPHKwkrP5nWkDtB+ZuqQzaK4Ri5IpgqtYF1CYpZgnK3mqLkmHRO17+8IA2/GQiGtoRm71PEPZY
DTapP86o13e9RU4IwP0FIAWubOiTYFlOu+aTaDRtHpoMuN+Q6uiMDA+XVRhNqmFiXUpYIqWQZHPN
g5hnBT+Bh1e/+lbUEdyNTAQLXz0oC3+MSf33twLGxwkj1dvxmsBOs5TKaTzIbx5q/EhDGj2TqCz3
1GkKTgmUudyowkx7uUaC9BtIHRJLhOZzYVchuNd+uga/tthglR//R7FFC8QHffdM4xoosUMvOi7F
3anD2AvrKXwsfc409x+wMl+/bih/V1fYxEw3ky+DvCipgI0epdGg9/iUbLB+A/EZ01RbOLKnHIef
H0AreZ6nrdy9Zej01nMa3czzrGOwGmpOVhgyQJ8LIBUFe+UJSeK2ri3ApvtB1PFUld/VQf4gAEAH
nbl+WjPedTe0JNqdoBH6A0qfsMf3HB3Pp/N7/+DCsU2DBstzQVm3CouRIH3OdpF2CbwnY0nwjpP7
Do0AduK+s8yOBsg8ragWMlhuvm23PfYQTAgVLZU8NnDgiagvQjs+rjWzvtL82dmYnFoxjxAMiF02
a5ffT3aPwYoIXkFlLpJn4lSvAVqXYPXxQNHwGNAxI8LJ7dLquZPK9qgvD/vaioDxfWPXSgHiwvdS
6jnst+2h+c82xKXrf/2z+DevG29rfvJEHPeI+KQbyv9ErOK6jvILqsMBNjSs119QUlmLG2Hl0Qi7
QiN5tb32yVJpaweq3ctijzLgSVsyMghSRly479AWDpRNXj3ODuIXUfm7hMKytyXeQVrMmC+p6N7v
jUjHCFi2tjhUNwl3gAeg+fscR2B5UCq48S/qQZB+0RdL/vEGdODOjts1+mJySg8p6jp9bN/piwny
RQvktYmP/PUSOpeL56k3bdZTZ2oa6yA14dZaTyR9Hsyqx8NKyDHtWAY3CRF8eMjP/ZoVZAHD1P1r
qgpt8A/PbTQdD8LkBuElWddkbtmTWikJuywCEsvbdgjE9nj/n9ENv5UO+MhIBhfuD5YkE4T7AmRR
qocdqwoQRcDmLr+et6Dc/x0qc+sUCzMIeI+U8Av+iEysRGoxxt+RCh2KYrUW1n99Ec8/GpukVQb4
/GSZPgUj5MtW+D8ue/sCZrco9swOG+r8crftR3pFWXILAZUpMxQtG8lEF5hkfK2hjjpiSBvbVIFH
e1scPJLN9A0VOPGG9I2Ar0bJCaRlKo/F21QgiGkSuWlFlXb1ELbN9sb7woANe5oUUSKtm8eZHg1A
wgoMVISpLoUwEpmQ1zm9hj41sE6QcihMzKWC6gYM1VV09KYNZcxjONb5x6pWTXjNsDuYG2vYuXT8
EUIfhJUjeg/OTgTVPHWzs++xeMeqYJcFbMBYovYxaEB/iHMVyGTOyJ1eb2gAhq8VtEMDItgkQaJf
3uQ5MvYBgAj6RIun9X+DLEghR2oSWdLUjzD4BALMTVojHxRxmTJIcWQhd+GxTh6s+6HtKwyfEXT0
3Llm+cC3iG1jIgsTq478V7mNXubpgai7CZVFAEU6dTeyUV2kAq2GprtE+hslDh5Gb9l6kNefzogD
8qjs49io0nOLaDRe1qQ2Wdi7i2igJg6bVT/GjY+QaXnAsWEvI5jeLifosugCo+s9pcyNZGltXJDY
ENmgBe0x1qBgYszeIqaoW+hqqf2z1KtNObvhvDsgac5xiZQjQutfrtA3odvnkIQaEtSRw0t6Sr5J
DVZljXP4aYY4k4MP1jLxGf0Roi2YIuRB/DZ4QANphrr4iWo2vIIjlpUl+5EQyS7ada0ZpdIA9Fhz
0HmZiNvYGj1rqob3/ZtMguQqds/fJ06IKlKCSZmfXy+Cv2sfd1QF2SlCJp1onlrFYWhnBuvBQhu4
w2+L1Fa7pWNT1cE950bSC+8nYdr2NXR6JDy4iRB+xKsiVhoQLvLh3qjxAOcz/GL5yAF+xnnU0d/Y
qiiVAQvi4Afa0hTEvpWd8pLCO4SkALaepowv0FGa861Dx2ndQNpsVyk4PYfKeczsbMbWz3IQIIuE
CTB3YWCdqR/tDMe9vYTD4wXP6jBTUyrNtv2BhkEknasJfvRZ/YzL+HSXQVnYyFyWdGSG9aHeZUJv
3WWD5C2YNULRO53OMy3MTpUfQJv77cn5NKENA5dFIiiPs1IQXdgJeWl7+jI14l7qomik8PfFgjok
HxILixMN6iX2yg5nvffI/5N3LqC3cmL4chZuiByv3+1vP4VIRO/bJkcZyFV/wH6UoCBH0pIPJ2BI
2+Iwe38S0xMD/CE5iD3dJW04ztlW+H5fs4319o4NEdrhOsN9HKO2fEUlb3RHew7SVMIB44CYkASc
YAlu2phgoyMi9mEL/BgknAjWoSvKPn7Slsi+FARUm428OeEMwJNt99Jeh4zy8HILqlCMeyl9K+zA
V6U1W7KN1+UjhZXsYm7OE9kukaKW/lhTkX/Gsbb8xc98mLpSjYnySFYnuMUQEQfcQhYCNsEOOGD1
a5wAbzsetShBiw2BRr9DXXNDkastZadH8G0QWPeCgBzK/3XxbUoUL/YJIstyZQjFtHm+vq7n0BAo
AK3tLMyFqPqtvNDtzQKBWdo9oBr+t8aFT20OX1yNYJT7+CSFdATM/wgShUTz6YJgb6kW1Pp2sXzJ
ecjodN8gss+mg1EwqGygXscGDR2PUuZX3MBxR/aXPjjpei7/sSVKQtQyM0EPVlxAYQifK4HbJfTI
EVhyTzRTSo4gFwnScaipxJ/By/tyel7YHg+Oux67SJSdfN6pnxbGSK0HHnuy4FWySKpvBn94uxZ0
B32qxzNVVrWRV0osKSBR/uF30C5DKc3eC6nfLbSovugc2rYRr4ZJlXlnHludyW3Q6A2rpth0yev5
jaMqP3MPyMN1zYwWU6FA2YegCctbB99gwM46tq8eAUmt9Uau835vfNc9DywTC3CTQ8xP82J3wVSb
Zi22qkDdCJzHx2AOaJPKj13WfmQQ6uAeTYPd4fNFR3ob+owRdhtAuntKHX2O1wFRNSzuy6WLdrka
1Cyij72M+z98wT8L3hik0au8nG/+6qWcQxmesM9cFzwb7+I2FfzzY/x6B4rJwdXtshHzF612MAla
JISW+YeSZ60zW2nMPObwqno+EoSQ0zPtK2Fw+yCx4RqNa6zkzYCi+driV/xBCAhinmEyCx1+TXIT
DKX5Jnucd4WFFTbCB7fierVpkViYTUs9c3O08wfw7GEydb3koVCzbJt+OTsHZuFvxwnIPjWJNosb
hYtZKaAkWM94D3ZLY9/Lemi38uwKp3tMA72VU6AF1itds9LNkHLfAebXlS8SeZKur+wVN8LCBmVK
9apukUE651Ry/MHhVHHuaSuchCz1uCFKdtWg3Abr5oBlNA7CjhUaaCkxVTTRhT21NtRiR342tf5B
KOAZ/rplne+85wvhvXvt3vGfp1ldFVmrJ7MDYKH/fTiMDJ4TS2FLSstLcBBsWf0Sa/vBMPhLcHvp
2Qz/AytsQ1pbtdHKUfvajUeLdQQ7caWiHfvkgoy3zvKAbgLz5OatV2yk0EkoQkbEiu4UcckXa871
yPpi4/UKrSf6bKcTn+4qCe3ob0hVRKEeaA/VacpJlCSikuzlbFF4Z+7pKJwgP6UsWCF3O/QABeem
vJ52Wsr6xJK4rFOZy+U4AUWOBNYT4yjwkluhM6g7QNBzclV08oW7MBa8aZRmTErCIhwVImIfnei7
Ku2xwVF6RFKg8UavqEfyxp2lyxLdgcm1REQcIidluWqB5o9U0mfHpVpT9b1L+q3t334B/TNFQTOo
yT5eNczpRWxt2nHp8bAIe5tMnpmYElesjmFX9MNQp54fCNp1IuRwfWP4zIpk63oSM7ZZIpGkD1PH
kdCsh/R7jSmYibfsjI0AWgnPF6QPNXALHEl7mXMZNa9U9rACFQgMXGDRC5yoSmoPwI1YqA+Fu+EQ
j5BFp7+fipGSqDpt7w+aq3dFBTD/FTuSBes8jAsz1mBt8spLGbD35ITRzKSlwyvc4kpcfVQWlpId
wW1gnwA/moNr5/T6+y4kskG4LejJ4QBDjJWCVHJ7wzmuv+YNvw5Cgul08pdn7abRQNcFHgFpJyuq
8uvJ7DM2vtX/votcCr3CVvDHUQCi6psIMO2ifqPNib4v8j2q2CBK32QkQJWF4IwCYSnZ1eP3rCxN
D/bs2fOm7/vlR4J3laQbZip8Q1/2vwTVG2h/Iy29QoKhkpuEvKltnj41fpp76Goly/MoB/7vpUYT
Fpf6zpKaYHaQGQpCNKC2wCKWonMtCQshkql8D9wYYSAwfG04750O0QJ6AAIg6jtI91RZaAqPM1xN
V7LinQlXCDZ5V1SdsMRFlmhw35k4k7vHC/YsSGOmSW4l71s393N9knLhOHVCJcVRCZvdcSoNMDLk
VS4y5TlAxJ4Lgqk8Nk8faGpWWV+N97hez9Bc2ANIQdayD12HBXIjObZIfrBk9MS7tJTVK07iKYlW
TfeghgKF4ZLPyxNuu+PGOwmerCLse8eOouAMLpQp40tnplcjeg0vQwN+4p7K5Hgj1DWWbasMdw1S
M3VWGigo8cHmQoVUkIyFFlxyC6aRBbWtp/zDsjqieXP4RITUt8IEMm9lpvhgDVuajFulto4ci2+G
MXWImtkkRKyheIrBeO5mR8L+1p+FpVBWuGczmnyKeUu3U1l56/XEb5TF8RRLdFyrbYGB0zvu6SZz
1x5D22EQNgdvSOgRqPKgYWLZJcNksNhahsreRZLbGIs3F2eXsMs9CPvxA/7R54lgGZ0GGFUwNb5e
ypw1M6yGwG5i3CmwYTh0XkOi4kM7DkVI7YuA4NO+VOOxWUWOvkkmXMEcf+satrR0xHPmIsu8NVoB
2Cn7X417TgBr73l/zHLU9SHOniRzsEAMPpp9CVhOaVxMZpki51rkELtHMJTBzZgsZ31ImIl+vsC/
VvBN7Zb+O4uO4Hev2CvRRI/SMMjboEHNlZxIdERxZJpnaHhKZnfPe5qLTJnAR1QuSKOHh8EBqG95
WoRlLyxyCXJWId3vW7IOO42zzbwSai/I+dAbnsdYQw7mPKCs9Rww+Df8lvXVTur/NLlYrCRgH5mN
a/3YsDKti19bwfMlYEPWfemqIIzFn8KsIrLUctq6TJ73vPbAZIm8vDSR4q4s0B+Q79/FjuSwhINQ
KAOCGaIQHGOLdIhSwUp1MknjTf4vw9pAdqif3f4/Meenl+ZusYI7cIpPhtqeWgn3X3di46xnjAO0
WtBuva1nx8CQdHc0Enc2HDfxGoa5yceGV93jEDLRrrE5jirrTHjth4kJwarATrvNXZp6R+wBtsek
GjHE5cpkOOlO1N1i6MXCRA4m+K/0ztbqSNgbZPvjwDZ/a272Z7uxLzVRP4UIOO+7aFnCFkxS6Kr5
DdO14EMmJPRknNdR+qXNaWfc8lnhNGKomauYCRhmODhjE2EsutmNx8IB/L6Wz0GkZGfqBRcCWqak
OuC1W8Z4ccPcqRmNGsdkAuXCTKBPWh4tJHQ+LSwQVgF1MlPEdqhSHXxnRufq4HuntO8bVLunDUmB
TdVPL8OcHiffFZ1zaXMZPjaG4K84Y1Cany8SUO7OQyzWPDZzZisIaBHtx5aezJMBU3zOu98M4pAb
803/JqKhbL2Wdsi6cARtZQ1iGFGX2bf2AxiYw5Enp26QnTjxLMeRkpSp94FaCRcwf5GH9vNYirZU
xp/H9RfICs5DE1azW/XS2gHG7dBdzqGAHzZRR/pMkP3Tg3tFVSrL1Pv66BLvCPQ2uEbN+5Ny8zXe
cvJ3C0uY/4rsbfnI27lxO+47P6DEa6rey9/jbZnPiGDLSf1ZDW3RoRY52BP5qXqhPEZvtcpDkMZi
BfjWhOLxdwbb+W3NK8zOpZksWjSSiUUjZMfZKLt+PpdsjJ3ugb87vAVkzyrU8QIJAVdRmD8S9cvk
5rrGCuy0sf8UuwYv1PO7bzXLfyX/Rz+DsqJQxaqSOSy2aXb8ogaWcqVRNvfKKMfy/ghpd93yUkTf
cXAWOA5I9Uny3S0xIYL7WJgusI82sIzsYBv7Ag3ewTNwqoM8w+TGFNdSsOzOb35CK4K4Ippez99w
IAJzyMdQLvqkhX4h1sVqgb3P74qXPnd641W35OKnvt7CmlJ4y9sf8RWRh4S2gXJ+heCGPWi1eQIa
/Ik+m8NZCSlJkbqxplXovJqMJoMKxZnTeQyDkjVsM0AjJg3fT+dOnVLnLbgRpX3m/vnKkkOT0dQ7
U7bkOYWbZOLnMRISCfYRy9kwJQgPMv78uqVb+T0INgSukWA+dgT8qdZ2pKEVXOwgxhcpG/5fwm2m
GOAdrGd/YqO2iYQu3inz6nRd1JeJAwPCbMkNYPJ6zAQsfw//J3N8sMBA0XeQ4d/L4AL2nRJ+8CB0
Gdm8t+SGKzBEiNPmEsHe6iwylPCWkwNi8soJqErgk4lLkGHeBB+q/B3Qj4asYRCOiCl6uB36Uo4h
Lzzh8hw4Qze+i47R0sr19DGsucQdz54sJt0abgKHttr5wLq6aNLQuLf0KDxWsTU7TsingVwqOmFo
sXbIbJRV3trMGhD8X0cwa7w40/RqKpphZXiGA9srev8QkjeyPAM7ByD30eDW2zjbCdYc+CAwcfP3
xZ3t0Dhv5zXhGvPGabWlqQTccxfLVthWgISL9Hvsm4Jsbl/LmVPn9fcgwCXv4AQm+W/E1tg+HugS
ZTja76cuVskVvIWsitacBvo5wGdsyjf1RR4MY6GAWIU52PukrtNOBVLKlzsPI+YZ16nMVfBX8TKQ
1ybVOY5+7vIim6xuvHQ9j1UsbVbCeZTsIP4+kcnEdlPZce9rf96DzbjwrfZ5CkfgRBtS/ugP5Ywj
sqVt1Chb3qjlD5MSWlc27XQCmkQ8Kxmn3Z7IeWSNIBmjErWXR0MbPHEIKCxGX3JoZIUAF1NfrxaZ
fW0JcvEI/bhBuWkssg3eJluICNz2r+vT2DQa0kV+fUP6VsP8vIIMpevN3eYkB3w0eLJFPgbNu9Tm
0kGyFi6VU5UYwOaCdY+IguEItpIveLlyEAMUpEchbr2NDq1ku+I1PQs63VqAM0H/PwAK09i5jeqV
0uZNy/wSUm8gn1TJjFCbzI8k/5k8R/FPiVX8Ac90IWS96VH64lViXrSQ0jERXp7Lvf+/36HZ/H7f
KLrrJQEzensBFz0RWbqrG+zWiSz+vYcPJ8rYY3OiOkrTOlBL0fW2Q2DBsgsUGXY3y7lhoeh8Xr1T
X1PSc1blm+8IqDFbjVdk68os1t2x4y2DE83ONk1OnD4sT8MNTEbkfoxgBOJvxEJvwDHiIf8u3pKY
Ud/DCRNeQSF8pddnp6UtYJ4PMZRQP8ZjMx3ogbBcEweEPJvaPKHIcBxSd1iWeKD8OGNWxdwdwQ9E
5ZakkVAlxdnysx5TtL4RgjXKIxAQabJ/9dAu9YsI8VEP5n0Nkmp/bDy//pFvDZv7TRJ1irHu3OGg
jIw/+J0CbXnOdkk7cDF+jiTQxKKIGMUEnp++SwsfSRGARk5muo6KnydYPi7+tql6kjkfegm6C0p/
Q+FnC+vXejivryrlIR4t5o9zmtPTqY4EpKUbOoq6jOyH5yoSSOCYB/Syr69dVUhahNWsH1NqtzCi
6srtMUicRYS5F608i5Hdm9nJAaIqYprwa7MfJk2yqRuC9hHUtqAAZlL3YjRHpZRI5O1CBehP3ocR
9AnmM1Hxaj7gcoRmo6mgcfEIi+s2eDwzWljToOfNUZH1wugAPqH2r9WOPTrGDgI8ei2IOZGP7rDh
7vorPlSPS1tGZ4r4m+cI3JEgpFrijW4uss5bTPNDBoP8JcWL1ClJ3h672lUFVM/HNjLVpGiUVc/T
LDJTRlbAPNPs2NBpPtioW7syi04enHE9WprJxaPf5wrEwZDPNvryp9TJiub8g0BkKYc+T3oIAoeS
iVVoa23k+2aYhbr7NTGqaHYZgGaXIy6mWEPBJbmUqFK9OKGBo5LLp17F4eAryTRt+4EBqxsbdiZp
gOsQzkTFK7vhAODP4MKSnpN1JvP0cZNC5w9OA28n/wREA5MUvwyNZS1gJk982fz/WFOAZK884nWT
QGNdWB7pdPl+ULh0ikz3HrIZWTHzJXbuvwV290dcGD02h1oN9+opDxRtTW0iIlWjsMj7JcYvEXS+
AVEeFerOzu7a/cFUgrMB2mnjq2TThCNN1Z5YXGAVNE+q6Syk6aSU6eOFE5xaVu0YZphr9qmBG6IF
OFrPWvkYnH0widq08+FXFTyZe4uvc7kTfW6d5jKhKOVgYipR7UBFd32jESprrFKhFKkF3uKWhhp7
RJnyF5TH13KEDzIYazFg51kqeG8boGKlqcmpOn2fheKgjFMY6CRJ5kDn93WetzBOCm1VXtT03OQG
1JeF2H42FyhTpBC6Bwv4tgzLMs18bjKztkha2s4uJqZL0I0i6hwNrH7fftp1LAbtj42eSeKDYiX+
qyPTL9Apunnt86hRMLUCzuUcKLLu1qKWU7dizNNS9zzvuTRoEYLy3QiZGp5llY/M0bj6lFvKB6HY
safmz2iAMfI6Osa3kD7zWSFlJa4TpmcaHYetJ2Px5Woy8oKkWbgCl7Qqu8YF7SL/mvsXI6z6E7jm
Z5gdnus5061/skRTDv3dfQJMOn6wf+A5YqgP9Dp+/grKL8HC7c1i8AVrCodwr9XQiFsoHxN4ykfv
b1gOdQKlnp1UB2fzBZgPVqEcmCTAWZ6f70R6tQrkPFxyF7CKPilBSuclbOkHE4UJz2taEas6aDsF
1sP3TH5BGJ8avrVqaJXacSPxLuYKo08yLxHjJe4I4u5REZB3Dk/uRCklje7dZa3Cijlq0iHk7PhY
Daqxwvd/LRuVrm3t91xXX3sOI4ftfEoA5YXTAy4PYnBF6zRr2bB2zh9tPiFouYck/4F2ri5J2Z2y
3ypPTY85AIP0540XfrSpCYqMAHPS2IJG2aQbeSe9T2mDsY5posG0vqFBPm1J5kjc+hPLPXQS5IFH
Na5LDtZfjHIWdjOGB7+oZuG9jkz4F/qKvH/ZLUOx4iUHGy8As7xLxV2KJbMe44X8FdaNy1+2jUWu
cfuY2LL5+FFSf4Wj9IV3K+rA/K+MEL2H+EW3YOqUdzkknFoY0nCXWDZgHSq5SK8hUJm8wq0GhZ5+
bb71QKkTxYKPSL+kNZbmMU1mjMq7Zlf/Y0WRimwyrLnlu6lT2MsxYc/q/QlSe0VY2mMxiAZS+wd5
YwkPCYlZesFWMeADfz+V7GVd7CCGgTXLqBhQmpj1OeffGCJ/AdQ7g2QH7d4+O2WVMjUHThAaBGSb
Jv4OJFqKhlmjc5X5oD9i4SDH0IbOGld429RcpQxHrHAbJ2DMZADuqQqgn+N44QVfNreafIoHSe0x
ACKI6e3s69xVzuY07fwA1tnSmMCYgarzRZTnVgYgyG9PPPPhXTocVbig2ne4wlTCmohp8xdWRPiU
xaoIKTkcDX6o1yKuO2eVPXA+YX8IvLLU0vnIg47fXTV41uTkaHwgpH32hA1kd4sXkHHeuQ2vOFSe
0bMhH+OzN8juPIP4Xi0L+LPFt9l9dgvZwdktGOp+KwTNX+CVHepqTJGImkw7SeHIpLDSVVH5/X05
azBt8T/+A5EmJ3T8vCNNZ7aLLZzskbta5erFEPi83Ap8dqRb/8A5OglLBIUPkgs9EFj3Hsz6b1T1
TFSpMkcMSrn5B95A92WcP3Gefk7eE+A460iOvWY1rX53tJr+I06jpMTJkd1q5CSoDgmLrZ81ojTS
7wf0pw58QkYZvcapNCP2Aq1yf3rGTeocPZQWmZomq2FNOpevNIyc9b48RLM7AZkqYWqACezdoWrK
GFP0SRqDVaSdCY+UIQiZS5lH5AgHmw87DDMbsOHLmxYsGnldxKUaXpUis5FmX2vRRDdUlvHwQmFi
HAhewUJY1MXqQ5u0Cv7kZ32wHqKuirtcJ4HPtXwiCd9bPRVbvKiKTBEDA/b4Rk60dluA+Tj5Ct5R
ilLx5/Ls+MADZ1eqAAccDI9aeTSFYOD2TKMc6s4wcm0nJd4XVWWl9DvdZKuvZrpC+XgBpr7KT9cg
ErNtWIqguIiRSMDVnYK8McmkzwZEEeJB9qZqTjRGf0bAzzppkRbwBg+u6ZO+IeVVEcXvRyCpAxzI
0BKXFa/3ZNiDMJQZPupKOHOzJM+kUVxynjNNkeGs016OiTqmzR6hxiW/H90i6m2YQHm8TkWzxcmL
ro53ROQggNcs5U5u0NNvoHKekePYJi1KFLeFh7mPZriJCIYvSNA8jpouxzfXHtEk8++hhHMKPfNz
MI8LnEuyFgvTyJvop+PterOg6CXu3PazpoP+lMoA0GcJqywd3ljEIrDaOfxpbioG2qoGOlDRcDv5
CN2JxY6SMzct6arbiei8COCo1v7iWiBV6KNNN75ZEk4QgrJaRndMhg/FGy59nDpxwighObFxbZte
cQMw8R46z4IJRXu7/eHvIClsG4OAYX/sZiOQZ2aK5CjwwacBhqHFYKLOrewGUCWoki7nO2K0MfHJ
GQldIut13WtpN6sH+7XEvqqdpdT5YzfO24J3Fh2jMQBRE/ey4WasByU8jAV/hiFGQIbhKrdQGSu5
8A4xSf5FVThZhftI064qp6sQYPd+WeWIm16TU9zgzN6EIDpF4f/79VTYDLnHrmBoVVe4T2E6djaD
O1V/HDgbTB8ruo2dJIKXcmaasuSY7OvOTKTkqJF8+nx0vvr/JO+1HSjl2YES4MqZv9rJT3Rknf9a
bCVfZK5yW1sz54ytswPzBT/lJd71S5GjTXwpRNYZlncyqce8a+7nOjTXtkozt/JS4wl5Zae6T2pZ
HH6GCtVCxI6lUMSvtmLf31+cEogYHzfNcVxpO1p2smRZtZtvKlati01BKrGt2TYnAPpsdTr9A3AZ
M5JkZUk704jSpkBMnkEQK0EFSKJrzEh69TXlnnVh++38pgLFJ8GXvWNr7UnAc0fdr2dyqHD6sEih
7RUiM66VGcO9HEvJzwzAKvCQFz2R8fF9aNLjX1bapmVqut3VzWAbpL55ooVnewI5kdeV5ckDq6XM
YScCDNFx3uPRn8YW3gVuj/m8cicMXfS4Ajd1YCGXjvJZd4O+DviVuE4/3dPr2iJuvUNznpKZRDVv
ZWy0gO5MJSYTpX55FPS9ya8JmHlxR/CNZgNlChFj+pVYGCjgGCKJY9gzcODPngQBBZwYdXrovAt1
C5yNsDTndSOWfu7TRXJk+mJ6caG7CNNjy8XtZN2qnM98SAQoEXX7KlKtvqI7oD/iGv+isnElNMVE
IwFslhwU8E4F7T/AxHIVidJzO5e7aL1afMS1sFXhsfCcdxbmKyTyx19ZH5fFh3TH+7BxroURv+8m
bm7t/LRginuZk3npdXS9p032wpH0oJwhzT4Mnvu6DdSWdMixOOUgWMRWpAt+VBOrg5Mlz9Be5Hh9
UvDCD6aRiOIH/y+KEsqo9Zz5YNCBjNXeaFQu2T5jr4MDZ1IjhMHsWhA2IhFEvD7nRnBZ0e+b5PT1
b29lmhZQ5cm4x8+AloszAlrDVdIbUb9iZ1kPm9Se/XtZr0IE3IsUCmTBxGjce55N2/SNyKw6PjiP
mh6vjz574ZghuvHL6pjRVk3IoaSnpIkofK0zagTztwOAm5x8ywAH0XN2OJSyMXpfwSwis5wXksEZ
1NRU+cFDVNuPObYAyWZwo0Z5EjYIyEkGI+JGwYqIoN202bDXsD3qcvFCgJMqKoVux1OIqOTzN7of
579TWy8FSFVNwfS0qR453KLAWKu70Wl3AVaTa9CiBeMWfb6luhkO1aVtNRMkf6ArcNWTdlyg4gKs
DbiQU3O7eEUtalRjrYjVQtcf40/GEUG4heqCeGgzQVD9vmJHVloKJMTZDJ2mxfXik06/DQksT3BX
JQQzTGXMydBJ0rVLf8hiBNuEIvp+ib0i4fJ6GbHOVdxFzr05HoWAIXKgLv+hSOJiopNsqTwtERlq
z/kygOm1Ymic+clrl/nH1Rd0jAzQGJH7kkohUGBUYhcwwOQnz+WhP01q+RpR3urV+bvhgFxmq/Jb
Gt/HH8rNvZ0oYYSlVsGBh+dHoKAV/il4kVxpCcQuvKRikrJ6HWOkp5Il7ZX+UrLNWgJNBoWVKa3t
RO36yvvOct+vlW9KJsW3il6jEczVwrVOS/GxqiULDpcqX/yDrziuSnxIcM7LVKACrEAttkK3p/A2
lSQjdNq44gLciVGNnRI/XIrRo2fPXkxn2zby7mHRWbw9QVaUqodzgacJPSQ+e883jDCvOujyYjGX
qvyHrqp6PtaIALEylx+qS+Zdnz0n56OiO8SqJcisLbzxup5nAxGkpwRYCIGJO09uutPZmVJ+yr5E
DAJf2Gt+CTxv8l+njoguSZUlWoALnGYIs/frax7iGMP2VucCybCqk0hqRmA64gkJJQNuv1NO/zse
O2nSB5wKICyUUgbWPyS0UZv7U4DKEXZph8tAtW0oZ+QdeOIvGcxCQwLeatRLeVBo6lBqfKKlg3kV
pYFjmA1glZBAFobAlelGffGaEHTOoRu5OzSHh6KvQo6wK5aZqH6+apuXrW103wIUbamLeA0125jF
a3Z2raBVUgCnY21NZvDB7QV6rqTewJiubPjWS8ORjlelqzv8qdB60AH8gGRWerrxEh1CwVCfi7qp
/vrI3YORwlyieNijhZpM5oAqufJBOuDENKWBD949GZxYXjwDacM+ToP2xNBFifA/EOtmhW8jX7LI
c5pi1ETLgBIfmOnMYU1hPzEQoYA7gZpEo83QhUOXWQRmpsg0yibo0TlfjUQ9vjCEt6zOke7EM/1V
g8edIVw29Z+UUqfTQ7GWFPKTtlSsSbgWzfAseD7uZZX9ugWO9CfcCD7U5AcVhXFakI+uwHrIrC6V
lcgR93vvrKB7WIUABnNnSqF64wH/DVXAV7/ZyF0ZGtuVgdHX488SMg46TtbS0o3xkFPV5ng3/6/Q
/5zR5lUykAO5LE8ZvSy1fmkej+G62cROEodJgCsROldRKowz8jLyH1IipLquj8Zn+w0+iS2JGoRE
PfEjGgcYfQACsCOgkAJ6opgTQKULhibejT85ZtWfaOoSJOc6a/3lgnO30mWN5xFO0L0POAT9OTh9
hxJG1xTi+Avn1IzTKwJ7U/S0VjfNs0GoL0Cb+cdxmQzP7f/DnlJs6ibIMjxZkOM0wiQzyWyEwO/+
iwxGAp2wQb0PImZoSrH9PzUoSk+81QllLm4kEXolcGuB0rp6CLcPd5Zi44G4ZZ+IdSZlqt0FvvlN
vJKhkcwGb5DjqNmpHhARpr9+MNgMyvA7J+bI1fyCf45muajuwgyI1uBTk+GWKSDog/xRG2BWQTWt
iAskWvjPwVcbCcVAcgurccVp+SIaUp2yt6+gxo6Bz/xdynzfz737zJLyAuyahU7pbOTH6V/ZXhOI
p74KI8RgUFQVyi0+r4McdYKkFYMxer9q41H3B/U/shV+FgPEuyBn9BChQCDe8WSbQUTAR8Wgz4JZ
OwUYT5rTFFANClnQQD/hTAACQP2E+Vs6z68ObJqY78vx+csxdoxjqwX4fCSVGRjapBD7AAOLg0yc
8s8Q9eu6tWZV9lglmvoRH3KE3YymivnqfJyagov/1LyVhxkVSLNpKrQAvzIB/Z+9o85SCiKztWb8
VUroXxjwzGnR2vC1uBdBeapQkLQSUstnm7F076iUVGLQZLSJ+wf37QCcG5ayFiIDJYrPSV2wavhz
6iq3QmCvVb0VvrOQ7K/hKuRENc2pGiALKQoWr0ZfFQft3y1+obGeUKbHzHZugvuHBCnXnHnPdsff
qLAVgcAhp0imeCA3y6y1yBmIik7cVgJ39r1MjsccD/URe0lI6oP1+G+VQR2aeRNNZXXqqpTiZnBx
0WEQvyXR9o8B0s33UyQKUfZA5PJ4au12GKEU/9Kg7iqNL5iKGaZYZZcJkOhi8my3FaasonBeIMOd
yAhiiD3l3FgTw8CLjszpAk7OuuTyVDx1hTqNzwjXAO6jGu0Zp4U0PClxDz1O2cZqENBaVUpGhp26
x6AIwzwkH1/OG5AUjnemvrVA5ARDoXibOv1weeZNG4931PsNHZutkQX5E0+eKRPJDr9uqdLYU61o
OOgOrdzeUmWCUuEN1VH7V5izsU+XiWfgZVIx5XhcYQafd3E6G8MXihCUv2LCIfjI1JpWpmrbJsHt
YpveRMPaFUqssneZ/Lss6KB84snuI0toxh+qgjBEP/QlaVB2MiodPXtSApzIzCAjBLEFJfLTUVKI
wWkJzza2WrlYUdjwO44XZEJxC5g5O8IX8SuXCfYab1i23f+cqpD6ZsCBYQH4MUNSnDzN90gGu5jq
i7D4o6QH4LXbCJldX1NS+tWWgip0yv4rwi8MoiupEmmCpReAeNvAhY/vhSnhFIrnxptQGypKbnZG
PCjfFnOwziWNtRug5o8AoVKfp7QMkLZ1g8wO1TM9rHQEKS2cOmoCiTefiRePqg5uI5h7d9TBCUWS
k/EaBPMzVZmg/252oyKuImFpyZonNkL9cqYKySz2eyhoR0+oBkl0fTGanHRqxSkxxUNjj0YXEqAc
s0/YdPB5sn1Z8Kl62BpTscOREz7BjfX1ReNi1bhUPggjGX9bqD1JJ7ky/ZfOwTYX59LXG2sSE1yl
Xexiv0KSuzfDAXBHpK+qmsrSTWx1pX+Q+4wMu0GncLBZQwzefnXmZWglSp5xipv3u48iHer1aPTu
IhS32Lq0MN7lwKApuwtqjn48IekhKJ1jcuTzqVnVbeGPYehFxVEZl0elLmNGFpaPOaNiKRrAam/Z
/6cFLbr7mxyLL/0x393cadddyWolWak7DnkA725V2C3zmtzY9tF78fiuP2dhiywMYiwd6xrHBHve
1NnNYGnJVEYT/ThZxaev46b8fjbGLPmnKm9braOAxIz3pet8Y4I1vM55Ihh+daVVvxfU2ApCyMef
WS7lquVw8s07hTs8ef8YfuAZkdXcqoah9t5gzmHoX8VrOk7JW72NJIeTb0TGOJLR/M9ZERJQu55J
SQDuK9v9Oi6kSpYYyV88b6Kq99eligyU2h5ORe8Fn4CSLgjxSeO/b7mszpAwSllUQ1TSO/NP6HQM
kWiOQW8P3Lx+L6YQQLsp77ROpvDeGuLhGNSFrrJr8376KvQhJ+7QoO/irzKsVYrUc3JFygEtv7RB
bfb5y+AYLiGS2mNwhc6D0DCxfdKTa2xdwfWJKTDMPIl3/hMVe1cTR3HDEQ6rXr1m/d5eCxW7MTJO
cwYrCXmg18xYTSS+oB2aWkXixGJi+8bj1MvOQLf397hNsXtLQedb8+eC1IXIUjMczL28vjcjdGcR
RbxdtQ6H+vU0XhA1KBbdtmbKy77erzRDqKtZlutcZ2fE1GcJdcgnpWqVqmKyVIsPG3Yd4t4n9Nmg
MxJkGFx+/g50X/I6UZvbojKCQcMpvNUD/3/DfNwIoz0rTLi/JgCUKVQgYK2dgDn2f0437F4bUVBQ
+O4g6Wzk4RGz1ocNTVs3AJHU59fiIzFMv5ZXuDVJzjGukGvWAPYPkturWSBvKAJ07Dp8+r319OU6
/qsUlALXee2fUW0oKSYxN9/ZzOQNyDmhaoyqSeCZqQ+vSjCKUx9IP1Jb0t+vgUY63x44ReRJkdZ8
LaM3ll3VK43M7wAZAE9Mzg1UkTzbawlSOhMQ7POGFK4z2tvLwsXNG95lHUH6VIl/0Owx46xXjk2A
IYgIIWABEV+zsJ9iXR5aod+79GXTcdoG3DGg8s5Hld0FA2QLxUbzqmF4axPqENBffXS2SIPfxTUN
SfNzygCUWsbdOicTWtTDiYmJbeXkg0+G80z7tQh77LmQx0g/oBNyTx6/R1O/VMjaoAHPA11oy/eW
Js8aHQTTr8ezpW47jFUZdb6VsNUzqARfbmn2OVwCc7VSsc1hMnJwWbeMCKOzDGfiBe8/zGKptGnU
oXuJrDTcsdbQgtmyFRoY5t34DMXVQ7gqRld8AOw7Pg4Gw4EYCjuOCud8fzv6pR6BmItgI2sENrJC
/YYBdxRkLdKLAky1DiXg3HwlY0G+qXT4zTZPofc5AUBIkd8fHezlbfDC/1TzWz7R3TvVyeLM1rJ6
H67cXvFKFGqZbVL16OAgmYaNe/RTXGgdYEFtiFf6sJbG6gSoLcxE/0QX645FxZCho9CyZOXxwt2N
IzzKlWeDYWqwINlYHTl4bZ31ixVkmEfP/lIuo7eecHqEjb4EAmYhKJj1OSiALOuixJ4zknUD2avq
Xsffmvoi/VhlZp9OaeBqU2MXJJBwcB0Fs6/IzoRJAKTbzqWJTj2Cffqt+6vdQt+sKkJfMztgX5bk
3X196CNBPc+lUbHM/yci3cvc911ymUJlR43reAXvS16bb6BZ8roseuH3Mmc59v6HFJX3RFOMCsXg
0ZvLQ57V9bCHRSxm3eCvQPCZ172YberP71b3B6+WEcKWRumGVTwhDzGYX+rFAn3jD0hMHb34QQz+
c2/5xD0stFJnKfrJxYwJFX8RPiT0M3tC6OdfIU6ZK3VuqJrk5Mb0MYO186OcTdfkcYa5gX6MKOjd
/4Tif+I3c8CTuKSoU1eX/HdgG3yokPcNhwsH6aqfNxATuAUmHGuR/9Jie+cXrFTBrLRk/94sOAwV
T7yL6Sx/jfbcpstw2fkI0WwqqpF/BlZGFCJdb4vfM26jzoRWe18QeJPccun6jodhQvcMdJOYBv5e
J89ce0TxZVAr66gR85OCCnHIngJ4Xzh9f7uoJ3aj62GRzQMdMGhqNUBkOy1qQGTwi3gmUwVX0HgT
35MxNePDTGrYGUA1CaYN/AAip5UPsbngdew0r52YaR6QQ5Sp2Lgay+dg2S5Op2khgMs9/2Pgc4XA
UszVSryYWjQconXkIcX5WlJ/VaSMlqSytPD/auBJYe2CQeOhpD/1lcYWspzxGg9ppYV0athPYSzu
snojLV1P1SHaa0OHFHYnPhjHeBijZfeGsmyo+U/xIPKPUtAYZKd4zlyRQOPSCZwOFyRH5t3GDn9F
PehbrKE6kme4dECvVHlVJIkMS+I5Udh8OMFuqzpqVKccezT0zuIAPuKenSOr/beAlevzzo7r5FrO
IOva2KDc4AsLVuLCIIiPDDlM55WMQXXun+YcSPvVtFIjMXddE+81rBBIID6u+qw37XN2tAoaFcrX
lcGHJ7sAjlMvNTx6syxmodbIXh4p/2BLF9E/6XgkwHk4iWbtCVbvoa4HscgWWsh6Er4DHkr3Db0n
1Q8lezc8CNCNbfy37anyU90SsEZmm20y+b5h8RX/KiwvtkIMMkP6LNak/Vvyv6FVMoSley71kfa+
TMGdVfpTkUiTvduKpbJBFhGuLFKgrDpXRy/+I+x7lUXJdV54eiOHu/dXGr3IM0e+tcCvD3FcXzTl
QD6HCMCwPmLsT+r5wf3Ru9tDRLasP+z95+31V20iPoKdLQ1DXARWH/0HirUuh1rHuEnOngIsLIOY
G16EB+1sEop8L826QtlAdVxD98CSVv8EIFhKOhoSM6PJsR81sOK5tObEqGOC+Zx7fwS1noRJiZCN
cto96DIKtmFJonn8WMqmMjYCas0av0PT0j6NaUtDM6DJ3kso73TtIvjT9QV5lWr5JwRtRq75muQv
PlrI6iHDNNxcvb9kQDMtgpXmie/tSZv76n7FkuLG8vJhwm/VkSOBd0fpThGSz/F0tdRDO8QJjVg1
n/0orhCUknYlelpvEgScqELtv3k9zpH4jQLVHvWonpSoUV8cXX1q68Inlk4W7Mid0nJ0+KEz1Ss2
5r1T78Rvw5n1kgz9TKVLueQ7a2v+Hl1+z0hn4+6trGuZn1NtYoMd9Wq3n4Jv5NOkfD3JPGtXRJP8
no62eQB7AeKwhmiDfG9oq9hblN3FFYRQ/sPElmedmgMWUrCpgdlA6F3jENplmhUUJelTrYYjqsYx
xSh38KBTDpAlhhyP8/AYXaAGjV9fVyF2XfcNIGeF3EdnSvFbIytffGCiLR5aALjkxouZm1UX/0qf
03/mKTuj0mG56UhGA/QMjeYPTh8uGQI3YQYDFp0p8ArmOCwA6YV7BN//Fsw3+mPpJNm+GYNunGLL
Y2WPg/0L4/90FbjRb8NhYYBpCdXkjd9u334Vnbz2qanNsNQiJByO155Rc7pKNoGIUY5L+rHBdFZ5
h7PkJcGLJOYfsZcIR3xoNxnLGsuJEc8RiyIuTKPc+GuGZO1kRMNO336ddcOzOx7K+2xkh49JiJUo
ACoXyVg/wgDbeT/q7rLZuQ9lWaRRhR4CZLhZCKXNJIToiXWQFVj5/GNzorxVoVexZ7+ptYXLVCbk
ziDn9gPYoa9dXV5SAfuCGbzb059ReSf19wIBGIA+gT9A29mu0mxM0Zk9+u0VxSV4Bz78KZBtj5y7
6sZd3fQqxz2CChPSKGJJOIcz4IBIDIC8wKO45s4vEh1UrnnWnY7bNEAN6jADigHZpZgYn/YXUy1x
iCZ1lcNwyEe5HSKNVDXzDgcYTkiJJdQOZBiEjxn1o52n3qNUXlqpsIFDOHw9x1Fdcu0n1jJgPmPk
sAC7AM2VR5dybXZ/EE1VE58wo/s9WzZjeQwGi0olnWaFJdUsSSPVP1cBXqthV7tmadbuRvJ5KaLG
yROmGDuKOlRGGElUYgmUFD9MlhsRuBIglCiGK/afSH1QBtuk6Jx763jL8c3H/EANi6Ej8egwugF0
GPZOVpcfwbX90XS+JEkPoM2ACNp9CeehztKaxBvFLxIwr+7CwLtjgj3Y/q8qANY1RsJLX07vIfby
m+D+gVAEHZ8fCmIkLAxtAVujFEDY6nVbe7NLbLEwr43N3hy5hldXefSvSzwkq4xjSS/VUIk7aWEx
2GyN3eDPzq9NiSL0Sv4Nnrx1mHFzdY+QpPnz18YYzZ1EP+Bocv6qzqoyh33+Ys2NxtsVhyoNN0CX
cdTQejiu/NShPLM+d0zMSHO1PGgsuxmrSPPlm1D+AErGMmN10ZJx7pvp972jEjT/UjXkf79KFRbb
D/FWUejkah7gq1gClCyCLm8N+XWHUODgGP7kVSN9QlI7UYMFIYeMpSxFMBfl+4Jqb+icRP+t5mIp
NPDJFjv6K4g+C9egdd6ruCQQLRINB77MFG0h++Y+dvs6es4lB8YR2BYQfOw1A5Xwk1kpxodx6vLK
zy3CEfjMXbgplCuy08ownPqEqFh/20OC6fz5kniU1VTRsKznSDZvFrSlh5TUk986LRE8AWOEa2QW
h0k770+D7m8rWT0Sl/7et9rtllNmSIZHuN42qUWqmn7itS0oknVgP5bY3ZbvFy4ZZLd/FODX2hxG
Fhd990IQtIz99x8XeTtSGrvXghr54u/cWYcJL732izxuHBEi1q9nQy6Cs+gA1S2RRFQ1/ouHtX4L
NwcNZxKP/zfsRXgJ0unAuXQSHGk/gYFuvpRt0AFkmlil9DZBlc9NdzdhJk4tTnb+f92MiX5+Vcko
VqrTGge3LWMRpj2X78jfkQz0sUTw+Pjr7ZxIgEjPK3bd70Ta9ZoZ46L/QGSWXxyEhq3HV+Tpf4oA
3xSZVaYEeZM7ul/20k7b95vpwhMMqTuttO1hrWJVGVDQFpl2HMzHgB41N2GXzksStLPeodVxCi4V
7P20qDyoaAjxz/IjGmuX16vEoMLzmzle2CwzLwFSyVsffLQyXWEnn5fdF60uwb4MWydYzQs2m0Lv
NEOxlcJ9f62B3k+KBm2gLwfGrhddk5ox/WKnBIz4IUQHtmyDBHeG+9Y++EkEMSYw15ucRKhmzSjk
V1V4lBZ4CDsKsqtwtA/hD0hID7GrdxBd+iCFtYKJdUSlBjSoez3xuHopLgpXA+aCggO2ymQIaqpw
pWeTrqzJbq46OUC2/sRrhvrNQLCPg2pfSVpo/OJodQnZhSvvn+ngsRwuh9jFqqLi9aLOm4DahlDA
3eZrkI//L/Ghw2jimve4bnw2Q7tje8fZUtIaikO/V3DbSrbONMSM4USMxknmmRvxrBA1kbAS+3CN
abjSACiOsIu9QavaKnpCSVsCsCl/pWiyEz5wWcgvWqiE+IrQVwaEtrqYTVQLptNXgSNGvmiY0wyB
L0dOZc5Gjgcxmgzo+ErCrvYsVwAhLpwmw8gERawe0IELLP5PMM8iDb3XCHtnJSsLhEWqj3IKBlKA
7aVKn9YVUXmXk+2e3D5zqUQThrC+u+PLNVakppvulobJ+ZfwFEoYcyPzGu/pqV/H3dziDmVni14y
s1ltDMyZQzWETqWD6fkm5Kekgtx8luBsjY+Wj31bWHYDvnXZuukhkmp8TggBF9k8jdtig6V3A86O
giSvZITLOctC17mddLraWH0m+o1DG4HoUKMVpXWOa7Zjo1MBZI5dnn4A42GNRw2+mMpeDYDJQnwM
4ojzw+bkKny+nloMorfHaEyFFgqmUuNsN3hvld9rDDRJvwaGjT1GKyfuAd0RYx+8ma7Eu9sPvH0c
/lTaJ1wtUTB+RktVrq5rhsdvDzBp52Qkd7CAU1Z1vs6aQuoYuxJR+BNV4ZyKMnPljBKGNTH/XcuB
/ADnHaFzmyYpbj0T5wIVWHRTmIVIqj5gN5jEQAgD522ics/2gQPhO/0chonmqbBlJAaRAsHvHtOB
h2vJyZe2pcjpEY/V9B3c8CdnuEn4cnNc+iEk664WijxU2xOStf8jIeXKp/amHlTQpcuaJiF8mGa7
h/s1jsyfXXGMX0lfXpgabhOcerAZADiI7ad1KsEiBgBJsOJb29h+Grx8WJRRbDkoF3D1h0H5cWyc
yLMf/Kp+z8iyfhB4Epi/KMuJRxQT1VoJlz2jWkK9jhhZg6uYlKsABGrOL48SVxr6RAD+roCpaXfT
SxceXuuHDG5UF55pEc79qd3+I68cAveBX2pMEzHQLakA7+UUTZzVH6hTeDqxx5vDgcaSbfRUA29U
JTVdum8sc0WQ7Vl05Yoiazo3kJBOqwTTfVkieF46xyP1ODX/wxKOpgzkg+EWRX0x1Zu0ffjWM43C
rAKmaqrJk2UkR+y/1m2rH5pxnNv6lxTD6JX0jD1SLwYuocddipBGzv1qbmNhVtgTkdeAKDFlGTQn
EerJgwMDNlwhdbNyql1OpoXKFCO3kNjUXiq0ziQTfXRewMIPo9SZ6Ti8H3QU1CULeBkzKb2H+GuQ
EtgX4gzd8YdQYyKre+oDbnBE+Gpupw4efE+7XpebHZcftR+fHcpFnrL8+gIaRn2AgLr//2BEuwAz
TStFv9PGj3RxzCIz8oBqwgzpSsogdm+Y6dFY4kj+OWTEy9HxYhq16LS6r4lpbTHOhpUs/+doLIYs
eu947QgPDSVkvOl8VzqM4XRzGYzXWUZ24Zv6yYw3ppuPgJlb833qk8u/yrA2Dtof+TtzZSTyKUAj
aegnVQn0bAjoPtk1so806VAkISofubsaNPSyMc18f+8mFo5NaNqZD9yZM9QNNAG0PTBAa1UWwe/Z
obbOkLbkewMxyh1qWVafjbeAykRrlIVw6TAhhtVmANEjq5qZsCLuetPi/d72q0V7bgP0OYGfx1ce
k1JkPPpxr+9DcowHUg++6MdGaSLnRQqviGQ5G62exhTMj96vGQePuT/O9OvRWBkmTO7EfOBroDwa
xvT6lpNN0vMEeEwlmbFye+1s8u6SbNBWAmVAR/fn/LhowCTJ6TwRZofmlXqnuFoTNmKyRi+z616p
ynezrc9EyTxTzpWj7c19g0d2zV5RwKwTdQOt4xZSbzPD9ArrjK5QWddsAKA7wlzszAQLdYFhbnME
43VrED6Lzk9tdPegsZ+CfoIKMlWE6FIm0ggY8VQxTtp4upZmwaR7cD/R8CPQaoEgS1BgxYaqIXzZ
l6yHXaIIc6JMWR2n6RX5KxkVlBd7r/9k1Mdc51nVKTwBrx/Ltij/uqHuldgEXM/K9K/s/B+r3X2z
LaDqkRcmufYZNEcZMr4sJqLO6LsLteviUzbltJv4xpUttY/PyujfTU6IxlTctHuDOQEwSEj5UAu+
GD4Er30vZ/VqTTZLg/Ats957IRqZ45aLx4szrdy2ha3Yk+5oY3KlQX0wfNXdOAB77z3AVJ6bDREn
Q0MufFH0o+QAaJxl3T/EistjzsKRddYYZ2VIIhV8/5BZEwqvEV73SBuTVUSAMpNymh2iQuAuwNq5
XUVBONprm10lgb7dBktPOXWoaky51o8HTc1Gj1JdL9gKxjP9jCQjVErKHumGf2Pb4qkHg3gLfEs0
78JmX/TfKmmhkEchFX37EjVqMnORmCPzNbjW+KfhtyFnH9FR4x9sTCakZltdAg+Wc3HHOq3Y2mnA
jhgoX5kJ6hrUBoGv/bj+c95ImcyThm9vbuVsphkbfbVmltfo+4vOP8DtT9QGlfhrzsHrtxYHQiWb
Zn+F4ZLtwQUwCKEivorNy6gVsowGKyX8xpUXmPEoBbyxrLu4fh7Ulig77fCX02kyIrwtjAISC/0H
ON/CQSQyCv4cTpQ0yVeVwUXSeUNQeRKnTMfjRFZ6znu7n4pZmXrjPiJq7TSqOj3V5lLDB/TNMmjV
ARyiIAPyNl5oLW3YlYFcsRtkStYZSXhkEgC36xDLCoxzkkhr7klykAsdD117CSlz2TyabFFQuuH8
jwUapQArJeYlpJQsukitqMtIptJ8Gwj/MmKBLC4ngTNTik3ZdYBiaRWa0MYIb8HRRoDa83rlBB5w
wR3Qc6+qKqo/wUuBHCqARHkhJ5nXuBahHlCyTZdxlDiqWlhEVWXFd3WfCsejDl6SrRb7bj627Rlt
JZMhyRjY95mRU1mFY0c/z0cS9DBkV8t9Ftr32LBn9Zh+2pDXyz6VtEtl1Zqo3d59u562/MKwretD
2GACJHXZfX0UfCQqvPYWwZlqPGTmkJUTGOETt3pZqVi7JtK1+dGTc8MHrByO4xFyMv7VAn3JuGRD
hTFQhAGcdLW5vf2N4RoziKEmdi9SoYdFvXi61S/UenR6ggMctJtbt2Yn/eW7z7N0UXjeva8l6m6j
i6C3MBUvoMkPmD0/H14rMGUvhMrbLPUK7PZrGfk6B6opge+hzqCB0yNeR2nl7ppf4SS4q9pQe/wW
3Ftb2/kRXvmkTb4DgEpC6zJzAUNSySDMpoqPmVahyWxbMhfZ4QU43gpK7TVwNueK3AqcpLaPaOs7
bhSb8zr4mh2EwcKOxi/zIVrCoRyrVPk9ZwOKRBBDMd6ml945CLm93DgNjTs2LZ1qH7WdatXe69hF
d26ty1Jus6GY9S81DRIICe8nJT9CfoMdCd8oLjubQaKwclCU5igTv3M28bjghOqGTOJoQzrMYuNi
PL/42bOH01+QzuqV+bJVh7fpch8R9KcfdaCqCLbCnbKEpDqzeR7omzJMpxYC+XtwR2bbLB7pXkLF
W+8hzFIUo+CT7Fszb/7NPv3wlOiN9edMtpOSU0k/b7wn5iq/NqIq0PH+jhDutQUP4AuoWLqwWVd8
b33G5B5bjjPbMHLSkojo19hZuH4YODroxoySgTV3/WRNeupy9B5lH5mrqkCvx5wWJOS3LqgqRtAg
Ex/PVwZCsw/Zdrn3tOwJVlDRn+aKNksLPUfwd2CDev41bxin325mX0qHjlaYi1XwFkkaGCo+K1iJ
ZvR56C8xrimG8ye/S9s0WL3EM0XSInkjaC4BbDikFraB7Z8gphrnUbHahtz/P96jes1+Lb79F70K
7c4Xjib9NEwXxsIlqIlTKNr6x7BFKlj2oLygk8PgiqXrwwLuxtWgi69nKSrJnpAWdXeuBuc3+eBQ
Qf97JlzeZqAPWnXfD0kLvqFWKhAMiWrbf+hmNGe4uRHOpnhtLSpoTee0veESLm3wMZqA566kGSZ1
nwQrRjPATAVigVS/wqPTL2Q4MuMO+gjleIhoHlagf14xb72CVbCXOWKUBuzmnM9MXKdpOxbowiyj
i92hgmP+x9o0ZP64BAzFo+MuVOWhFl1Jb4P0vUOzNzRGPJ+Kh1ILHqFHo8AhMjGjxv2Ea9/XL2ZN
t88w2WKmnPeLGTDb9+txVg0du/EO2sVLMRX+KpR5J8j/XE8aikS3AkhfhcC84m59ybs3Bjnw/r4d
yjuK5pY9OYW0y0Iv5M4TfJ542AAWxuMzVgcid67zqesRGtjggiIc5QBjO2knQD8xwsF8hDfZ2zSp
9H+5/GO02R+vlrsEXVhoKFvqADlw+qfN2q0ShUfuIvJhMxTTau2Ws/tNWYcFJ9pLkVn8viIfwTu1
e+z+iv+gvIABEuVfrW3AXBR2mxi7/pP+TRNMmNcczDIafZvQwtC0eFj26C4xfRBYIlECQopXJk0B
/NqcekgQpulPL38TkcyeEh5yor1NdK5V6AG/ilNw/Qm6+4MXqcAweKYeqFgX/89MezlYHMEoICTn
PdwI5WzkYUFn72DIxUYeijjsFLjPUrjNg1E24Y4J+1z5Q9yPndOxAc6pOR66zbDxe4lIqakJ5p2l
U6491+58PrxkYf5wSUWkJLaEsaQvl8eJfru5LTHhAdOQ1yUTWgJZiQqF6XrsTuJgSeWXuCnhLrdi
495dOolteGdMDQpfILbWNJnnGjutTtKNHk9bTdaiGmucYD5PB2kh46YyckHBLJF1BF6MZq5r7zKP
vS4qxvrY7xDD9ui0IuSJM974bAdk60qMTuUJzvyBptitK2MlLNR/QtP0dV2w66kODC4uz6L7WBIu
WFqeWsKEZCFKVSRWRKcNkEhMkYuYTJC8JS/TvfGE0v/nm8nZylgI51NVQbNYA6fE9pbcBcfiOMyW
+lpmUYvpUWIxKf2JDckv3DRBCGTFOViIDhfjaFOX8CFQy0bSEgd7HRlIP9aELMGKsrv5P7H6Neda
YcUn2VrVXizc5XtaZA68KJdJU1h04DZU3mJ3Ztb2IiPcsOPZj6tF5yRJL99DEZzslTWE/5PECQxL
/ZEdrBmYMndty1TZbe/FQlXbAmUO/FiH7xEowG0a9qU99m/c3bxPJP7Rvkg/dCuyi/igq3ZR+1Ow
FaCm/wUuMQujyD0FCmYKi4HAnLUdS+dA3eXYiACEbsMYzt4RgoKS9jwkQtgwei1jjXxsMfi3zjeJ
GlqyLQewAgybslMjPkuPBE/xhE0+5VUdk6alHsMmdOoa0pEo/x0zfP5j+xmYZ4fqIpggNrEWwp4W
Cnb1/jfC74glUS67Bd/I/9xV+BY82kbGwKd53lbDv7o3Qz4tjh166l3rjZ+7BaShy2pzSA1KLL7W
YtY/r7W+1Efo6c9myiwkoCpfZIS4Ovh607N72HssSaJzUiTwSYQYRC1+6Qew20XJ/RHGlPPEm4oX
QFmwUVHDJLeBTTCG3TnkfkzlH6Xs8jwt4yPAUC8nbcYb3NVv+gwDqPN120bp7ioEZrBX6ot5+zCI
v00GDcR1UShN6V+AoOVD2KgNzNzqq7ZifOW1Y8H+6BPJComokmNVicsnmQfjNcwm6j8dog95Q43Y
9Wtogjso3j7Li0MA8nLE9zgrlt6zGc7NH7fvG7rwgbRCzEoP9aGlS6qDtphVeuzAXv3cvFTnh9gL
uwfn2ufWQDJSR1Rs5HhtixoTaDPFHKCZqhs8bQE42k7nAX9LZ1xvWTfOAJM7yKd9EMOmC7UJc5JI
CXfcEhTWS3d/ksajevdJWhxzNrvLV392IKzlMRMz8w4gxDJSrEWb6r/1iCT+dasMCknmVRNZKfgD
NrOMrlYcqduH+3LpgQL5nN1sgnDenNgYq2TYur/zMcrvqwHuto7NxvUrI/EHjmamW2913TWY89TU
P4vMnyZQ0SUJuYn+N36eOOLVIxXdSjelRUwpXdDLCZ/LnJQWzD0sa4hq+3KhdYG00PVnNJZlRswq
n8S4PEgMfbdI4Mm9j3cces22UZ+8z93Wgz+2p7GEdoGD4dmD7qoBeoj+YLLfalNHCAR9qmZTa0Ng
2qNd14KPWdfSoRiSW2rOhBa9AVeYQQx3lpIEspoPqokn5CNjTPYbjWhqf64niZd5YhZl5fVdTHcd
hWpu9nNZkdHcx8jIOzgdz+Y9TmV9VJUGFPO5kFrR31y0/F1kTalKG5QdVl/0HyjWU0Eu7kWY26yQ
L0KquSCDx09sZ9bCbsTx0uQvh9E//63AdauNRWPJ2+5mo0JSaqgNVvVzjj8UmVZMdfpmUAFyUqLF
y4hoTm1dm84NdmbBH8Fk/PAMZc46CQy4wDOjerVoFangTFR9X2r5XUqJMAWRK9+i2NThdUghVITp
rmrSBzT7bgGamhnbWxwTv2NwmTpN+NFP5Vrc3DDySDFj+6zQjYwLez9mi5AdS3Or19gnc6m+pTYh
ViC5xycHTiybrCnlt2aFnjqhZCk7tGOfKWh3mxoBKpGBFfQUQ6XbnA2pv1OEvREOMQwzyZdL4U3b
2w8YT15SWsg2XnSfFPNT56+prTuUz27bdV+ueswekhIX8CNJqfcmxSavkb7nJL1ZHc23NyAZv6Q6
xGmzJPAvNHxRl6TgM33ECx1iZRxnrOf10ntCB47ck2lcdy0Ajc5lSd95TZHcrfavHjMoZ66CmtFk
4A+oRP+cBgyMRegU156UppT0NoxgdonHaMlwypxtfONqmxt4NQIHvWSDGTnZxDwRYwaOby2DVarv
+2mjYCLBObTxzL/WKpgvRY7WQI8ZUK8fs/mbc497IEB5SWMF0PjCZ+XxPaMnI/7DEStewlkZwcHS
/mlaoQiLaWiqe0Cy9QVHcSE3k2Vx45dAfAqUpcTvni2j5oMuwM/LnCA0OkVuzYbeyMD7NbazTzhC
vcViEcXWwfL0Xiw+wtWfY0v88eZ/eoRU3ITG9Btj6yI4wW3KyXV6m0VhMY1WEWpsrCO1D9iF+JAD
+RGsi8Uk/sPZHyv3RVFcVIL08SEbYwWQIMGNzBTst/oL2PeCxAEI6Qvdq30IAAsTknoYj1WLBvHq
owdkMENG8NE0tPCUnFDuYbie/uO2gNXL+EOHye8+7M6g+hlmjeY+VBrur6fneqrn6mMz9GLKsbss
la+9DwVFokdrEp/0NkeIU01tJfyts4XmYAw0aXQKmspKWT0YjOT8Y6ray6KaGoJ1SdP9Jiepqsum
cPl3SRibdFUtyMUJC56gqxW+y7RnRHgNmksQVkP0eXvHk8HDUYq7iPL41UGJgrKpIVOTCTUKIUvz
j5U9AsT4bWlRWAgMdq0XjC97uDhON49lt8N4Mr+Ca/PLszpLtLrw5mS6UgeIjzdCowmrw7vpePhA
+20MnenlQB3B7J7rhpGhxQ/pfNIGpWOWXummcusGymg0BBERPjRXzfa/PTwOaK7uCLFj4sz8G2sZ
MXbvFtpOZ2okZ9EX9zycqBRAj10Dg0yDtR2xk0ra/tczYJQw8exlNp0bPoLurEnuRXoj5XVuJpZP
L/YTaQvpiILCbjglWIak5SV2r5qmsxGjEtIJjyvRb9amVF2aY2mL3K/ZWqvV52lHUDXmurbClupL
q5LZ59SOLWLAQKwOlt79StSOiax95WZsBOe70D3XBKd4ULpPifeuneqMNgiR02us6zzplRzmdXCV
CqAaPxuZceYh/qW6dyq5RtOh2Xox/yk+yx+OV3AMFfKjP2kW7XmnBlDsXhDOreFUnpofM+65YBx1
hjHURSwH1Jh+Kz8mCB0PLKnglU79xEnLuiz7WrD59vl1qYKeTqbDmBMg+tH0KvNp+8capU8/31eZ
cdZy/TA6ho2eR4W7ELktsAnRwg2Qa0UunwrIkhh5bLTmCQuevBSPhF8ZS/tp+Vimrqmdz+53D571
NHx1NiPV0daCWjdZ72bgslHhOmT0ms+9Cs3O+9v2zFBH+2Y+5FZW8IVQ84qhzmwdosNJABPa+oZS
a72TaHXrQgxsIDgGyM+2bchZe6nivSlJ5PlfWtuVVYSEr+hjgW9beCbToyQrlyiynr/1kCbcWON9
bA3VXJZu0eHYa4zA5N8f2GPYRTAW+wudOuf7dEDFLGF2LX+3T1l9kDLCcIxJOj6IvzyS3LdM3uut
ARsEkongJMttFiQkjsGqkdeV9K0w96/Ty/ifrEq6gwFpb+MMfjFpPGMzJ7IOXHXfvm8/H6JyuG24
OhvgakQ1bSuT8EofxR+IkEJp2z1P/E3MMmwLr33J7He76rke3A4BgXhhHGmogeJN+gnpE9LAGMsd
C42bbLiGSPGa4K7vCLXRGcsZVAosVo72StQv+YkOedcORBqG1zUgdPUV/6AnAew16zmnq0+KvGz0
cwISKyNkqNbpJVNauwd7USKk0g6y6Sqb9ncHaAO1LrQu4NFjDHQh3gAJ/+Tr4wMmm6eq2q+r0QRv
3zbrg3eftBf2ygWpB+dZC5FBPyXodBv5QXTrTGlItaLSD+BlY/u8BzH2k+Gh3DFl9HxL5zWXyAZR
RJPLtKuKabgdziWOKMNBrjfHyeUrolSVWgyZJNpnEW9Afkc3ky2kGn2Q2G0NH17ces0ftDBeH074
piZXRbvhN61PGptNXaI35oXJlvja8HThxpI4HY6DGXMD3uOJW3+foeUo3kzANx08CQg1CaCwxdB0
H7HmRqhg3UngAX+G95dqu0d+CEGZoSNeTeWYEBnEB2e91B3/VaHcJsPZGKQTADDW2S5WkY3sKO8m
50WvZbgFCeg7NxMlMjK8bA7kQvbhi9IG8AzPO39hB+L1tigvv2kj955Y/7Y8KjXGpUVX8lhWYKpu
9alQl44ej0xvpqrXowePQ9Q1Hu9UHeLltcV61buqqVE5ljtrjLOXBHUzKcpoG6lXiV67Ms1vDUul
SYk4pMaqaXX2Pnd0QkVvEsYd6Px22mu8ZIH1P4XyV6L36hxJgnNgdV3md9cZa9rksqcK5UH7YPP7
Hl4mULtV8iHefQidCXpR+c50yXzrgVNwBDZJBhiDLneXEGJT16TivGLJOhccwolyQnlLF4NQ2PWg
64yKPqATGN5+WOID0MnYhhNIN+OwmpLF8nj7hjjEIk1/hh46YGyagM5FJF4gDMkUHeUiZoh2SBsc
BdVPKx//8/Fp72zvjhyadM5LupJK/ZFGIjwKtdZa1xCXyyRvNkEoqRxq0cHeHJg4lycwFnkJ+Xtp
YuV1KxrVNcDg84gQ7jn9yNaOQlc+uTAQ7SZl1I5vTS4njMBfdI6YAKEJ/yYhw6TRvFOzN5faK0fy
6C0k0nmpTKL38/gNKyTD3StjE5V6/BrQNr8C2qS/of0wHvi3kD5ian7IrSr4hq6vn8GVYF3ZvNH5
H6wV46IaFi5EMROXtklzgsvn4iz+6dvBwv80F/HHvx92GYicBdhYdbIvMrKeKofN9O+3i/hWsjFt
6rNOVM/VJuuIOKLpoIjqPbdlUrfNOfn5wPYEmNjtzyQaeNDcjHLB01sQZEzr+YfxJVqs4TiQuszW
gqyAlX32C6hdCLA3nLRXf3ZR0v0MwgkoX63huuniyRI7GWt4vH6W1kQZLlA9/Pf2RB1zX1Jt0JJN
05XuGTUbe1JzWNKD5IBI4gv+NH5jxBHpa1HTI9H5T+fwfzRRosy2XIGBrtPQdbu0QoSMYGJ2xhpt
/emBzVg9WkvGfnrb3i4RKgDkG6Isl0vjHLA1uR86CWCWtD/TbcQscfnOGYpKT1YsT+H5i89jvsvj
WFcdoRZaxmc3jV5mZDmvkctEEfD7cBYRn0t0nLy5t6U0SDHSDuh3nEGJKJi3RgRpTg788KIA3acK
6pj+uO/iW7vgZGJDd7364B/eB68GcO4avquQFXbxrlmYQikl+CB3Bs0hcmWnneoDQNzT2MI340jB
v4vU+pyLUcA5pxyJQCpXdw4pTaA7yRlLAH4RraJazHrajWmHGqIKcyCS9nxLW8aFNPctmm5o/CUN
Gwm4Rd5BnIqjwzSamkxbVXH52Ket6AJvTeFVkRqkwhxNJk57KiNqc7YhrkTRtkv/TVpJMS/w4AfH
ZfdEmGaLvUwuCbDLyYXxLmydNLp+MxiYQ8RQYs/Nn+PqH3ZmbN2Ed6He8PJUFO5vCZqMHa4+9jiD
C0EVVcsr2FfYafzkJCLdKtlRTEmPntvJYs3Ynrp50SfgFZJO7DfHzcJK0A0/AYu6/Dg/y8ojCGxQ
kDJZHZNVncf4EmcqMq8CHQNzFmepejRN5/hKgevEGPVLBRPyu8AvDx8Jw9jJ/0wzjX5IjSV42B+o
iT30Kw6qoFQkjURdxdrZkMfQlJfDXmF2hgoZnLKTRbZuGjtnHp4AzM7WVL9nSnFFvxtgDo4P6KD+
ROAn95R3ddjnTOjNkSt6TmwRsy2N27xqdCvhSXj4pUYzRfjSwrER2j4n+63PCkPP0qf7q85bUGEC
VyP5nh4r6gLlyw36egHLN9gj+jDL10tPmf7uz2/vWYABwXnI2t7qO3WoPDazvJpMwP6lD9deNcg8
WKz1oZB4KpdWSi3X1faZJpblUIKh+VQvXwtozysqeqnWyEWBjkQ1j+KJLx+2ZneHHvS1YlNkaBJZ
G84b/nedPOIPYCXhSUxisuG2vLACGru+PBD0XGmJfpfRFUJ67R72w4BWsHhnSIivVu2O6JJQkutC
yjxBF65xmMjDaPTqSh+kKnPNrBpe8UMi/YUljpEhzSCrlRGtyliso++AJnTyqb09KcpoIs0cJYwE
wEhxmjnntV50cJbEC4XjSVdVIXradmIYqJtq6/F4bpnl9Po/QnA/T4yt7cOzicRq0XCpqXIPLPdB
JfuqU7UMU7+7gkNL+sM4DlHfhnOhw/JIPSeBWm0slqTT+qappfO+K8aJqWwn/mDEgUE2tkEFQ0af
WvmtD+KzZOZMRd82yzM1AzWOMeiJSMW/KwJwpoYD5G0mJdgOjxmHqjMdgQzf0gTyBXKqkPUrnZzV
Of8tTSjaxQ5QK7fKpi1jymjuvEbwGNztAOeMs/LMiMy98F/hgbqfw//nQbMtZLfcf2oDz9c1baPo
JGL/Y51M0W6X6UIAt0zzxgsVd6hXkT8txNYjBtTJxhJk/Rxem/SvW0aNgAaUgUL1k1CGdsYzg7TV
9zzFHQaMKjyF3OA5QEvjm3s1Fi1CMSqS6a3h2yRIUoTB/QRiT0/wwmWyBbY7HZpGrhuNdk+Fkn1i
il3v/axvEwSDV6Fc5zCs0bn5XtDEuLadIRoF/90sHWdpLRkcYE9xQUdH18EYTHnWz4rDzqaTiO8E
T/qjB79hnikZ+uE6+I3zcJHhZS2Ze1SDpTTtgfqXoF4eiZV5lWW51HPt0ltsOqxxO+OvnVzwlPAF
EJOl9Nm/EKSKm9CIkASod+0k91Orga1crm4Kz3cE8MQgViO5tFaAcq1tle4hJTcwhqGHFP8neXTo
6BqPo/5mDFLcrXPxbdmhHy4nP8N1eshO9NHUqLURF8fw//c762hyttD4fcxMJ6cWIOxV89NVNIam
z2/fqNEyBjmnEyx1/Tn3xvW1uE3p9fS5GbUnJEpbZTeepGuhw8stCvg2v5Ah0Q3CI3zy3liPPGVT
owWvFJy1dNwqte4hdzUpOpOKYmv/cNAWybT/pWIuPYe3opqj6Caul/IcwyEwtbN9GNXb2z3XFlIa
qYKflDQ5Flkiw7ZlsbDl0UVtmvQfE7bm9UjpBdQdzmS+05dAdowRWOMi3fvmX1YBqRjGo+OSEuZx
ca5Iuf2ONNxcjLvL6RUL3o2B2cHYVVLupijQJXoBXq89+37cZcJ2/jLAv/28uk9fvfIw4f2pVJjw
EGQJPkmcBQX81jEnH/IXinb0PvLerRG7yhsZr+3NjoSqiwi/yLwua4kts+n0YsMvDWGE63dIGDI6
gIIsEAI40P7tj02HkRo2W5v3GOguvkhbT/GNfLW7J+nw6jy7DtF3yamxzJWwtL9F6c0vwM3t1750
YhrFNkdMdL0xXBnkcm6dQuHulQHldoMYgZRiT2NJMHGIEks08Js2yrl7vPyaaw2O7aZyxX891TAI
HsLohFl/moIaqVIV0Yg7dOdaGH/d5f3N+UQ0MNyU6dubzxGCfVvxEpsn2n/CpSm/s5sStcaMQBgq
1HFCtFqwm0FaBwY1obHf9FkyWqroKewDqQspIN0Chz7WeYRiewBoMNUWpgcL4u/NWOGRovxAphB/
VtD5IqUTeMsigs9S2XB5yUyPZ7m/ShoW8ERa3Lz+GESg2CDbeFKOfFl5D9xZl2v3kBmkFmfIuTVO
COZ3TWs6/LTspAPRz+QuZk86u6m6xp3+knT5wyYWF2OHVJuqvPwAbJ6W/PEvgEyKZK0D2Sj/Qev6
2BCouAxhxgtG4NOZe9/6w6yC6x2CMv70KPyLsAoD/v0nD7WrsaPRAGz5vfRU85Scv2LzptW35skR
pUK432O3irdSBjZ0g8L/9yVSRfwXnv/b5/M56ZhUi0WtHortzsqFqcBtasVmcZzE8Mdo8HZ5TjAB
EIzRD+PvCcp4lX/r5l3vRj1gLW52AcuCd3K3sgBo3WLISlSf2VEuMFdqNy7I6wCcJGpww877qBgh
s5N+fF/nR2BYdtzDF112g1xOMlRk1WY+2yUXBisqISZA3UTRk4KJRUjr/KkV0la+d1DkPAcAJJph
n1lqn3DDrt5uETw5Q1NrqeOxl9Nys+kvz/bt+BnH5GtSkIa/ylbumtM1z1vt0LOhHdJ6eej30dlV
+cBPB1VlY/QqoeHQxT8fUMUX5sbT1tRrYJzy/Zwcan1/GQXHrUmB7SqAn1iJQggfvA1dVMT6jJBO
w1w5lJM/YtpT4PuDyl0Kiy9dNM249D6SM417FF7/Dnf1xWUNVJkc2NY/bkepcLNzy3nHNGnAudv6
ENUNbNJPyGXg933La8Q7GUt/zcwzCmmlOc4BzHw7sYGmyIzUjBDdEQVK1ytZSdNt2sNoDQRKDd6j
Kv0ztgKx0VPVIRTtAQ54e/yYZaJzRnDR3/vtZxxnmy0gs2Dc06suoVPDv4c9FmrQwppbz1s7mNrw
OEjx6dCnVt3aHu78i9HcvXnkM7HrVJuzywQlDNXrDRM1DuRLMqRDKBFzMNFsQpx4kVDcn/4gQp+8
ZgDL6bSk0Wel4oaJK5dEOqkeO/U4R9xZtwTn3ZdlaU4kmf+9Bb1SpSBP1DIeaaANn7aKcIWhpIDm
SgLNqWrvVhlpOvkO71Y39dQ1IOXWF4Cd9DVwySHfEBzH1u1D+DhDdVfZr3ckZkefGdjBnlVk69j/
A+waYqN6eh9z0rGBOW+fSQE4U+brbJDNHHrkj2XboW8kJYhcMryknTMbHsTAAk91HtTqbDDs6JUO
YxlmRnsDEn7tszSfDB7g2PB+4Vg5UxuVnKlTB7k6L8igxAmnWpO02bRGInS+pHXB20y69Qd7/Y32
3NXzzQuod/D8OkpWYdwFGpQRv5DMGFLA7It9IBpyXTzi3MOqSnQYGJSJl7+mtBiuNw9Zb/e2Eejl
B7ObR7e6HatzsQiN5fWU6/sj6VVQzyWhIYPrQvsDOVG7j/cTMOMu4/aUKGjjt1j1ZobUAgMs6/Pj
ICo1kI9UvtJN2/tZ7QPZqDTL3rE5bMwE0hOUmnHvxPQF9kQEUkDXhMdj/AXvRKeYh9CWtFrahtr6
bSkQCoZtCAcko9aoiH+lxKS0l52yLj16sSB1ph+hCrRvN2juEZsCnKoe6aUBwufqr3po9Pf04l9e
G8COG/gznP422CrEm2Q5U6zTH5jvRZPkPyhsEK5ikUjYgTrJ6iesnPpSM2Rk2F0+F3TaQv2tB7qW
3P2iKKgMw6iXc9niYG1MPJlKquIRmH9MlCwAzeJEPL7RBQGUXI82kiTitozZi0rmKSNgvVvXBAvh
TQADHNJ6jb+EpQOW8BRb/CddzNLbOD4mqcUC+0gB6jBNvxz3V7607a8tTfrLmT9Ft3aI1o/OR+kl
2YyKkDBSmTeXy2Q0yFoTXuJQwn+Cre1uUG+XNETjHafKy7+xDfjPkBT3dRPhaa2xW2lYirIudPw/
Rubk6DdSA4iYas8kWgvMuQI9qP4gByVm70MtzIuG7Ec8fmSGMeD+yDAuIeLnY6ocCGaAhl0LOoP9
PkN+F5RDOBiDzFzBlho2O2950PDXJ5Vv5W6Tdj9k1HN2Po256WX5tMh3BpY1w2saXXUd0W1K+yXK
I/gr7f7Ukw0VRe2qzNEbSK2CUUuGjy+iavfgrrwJ6AWc00DPNspPJJg0JEYy9gijqUcSI03waXF1
0zw9CKTCqsPEqlwPLHJVbTFwdjwrhGNyPvX32CyUS99FJbFcYQ61/j4t2OFXEzYg6cplMkMB9zn1
haHpO6Yb2VPoNbeC6k/OVvKzEyV+SjIhkSibt1d5oT+r3Ab6MgJq4BIUpYY2ql7c6UMwp9ZAouyJ
pgL2dytKuP6PPYIDoiXXW5D6l1QTxzn29GWTF1xVfzyZRgPNLNMTNOEzhctCEc2PtFN3tVYVBunC
oKwCjIyH1TcmsXkQmlk2YLsglCeM+Zlp7VFnZSXnQ8jrYrnwY7jijumL+QCXjDpQGIiAJvhzOIRN
kMagsNjrDAetoCkwQRLNeK3hulENv0TF9efLWDYkUVqIopRDJaaA3ak3RvsITNy93T4ZwfEWgJ3+
O4WilxJ29DAkN81uBGVsMqw86WYbDSdOf9EROzr5/88Zhu7iDYvf6XRTYLki7yl1VZOiHvL23Q8u
bkasLXm+86zoetn9mnLSGi/XPFmaYXnNKLxv0cujx6i9ijC6HfZS9IBqsIsdtZbbvivZ+6Ooza2m
hn4zW+Uy1oOx1HsNgpT5BkKzwMGixrYLNDEleVvccQMKOi/LevZK0tjHb5qVqWAUrKx9PnQYrHg/
AJCXY3U6ySEPv4mI/SNU3o4yWJW5e80I0z+H0D+iHr5XX8wNcwybvmhbZWKIS6VFEx87G4as+AiK
NFjNmSGuB+GdCeKuoI5klxjT3ODHy0naUKtyTuF12eZ94OjpR0V5NR69M7xciwLrqAI1SgShj55N
47LTPqR+q+xTef/2ftHkbZWhfWuz32/lxgENEr1LsC1u6QI5SpfUcOfciJE1wBvOSs4QofLk1yRu
HEtOdG+l07XEu2reARYovzd+HlQkFN5wlGKPNozknPQqCWO5hquWZ0zEu/Uz0ao3+Jhig2Xy/+hJ
n119Suwp4q5DG9tILA25FwEFbnI3D4nl6lxtx6ioD+1lMLg+Xe/aUuh+eWbMGMFJ33+MuVat5YEm
b/gENYYVX6QT7WKHksHYmWu0GaERILTy2JYhnEZO7GsEwXP2KWDJlCn+ESA0ubFoGOEqrkM1bdwJ
M8h8hKR2mDrCSFxTfCQ+GhMGNPQjfRV5JSssf5pANQnJHD/kV2TMmcLC7gTaxefIR3SNmSp9+lQ2
2gXndFCGH8n0oS13P3EBxFcrIndMysNFwMJxSkV1TOp56vnrenQ+efU/wOVejcm9GlBVrZR6EPUf
CSS3zlkZQAHTuwiZG3praZ5JaicNYAN3Na0CwDIjyVvbV3AsErnVtOJTIaYeO9ZRLe3p626zqoxc
JAZJeYyW1F9DYkuvN6IW3UhzeJFJcpXvod3MiIy6K9r2Fb2hx2wikYgmvixQTsbdu1iFMDbkC0eR
ai8dUx/zTKz/dCbn1KQ+KHv0XdZyG362HZ3gIX6Hgg62A2A30001ZbHKZF3SIcUA2X1ESvd1PU4Y
Axz1BcKVoTSm4yqsgNH4a+pyrm1hIbYa4vfKgYwC3I2dYDOWh70/2NuIcZJHGCcs78ibmF/fiq3x
3RPGRCrsspVi2ynA9s8idrdcwGy8LmTmkG1dp3KoEwLHGS4Jiy+gS/XjM92gpFUXXfjdGj/vR90P
i49rCsPuSWd0UXyWNLXYEKVXA7nUu420W/eC05NjKV3EJdfxHV0FddkUtdRq7io8NZwvMHP0GwFc
tRn7xus3lP6t/bi/jrRmSqW4T98AWsbBWuP549texvoCRuvqlr5Rtlz7J3hw/ctYtok8+p9Vv2Ay
4dR9djYSV6BlzOnO9aQF0C4zXj+6u53WSsf6BV5y7Pqu8rGEE3cqLbsqPJMEs2mXIbTxUv9bU0F5
GHchYtOUEuEPNIox0d5LW+G1o1axzzNs2ZpadcVkpB9fTpIC4BmQFkTgD/jhT03K3I6ozdBFOLPR
+wQSiAYz/+4Xkvc8jsGfRsKYSONSrTaNdouXFGhHqwr+QKBTHiS/7VJ1mPWXfSSc4qEHK+NrCnKa
RflDhfSFwcj4ID5pf7TZREi6JpdpSbmBhT1SpA+qq05FC0c4lq5vj0nPnGmVms47h8NFoT9l4j9u
OtCYKDG6Y25x5UO3w6vOc6GR+4CHNazpYGYwOxbnnarTEKWO+CDcuSMwDAkwAu/lRaKqd3ousf65
eAyyjGVcphhPtxErCh3oSfUgGV4Xgdmg71pLkc32eNK4fYnyafevpGLZt8WAaCh0jM/vG529945j
4nb8VWpFCs3fqYiBq2XzmNOvavmnTMGTayU09WDWFtbgwWWkpsZxyChy6/7V1pEqvMqO54+T9kvU
JiutSH0hKb9QKE+/AFazHDaEfZEGmWVJsI4umUoCGGcnMPmNn4CV3pUSUE9px7FVY3NJtwKZaViW
KevMZQtFK3aMk4sY06yB5At7VoWUUDAbeeI5tgg0zLYw69uWw9+MOCQC+mDccbyB3i9ZS97dckdy
k8sNbd1UNSPimm6fjAsr0IC1P57i3i9D1gxZ25gY9cJJVEtQvYWEmE5KM8TrWSIHHqmR3ZaaBNrW
aExxUopc8oeQbSjCqwlbY6et6a3fI4s5Mof32xbX7+x5DDf7xoO/HE8eQeatWnHM37C2oE8Sj85L
hOh45vWEPWomIMeanMrRoLbI+5MN2Q6GJNXAJLKRSl0W7Ho7MX+f8Ia8y9eXdIDOzM36NC8ebupq
h5RP0L1Ik0/ncJhfVVl2pt857ctokApVKGt15RQT9vG+iJOpXC6iS4WvRClUTFUi2b0mq75aiNnQ
7GHyb2mRPE/lwiiqNkrzgbTJY8J0n7wMwuu7P0DFNLWaZ7lMFEtzh9AZ29DR1buc/cIC7BD/05Ro
s44zHz9DJRAbP0BwKQEu8mNjr69NAx7oWP3zDrbczlMzI6iL5ZHsdeACv5FINKgQpEAnGOwRm4lI
WWQDL61rvMSKjTcaAUMO9fbEqqaDL9NMXHJO5C3kI//eFEf9T+ezrJa+mGcAIOdTL1RPUIR6cXMi
3hDpbK4g0KFRtPh1ULys9C4Usp5kmVTxd94/ktDNqSm3ziYCq4Elz1N4ZBBRqV0JhzL/Ou/n5BI/
y2hCd6fjezHtR1VZPRa1xIK7+NsINxPEVDvGvruumiMSIy0tulPhmqr+g+jHVdvbpeNydfoPWljd
PoW7di+nIF8lzPs4oOGPCXgfiRlhiP4HcnPJ+/xTtAVr9Xu6mnoll+fSsL2x/G+HVRe0dKcKKWnG
Lv4NwLHeRzigWFau+qd7cIZKa8t6fxjLExqCafU1vf0NxJd0YRiFFQc36RrOuMyp5ippuIKAzzo/
T2ORtNiIEkIlT/YQtK5rTRm5v9DVxNd5VT7crmEBuktABfOGa5mPQPwGMmFhAZ8IaeA+sSRzhTPa
okKsfCgpUatzsmLP4Gj8YJVBnrtCsCKkqP1RZ5nCydmyRM2Fg0Gq70cRc0TLLGD95OfvGbXo21C1
WqwqlNE8X++yNXUWIGaiXYsqW8n7FajGaqEpzxZahGEwDt2deDFar3nZ4rcYnTbLvS5W2knaJSgx
8JWhCFwBQWd5ySFyZcwdj5W4CgNg7in8ecUZPsmPMTWOASGkWFhOjcxWaOWN2b1tgqJ+p5Tw1/t2
oW5kIIuyUjsx9oGjgzJYlHD7yM9TVwGOrd5MC/CIsvP0Z6p4JYMG4MniTppNyoiuAKIIwsPBC5OE
fqN3cJ4b5v1OtccuPx+LwJLqiiOHj57pWxHF9W9cpOEI7a9SzQD9qKLO9ui6Bxf3By1kLHQFV/R3
b6n5199hw4qtQyC5R4l1eDDMtztzGhpvvhJL+TPZJBpbtFtaOGx9Zy6192BJoAb9DBYrIMJpDVju
ewba/6LvAp/NrDZk1zpNQzx+vki9UIFY7qA7QrEkLy15k/hgukWPMV+jYDbBlRhWHK/XaWc0ZwUa
N0h/Iceduy06OtJHl73gn8jcthN6x7xLzAINW2J6RwDUIEkvcs17M9sYvUaOG9BlMEQ0udz4+1fP
S+6RcQ0qdIDGZGRkp2TU2ki0Tcuu4Bptz+RcXiQSaxMmigTCPqeTgA4HYAYHk3mOgDV5vMHAlWFX
siedveYrIbhmBFQggkkUh4n4pmvVM2dQB0wgyv+Ap26up1AKjde47rYWGh5jChmtbM65ZMaphI2h
sqsa5EkSMYieqejinfG+F0PlCvktK3sZxtVZje8/nIYarucvt7c8PkBCPMofzOrS7lH1EzIDxPZz
mUriBq/IPAW/LAFwG+25yP9vo/gkfGETnjd6ScJUmwdqDtQRgo7tRnM6vEvY0KxuWudAhLyVqUDe
QwJ9HKAGzAhm/MDoo2j4Mn+KNi6wBSC5Wbf7yEHHXYzCVZb5G60b5qhqi6nA4oFWrG3T8Kk4IDUc
jNYZoYoGcjRVT+g0m4CPV/mNA9HVQlBi5BLUnlenu3EucMmVTeZdZIP3Gh13vQy3ExK4W9c1RebX
Lr98cWn8omlWslDABGKQUhVz2lm/yoytbGr2wqjCzmksBHn5mqXb1YbpfstLhw8lEJvIhuGkCBZ3
0hs/Y778aC/WbuREGag54EqFwuVhM1w+a4qzDvo2SIZKAQ6YeTuflQVO1gpn2bpaj4tLAR0Y1qaR
+2fHj1wbXyCw4A4PIa1WpsxLtDCNw1rXvNegpPsZ3iQM5xujQUkd8CF6fmSNErwvZEdhjjE/9Ssq
bqJzA+VOmtBdoFZvGhkCXjF2j/4F2q8Lghr4HZPAGncIL2tMWhgytx4mc7chAHp3Y/LYIJQNYbCa
DVw9dgWlt7lhV5S+AlQgqmkUZkf+Up4l/jf/q46JAcK/YAuuugfzT31GiQpMvuhM1q33fJiKu1Da
Rt6F1ghwf4OJyS3hIxrHyGMrZcmTh9JgQKmANjizGLrdKT1W0Bs7UTEshbGFeNxPQD3Omd29KpNF
LCyQOirqdCa4ggLyWBvDR72RN/L8pTSB5RuGR1mTTyhb47QRgXzoHA4093XHtOC3ODQssVByOIpZ
tf4uxmKnezCmO0kMzT0Xz6OdYeIulNxdc4hJpsmM3B3/8VM2nIcMGYIgJxReZyqWom+BqvXfXfjt
ESE6wQem7lxHKgqTg1otSN7iYGAPn5DSxpA+KoI0O3Fb6TNX8iXCgTsn5P9nlkU7T3Y2bJ+REMOO
/XxNp1YkXDvrnsndRbf3rW9mGyVX/1yQCsqkHqJY/6T4v/JgMxyBU1tLIuzm9BKdBCTvzVvUacXk
W0Nme1tMq9c3vJ1MWm7LfEX0vzJcDRw27u3EXutWS4yEUH5C/ZtClSSgbj2sj8G++rLZm3SZegPV
5N1/oae1AShG0lYNT2PPp2Q67lPX05e/TdpgcjNE3XBQY+8IpDzSmnpskQ42cZ9vE7GpANGms9j7
LS9xrypgOitechSaS8CnEL6w6cnw5g2aBdDxL6yZJtGuS4xrQSdMWQWO2RsvbWTIzHljmTjoXc5l
8O5aYh6SNkjXeDzq3WI7Xvy31+MuwlyxNC2WXUofPOs85fEEAAUW8oIB/LBlnvgpX5Bd0hVuLDyM
BRdjyrBbwV4I0S5Dh+4P0hxPqLJPbtQPm2b249c77NiUhvIaEGULyNAyhbEZOr9BQgvUDYFRigEo
1ZLPAEfg2DMwbgpsxP9heYARA5T36ivrWzBJhER4XPxybPQ6r/y1ejfu7PErKZ62pK0bOEl4d6px
4D1hAXrezHMKpRIiANMHfhWitdlkTlw6ruEZu9wpgl9jQYe1cw4iKu8yLrhxTPx4g7BHrP1w22P2
GBHXZh0qKUDmftv/Jn8FlIIA+knbxRQOJIgxMfeH++7kgT6OqGcIsKcPnI8YTYbFxWqFliA+oMZ+
VJicWc7Q/GOIfLwnjOT3hUnvaMTuE2zMGWbq1nxgTOijZXZAKi54DfVXHSwa8K7RTEy4yLwFOnfD
3nY+rb5sBIGu49Nv3ZXLkWQnkg7AC7ngV0cTfZ74eC9nBqDvAk58MRZoC1LPE9vbTQhsG6z/2Eaa
mX0TGicka1WLcKdUckYmzENQAgjr+ae1xIKfnNPDKJouxy675lWGiTEsKQ9gGfE6zvJCYSwxsdWw
8Q3HjYdpWmis9yvkt/k5sWs7cNY0hfkQarW3l+AqcfLR2YbwSm4qySEssAoVlK63YlKnXfjIryYl
lF40bo7DstaWIJW/FxRavTa0ltetBVmtFJk2UtXK0DzLSqBKDRkYsyeDh/mwI7Us93Z6i2ju8+c0
LC7ZPRHP/fhlTn5zcteiO3PFAZDYO8LFZ+2b03DePXwnWIetULkgP1MsK1BCfngW+38dthDF6nOB
CR9FDJTGmd6VUAK4L+qQgfr/kvd3DxpZzDPafNxwVA8jeGypyDIESOY2Xs4QtDXknwQ4tkt1cxlI
TGYlR1CZhPpvX5NS4SCufyJ+xWa5qeSYgAbJaClLKf5twtRdcLI8GSBZTJdkxUJx/ry3NSTbbPoZ
m0heLgAkJZZiiigCGEmS4UQdEivOfikYOqJb97vaRHDa+XAFWRIPhh5REoMtyYiSPRQ5LhOFH13V
NZhRgq1I4U+PaYHlex11awlASFNXAecXH7IK+Q3XslAfma2kijKo5zDS7DQvAw0N+u5HbMxk7N7y
bJkigLBjdDTyeDlq7Y+4BvZ+kl0VvZ7JqCygn2+gK/TGXx+E0W61I586eh5SyivNTKSeTNlBqrcR
AUeKIa9WTBw1MtOeiMsoE6UbltJB+D2CsK7UPdHxgnSXC2Zu9VZ7503O6GhtuItD9wAMEULAW7Wb
DVUJ+AL2wylX4WtJ0SdknCMGlgLnmqZEKOVn/K4mv9cNOwhpGL9ry+GsDJoT3K0L5meZ/tGpZnek
QroeXYCOEYJOKAAxm3ybMoAvUQnKk0KzqF09GwRAMtZsHK+aiXUVKQaiCrsL96xBpd4XtSepWSxS
boHZGGSKom/AD+aW+fRjZj1DO+lk2b75kbF2gDLYRQZITpmppe3Z/SPUlIUW2NdTwuXWXRC839XO
89Q6GeOjpPKxtPEv7jy66emRHKjvM6ZkG+yqzcmkTH4Fb3o2Y0glP2a9EgNssp/B4kZN3MgVH1I9
FAc2uUdssNpI1um26ISTFLOmvPnymvsWCkYLkQdbqS52FQu9ZRafOt6YMLNGIefyIxPnww6Db4IO
CY/i9PGJQfTlE1SW3YCZ2AIl0DeOMx+mvY65acNcKgxwbqkJDfqJPDoDQDWIuutgP6gsnxXvJdPd
GSp+7mTnHlZqpnd7rDQ1DCy+A4ogGpYWEsENa2CzQRhfSNKPSXfJDiROpJnN4GYoS+IYTFVR37Ft
H7UWrho3P3Fp/xG99eO/9KEWpIKgC7QWWWFrjMv08DrfTtE6/g2IHanM7Apn6ouNUPzd635iZ4qW
BP+Uca2qqL3+Q1pzHWdu7Z9O12P1FskyKV7gO+IpQBwTC5IPnVwXYe3GSYtBnVmwoSospcAyqeYn
u3LD4KDzPzMH8unQxgMtKdtocAKAp/ZRUybPtM7JMh1dIyF0qsoCV1XRq6rFeAxTy0ox6EiwBduS
/BltsszLkP0b2sPP4uEgvws1tjaPsw14AgNSeJixyBrBr1PHSNMlRnoj5ExMbPDWT1ueNpKZQLHj
8lGNlVFk/bn2RdNm9GTroJCr+ablgdXKEDmItBQQ/7ChIhBD70hFthclWzxL7rG96ItA6ybOU/yf
bYBQGk4rVDBJpf+6uQu566EIlj/P0IApUrBoQRt5aiq70T40juWfvIEkMWerE2YlamT65vZXj2Oa
Ok5SlpeuPdmgf+EH8WqCj9HPOXKACwNY1LN6c7BpNbZ12Ru4FQ4DoYmQh/l4kX2BP6yysEvix5nT
TpRyOkUsV+oiAGXVKXXWCKfUBlrsn1kL7iO2mm8UmWjPASVjT8zCgrAxXX2/4aSPqvM4bRiBnyfg
wT98VTH99ESvIXA7/vVKLd6KvHfi04urjygFpgLrIRE7PilBKQmuqiaKf4zn46na5RLsEURssObZ
XqIcWFfY6dCFKnjmkVNT1/ylaj61AI8VU0j+uk1t7INA8bWqPSCZkKprNiX88Bgwsa5oeCCkMlh/
51bkO/6pX8gaxaeI6QA0wzXLSKBv84WcM/ulWfqW5shYtYv6ZChQHTdPvu4nWEut71E77pmTnv/7
ORHbkK348L93pHn7GAIdpFQgqFzLLDs0kO4Y6IUz1rMVXGw6FHEg2Rw1LnI49CCbBmA/1HLch8P+
HKjBqLi5W9jiNqH4A9OFK8MqdGzUbS7Mt4x24oW2AnMupmbjpkRE/XfoIapGKZlNDCsYeTb2fT/B
EjshJ2DayAiquQB6GnENF15FixZ4HeIysr5ZB+H/1Nyq8RZXqA44yaGvKE7FNxWdsm0IHdsBr/lZ
wOfjRCt5uHMCQKdYgMAnjAPzWpOsDvnKuffDMn3Q+Kfuyv4zhUE3m06MgtgFe10Iu/OszkRdA/8e
u6a8fUCU2tmpntXroamSZYbEwKqNuSaeFIdMPSf4EUONctRJD7zBABV5le/J7P2Ai2woqfShd8hk
XxyXN5RU91Ndaf9dIF2WitK4Ag+ex4crCIvWAYHw8SFVQLvvJ3GjpGO1O7y/JRhD4NMHah5HTHWe
uBkzJ04Yik1BTds5w1fcvt9M5jbrJ1dj2MvzaYwV3IEjeZEJEWZQ4DkBesI2RbyOp3zE78vaN5Nq
Mz/ugff58M7Iig/NGeqSFYWdhA2U4TSFeyFp15JJ5/+mO+Pk/7OixR38rCkUDF1BVKc1IIA53Bch
8V57LHR2J4uszXKpKVYkDsenynTGtg6ZFN1znhSm53nfJNWHLxn9HPqQ8IzZxq6/QsntgqwHCyfA
nNIZjkbEdIaWu32QaWk443FAwuYNnrsX29nOoq6DVTeqiSh5abPJL721aPysvPWWiqarMwaky+YX
a9mxnrJRlEz0m8bDqbiKSpat8ciLUDtOlb/5HKdY2QvNWU2YYOG++8ujcRegvXlyxBhj2fBgfpN7
0ay/sC/x6aocHYoDmbqBqTc1vrfvRL2tPFLt3iMQY06m0GIhBr9G7ZLtFAMcll9S9eSkv8IKgdBf
cQNPYrFB7w+ZtAiwqogPulrHEt5kwEwags8GyqYHt4GpiELNaSbwxpH82X7XsNMCRB8gyGbutyvO
++JROG/EUCmKx0N3dqoLKHLhIu8eEmH7WMCFB6LO25vqind3PW/Cj0p8VWmwSD+yftVLVqEhCPL8
28u6Q+vGk5i9oa/YHfLLhJRue2XNITqwE58rwaDMr6ghuLYTqj4e53y2bl6Qk2w0FpQzu+49FmTi
dzvijf0E5Ybozh/lmfVh2wdksTb1Nucqv3VexApNn66mDM9aNmrjp2UT3D6cSC7jNJI3Y/TXCjV/
nOIrI25gqD2+XJVQG/rIKbdinHpWBe/w4IMBwwcrTBEhLN6MXxU31GQFHtmz47Qamh4ZRq3HHZTg
vgteilUgVUUhnoGt8XhwNCIDHgkckKJTayJF1d3mRDahoTgf5//Tn0dInyZkVpnk8CGxYc582giw
O+7t2RNCBMKSG0HlagAFWkUNekcsu9AWPJ9xN/7F2GfTWz2WzEzemw6iq3uUNosIQOErce7sikCY
u8OZtbQKfTjbp0i5/Ib/w0WHwuK3n52SmHUVHiNgEjRZjPLSABOyMk23XH4+LrrKETSYYNnP9grp
biJJpAn4+bSdl/s9DdwGnKnbXVM9X3xiXG+gTLzYJuC0YEOTJV6mOQc2UPBvlK8jgr49/3PMec4b
N796PO2yv0p1KRS7B7L4J1SWu8/yzVkFDqk6o2MbzCKIjD72GueDOwz+Y5yXIQz/81noG0/xendD
RymY1uV/xFBJpTJhMM0t/MqZ6WwvfJdpy8PHFGZY3sknMTv+d6mdSgDHpcxe0vh/KVDCBEuL6c0Z
RQp8vZEHLYdU53wIb+RKHUpWj+WCTU+Z9g7+LFIUb3lI26WLHVeFf0m5CfJdcNy7R03LWs2P9sGE
z7QRIzsOydqVqBaP9ZcRvvUQlloMPYG16us1/hn/U3SkzrL2jqVCnEPjPH05mvXDvQT3wLSATgWL
yyImVloAw0PxsrvAalyUCXP+LbbYsv+ep0ZaopWQkln35M9RvHo8qyPe+nHo1gZQ4SvduC6lduiW
zW2Mq5GUOoD36xKkI5IeOaO+XRLm6CYChTyvTfLP/gB/NvIhRXiJl8584joIYXwErsDRxNcjZ9sR
XEKKLXSx0t3vY7SWiScjW+LCIzpR0QcLPVaRoZIEohAFXxxp2R6lr/hrgGqRQaUTDHM2o5+OlpKf
TRz/aNWOaqgFAEFYmMHOjlPcwEvTNThHyKNx3hdcn+Z75XaRaOFBAfD5sOoreW+E9G3UiVtNBKD6
1BU1bAe7xg2Cak5hWevvI2cEPYWfnw6NJnPcO78ksOCykkKYoS0HoIe+exDmlhYijpEsT8w4pPMD
jd/pzhuu8qNOpuuFT1v7fb+48i9Nepo8xOq7AlTGnH2VgWmttlebmh3J7LR0AUR3df9AmMNEhKso
Uig59xshGGSBBfaFiEscrUu+WvLq+pPRCAebokvEe8Cs0exJqS0nTN/nBWSp384q2vJf+YYr5txf
anYKSrLvUFHlWRMwnaTl52xYETqdk0FDFRtCiXXDBS1c4vB80pImCZ5YRQkneqL3B9CaDqF2co46
UJaudVspkS5+Gx9ql00tdfTAbNVTLYO2QpO54iCi2Jl9OreaHwnoTkrbOo5dNtdRu/GoS7o4pxIY
7Jy6kP8uP/F7rmh1xcGTQ5G6UQNw52JcwTSmgCj7AkYswWIxE3HNsxX7CqfcNYwzGPHnnD0PT7et
DUVUwcyOvLQK3Sch+j+MVbDaf/aXEYUuD8zojg+ksLPiyekTw9k5N0DEihBsOPtmHvJM5imlOn1U
J4+dotCN1SN80eASuPeaY0/ZS0lwATPVQ7LYow2VT19ygrJ+Gm8qwaxnF0BdLLD7sxzp5KeRGg7F
5swKjNltdUf79zzWbloHzGz+8n83Acwd5EiHrWSxSCEj8tX0ub7KsjbeCPnyMgl27dAF0Z2TKDEO
ZgK8g9seYjBOpaFzIbK/WkWYIoBO0G/47L6+P8lu/BV9r/MpAT7iWMpuUa/LcD52LI7JEa7ED44+
SPbVgH1MKWtrW6sYwjStB085whNm0R8UhMp7ftxKk+UFGo75kMyN432bwoz1Yb0YOmaIk2enFzMF
TtGywVfQdPR3hawxGjh34vN4FCoCjgAYnTWauqo4uQxfc+tzjqXfaEyHeAImPQxwkA6myBzDtX5o
7Aa1x7T7Hx0Stvs0afUFHjCQ5li2yJVd2qhuItTHcy8GfirCbZWM6qtQ5P/nKrVqtKptUNV8Wus3
G/EuBu7yrIZlIXE6r7dQCXZvWvXraTecyzHxvwPVgmB1BibSZEN3O6IF7w08XEcmlwJnGgkwwePA
TrRwSF+3kzQfZbRqotOtfsj9ll+D++4aCnQ7s8ldmwKcoQoATC6DWh73NC2ZbLNLFLNor/+6/K0Y
/bmpEvu4TdWMUhti45f3wF9+AekVHG0nm5ot3lTpb92sqlA+wdYV6yUQDcvd/huk8inhkywT6tpY
vw9afTXnLP/rl6K6llvuMmGYlHQWBQbjbsTJW0gWAUIixNDJcO0QhzE18upfwf5h8gWKb1srb6U1
eiRJDCKdjdV//vS5WhOgdcJqraQsnMF5ODVoTIDc03iDiUC6dW1VCPw6I2yqyP8Wn1mWLPKGRwjk
kA0RxdAKfEe++e6Cl7VVfMPF8pCFBRqdWAL2IrMxS26XNNO4wiz+zbyvZWOIV2JRL5SnAmmHM+cs
PRbuR5nCFE4/eLIyJtoWAHZm3k+bwVDI7qjYxJ4g+09KGdqNWE/8V9JzbXDgpYiSgaJUbJb2Fvx2
x/aDjXS50mkspHS2Z+6uZB1qJumkL2mV2IDYcISf2UZc+3zUp6rB48V5kEAiOrzEy2EGI8M2Hl2u
XQqzxrV1GH+NcV4APP7CmSV8vFH68v185jXFpdpxufzUP0ePYTOP1xltPeOODLytDkhdFM6IZQyy
2Avp/WixhxkLCdEYbvqq2KGxOKIIPrt5IztJJiO+lIP3oF7APWaZRzs280Mu1AISiKAyvDdhaHSx
P+3n5+Eoy4cfDPqNOCMN1Z67hrhVk1mlhtvQ+arudG1NTbqIeA8BxzJBYBmvW3v30ZoLurimp6qR
p2+NHm53Fv7FLGpQcu2ZSDH6J864HwJWAxdxH4UdD7FGIwKmp3oGs7rkQo9UD77nzD+feibv+xS+
/nrhFlYmGk8ZERaCj3gnjXFoye1YH9dHIpgxftBlDU9y88IABRMaCl+AbLWSSTxXfGHQ5HWCY2d7
yyXcIgiW//5f5/x2sWQwA0KhFoxli7zqP4jXguJfAxVzrtWjegHoWDQt8b+c/5URgCmCBlu0Fpq5
oe+Q8GTB2FXX6zxTpG+wuOYUy4n5bUDOM4Od7VrRHTbWGut363EoHNFYF8IzxIwufABE5rLO/dag
YNdzVMaJg/3BxmfqnFnet1PFngaGQaQNBOPpwUWFXwxs9fydFx+T8QFn0ghtiYGIiTcfm6ub54OY
YmNqRBkRxFb8Ma2068YFSEEcw2+8RuDTQbH2paFsZMOtCdRQ2X3xhlScAiZW/zN+ttqeeLds83MC
KN71DbjTxZVgOdy7/Vu0XYkGiY4RPrxPv3iJ0pd+C/68h+twdIojciya213O/GGJy0aOXxlzh1Bz
PjXGyvrxB17nqnPSTAZsjWClXAJTfaG2Rk8k3jO8aHqNeB9ddovm6rdNG45hRvnxlxOtAJk+vAaZ
bAMm4Dkq9Re3c5S2ugo3XdI2izocTz7KGIz/2ndq9R95pFGNews4PT190Pep21mE6iqhOkNbkF4x
ImatrTz4+mPwfpmKA0ZAVM6evlIsMZWgcIVWk5dHY2YlumpodG+0I7pn9PlNF2dKmxkYdnHEljmr
bTAiDsXQVA1mxpQuXnM7Lk/TwK6YgGeVkbbGxLuTQO5rvq9xCReE6hgC3CNBzUn6Mo0e8kVTvXJK
rpv5YxdHhMlBh+fIDGSN6u3/1VJKpvSUKwkWAVhqtk3muuN6fxuBkPOPnLM/4F30hpFRCZFchi03
j6zKWzzL+6Us+FOXt8OanogfJas+x6/t2mZdZ6Lgl1f/nWeG8DG8HvWZYiPjB3PpDquNANJ6/EEC
rxZgPt3SbdPkK6l0tFLQiabqapfZvgM/H9y93I+VfBRz3B71sXKMk2ZSSPg94jmIFQr3b0OHMyU9
AHgCGPujt+EQdlc1qjRBXIZDJvXJzOPz2sD6mBuwMtRA60epQCZSZyN3VGaw3+i+u19GUBt4/LyQ
HSZ7lvsR1oJPoelirjsqSd4yOCMqumZl8yVtzcjQ9457ZRPFB8C3Tp0FS+aef0psZfK8FaVHVjzF
OAq6qcTSdS0Bb2BREtCJNZVrBbDUB0aVgA0h34FCcd5OwMmXyH4JvRnqIRhPdeLf+w+kU2uf4+ym
7mMhocUbrxKgPwasIRvIOlkBU/zsKwiBt765SwIOo43fjwDKKkbzQjntaDrj1WTkTLULCuccmbga
NNm28pQAeUmlChxWh3wxVjYtHxI7vk2OMdXlUFElxlrzQgtFmNAc37lgvbw9P/Z0tgr0gLNEH8Pi
kxlzWT4P/GZhM+j5zkI/AGZSfusi4L1Z76bwAfKFhx3+VuvoNzrYPtslMvfH5+rb0Zm709i7hLNQ
+WcEoVM5PzPZwnKit4oQc8NbFzKRXp9ioI9WWHhtK8cSzEx6x0MnqMfeOBE/YlbNpLQtQ+6I3PUZ
0s/SXv4uiLkITRAV8uPDDH8I2TOBePPfmbYsLXwv3aKY78vNt8PsB29E1XK1cRHwF2gn6WyJX45d
Yqo3SFP1HM9iywHniHDoM2K2ypWcnzYMYUXeek34GMcCvFqoghcNe0UGGaZrDA5iFd/YRRPmVVhi
V3LsjTyw5tLZh47xxgXYYaW45a+KUueQEm8vdylWtFCYsN36DRqGrjVtbM6DKAAsc4V2tyHaJ+Db
gbSXvVp7KMqv1PWtDdWzoD80g0nf8romiajAOtP7b20oCDk7/2phad9lxM4Zb5lxoM27exY3UKVh
6IDUl7ckTYIk8annUWL/IpCkJdoSRcuCh7xnU37bm9eLjQmo2MwU8nL1TFTRG50vkmRFx0AjQwwW
ToQV04UFjngjsUu9DJOYyeljlGKcfl5WygLH+WNAFFKFH8UNJiSRb9n5l9Sfs7INPVQiTRvCzZBg
udIfiEeaLJ06LQ7Y0C4Xdc4ks1S6SZPHHCTAz1PyAIuhWwPAC6DLuBXJG2Z5P3IgjQ7C0lAIOjXN
Ve0DAkkiM3gJFvqP6UAvS4F7baUgWXtRgxkBQo6dzMkVmGZfcQS0wsrypTGMeJrzxZqrEiZEQJtf
/GLSnXYMOlSX5CAKd1QdAi9sOyKOm9ZV0RvJOgqZglMemx+VDnaEtgAkibSSLphlaSveQd9Ul+TL
3+DtLKnbTCgD9Q4ooFX1x9ftyYuv1xKLzRTqMkT3u2KDqhMHKIP9oqoOf/LyOnB6aZv6G1hoKVm9
yyLyBhdGFXPm9WjEeCuLTbeKLyye3bQxC2IJ4bIMAmHOwRfTuDWnyYSPNZaXnFDmphfCCyKI1JPH
mT/Ci00mqGRiE2av+K+riEcgtMMxwP+d6gMQOK0efHIWFuaStO3yRnus79dle8BT3YVkPZJ6brXT
uXcbnLLnvBlEwb2qxybA84Ag22KFH+gr2WNoDJvoVrrrkZTrTFtwtWoVPYH5xwRNF7sZdpRF7fpU
w1QZI2l3F0wCKNioJ9ue4LHbSqW5EkZxGVvrV7hOk3407shBzggIwBFwzY2ChWfTPHCcA2zADA9D
34ri1oahvze5Awwz2/GB55yaL+FiVYjvLv8iypVrD31q7PLke68rKRiXe6dps4kuyVsOuYHDNITV
/Jc+/UDf/XqBG6vpMFm5ZAvsTMbo2LoNkN4JjQTbkrPXsyi4F8sLvOxbVmzXWuwFgvmhHFvCQDX8
dDI6mIV87QQbtoqzAHCO4CRcguSxp408+QmBiuKxK9TLNsl+mHFnaaec9xURwgZ6RnIvcTXuyCTs
fkv9QBt57Uc0YZ4slgcwyM26GcLbJtJHD5NjRNRIF/KUGlejgto5jWw1PqgYkXxGbiTDValmLVFH
ZCQDT7kYTtx8ARoKtBB605RSov6a/ipg/ruiJlascoGox9eDKJZJQF1cgasH9NtN4gKfE9A/AkMt
0juHQyxN4hz1sY5wRupPG7oOyhNNimEmUWidETNlUJTbTbbHDicFbC7fq7d+1Hen0VVcnT0avTHb
0AyNZ9Uja1pmQPdj2bNWTYAEsY6WSR+PcvVLqOfhtoaDKU5FAQNLOMHSypKNd4l1Z5zZsxQdjMV2
tjaZotb3dRpdLI9AgUMXm9BlPCO/nGn7JCtn8iu738svPgT2z2x+O2DDnh1+pyxH82LiD2qwTD2M
0HLq4YpWbWZeg/40XEEg7tIa98r4mdaj8OOevVCslDDHvMkwQFPe6yLPBQjhs8diPKPsJpIHywOe
utzRTgTFWIx/h2dcqXoAxFr1FXpJQSWaZqZj6o18fj0+mJQeliIO7DGepPTiLpIjVcQ257ma35+3
1pFa0m0OZxF+w9kbCIaIpTjk6tvfgxURK+ixoQZJrYz0oo6V5deHVBadhOcY/EwIh5XKKu94Huf8
fSKCj5zFgDQO9nGhxZYEq1uu3tUtaJKsRvPdED3wfBOJitsdANcJe+XHOXoiqHLYePC/cMGEh4lF
dSyCFeIFIxSMlwhBd9cNkylbyN/+4B8I+6mJWuNpaQcBJJIadbLV9PPVgLwjz2bOmlQ1mMPH6rrn
RTBFny0HPUVdyU9yUqB9Fo1xcrOKbPKTfY/UgudoGjZriXe3aBREDjxPdvNrYV+HdiWVqOSVoZa4
XzP3UBIWEqjNuwV9Fn+f4p2FAuRwA1XxVvb4cZpg4t+MwgzAytBpX24M4oBSFUC6ejTFe1OpzDeP
U35J3TTkZpaPuJSRq8OFXmap/U6aeFumPDrGaG9isIjkht7zDIjRc7BTXGySVbltkyPTs0AGkJ3e
pABjNdTTTrkWoeWQ7Df1dzAMmoNM8D0xzCe7qYesdqQfoudeiEQg5igGUXByKfMRN9s8KS9nzavx
GjSu5NZfL+xLCtahzDFYD9FEyrsjT/AJkURNUcXhyOvH4dNQk00D82VoAOhttmfNS8o45LTomzLS
6GErd7cYeiru+/QFhJF3skOA4kJPucx6pzMwhw9Q1gzoxlxFd3M3/CCx2pMHwNP3Nb5Q8n6malML
OVfDRlJZqGCK888mYqqwA7/e44DvtAZGfL9ar9D1vcU2A6JXLTYQIXNZyK5c0tfITnGS9a4lwqD3
TIKVhIopoNXgI7ciNobPOt6R5Q8COxIFgIPC8pg9jkOfjxcAjqxlBBus36m3d9ddATk/F8AeJ5Up
Waxrha1xjlQzUR/bTRxg+FROuLKb4+pTihIp3sWiffOfJmrbRlnNH97m8ZJvdO/vGMpRYvbX6YN1
KIOb/wTQYRSUMIciFRA3vKo6Q9upC4TBI4JMvnarfGTt64daeSseT+Da2x9jEnz2LogUe0n/p+ci
wRbkDSAixfWZiGaFQP3cdOOaGy17ijyO61rfqtBz6fnWpfVt2kiD82Th192WwPzZ+Xs+mOfPmeVB
nr+6+mJOHDcXUt6RISL2LYEQeeFNixCBhUek4jWqbh5o7kPCp73t2+TEFMpAqfDbLXVlNLjAejQ0
Iy32F1WEnoNmLjf3KFJYUaz6D32QqZXP5ZSwh2+bebxshXmBODNNSFZgBzkwFUcprRQDh7qAItNU
AjRaiqDzW37ueY2YtoNbGZf2TEUvjgg7fRHMacFIPuYm4WmFq4ggitQ7Vm0Kyjt4vcS60lMNVPJ/
AKCmOBAWIO0ovNHBbyMHYCPEck4UXiMvuzxfNhke14qj0I5F5g/LrqykiblzOVFvcNjXxGKP9LvD
64NKYvvGxvwBL2yH9cSQJx55Dp7i65JFupjvlyb67tq8xbaGQjfqEjeLbKjbrVgoPmA7103Mx5kp
e85+EKpL8OGr74oA75BgNc/P1js2uDKp/fKw+2qN0B2oAYACn03eTC7LGojlBGsrvEpT7IozFTwF
UBiHHbBmUfTWvoNb0cu1fUf1hdQXLAUH4cSMyLTBe1EQIbOhu9AA6/b4HwhJeh3M8qZtT7eOiYoR
3Q1fpNc1VcK7+VCkA1ZYxLh5nSgpsoTFIWFLJuMecl0WBAM18jQaiIiVNaXO/8/ORYVTrFJUm5CB
s0B4bIe8V4Lzsv0ouBQo4KV1rCjiszpt5W+ZcXsp3NFs2V0Z4GHgupWNT/8vaFl0LbpxSVwvDsY7
Tumcb47TfPPe7rNcBn0SdguNGVHt77bdTfDTeW0Gg/6l2QgGJK1YsGhevmxkLn9up7hPjAaX2huj
ISufFFvrXw/1Ufh2Ue3JMVFRWyzXdHvPatVVSasg/9M2tUxBOs13jhdvp9hT2F3EJYhYy4QKABST
HWCjY2uy07deO2KQ3cxN16VaOH/jUoXd+Hr84nIcnw2rAxgvHjOD4gPyqJBF86xL/Tw/nJsAD8NY
dYOZqgAG9/YwVXW7kyuhCF/sT5GVDcXDQSMjW5fmrH0OFNhFuevdu+tHzJnzmYvnhT6b4gsIzld0
ezJo1cy6wBoVe3dshCHPGQMk7Y+df+LTqauOt9nMtlYBq3WvrqA4supH56ZtnUqKIjy9xq+2b3GM
4obcRb1UKRO24Rqx2oPYt3cbyFs/TQRhp/t5jvyEMVxf7Q4Gi61CwsRGIjR+dwTbi/qtvJKnp70P
ZCgopwjrXO9F3JfQ7gnartH1YMNvpUoULPHMw0MJJljCf5plGIrucS20joVlkafKfcr82aNH7BG9
PxIDbpYlT5x+kt23lTIY9Me6xoZR1DpLqHu3ewvriIcrftPNFQkrMG7swzjImibLHZlWvO3JHDVA
/J+aJPm7oXKZiwR0Un2PsJcNhe4zoltKq3nJeZTu6jWNLc+Yg34iufsRLJL+QZ6Vy6+kA76b22ZZ
tfAXztyE//BknM8+dbbAh0oIviSjTXQ5erNbqjtyhtK0b94WYvhR9eYkJMZbqw+IwHEk16EIFjbt
vNkeOC3Tsx0myTWt4O2dxEa/JjDZGPgvepEgYftXDb6QMBEbS4RjrxQPm0EgV0jcxqxaXaEyXdZq
/2X61Phv7QG6CUFtoHlugC+YleC/OVtcA/1S4yLGicB445AVbMt2wSml+yMNan4iofRhbu5HLGoC
wzexKKVC0LRzxKpMk/ZuzVHEELuOH0G3Og1ek/9QlLU9vCeAAS1lJzjFi/wu7pEQb4CuTnSdXUsu
dVc8CQl1dZQbXkWCS5tnbSjvuzL7JvTnQGrsSkmUDQBSzA1MhwropDngl4OmI0fJBnk7dONOrO8X
z7YcLMS89LNlbao+97NdWufBEdUaIsZO94ZGgxoVn53V0Gr3L2W5dME7dv/mmXuqf5VEqyIW7y6T
WNJlpqOlYCWR6lg63lnTWvS8Is8yVP/Qus8mtk74TEEkRQkkKcKKm4hWK5lKr1wXuaEGdwTnJtFC
oea1CvvEWBJAJeaMr71nOYbW/YDJToLDaMjuIpSqAlMNnumtItR/kErdXSAkGj0VoacNgkffPz/U
n0N+4nrT229zC1R7qltS6ElRDWNEwWazD6nhwnBk5EPsrBwxvGBhqw1pG98ESlVQZd2PLTOE3K1X
OgV8UjNOa9cPg5/d1+242U4MXNoBr8cudn/GB+ikpbEbITaMvQ/TQ6L3NtcQHbqeeE2QLqV04O8a
f+120o1F+OwvPf8gXdjKhS/wKeLozVlB+cVAfjZrbK2RzyUAGsBe3o9K+Gnbs+Jcio4FQ5he84cR
fqpqIlO+2FSt0j3fJ0LrXB7IP36dDvoEnnOJZblIhwYY0sSk837RCXgmA8Lfm5KcpEaSUxO9gM7S
x3pEAKuo9o8In24owPU/C+MsbhnT/tFYJfAROurzUGOv1T7TkqFhSfK/Bq1+YIsdcnhuHb3m4mhn
WPSF+gk5hEYPOW1bdsYXBYwqW5DXWaw1klC/jAkiq284opBJ55R62DUnoqaQ4J/u9rHo6E5vHQBe
5jFeSWRPd1trLm5RlPBwua2ELenIbOTtsFsU6s8WmGMKj3NNBrXS2KktQCWc8OsGipfrH7aasoRQ
BjTp5LDKrJeLx110Qu1B80ExvRnsgn8asfiA/36hLwyT3Gw9GGSMkm0bmroD6qbqs2hL3a8BYaip
2i9NaKJ4ib6+34WUF8JtK4w4E6K90NoPdb2yAQ09AaupP55bJg/KvsVof4gL8CayOiimupx8UvjH
hbJwsxpbLn9Wih6Rz8Dr0Fa8fDmrG8xN9ki7rxUzbzJOLw+Q5mbzuXbZilPO60kJgQVO6snQJ6LM
4Bxdm8Jd1HijGHw0n5VVTAIiXceUP9GJO93zzUke3iW4kYX9SyYlmzVirAfHU4P6h5sheZuXj/0x
0nrxvMzqzGkjB2ruUYnbPXfETCCM+M50iGGTPCUoI7N+nQa3hVJGT2Vep5TTjQDUHYr6grsUgmd8
a3+xT+MzhokrivQdidNqod0uptT3hQjocWoG57PfSvpfaAdel8ZfoIM82alrehdR+UE8rhb2oi0+
hUON+jK/O+vJ5s72Pe36bDGmJTKwco1i5k4ZwLqbfviQncArQ6YQkXnhvWL1oEgO7Ee3+h3tQ0rP
LuYSVVmetBt8FRv2coRjqJ/o5uxj2s0n7gmr8lwqkwJAzWayhnyerJHRBnekNbdLT4vRKQPy98xg
5fsNhfqDeW9gw+zB3r7Cy6vc2N9JewfHRjWRoPDhpiUcNjZZ/jI08ObUz2WBahg6AYdpO8Xe33bV
Y4zMI9o8KcSmPIFsdijRVar5JicY41QTaz5Ox4idT9bWsPf1cMZ1NBrrAg8STotvXTO3IKWk/Jde
k3JnkLgZkw4l3fZliKYOQdqYtm8nnfINgpN+U1DtJlIMTCPVZvywvDKSBbnkDT15eOJDKViundxx
f0INAfQcK5qoxb7ZdMvWe7MmHFn+cHDoeVZ0Y9Zp6yeMTZrV/RUk4OYbByRDFLjavlshKvsPpYX7
MfUbnuKubDEmb3gHq80YhLNFlTowbe3qgNEnzs/0trjFrHiJbHWe2bAV27h/ZTy4T6UPDEs1fQXK
J2NF7KebwPZAfL6Nng6RJpK9o+uTwk7qiBZlOC/tWpKc15z6FpF8lOWFXfs7/D7XiQERhKD4r46/
+rd3kT9IDeEf+BOZPmsuPKidSJ5V9u76CRlgwFBDHY2yVZPTDnVNYjfFQ5N4Dj338XIi7fMU9uwb
7UXKK2ZxGfZ2qWuuhfw7WOSnZdD7Ti+Ul/KVHp7VHEHWnmEstalFNZDy/uUnxlbFAl3uzd+wlKx9
lB7LPLtCDR8xdalP79UZiQ9ksYDf+JtrX6VOBgWfnmm4HDT0ynMhESSfAJ6qPNcWDamXv3tc5TWl
cWlx0NJOtUFwX9RtEB6no6vN5D7QXzGPOjT1JMkhRTeUjqS1TARN09TVGasW19PcjNFjfjHQ9Zjv
7ZDVE6qe2QxCKm7gcseVinpburrTabybdbKwhi4OItDtMRvRIAWCUl/jTx/gjBVczZNQp5o83jZY
HdrZS9PUen6DIaX38Y0HRkJqA8hHFpiUoYbG3wgmLQZs6sv/lxYvmi574RAGEoVklm050tFKQFWP
Fd0+NjVGl0QVat3iRj31YPTdkBtyYIgJGlOdgTsPdp6LIGeG4KZLLt6xV34cKr1EqKssUliLJ1fP
P4SGoYQh1V4ZF1bL5RsR45xPMOXAu5Iq6/rPWIxrUcNH31mnCWhiccncOwpriFy9XLBhd+oliscY
h/f/OqzOgC65/4v95HSIGc2fFEvgUP6cl0xHhVwtYnLE2c1nTi6UpKFiqno8fKbqL6yCjMSJB6vP
8h4yliH1QmG6oTbeEED5rEAQw8fsmE9oF1nK6va3AqPLT/c4XEeo1wArU+PL6Ap4SvtWY2lhJHht
+JFdIZzkPopTRUHntuOt/oyY8AYsHP8txrcHpasIU/4v3O5HmgEfytdjInoIYZ3K/5ExBcUXIznr
BBJq05itFzdZ7N6uSPtU8kU9TYp22NX+u15QnYlspnuGCUjAW8J1JUZAbSz218Ipj8VdgGQm4sH6
6X5tTFKvsyHcuw+PhaD04RNCE6qk6jcwuoPXi1W3Ep4T3Y95vvkHwE9znqzaYlmaTefQPMkSBDof
gQedBhJYyhvaZKNgexejyuoaG+pVp87GcxZoN5srmq94GjJ2MGhzeWwbbBOu2vhA49KlqrEG1WK/
mHqATTI8IjhaCPkV7NgSYzeA96c+3lbDbsR62MAVOIPcIWvKquWDd2BSNmiUX40e49kzbWzm4Jk1
ISXnQdG4gL0Udid6GjHqgsjvoTJKfKlLowwieWzHQd8ZabpO91CpEUhw7hh52CTkuxbXM3IQfudo
+XbQ6B4Lg8W/K4pyYoba2viKgDE14NvoRARMeQHfzYi4GH/mOPUznNTZ2U4NyQWqGY6OEeAnYBlA
lNNPQsVJy+gHb47GXASuOXQIa3PUc7+UntRjAUMfdt/YUk+S0hXqzhaQlBoFwJ41ao++pvok9J3M
9o9SO87z4JgblMRZned9LYFdZF7cDyC08PkJBELLCXLYQGF9ySNk9BAov0JQmsxrak9oUJpZwFW7
zrzHwC9T/OWEwI6HblpHYQiSSvhjGfNlVXZBZXRVKKqCSXcgUau/tHABu+kDIFrMCS3O8Ym94VLw
vgcHPJA3shhj4wj55lhaSyNUyXK2PgfYEputSnZeDRlSWEbCq6hJG62VPBsWXNr1y1cEDjFI1lKb
DSRc2RfnPiNuT2d0JLcOYpf3Of5ZnEAk2tWh6yxUyQqpTVuAP1ux2rUIEs1TkfUVPQR07lZjr2KM
j/GbcyvumfXjtOuNSX/ZBN+dVyBeIKtyj5No9tckMQjnsgC80vgOPseOGSbBpafi1ZGastpAS4/B
NHBbsU0y+Neq/NgWTqNjnwXE4pazBIvB65K8Mwi0xhlLgrF5rUJmFLWH6G7iO61nga5/6ODsWL9C
Jg997fMKkt41GhfvYv6Px5NXARuOxml3A9KRvEDCeanvuC3c3xKb/UhR18qzubeHkwQyCeYyytzi
MD5rOQnnEGFXaAjYrw0r+BKAa4ACiJJEuwH2pI0rwJOyyJybrkDqjczpBdScRbVu4A+/8kMNI0Qi
hXRVmRRB0Fo629MbPw20PeVpRdmjMaRP/8DRI5+sBOUGzXFmE9iUEpiwr1LPPIN6b7+FC0AwXJnX
a+1/uQdecA1KKun7TiG0yxFfQ9ks7EYBSqlIuvyZJ76Uai+dB+ifplcrkOdHmIz+1nU8DHIHVJn9
2Bo0rGUoH25VgVMwbvdSnsfWAqpsIiZiKDOQJSKQPOqRG3ZdtFGcwA/+jSw7HKXpN5kZIvjoMdeu
dqyzvYgQdUbhBo8GowHS+80QgKD27elIbTSJyddPGRA6ZduoIxwmVXO1R5jnrJsBDHlDD6pxcYkx
umxnstgdgEsH10qK6T7PZwP26S4QLjbFCWf4+zMhDccvexgoGsAaT/XO5AplpU2k17D4jlFHH8BC
RmIbvzXtqGJF4c5oYbph2qrBG8A9mqCXsfcXMXKr08KchKhXlOUsTtC5Nnl69+26KlFGfqEXUBBt
/+WH9TDDWi0sNfzXe85Bc0F4KNywasd5HnEqqCBEGI9H1p3B8XFIQfgQEn+q91eV5WTxdsaVibhR
GZnw24hwvNSyJgQX+Fv7nhhLBt7FaDt7CcPiSki3DI0ifsb+csMdX0PhUcanTfEJjBCkMg+07G2n
/UCq/u/1RDBt6M2twapSPR+nb8hOygFgcxGNSwyke+kOgLIWIDmk7ifSMEfx2mi5kx14C4lsqUMM
WuGL6jgVqMDCewNKNOYe7pWQdQyGvJFM5swZDkMmlTIz3xN4D8Q7pFq6FxB1QVmBKxdhIWMzNRBA
+Cx7cE6STYMWgXXV9NJqAX2PVQDYEBuBC8ZKtmuFRNkLYdlyf9B/SHQ/abmAtfZu1m8rEQHH1XxQ
n6La9ld6bpVQfsSzpMWjotu6ens/jg8FNnyh+aPtRrjtYPM6eqjhQrsij8w0iwPTFmXKzjhfeZlk
sbMq2/g0bc97SBBeaiTLEtHylCM2AhOQceR96ToKH1+BQX/36cdZKu/HnbujztElKT5VgZnP2tka
mYtgkTNBP0pldbGsormscamFCXYw6H2KAYV+8jWi+arOICMYGYeR4qqdjFvDRoQ+H/UmK8AuZ+J/
9Tl0WVDivb+oJR/v8zvkSqN+NqWjVx5fUn1NNxjow5XnXnlZ1ZEXo/vcNKmGzuLQ1rF+Qz6i4lD2
D73AcpCo/w7bk/+FC1PWhgVndTEoH+KMHEQVb5ndSmgysWKppkT+jd+txEWLE0b3bztH2FnIQpkG
G/mE0CoZGXwsX0OviDfp1pKWeswgjK4R/vR5cX93jrA/TmIOmSDbBFMhQ3lM8JyHMapqkMAIPaw1
73mOm/ihT3UIFLX8wXRPoh8bQQSEd4fLx4PPR5BsxTMnZPohab3rCUDP0d2sEMyJMBHCMk/8m6M7
ZimRTa8NBnKGegSpar+IL+uPu2Eps5bc69TiS+7kno/EdyYmmV9BwGsymb1QhmaBrFXFvaCbXYRH
7+5nFpOcjq0CBv6rFV/AWgr4Zz4vT0AMmdxxcbyaDQkyUpvmLkm/llKF8Uai2iYcjwt/MuEGSLY8
98zRAbh/TJn/IdzYiqk8FC9u5mepd5nLkjUG8m6ttDmsswTIfgV6OCA3AI9Xdk0ZIRsEDv3XEG13
afBrUUxSuCNKFPkWA/V+M0MoZS/YpafZz4CwM2Wzq+yGUb2zgwM0cZD6KDC41LpZqAloDObC/jS7
QrvsrdL4oyEjXQx3u9TCgIPbcqS2AvgWlGMgWiSTVE+sQaYOE5ktTbhtNIEpIl/HzFxUIA6yul3v
7hNYhspFDkA57TwkY9oxbaexsJbghRY0UHUfUHdf+nSXia+EtOQNNRudb5mXKrhONLznXboO898Z
IM3RXwD7qjttLH+Y7DO/y5tD+ZSoNuAXvtU6hg/iq7Kdr5mIalE7f0YAm0XDuRZWO18Sr+JKmacd
ZNqgtTI6AbeIqp+1xVeYDuwPuMlLIpqYFgtGHWVCjJuJztlTTlh8H/42cRqp9yZBY27l3Sazpjj2
ZyLLr2salQNaH9If4u4flK6t/PCAtmPyEiinOW852mMzbWTLo6K+/cQce1bfSraKplZGTeu6LibE
DYyUxl3478PG+loHZwUmvKlOpgs5AvpYBVNaM8bSYcBOPCsCynvXxOSPrRIX0567pu88FK2p0tSU
dNOO0yCThuAWZ1niw63VWToPA5U8rBzCuZXPUrumw/c4Gk9/Upd2rVHApXSLEN2FQ3OtHBxAUxfY
O6Zea/8hV2q/OwmTPbKYtvHlGUzWfK8+UHKEuHzOYvBs5BXn3oD732czMuE4/VwEkva4ABLfvvES
84zDwWaAk7g1PkJuFdFtrige1wbNgo+eodr1FIDjdwn4XWk1H5/YgBb1Ayr5LKeC4OfFIuOA321a
T/cdOh4IRqX3M51uekUnbQuAoK/dLk68Ic6VLPfTeD1fRlx6DSnRmWPvU03gYYSX3svK1gii01tG
U3DcGEzEfeyCdS2LZELq40c8krwsFcSOS+OpP87zibs4Ogky2GnbBg20mrZPE4RebrIPO46sGyYf
GZd0N4NHjn7N72gDuY6R6utXaQNmDpuxPyJOGr26qL0s2wy8cJEU7ObHzcRhAEsGZC6dygGCCuF/
6v4U9qZ2CBwbt3wWkCNKKUZ7s6IIf+jGwM8PdTznNoUnrwR/Q4sFqwEHVmbv9uz7bPf7q97ZGQF6
TRq24ZbkMN+X2rJaAxQxyLeYf9Wt1X3qmHG2fKMF29t6tuoCy15V8blziHk2eBTEpVF72CQBz5oC
aubJ1VkgrdlKodKMjdHv+VKA+ocKcGdp9ubb4kp4FQYVFClT9VDGqB+B+OWaVafhdqsXUXCWJ0Sa
XXX1l5+8nATJezy0y3o0m23Y+hKtf++YIYmA/4NJcaeZhMxwvJDlzK1OkUM3Ube33+dUJVXZJO1+
37jZWfQA0nXBiNzHnGc9vm0DG4bdBv4soj9fwDN/nhDdzSeCOLaPqyJqA39rDU1F8G2nGvx85P05
q/jHf8XxkjuP9YnE49rmPJtrpcXdx9W3QiOO3snPEjGR0P7GWqtVACVqUnHIBFH8PtzZ8qg1vS6p
iSo/ZWrVJsnZvf2c5dQoLcL083n002LWzh7F/mHYEF+ZBVplFXA8peGonWuGPqxrqx94W0u/DF2E
CpuBTLdW4LVlCh5AeDEnRS2HPajhtuxpzOgsU5dIGaDky13/G1m+EstlY5lMfL7rw9HXqWlwowle
Z60gXGr0Q2XMr7tadZULBG6Ln/AiHctf60OC9CUKd10CibXWoitIQkoo1sq+uwIs7Iuz8kLed8mG
j9tCszmaApftsLz8iDHq5T0+5Jq400AWlus9qjV7SjMe8xlGP+oAhMfcUw+9kRP+0RVcX0Uyx3qL
KXUBfN7zU+27LOnKwDso8IhocbyK+wR/l0jB8rV7jZvSsk2YmlRAjZFNb+Dk7gQPOUr1Xkr9SUDT
1RYgEgFBfS6qlTudA85T7nmPYoIUQBlPISWfdVrDo2tu8lhBi03qLx00PHEj6418HWbcUQlhctGK
OEhnp5z6h7NtUaLEUCnNeM2d9IuR5Y8PzlDf4ozODynnskPEG8ZyDVbgQhmXBf+hpHLhI/Ml9WL6
HSbpuHfltFTNDKNJNTiNEHpmZnas8N+emTTxtN7gNvfPW4uc9SfZrXE5dw8ycPRxrSiCYWpPtTjg
tmskHiduyHacL78tw9HYqgW3yUeqvT4qrIBrRYHNm9ztzTgRPqTXQO0PcExCLdpz3X9t3ESArI8F
ztf0izLrzTIVXX3SQtkL/kVLpWm4hh5lxENhwSBaGKjm+szAkqTLfUj6egO/R+21uw9+E3IxzyVV
6oWTUWm1phzEzM3tDK8wOkXUnCVXf0UkywxmYXf3Vjs63XpCJkXqDPdIxuSVF1PqZqqhIKBGufUz
1OqlC7IS8MiTFFoejEQgkmDegmsVNJ1AP0NszwfnuRNcuWqnTNuT6hhMNkl2Vop41knNIhq7P8H9
36y6BVMbo4YeYNc+x2LCsyoLari55+XbRreQG7y8NQGr935bj5pHoCpypins6SWo2tBVckrWfT1R
QRk5BEHuQfvjBERf9gsipube+ANdOX2awNdMzof5QzrVCuwDAAC9ijqZKSj8/gHxHdVoNjlkuRBi
jmPKuReaLLVfvj9sm6lVfaoCjgr5HT1ak3kMn/S8+U0bHYGg5WMRibS11LZWTyflfN2hG/0Yh+Oa
bhCOGZtcv+qW0MPbJEh+XbT4FIYfBjnVtJ8GK0tIw7DorGlQos6NKRrtVDIZxOKiPSFKA/nh28XJ
nTOFq055Vhr7+VqRJgBXFeqj1IQspwfOys1wPwk3ftynLjKXWFD8+xKkKArxUUGe2ZnTGDswaAj+
YcoXiC2UatJSg5Wls0zEboC/6UFnqt65sWOXhoTehJUVKIoVrDomtDOUGRzCgc4XZWzUvmO47RUc
PQiJH5SKPlJK5gyD+3fRsRLFOhJiIbnx6AvdIf66L/zL8lM8gvehPdUSoKZIigTfKJRi7XMQAwL7
LbZs5mR0l43eBmo0eNliqG3aG5PKA7K2ATCFuDyUaNCQl/059RDdjAWB9Pz/Z93wY5rjxRa4nQbe
o7SR7+yG+ELKnXi1CJPX4Vwxo8XkTU/3woZLr6rGzT6S1/BKFH/MRYGgb2UesHHBlq4MO4/J14Jg
kscbST3uMzN3enxgjRu1syoj9o8yt+p4POEByfD3YuarqEmcirwcA9rdvsyR4xFK+30REujvAfLo
qNMg9qzHZ8EQPaptvMoJPOHqtAWJTPq8ECWe5GFZi13l0/e0/0A1lJ85FI6+oXZ0NisMqV9pURxp
xXBtUqGNCt2E83ua8eTF25ykp2iFPvEYaHWbJWazBpN89iMW/YxzvkMKXa+t2ZMnraM2Uk6q6TB+
PTiByOC3BJ0sVMZ1iIaZ5ldlduvgCF1o1U6UL5/Iie5vKW38ALFFPB8WVTeIhJH2Nw+QCgFqBnur
KroVAhPi5uR+MMyxuI+QbuGAOrTQuLu+PLxq64cPo3iYJYZbUNI76055CzhqAn8S6AHtgsJFwGoU
d5TWKIC+0r1r/dqE/zXLE6AgU3ZWA0flt3VDIAnKVjTrSFehq9Eh+Phxx/7sLmvv9stTnsmZniAe
xEnXuKbhYVNd6oaBws+GcupqrceN2f5h9wZmPhgyg3I866lqnzxym8soxxwD85xKiwsLVp6CDihW
iSO8gfc3kWNHXD6jnA/Ko+o/rlQZU96yu9jy0LQsNJEy830zbwHj46jzCrLThIV2uy9nD9cSjKoP
tWHKmtl3YKO0hROhYWDFhsrmMMzqDlnyYEzM+vGV8lT9hzJXSx/d+xgwtVHPLt69oW/GXoPkEEmz
2c47D1oREZfiIp53eSu43M77xC5zxwJsQLdbT7EoBIuw8blXAV4IEs2mf/DZ1WWw5BBFIPIIaI2L
o8jA28+BfcofxRyIdsLB9pVUuEqvXe5j52jmofXK6LhsJrX6VVZF0iEA0EVkw6jwVcOIWHysPbuH
RSHu8av1PggBFbuOV31sI9z0CsdZOs8B+G27Nio2vz7nZ06kVMdVs+wgoOXetEc5ampmowEzN56x
aUc4UVL4eetMjTqjEhb8JSzf12Oq8HvArT7qpPZwk0OuIQQa3qNcUZLux50a7f6STskzmpAQ5+g9
02SDO+waXSqb9Gj8aUBwnizMuuiKGsFdw37+WIJLjMh9f6yx5HtR4o9bs0/qnLQdly/AIQbQm4Da
dgbN6nzqu0eFtg6eyqRu8E/0S+/N+cR+5LfnQ1Nl6stnswfuxJ6ajXKeGMs+OIVvuwT/Hcx/FW6n
QcLEc54pXJiD5jxZ1MjGo8LwHEocytTbEt3AAOOn3aVKHishlisCkR2+6kU3mgN4mu9brAmXfuIW
/AWRJSHlyXLDdirbUggNc0A6fn3yy9lGLQ8lZPW58uBuK0Q2lhY/b7yTsK9CyPp51nAi7QQx+q8/
PfIC2Syy2ZgZpddqWF6gRcMav8mPn2OKQtV+EGHF/6GgHsKTo7Ir/o9hGyNiAwFSVp6IFM7t+ick
5Oc8AkytcvydC1Ct/zzXpAByBOLwDHmhcVV3cpYX09YrRXXuyu2EZlRBEdmL1Mgmcm1jO6hLIMNw
AyG+WjoEnlR1Hbr34uUnf/wczyghFbbjh6sotXckkfTJS8BYwkFlZEHzuXRcEZdwlFc/OFV6opk7
plIHxh9/U/hxlBkWqpokFnijlVtCB/efcdSr76dxWkU5t2GZW3RVKwVqkBUIWXXrlAqhUGkHuB/l
PgCESwEAudEvRXkvU7xyveHO5CxagqtHxzXPk3Fnkddmt3yWhXjuaKnhc5PJaAUAZHXgYyuJFeSx
8kxpLnMogwbcA1xSjRMASu26ADP8cvWFbd9vdILojcTAaFqO5vpxp/7lKvot7OMFSNckSAlbY+vH
1gGEw8OSCOfbBoJz4sy3t82ycqOKE4RhP43/W/6g+oOjqZSqi/p8cdyX/IO/BWWc/h5FUS+VYt35
A4xIEMMs7ych4RHU81EJqOX6BJe9cignkSwMUs5aYNGr26OfYspp3RdmvXvAZamSnEc5v9CVrtbw
zY58olDLNn7DxH32g+RTyTqUdThCXSEyRGqc9/8KeW7lOfa1rMPzgoJj5QhMKZJ1B3xgYO0miomM
83kVPbVa9SK+SB6yIcbnhfPNeT7CqO433zfMy0jNDYaCX8/LsHZ2Ju0nrHTF8sL/XgFcoRwof41j
WcnNpqu85Ama0889GX8rNa2nCSDtQj1bsrzCCRnzXObqTcH26y3/ZYOwgamxVLpkZtPcaJ03Esdf
35F1eHLT81oXGNAtcFITN5eVsr2ghpQwhq3Wf/7THSOeljzMspECg3HgfVyNUcPnfYjiJKfsZL7f
FtBZBmVUY55HbNb7o+L4y1J4ohODnmz12KS87iNGbYy2mAwBt25IBeD7qrKpvuBm8B1PGXWnKV9x
cnyffglzMutPzEdnWOk5Hzxr6HeQPaaYPshXOxxMa+Pln/naHFAqgEc+hrkr15Ux3A91OK4gaZYi
wWe+e/MNoBGl5WMnp3nOZVZlrYNkwoM4RoYRX29juHEYTRQvDPz/QYcPo7lO6cOTlwufFNW7HkH4
2D4lE8unwAQAIDkIAzJgyxbAMlxtICpy5fuGi0qHY7z2r/JnlqiQp9YG3Jn+FeTVh2aesYn2LpZ/
WC82IFisq2UszKWa/AdQ4mN3KEVzwNYXYspHRfcuKvo3G61v+n8zcqV7kKwYwucMePVJVLmJdSmo
rJ1eMiDu6zvaq8FLpGmYeFaTJ4riCTCujdsx+GoUkHsybHS3snJ6dhc9gd+f/Jr7JSFWYWnXwFay
+TbQ0preJUIZaZ4GzQWahI33k+H4Ca9XCs9kDySAMKO7Nr1LKQGnAbLAvBzOFdxEHPQ7KetEB+Sg
QqyDL5bMorEnQ+443+fesPnNnZvh6vb1IwLNlFJ80K7Ou/34C84u8i0Fq7W5hwIXyKPopjNP5ggI
H1ANTVExuouD+VytHTdEVfLTfuxNuZrTjXR5ugifmbUATStjFiTEBBwy8SLpUsiyWXBendYFPfAY
R1LFjoc9nwLxhpp8Lrbqql7BUbnFZyReN5RlGzDKSON9BOK3XWd4vesZnVuVnvHExd98ivqRUKxL
eRO+8ZCGXKnlKFzKevnhaOcqkE3KrPE1MzEmz6V3VH8oyKwoTuNyceLI4OSfLAQ0JILUMPz2gCKK
GtM4uOKGtyCJQeU639LG+eqUey7QnhH5X8ZYxtBVQfs3WCoOZ+7zAcq1IQFstmLur/pdZSs1CbtQ
Eg3pI+/JiYyuxI+irvIWdbaf0NrhAPMmXfSX93aUypIhIeBK2IyZQpSZYt5qljIEN9fYYjP44fD7
slnFzFMHvMuZ3fhHhACVbvRAYjgvXQBGxioJ4P7UMtp0zOPo5F9Z4dkGvP055BC0p0pSyy+Wfoxz
r70NfNov/pftxIyGrBLyfnCJXffF0nH9fCNwut3RV49fboWKSLlL9H1wbEobVoaTGvx9MsloLO/8
PewDtrBNDuVT24oJeZ6Ys45FkF/YjpRdPIeZXuzEiQMxSEJqlLeeSy0XaLtQ2dQXemZtYU9vF/IL
JwiO+mtZI5p0aulQQHX0/lF1tf5Kdd/jUVuMXbbHnL2b9MI/WsrlAZgHNfOZy8mEbp3TQOqL8oqb
N/P537NgYr7R7L5XZHq4fz1Rj0cNzDEZQDQM621WISjLj7/j8Lyn1nbAWI9wTsmgRoqOUrWvEe40
SXFVk1dvRDnRoPZWO5NHJXb1wZ0slynpvkm+ZDrelkVNclW2tlkUqbz2y0zE/CXe8Fx8ClqqQx25
j4+WeJY1Z3DxY2ryjx+cZwuHQtR2LWaWNtmDk1pn6jAFZSwczjYHD1AujvNSjYEOstQ6860eCb8W
H5TNpL4kkmG1kqSbcJl1y6i4rRMm8vsQXkxYwftgWBvN7rdLhPBGLS106X3Zw0oWUT/1MTUmx8bt
SUYNR7lALmfKeBd9f6tr2HooxyFvsFT4GbtNhSD0zaKjWZs0wCbnrZvF9haOdM1ykHCAR7DCnnVV
dFJn50LxgOOzY45/Ozw2FzCYALvOmmKaPvxgs/OK7LOMMwIqe1rgU1dun0Zdnr9gUVQtpJNLSDFo
AelrDysOfO5IeNFMqVA0VWrHnsZNKlTtgATw++pbcLhiB1c+UaUXopEw9H9Vj1l5migB4i+c/+N6
VdNvcZoo9U7UvUDY2SMsTV7S6RLRzrsJK2jJx84rZwTk6PINaCjXw2yqwTizf/oIEIt7lSWfjcma
4d5xu73ywfXcqyFbVK7GF/+tUed3fxEC2y5wHqFOuHzDduKY482wkw3crgil8FwzcEWbyKHQs9qk
0H4WbrCmux67NRG37JDjYcs8vwPK872SsgrRwHuveSZ3Bp+qL8vaNpvNeOEmQSNBMUhQCy2m2Jb9
rBq3+IBQt+mtB8fSMeGqD2yNxYlDROxyMtkuU7rXgM5HJyGAIH08riMugO7n26STzYSvzWY3f4MP
Yq66/OXoW8Xbc4/zXnfUYqC6QyKVHBZgAWMbmU+w6GN/RLTMITvXiBowUoHm+O3oDBehlVmF+25d
sOk5Y6/XHDuQqikwmOJ245cgqAquOYlo0xOB3V8Hnd/9OZ4p4sv1a02I+Ivn1qPG3qngfqHF/K1c
zEyNubnOBeF1GtNXY6xFpa8dXFh+OrxGn7Wou9yMQSAWTSduEAcBrolb4enlJ0/l0zNs3Ve4kgWo
Nfll5jcUOym0jNz7u3o5Mn+DrPUxKCwDimqzhvsT00PjeTnjPIVpoZWrubByRhwISeEznZJ5tBCx
UNyQTocpDiGleWdJtO0SyLbe+vyUrCVw0gbIzKU3TfdeQk6asTrlCe3lF1af6s0aSlqwDxgV3KTk
w/q09WHPUe24zZkrNKZ3ycUZMbdixkMR9t96I6Yi5ItzdzRliSYXPtPrZ1JPaXpNfAFONLP4jPGi
yTaMh517+dWpoDZT5uwpoZvx9UoTKB3ng+VuyovMOumAqKusCdWqOjaPrXzMeEFjJ0Zk8I5wJsPS
MZfCSwxaT+ZiSxMXwZ+qhchOpSVitngrzByYKhiq4Bgvg1UwS3SpMOOZbBI1eO9yqqUdSi+USYNE
P9guepJCOOk+dPCYImXbaIevwdQf6Gq3Lx+Hn21/SgzefrXD5iKf7VRRmDY4o6vWq5x5M7RZD5hl
v8hpNirEGhMr+ogddzB5jEscCfLM9U9kYUtoUNoLq+6ykwjHUcu/3pXc+OC2+RQzkvfxRD8Pbf8+
pyDjBn12dGioJIKFeJs9IrWZz6shmqlhAbQh/b3fht7HAZa7Xqt3K+/UZPV/gn2Rzv8fKDMDMdgi
yw2oY1IN9cAEQBOmdNkAwZWRI11aq/K2/bLc/gpGu8/CVOpU9azgDZdBdNR4DHYE1Ch2EVfg0G1r
E/H2GHEyBtCHIAwb7XCeWa1lgpGrZSUSdxmECYtGh9auMs9UB2owb6smGHVr8Eaicgj9/664MchL
WJaed7xeDiUlM/7hDMVe2cLeLt+5uE74GINGBOUxLU4++XVO8qEZP/0D21T86RFsCmuqgMs7o1R1
hfe/LDHAbSH1Lh4/oJJCY10XL3ZEhcow5JHbw5g2PhXP6dmhHEqs0d+twO+rSty3nidO4qgXjJ20
Jthzp9u6LpbKyzZeJDY5Jk0oQCWNEhLC2IvVZOD5ZY94gg18X6rs7lziS+CPz6RCYisAgWPM5dkA
3Ww93Ur40b6iIVLzwTZFOG7HLe4nuegnJK+WwtzfNLSrTWcElp82N99dlM3qw0Xs0RRiwbVUWIih
UShQpuhkEBS+BsDTFkKlb2ahITu8xLiVRUmaHk1imbIRwp2Io9XcjcWaMAjERRX4VbseiFk5dNj8
PG5HgUxRUaG+i0nI0mnivsNIozydEVUZiR2VD7y2FTb6A5QJLme5nAzLBne4zjTbOLloCEIla6F/
/lajBaXK4Pl2YBpXcvBA/YqYQa9hrZPjxlq4NmGDSkLLtHenbgNvH67IrOJj01o2uPcNtucvkkMX
elyu9/MPCwiFRnYPblGchblXvlZZWeSSK76zqY8txWaVw4SzNIvGqJK1M1wfXu+lueK1fbfkAtja
U3CQicWaLLyt0vkeZJQmmUMRrNERUChze8k552F4BqCmTieL8tL0vhe3QTODNKs8fqV+uGzmfmWY
GSnxyKzuGMZF68x9YRCaCH63CIWS+k6fWw9CHD+0Cz4OMH3QoDklDcdWCPzjZlJtPvE4ojQeClPJ
N6B+Fi7021RBKC9tX+ij4Aoy227grBV51MSFwOdyz8hb7Gpi/Skuiut2/xTnyZJpD/RS2eVernDv
6/S7KGMKafGmL8XkPmrXHoa6XMT7bdS0cXFn7I6FLEcCUVJ/B69ASYiHECewr6+E7yyFRpV678Ug
phYGnaj2S45qOnJbrF7WTiNmNe/GtLxwW0vEdeXzAqVpQ18XwV38ghvXG/3RE+V3aY8R5oTHfqMX
B1RpfynDWvHny1EPsec0od6WYcc6eBdp7fJFmaCSWSi1LsBenrJ5zRAGwgGcDuOCU1VmKkdVhBz9
v2QYbs76oD6gYEm7c7fkz6ZmGaufaE7gtaWCFWVfOse43LEea49odYesnCfzoBM65+qNIvvw4Hd8
fuYVjAHSnr+bMwDHCi+b0eDrzlrSP40e0xqfjb8H7kpxfzhxp0WKleil0iYE9CqpQtHQvwa7zlZ3
/gxr554cONZgkSsIcoXlBC5uPdvZc3s0/+0nStrtjeozcQ7R68XjOmkIjZGaW8jHvNu/1ytjHoUW
MkjiypfjSCdrU9LpCRYDU3XofQWgr7fNnpkSv9Ij+fchvWWshFKRBivgwNQ7it64UWw/BsfWEoB+
ae2gDoHngQiBwlDpUePSslM5MtHyOaY3O86Y0zFc4OBfnblEvBkEdX6Yqhu+DWcv009nAQLNboC3
ucc+6K/QXubd5Q/X2x/WBo1lOy7GTWyqPO7AjWRuthjRMHSQX28kytchY0IVdgor2HnzDEOJXDG+
bMoBRmTlkXUsNPj0zsV9Tyziv7PLazFIRIdgTTluDmO1XI25QbAZays4q4wk0ykHdLfprv8o6MOH
iPFAsf+co/L3NvNvV25SgI2R3FdvMU7xbd2oXuUzr29hIJNl7474vWnS1nRS2YuYoU+Fd5amKKgZ
CRQD97uocFhGityPqCZ7PgussM6zRphEuvsDKC2w30eA9nckuuN4RMdlEtfhXadDrc0Px2ZiPM9G
alRpid1/8O6xHdPA1WzuiIyycc/m4ha33lPW+pOuq1ABparW4cMgF64LZWxvh/jGERu3ErISdGOm
JcwY2BEvzMDZiV/r4Xesmp3ce6zPazHDZQ4VZ/AoV3D54YXo4ZUUYNTuglsMkCoKWqDWUZc8zkOF
2iWRHwy6o5zAJcFtxI4riutAPJ/gPHiogSQnOSqjcqTo9BKq6GjUVMoCkWiQVyogzWEAomiDUY4a
/2ZrP+3a13g5nKX0kN5O3DyqBqZTxJpPnjgly3IA08pdFU0nPyvAeS/cEWoMOhWrH+bsRMb3lnl+
Ur0VSmvbym9c8mAsqxd/rZ35h8vBUiOfxcdr0hz4ajIFVv97GgXVb8iEnklTwOPTBhEEs4OL6BqQ
ewiuswoJZPuGgEtxpLAOj9xsjuGptFQ4CE2e6ibWC2MTj9WWH107l8SlXs1NRhBCdBNTHaAZs2Z8
bMnft29nkcRxB0qrFxcswljgZigaqn+yNb8E68+TALR17diXs4wLyC7vDnyXVRfEsbXxYPD4KBAi
PA77cCzrNzO3O+a1Ue8XQM77PBU60yb8CNVnGQeIsuKdXHdkKVrZImzf7mzl84Pb/VJKJfKhkV5z
HBvBtSS0gzoIcoCgf1dSPggcvCj1DYssVh9WBf5qyJHHPSwwCZqY/Xd5t0qzxqV/h+YkbTiF3pwO
C2c062Tt6fEgYu0Pq8CVH/270B8mnl/Y3Fmx9yHJDw4+T7fP84DdfQ6JlWKg7QvSZ55cZi3AsP5N
B6s+7F2TFUSWv1tKE5/qYL4X0VEVzlGzbzLVdRqhZ6+H0GsWbfzkJ1446OD9qqlr8yqEoBcYIxNZ
EGNqKHjDiapdNKbtMHQliKsyM644I5Pi83qDb8En3DYRFgXpxZgPG33azCBITsXxlNv0kid9KzR9
uuvZBe61DSYOmHV8hzp2yo6TGz8Hxr9r8RqCpGPnYkn5GU7z3//7hUGLYIWyHpDk6O2wq8eyM7KU
WiS0Eu8Crfo+vcg2I62S9z01M2db3XiwHUBnZn4yflTOryFTwaytsJhYX0cfUR3Smypd4iIhc1Jb
zvKsIgfkJhasU48tuoKtt9AnWvYO28yuHTIEXpj1RLTxeytCiQNyKmQt8kS3YRRKhgkdE0RXArLJ
5FbCwVZ9X1cS+r60YvX2ei/5uGwPYwkXYbymz4mT37GAIfC9LWZo3HOLhZ60wfAwVUD+qLbT5ucU
YdzpArN5w21NMzm/I+IV91McOAjK/ggMl68j+drwQYXBAHQo5uPiQUFrSsYB1PNB5RsD0rwGkHch
94IuiHDCzdTvx0ozdnm1IvZxn9kKgGvUyWLlyAR7BYgzWy115cg2gvJybCqLfpE9ZMJg60x1WxRr
VSQG9xJvuLwy7SEGvyJf0n80hL82L7Lg2m69tptoYUWxlVjxgHdcRT0DU63dwGmv6ePDr+CGGOWE
DekRP5gQ1vYljycTlWcSs89Rzsa/zSzmNIDFWLUOQQFatH7r2PxdUPWjMG9Z6/B8m7Zz1h73ygq2
6N+Tbkiwqo7dvm6hzjIx6xURaBsp6pSGO85cKVvlUhhRZLhbXNNKRWYYPU30dLgFGS9D+5CTJI4B
1QGDFkhTo3Zu4H/S1UFdc1NX2Y05wrGRsqKtXpGQvyWD8XEti4J1AxFWJn8TT2iDKdmWHJ4Yqk3d
JCQijqBoTWMq1OBRJaGBZV+SsSv4QtKbFtSL1C67xYB+wRYz3OfiYxkDhicCo3M9TZxegbZQqLGM
8O8gcUhiznpA2IsMbdzcTJgupqnJ/CSXkjDRliqO74xKf7rNF67t2MHuU4yAwA0/UX2UxFQiruZi
4+WxRs21UXVZBtdYZhflItnUXskFVl0GeQYgc2HugGMUVOgouKxPZDkwD6Izy9GSiJs5RQuSTnh8
UMTcrNlGZM5k3pxXHlbR9q8XREmLQRGLUopD/Uqjx50SykdevO5m3+iswrjAIiFvXNECNK+78RhJ
/JzfX15CNy13Wkz7D+WQqoaTURx4vfUvXg4EXiLcB+oeNQW1KqUMPgO+htohAJMgNZZC21m31QWe
Ur8weVhj+RcEGEIUaZhPu5yPfZ+PLWHqpcfsLKVpo4OaBFbXTkaW4YYA87o+706xolhyD3WCheue
43k73U9tI/2NuI8azln9AgsE/JMPtxbW/uXcl0wxNMlfn9VckmPVOmh+2XKvN7++JfVyvT0TbAW5
HdTQ/H2xJsQXF5WhK+y7CGgQd55PiASXxQNRKlfs0u9d6xsyEc/QDnsl1dRGK7a0eTiE4QgjnjFp
ipFAGohd4hIrTxxUX0lvj/fzt99MZB50iF8polpXKKQrlM6y6xpageGe5wBIERpY32JQO9BorVGW
l/NLkHiF1/U3hwL7Odztn5QX1j4Lu/0MXoam8JcvyQjhY0EW7B3LqHsunckcmig4rPsYeIriPt8b
TPedAIV2B+y66tKUcb8y6oNLpf5rzHoQqLRmYEm+yVs2PD/5Dnw4VaJ0Xut1nu8O2wrHZTwCdmMe
cmREhHXPfDIAD1AgD+O9XGYun3PkBrj9Z3fSPVj/Vkt6469gkNnHZ7LzNyJdBjdf5g1FclhEgKjC
keH8wYBorGsm7ZPrcLz8Aey7ARtZ1lVuC6vP8FzQmxttY/tZDZryFSwi8YoFVFprzWC7dR3+U9L2
GmnTXZcVLXK+TqkIpKTlZCmlYKOuLJrXgCnTPMItSGPHZioTyWEAVQ78uiOSiUOha74mLUp564Z4
CvuO1radGuIMzDEeXSEVCbradBA0KtI/5Uf4IFM74HXgs6orTVFTh3KI8+uM9na3E0jnHq3o0Lyo
aas+kPzv3lmSW7EZxXiqy+aAzTN9u/PZzsF+bfLA7RXy/QQII5t/czs5eGOora4vPZIPbirEia/J
hytqi9tkSdUI7zACuCwyo5ZwpYTzGo59LZEK6/W2mRi5Ti65SqzZXUHKV4z4ZbN31ABdHo+S3I4N
jMWlQZWspci7NEn+EFOShIF5+Ja3v0zUGe2QPNN7mNgas9DOkJtJvDCnh12nF0ITlnQtZqsGoZhV
+Pn3TFecD7Ffx0MqOqMwL5b4WdPovhvcGBfz65fix1ND+Ze48YaZ6D1vp0lLynARq7eDx/zjd3GP
rG66tmKf4/KfWgYajAKCjtIM1myiV7Yw3sRsfDY3vHt+8VI2+CCcVxGxDoQyEvpwYToKcAeojJMw
WOQJUWbHWRhkFD/utt7bVRXnvv3LcKNImmtiVqwDJDdLMpf+UOPPgb2+hhYCjqsMs8XDjJlSBnFz
vX6IDiOx9rY2AgGl49CayBAYEC0T6V1oGmo3+Rqy8U8o0p0T/Vt23pI0e7GM4aKz+Lfv1bBfUjI+
ufluE4PU3kEG+Lp8nGzS9jlG9w3XwPlyMVrqguzjNVgVrvL/koX+1ZBkozGQi0Lwuqms9Coo26l7
dsZIA8qE8BJBYIeusG30ybiY022LUpTA/hCE6asb3k/P51P1WjSmSCiW9g/EfwnFCmnRwmraZjLi
c0copfqH3R2A5JaqXSH2APzRNJYGD/FnDtGWu2ggSuokGZWyKkGYfq0zN/4SexJkKqlYxYpSQS8r
dhaEFdJLFpdk5Rbp62IM/ooJnzsv4Aj9pz8ukZCgfF21GIIcFC+XIPsB293/RiCt5WDxfVk6ItKc
q/pgjG94ijqZSRIehMqla6uivLxEUTVAYxXjOSLt86p24YTzjZH0LnwJVIYmb0jqyT8pA1Qe/CpT
YnUBAsJ6qK7JN4TF70Jf7ObyO/4Lq+oLT3Pet3eBjgj2Cm4x1I5+MYxRbjwVSP4ibi5Wr9gnM7Go
/oTi9ml2SBBPUnxNGpMIrZoPsgD9e9QAgHfItIOlsUHcR2qMlNXdJD8DzGhCVrxzhlQyIOJ+InNB
8QvKTlKFZwZskFbcscLGuPDUfnltzjergAi5SjZTph9/RbWAkpB13dsacSCpI3NraiB6Orx3iX0X
kvPByuY/u89bdB7L7wLkLYQLjG+XLVC4HU4ESMxS3jgQjIMAucxv53cNitzgi75LgIa3XnU82AYS
nWW7RdTc8FwAsPhu5q9CSsq/bwh5G5ui8odLK4To+DmIzbaM2JuPl8kc1WsbF55eTPfl6fpBUI3R
+fnDteoizQjxtp5RstxpAUHruun5IOKqBDO8u5Sy41cF+NUC20xv+qs+sTsMGN8deu3IMhySioMZ
OK5FPFfFxkI1b2NtKSIrdir6pXmrG/PB6kKeOFihVB9la6COJT1csoZegvdNYpWyqd8CVawC8n9Y
ku0IOvJunCtCyzdY8rRGqSO+EoL0eF+8VJveP3Y0V6raduPEj3LBxLtDTqLxpEUCidrcMm+P3EHH
f8xcyzIZjTe7AghBZYs3k75NOxJGrJawT3j1ydkyPwOZ6+jeSNuHbTZw/TLZWHUBbE8hoMEcU6No
C7yjVG+amnlE1EYH6D+lvoLB4th/2rxpDwJeB+XC34aXiOgzKrq3I5Iv5eFawdaiLE2n8OScDYxh
pYQE93LkFb2wzTJgbhNXGGnbtAkIrZHA2/pdvlo0TSOQjBBJJ35ovuDAMrxaaF4HDnXcoB3Hoh/B
+A2MVjQES7b+ij4ZlXxtzuz0Ur2IHgYGMqpjbbBQNLFdmAqemySqCX+JeN3ty6Ggwn5sfXyqjxfh
N35wXoEvmP0hwTxRZ9Ijhd/u6WAMHoFqkgnQLiS13GpPF+3B+tbO2bO2NZo/xxyMLxxoyUpFFDBx
iD4ee8wFgnohL9CmdX84ta6lPNpAaj+teLZwf+U2AOfykUPgz+kbsQ+JdzOoSJ7lkRe24syhjeFo
MXk0bOs30dt5iz1jI/iLXLRWRlP5e01uq9uCgqp70o/EborvIRMR/23gimafPauOvF1Jt8X3BP8D
UF8iBUVPbspF8nNC85WdS/GxILidWGVyJEyfyRQ8jpMkvSWwdB5w1M23Z0bwdYUPkhk3P1571ttF
uX9Cr9lU5ZeZ9oNS1BNGOYjM/Qna0vsHAJR70mBYep7rCb52G1GkAymqm/wo7vrPo0XHFs2KCVGn
ACn9QrIaSeKGITXiN7styp1VzBEKWvRJd71AESPa4kp5nbx9WNWgmi1P4GudIDX01srsSvjylHsC
kd7PO6mJLAVnmwkvzrMjJtJAClsDFQYgWqLCw0LK2BJ+Cr4TKhSKlIV6WmAAzbixry1K/PIcKL53
l9GKiAvQNdE+uTb4CdueNSyCWrrGFHsUz6jOIxbIwD1QlLzxEhv8G4QTdRoYsO4+zQHau2OXtOcs
vEDJOBJc5Ks6sjNu3XN57Mr0C6+U/5Zmm2mN0+SYvqaEnxVEzir4j50ZGajsc0mrTJHxAqRkX++v
64gOoXZM2MxPekexyk8TnQIB/gYFwIe+Eywo2AyNKu6+R5u8IxRmiGWG5CohG6n/ziGiyxVtxUoI
9WLYgcROoikryy//yTP0c2OKRnA2vjIsrRCn3tztbnGwSaX+vTD0bexGK/VLkTcIYyAUur4Fn7s7
c5peymn0bppxmm7VWCYX6QImE6SV3tfpHlpZh1Fr5o16Q49YpTc916zHVYEIcze1y9jWNXbLn61u
ju9doR8LbG7Mliz5jufitM0GEIQ/jaxQPlzZxmRORz9EYQcnlFpr4N8pj1f4iTr1hyw8/UskAov9
eclHkZmubTZI6uH7fcfP23IxDZv8hHmeOvksO7EZaE4//TkLkdyPOgNGImf2Zxm/yyNZa20ezWca
w1XF1xyWl5z/SCJKXm3NCd1HN2l64aeaEyFMamPsz9+g8sxxy7q00VIBEnaj02Joxkx7LbzNv+ms
j8wNIT3TB//LNWVhQgRb/ZzkwQaCxppWyUeze1o824ykLCnSmpGaUkpJDf/zDUimkJW6cwH5N+5n
zhkwVcp+e8RhmUyAa2Zz97RVq8MLzXM5UABLTym81gAzLvKme8bHRyDNoCFpEBDk9HQS5DlBGDS9
gAs3C5nvSKBGvyrK4kHIlkTSiiWHH93OytOYIVCJcQPxpKhKIhcLjAeEgf24LVXAKb+jgEq7dKqc
nQzITajx2ZZ57wkBCjIP2FVpSy4BPBbXQjlqBev1lYH4GPaVxmoONavDq5HUV36wa76Xmj/yaQQ5
ai/Ww4bm+icp1crQ/R6Bh+uRx7LPlyZfat96ppgabFf5b6W+m4BnNLRYeC4jPON8YmMD6RcLjbC5
sUSzOeuRPWL/B0i9kmsOTdu8rJDUmlrqzbgsN2tt+p+x0AZ31TdedVDIAAr1fNkdsvwApuZq4k1w
4UoBL801TKIjlsR7UoEI3ZuFD1bkGPWnp2+0fCgsZ74IhO1EuZq15/26yeGPYG0GZvDbgF+9JZZz
pnY+ztmbLQ32xSB8Ina04IjBocK0zZJ809DJEalyyyrgQSr2PCiOkOlHJib1gkUqmwE6ob8mJvrl
c96eJI92PhNiUglYqE65LPMYtuqTFjNN3BK3DvksER5H8HVDokQ7o6SsdSG9njTLL0XEolGsMhXP
fmqpPMs4D5AFmQ9K7iIhOQukJXAlK8xiuGGo8qG1dpGJLCJRCOthjh5j4xyiids99RjS2aoY5WeO
9Qx/MuC00oagZuZ4laNIYnyErHSm2lhuLVrkXAN0vEJuRNId4lq6pFgJUBSOIJNSDgl+rH7JImJK
ZNFhjHSbSbskQJhV2hLfNiuD0sBHhVmG37DpqqgTctjuLlOUurdu/8rG6UB+7jvwhuJtnFjVbBmo
ieov+/yP2b/4GsBDuIkBLnkU85IxSDIBeBgqiZWmrw1xJSJQ0acEPEkvxFv3N6OeDNrNdE/bwvll
AHNBV9UQwnm+y7mVJbY6/LezgOMYHkzlHlvJIIC+mFpbyW4d2EBLveWl1m2SwbYMgfSCQV93ApkU
z8R6sgLZQ+mCl8jFQX9oDRZFnwmUiLbv5ma6NspN9FKXQyalAHtmn3kchjRSKKsB3y8wkFBJlu3g
RQ7dCuwjpXI0SAVW8KQCLdw8OXyr42vP72b3hMzn6mBmP+UF4M11NUNDQFxmY7vVLh9buR+zKQ4T
Mc4zh6T2UhIalYrDAz6xTfFEMl7/yzvOwfCjx7a78d+mOCzOzOMC6r463C+g+/051GKaw7ZkAk5A
PJzcYHyffCuSKrSA44Ho5f7tdF7s4wyYWoEKhnNA6OhlESgsRsGAf9PzmC6tqq2JEXGut6tGJgwD
eLPGRXrC/vFaypSrUOItlGi09RLpCI3uvSeUFNXmuyyz0+1gGTEmmU1SfG8HOMfKC/6k/AStHuSx
U8GQ7yDoVdD7+xYnN3jFHZ5k4BsAB6fGKn6muxyvITV5iLMP99Yt8rOGPsri62FvqF4hHQC42HyB
L6RjgchVB1BH+DbJl13Zk67GJDlD+b0x+VgQwe/CMWRyLKxFkN0Q6yq/xPaHhDcIH0BvtIuOnivB
FL3qY1mjOoP4sTDGON6aVeLN2mah0bEv9JF5BdiDONpHRaoJMIWXtu/MgV7cMAXiHuU2JxYVJt2l
PRwYB983XjHkkJdQwEivHZxa0tndNXfpnK8vwWc6fFFce8JsMzW4WWaQLpHlZaOJ8DnEOWJ/2yCg
TX7tIKY+V0q0y8lygCMnFkdM57tNs4hVYdYgB4M58ed6S4bSZ5Yu7TtT2jq5mnUphXuYzX5pRsvI
GcEDw+rOFlq+ppqmePtfZ8eDMFbyF9lA5HDh0BgMvRxKQBSpkC1BZ9ovZyupZ8VzP6rkBjSGvNMt
++IBxAZ9YMLfcAcXErXT5S4Ky19ks4UQe5J5XrGLLNE2MmMOQcC+WI9h5Ss2tcbbvInR7dHb8wrL
nwah0KTX1lPveG/Zu3znLVYeDn9R0RuQ7CYFUTSlwFYma4Ld8ocZGBjUhJHm6k3xOzKZRGFoO18E
YGOo9AhCc/lNVu1FgZeV+QaAZFc3+iSK5gYo4DaPkAulHfygV7OTKkIPP6GQOt+CejoxExlgFZfQ
izOPl8HqNnJmsaYYpiKWZRxuYaP7Zf5dNc3lIKM9+mymBKuPbMZRjPDsOvorUUK4p2pMgmwpniug
ztpIR1rp3hWsVjPH6W+E67nlehtz3VkQ03DffGmHZ+cyXOAUY76HGrqiDdMRdUHPaqe7rBjX3d6z
QlEWKedw2zSqqWYhYkV1xZPLd/l89QHmNUf81iG6Ot/RUEtIRpKbJLk6mEeI/ew29Ad8nN5lR6Sw
BBNvLsvn+ts5hLGRWe01JNSYJqBMqdBZBrX9RVUiwrgC/fmPrl19sVxZsr3YL2ZhtK49VVRUCsED
qIQEyqgCk9lcYkk+MoH2jSHb/zoetg2dE5kEgaq6OGy2Fs4bLrlxP54Ym0isMk+j2YbCNOHNRcqy
q/SCak7AWVPup5m2yJte2jL+iNFxy5suCaesgj6Y26quPRyp0Eu5+2gMecB/KR1gzh8hSXSjic6Z
F/lAOSodSbAypdDiI4J8F+0JAGe/S++qwEC/IGp9yRKYSSQTUHmOD+JxJVt9wKSnWFrWyaqZy+77
uYhsulprYi5Qncuqf1V0na7BaIkKTQ+TUy7bOBU2EKmrn0NzDh7+P7GSmIAkMKgYL9QoEq4ln/Kb
Y5wfCHtY0W4NRMu4kbQemxQqvxg/e/rQwjaRi6OIwyhbM02+BJ3Y3Dz8uaLE5tLYkc5DMPjA8ODD
8/3QqosIxZ7HFr7yRO5xEWaUbLuJycve+HlM0cikuwQ4Op+iPZ0jAn+5ZRC+sPCV4iAMUyiTuOkK
goCdpjkIubMorodIFrNgVBZo3yYvDM6MapbiE3OeVxybHw9x1scWw7TdaeEn7v+Mabth0Iv1wWJL
g0UQ4nNtaV3BtB3zWQNPYw2UVVwTf2pQhbGnD4xjCXeDf/ZrHxkmUXg5JB5aaoJzNAA7CV/mB7y4
CJa80h1ASRQMBGagg4av2KaHzLQdwkpknx3IH9L/qPwdWf/HkV0GpNS+Vd5BYMGWt0R7sKHod8tn
DQJU/OAxiy41FBsAbcL3gmTxRDHGIUUCToZWhnm4LLlYYpQAoxwyaQGOPEis/tmkl0kZK23MK9l+
Dx7MqV13aimA/Io0duPWGqbzu8KtTGCk+8K+91i9REQUT3YF7TIFTonHURxM9dvQt36M8dxI0p/b
rwOBlv/l5Kr8ParXVKbTHoCjQiIdEgVyw+nnYgUBeZ6oCs77ZVVr4A6POtxNcLnUCdQZP5oOY4fx
ILg4YYaaMv11Cu4UGix38EcFabeUrtfEyJqf7Uy+fnMlu9TXRtGJfSPIKDrC9u0CaaYnNWq6RQDY
ovuT+LbzXRv75W4ZCV+r/oXac35IzcZE76W2VMH2+yBvFKLw+f0kBDjHGcPLi+A22Dj5S8D383vm
5/hBWrJp9WYwuIsW9U9J+ZymTHiorI+WDvsCYxjM1iIQbG1ZSY1xUjaEzSmyZlY2qbVOsie9PKBn
Fnj8oOAR8l177/u+MZweh9I1/f5rwUa0XA0DRFybzx5oBBhuMETii9PGx9vkx/TFbiK8Ggl0tK/3
fOCkijZL0vb60GtDn0/kNW0wDy1qZ/sZhrA80PB/FfwYiXN2MT58kfY6z0ulDkuXJV5pb0Cx/TpX
zq8eFJjKQKPf4CaWNkwJiI/Xs18kO567RaPlivFm5ZnmZV0Lzawc00CMgImU/Pqh0tpm+ym+pxIf
Bs9UZnEtakZAdkFbRpjDDqMryubrt87j6KVQsWnNtiRle/yFZQ9nEUdeYBIp/i5F8u9EjW7IKu5L
BJDs1AcHTt0+gygW1Ka0YldpGSPa0FlFLY6HAsf2TbRxAb15/4ODGInRKz9sfo210xzOB+BJE5dF
yYCu76XquVHqzzxWT5ox2NZkFRziM6C8RB/bN9MVWfSUxeD3hS7qrQQJmZXm6mr7hTFgW9XQvBb8
+WkNBfidpvaZX3KwmtvzUbf43ahQfQaij7We1Ps0oyAQ+MkNYa4CJFbX7yiQUwhu4YHUXKAdauSH
fmAEMs+XkzAnLdmdHwzdNrOVo5sqofSR+/9+/bbpjrV2KUt3pdBiODdT7BAGQF3kX20DbF40iAvi
kL6lHdcuPz1ww0NydRssECsVdnAQonCA/C/PsDO7k+PBUExTzpkzTQNGRIaOle0iWjgK/JQYMin3
mvshdgS8F/yCVeMpwdSgPQpSJ1HZWyXhn0W14lNMX0tLt9KrJnbttskoNJWzOmYnk7Y041bWA1tg
shJeMJkTsaOX9ozizJRmKeJYRKqT5+AhPbvlZpwsCMhdGE/DkNYsZt+AJP8+6rBda8DDQoDEX4KG
vPNVP+70gBCPtVL1ggIAGy9MS/6pfy3DcKadgD6lYHA1ELvcKjoef0pz/C6m3FMm9fgbgn0AcsG9
FszArmCZHJj9cQBNm3VCHkfwSbZYKoclVghyZjPGAPh78lVy7mLVP11G3APva3itzMQsW4qVGREg
93zoc1Hx++6l1QAyw++h/ArWFvuuQIsXPk7IR/T2Z67i1DHX2WRb59zTxStjYb1h0vY3y7LMDEoA
/q2vczqVlMLHnPeEvcNNTxKavfKvEwStDS9cHx4m7YPtY7uKY1XofnDIl+5aQAmw/FiJy8MbOvbD
WD8fFTMsSrfUbMnI4lrENA7Hrnh00MzGwKxVmKB6UQEZXSdB/sSmeJM0nVQ6tBK9FDmY1KiI2lPb
p9GiNUmbfXU5WEzxWqyTmJ3/zIhm9CtIdAZhenTdivXCxYYWVz5dGPGuvpV26fwJ570cNmVZYilL
9KgMnKVZoydYX8YyGNBhbGVrfyoCx9UFC4vJjbzFAiR6nGAfIALmA5exqDkzUaZufDp9/bomKFqu
OhXcwNTTegCTpC1jY/BhLIhlRw0d74HAQPs8c+xsfUje2CW1z8Y+rIAIXHzYW22S3SuWhzV++3L8
FgX54yuKT6bzNLNQao3pftejkcIPilCdCBR19DuoXS6PFHpLNOReH7sB9NP2TCznvV8dkvcHxi/7
ybGDn+B2j+z2lTp3lKjbzNxs26jvU5Lvj/wxijL2WgoqBiiHxBTZEn3cgpFMaQ1yiR0Y3CTJLE0+
blEWg+8mTbOGC+/A83Hov7GcR5dwxaEVj9bp0FEzs5VGB8pTvvGSx2cSMPqXVfoHMr4Ck5eejqWP
7D5Cn/a0Sa7TgqLZ6C95sLztYW3k4GFNPpwUfhNAT6ZmVYEqp4j4smLtRGSnpS1ojAAR6gtjTM1k
zdNOyt2SVo/KaDvnEE2CyERA/0ouCAUxPbDpkVTGwBXNqkhekhUSr31cMI/NxuNrsDEMRvuZYuhK
RhzbLynycI2J0EjnKvckawIB2NSlbZCL7RaNewptyarK3dG30Bca5sns/WvISa9vNvuHiVxzWrRH
uyxp23rmRyZLqDW0IkjO2nvOh6ri+wtrD5/yslqvlnOLIiOjkmPQBNDt2i1cjXOC5DNxoLLTmCzh
/06AEc4xn6cf5aki2ZkruztTaql0bANdE8wKBGyni8XsTcZhE7pi2FNWE1fFFTlHfHbxwAmMTuWK
jDpshFGvAgJb5V8lahI2upP2jNFWd0d6iVSUz/p9Rhb3nXgsjjMPECGWcVRMD9CvO0gyOfvZhMCa
02r0qHICeECpdJ2jH2LdKM9R+DW4Jhj0xfOARfVGauAZ0BCIkL97LRgkdFoyNlNtNDkTDBn1dXxV
rfmtOYrJUb9oD9lz++/1ROuH3iGOZEic6hCdbH98nAopVFjT3YNWPZTOK8O/LYCs/MsxmZAJTJT3
TfONZGn0tz4pYimW6jjBLfTIS+1U8pQxQdRNBSijKaZ08LiOi3QdH3nlrbn1olqJRZta302Qoqhe
pISe2Tjx6tfB5AOxEqN1ZDWxixoL3VtVB3x0fnF3ETdCRvvjPH3NA64IURNTIGRe7imiNLOcRBaY
Ybl0nje5R97LVkCDyBlr40baPoyed4rVefoKjqLpv+HvGJ3M4MuoxXzd7xauTqY78/l0XZklPmZM
0psu/hmLJf74aNw3J5q67ZNYC0JVVwaLfxaDjp4bez/Bo1neoqxcEURgqsFJ7gJLSClRWmF6PPaL
QrKTDbeJ+mVE/oYRrY+WpxPhEr4VR0Joq9aK3ewxz/euxZE2bgSQF9RanfzUgEROnsF8m17BqXmW
jvJJ1PKOFI9q5Lc9qm7WaFad03MFe4lRSjGGzglKtY05YuyB3h2hfu45plQl+QlCumanos7PlUNs
avVn0mA7xJcm0m/+cdEUA9nGU0AZaBo2VqHhouMn3rGUDUHw1Fu0yD+gCqbRMia0pOyuAlkj2pth
RYNu32Qa/Ob0uQgSCu95inL91jD+Z6QPfFH+N7rOyti3sMG2hVdeA19ip//P8oIFj1Ij1Sb6auTM
Lm4PxVDvV4Mpp/JNYbfoLYmmaFBmY08fLjWMa6fyS6uFkJQHmwUOeJd66O8enFXIWgpFxNasD/nt
Ta8y/TmpPimiWsEP+LlzFK7jh+adsPmBKvURarapuiRIQSWHRHvrN/VXQ8FeE/AqMqS6ILO9LU6Z
cTmJNs/RqQKSvBOjzMmR2gMqJCtHh8xH8sxcnXB6WmXZhiIWepXZfUiFQgJfEgef44XN3DuFBZmS
dofZlsua7xIrL80Sndo5FlSpPFHOxKbsH2U9cbTNiesS/z2oucSjCVujmBjp1R809711e56z8gXR
KxTXKotM5ArdMz7XMIpTcuNjfllGkJJOpARKdlv1K9nGKPF5vCDDO0ScAK6SDI4/1vXCr3261D10
UcULT/GtJFq4U8OWsRqYyTQ19+aheIlFMX9MFjoz7q4JCrXcOqQMD6yqF3AZgy0bJrLP6zphqh1h
qEb7QJeZAZX3Aq5Ow4pBXZWa5Br6CJYYSkeLLzDD9WslVY1ckGNz3fFbD4tdbSVp5aLeFxU4wiuk
5Ulgcu6H/+D7Lk0i5mY7sjDqP0eWSdKKn+A7/OeMR3+tFgqj0t3N1UDuz13ugI5033QFZ4pFZEUa
CejI8m2EoZORc0oVGAVMiZ5q6irJYCgMUiy3+xF5iCpJLUR+pfpI4oSnWAq2FWOI7Hv6/Q2DrZV3
ihiPSASgetDo8NSIzPeuDmBKt5Uy+c4jHQy2Hy8acEsTLw3AsD3bZFrkt8llVQg3WUmpTRFqdlJW
NNhaSuu8raSHQTt1L4ohb6VdXAZ+ftsxO0MWxbeIM54/23Jb3wXR9RbgNzV6mIZ09fzagZMEc2Fn
cJ6P8y498Dg7O9cQrmO9asPVMai0LKQdZ510czP58IILlzkBt7Lb2P1eiKN8/dqX8z0mPES4uCGj
erk668T71Dn7fnLHRoKUjdGFyhh0e7OnwkiHWiIaGzT1sCM+MckLCaAF5Mr/IJiyKbHZpzJifWFx
N5KXuOskLbVUPebj1TksV7OU5VydXzNDg7yayonSgSi8RuFpY3gk8e6jfK7+MoloFrawd3axAvFV
XtmiV8Tn4vyHc+p2Am6S0l664a2X2NDWpEFFjtubzel6NoNvD370tZRP4OTCGX2Q6bQZgcDTmCQd
ucqXwHC+TF3d4HSD8tlTclpsP/vag4ovcDPRqWvaUv73/R3kiquVzqkuUX6lR4CW9DbwY+JeX9ef
yoFiwe7ctkt5C8OgvRzoeygXxr7b6fNc4Gm6MNnJ5/ubMenpAaEhuJMqKAEtKYp+x+FVn4+eRJtj
BI9I2ciaxtwXZ4pFbxLlhG4JTo06pvphg1IMke7dM82lcYNwpnFN/DLU668HYA5Yoe2zi4S1ATnj
L4g6fs/WY5AuzGTXvnHZy03dQfxhD0tCqMUCaroRzbMJ/eGOQGXuXkdAyuRc7MUBjbHFy0kZxkc2
8pGvoeah+8mwDtH0CTs56GvpAAF/5Y7FU1Uw12UD7ZLz30gV8wdBjI1tf0DoxmuS0T5QcPvwFLOt
ouQvD5IggMS2w2wTbi9cN0FsBlTvW2K2pZYtADAQIUT1HSEm6cKU9uXvnFrEvkTwqz8hWa5EsVKm
Um/2928OdDKv56ddUYiCan27nR94FDfgrWrkKL4o8fdTGA3rOZcj0fAiQAZ8TpPLdHbCYYmptONo
0kKKcKOIPnwwGWrTZlHsKbYi/azgHz/cdsbSsF1iHoFTmbXThmVH+h9c847KcaAydLpjkXeF1vs+
zPLDsNHg81NnL6x6ll7b+TrsmqfEsCnvG8cnEwreLsy4bypXKJ3rztyotN+wKLUBWm3Yh36uolWn
aA/ey/j4vgVWzPRIe5tGOOxO59nygNJyNbnsgaIgOhztitdXoptCiZA8UTESEpWti32jpOCFJu1x
C+nrHkhR1ErMsjenJ/dW4zuI6KmrZWjAdqCz1rvOZ+IAww2fBwqoSqU1VuY3CFCBGLPvalcCm6WS
bwMvFPD3/HZWuVaPdtNudaYbo1lfZFl/3FKXofAeeaIEaJOZrX7HJWA3ToqiPgvVTNWloWiSDd8n
mxPxv1C3T8EIrSjQtibAouOdcjxgcRHKjyVs2J4y7GoRnjzQC7s688JGFrqSeltfVzqLgfZPc9Xx
XE4zx1SHJXa7mCy0Y6DCfwil6CKnzi1GNYG3ZcRf3ttKzzymRPQPxl1W0h10oh1rNaVeBwXTQDGT
1g1DCCMW3dUQgKyJ96xOL4lr5jH/Hv6vyojzQvAMwtcd8z29OeYgSkmde2ysz3fIcS9vcJkKrdtE
gsbEGBN/ngK35Iaq30IxoLA+OIivoQXx62Oub+P7wCvJqaT7M04h5HAS/FvKOZTo/UsWJ2IT2pgq
8/5eEAgEbrBYbH6nsr1kKd9SxTyE0FJZzBIaLGgcebDpFdy3y3V7qdYE/R7TnYKPBG0L44gULQ0j
dOpwkEkSsIZgnWJkrhn3GMeMphyRtYo8nW78QwMIAvO0680a/ITSyrpk8UOEtiKdKovRoHJHFuOi
dk5aTWQ/M9d1e3xKdq/JD2H3WkNkCc6J4ds6h9kkw/6Je+odMthghtIw/Mnw/7svm4MD9BSMq+Tn
1ptyvVlAhjd31p6j1+NJaPH/fEAAXdmFEYGon9GeR50O576CpM7RuyIt491t+lGX1xsEKg5FrhF4
4hdz+tHnyrOA2NbeLvjMOLkVOtj3U9iuyBWyPK7CmaJhdHd0ghnODN7O6nZ0fJLkqPtj5HEcehDU
fFZSLp4YJ0kcMExJn50uY7PpbXDqqpkQ+WxipLuWxu+qn40u2VMPH9Qf4nc8MvzqT3Ko9Ea+WZMu
6HnoG+V/gXX3tdTUoKc0DuBnr+ZNPtCT6CXSaSTTq8w7UfIgsYnpEV70lwLXYQ9MygaN94zTiESn
2R1+fWUiL2iK1vVgo2jzgfpEMv8UaPe1i8oaAbLccNHGNvL1xsmWT43Fb87kddu6enx2enRx0xGp
bKtXZjkBV0XdiL6wf8emhZisNsnprS5sBRm0pIvzPi0kSRqZ48mtdV3M61ddZnW3zSohMY5U6AVG
tPmFcLkA0yvb35hJ96O9kG/3pq7txZK4l4piS8BOC9B6iisS+ACkh6beXAh4JuUdk/uXNB7Jj0Fr
McRXRAFkbq7vC9O6IlJ9M/7jYCAGghmK+DhtvNwLnyW70DwhwSlFGBcbM5pimMVc1LKzWq1NrkYc
oZMskqogYW7okLWBrSGK4m7DnA2gmZayfzmM7oUuc2FmCoig7fqLelCvP48sUiXv73yP5Yt+BRRx
OigFtxYvrqNtnuGFYtZgeKIGSr5L+cCQhyWpoLdpX1Q1Ul+2aKgjZ+zuOmPu0uUnkkHgGurRDwy6
A3dEetDyQuyK9q6AIw0GuRkXXIbfp8aGi84JzuD1cd46AEa7UIB6r9EiqKqxKePSGEwd4PU8EuAK
87fWIf06s2YDZih5ef+wCTfC6lKPX1MlJaTYkJoZTaJeCESOjL71p8iUyEOetSpn8dQfGac3XlOl
jQ4VZTfmlTUnIdDLPh6PGqiZu5H+I6sFvP8N8Pm9F3ZFXSjJwMMprO2pMgjC0j6QdYzdMApnn19Q
HzlDlRbQuxFyuvqkRuaEZWRV75m2CBoC60vjxUse0PCF9SE6Wjhza2fJ/wttNTHqTKbBdQUFpyVx
3a/aQ2ULZGEnf6Gt6vHefsLlFsfHgyAjQf/pqky0tFQdQffIBLnoooj0K3MMeHgxwHuaYQEw7BYA
qD5NxPwtr/tiAfYHtUMuayaHnk8GPdZAGa6PUj00YoeZotVHWAqkucTwV+hzJNa5FqFu5E8Qmfct
CKmy1ck9/fKsaHwVEJzbSi0sZ2H3lvsoh7wlffO4UA6U8Dn9zIOXScXCDbIqNJAjQ6nYBmsz7JXJ
jfTBWVY/o5pARfNtukvsjgfa2J3RmBvXNw67MSJpRL4q7mMIvq0O6JvNZUxNlTS44libpxiF8E2n
SW4GzFhhlcs/Cog8v0mrDQrI8lQL6oXYaKAxW7uS7RknvIyhFJMatFPvQ0qdOd+Gga295pfIXO7y
2OjCWyHVpj8W8Pl1DhxaeVsfTERrDoiEjTChp+oWMzk7X69kNMoGgW4iFiowz6Y8U5Us4JzxfqaX
GBW/2LwHVSn33ER3VKOCWXw2TFWa43I2AegmHgriH/GRiu5oG3/lS01fvHRcBfeON0Yy/RsYoYQc
NNvWOEo9JdRA9yZ+xUCmhCgu12waDR5uEATde+N86KqdZkCyUWZ4agNqbxHbLWLO7m/JalSlYhfD
1l1mmIZkETX5HCTMfMUNEP0JOBcuVxqkSqcczzDCrnvGjQ5WcIClRYGiLE9+fNo1FmhGrTl3Z+7q
DApV1KNSjugIkNSMUYETKXpA/MmlF10fdqVNr2Mm/Uolzg02Ry0dDNJdQHpNLlom/vd9Go6l5Uci
JnTVMhiPMZblk5RjgPX3wB5EQqzd4gDUUjF4WV6RCP38fpV0mAVOHFOpnzyNDmOxWDH1Q0avUTjn
EN6nfx8VV3UmgeP5oQXcGyTXxYeY3eAMOKiULb9QpuwJVuZoUjih/sH1eSes+MWt8bgNcKTFwyCX
kdEGxRiJcWvZTZ412jJGyMek/MahBBDKtA7WffW7lYU2r1jRggKd1oufM+gkif+2/XvslvQunPLU
Ynydi0k+umxwFcf2xdW6UfTfl1uRbzFtGIpvcBxVYItBuUHycLdJ4qbLViLUCrPHeDkKkA1kWnuU
Oa8j4LksP1m7++xs/yPSPKkFJeZNw9re4DzCMATNqYAHEIJRuDOB762vwKsorneH9uM5XYMZQo9V
KzcFAE2K0sB1Xdl0sPGpLfYEGqdd8HLvL3VEo70OJ2dWGoJQyjREOdVQy4VCfujhH+MZUTnI3BcH
1TGpDTWnwatJD97PJ6v9ZDkMxsOyjo9vnynx3glIKyb7Qsd8WpbXcfEwNph5vd+QpA2NS14Fzxm1
172SR5up9pGVqypRB/ZH8qjFonLaDrCXxvnvpLMOPx0CmgEhh6gTe0juH1o97Rh1bjAVPBYSoKpM
lzsFUMEopL32h/56sAnFs76QCG+UIwx0W7b4tGTJSaiOuid+0qgUra2w3P0pE2ErOrfVotxIqM9c
wlv6Pul2iUywE+kUAYNSMIR1Rw9hVf+KpvJkHmpiOp/XF2qALzRapSoOkSb2vyEMrb7pSyjJSGyJ
Rv/LLXvFd+BrmvgSGjgH2MAK/m5Qu9hkGlsPo4SOA+UaKFQxp9IS0DM5YBlYbeKAh0iCCtAkDMD3
wQXwQf7tnxEzkRD9bB45ghiAVJ5hqFZ1GFXd5N4twZ/ffbnC7ef+FtEoHKxnTPEqniXtOhobLASx
RJfWNf5cw9LSFbg4sE3yCNyK9WFIMbPLSImDEjAAVLt9kw6NYA7YEavmARcTJxo2UcnFeFtKAQD/
pIm8agt0dXiThjMo6TbDPsmnso/vYtOFuxawxXHYu+kT4eoLJS3HhI0U06nrbZZz8rdZxj+ji3km
1rTtGjGhNf0x+nZO9n2lK7ruJl9tJeaztv3z1WS6G49aIMvwU41x2gOYBZW4MNljpPWD4tFB8UMQ
WOfBgQmBYlsnXkUjO5Er+XWpQMjiIq/zixvEVXflLGzoNxYxEtuNCwmlrsTAenFYk+6TuMlZCG/6
kMnakCFUFt7K2elVpjPjl1YfY4y08yMipYZdHao6rjMM4cWJoxMT0efWy6f3o/R/4N52SRpDApFs
0Ltk/1CuDoTApW8s6bZKRABYzkf0kNngjvUweK0DZ5V/dx34IzmbI1+CgpTPmg5P8tuBFV8EYeHt
SK0trUXOzEdG0slYzjsZjGzLBKN2Y8O2uTdZpAFFjQeitd0RQ+jmnXS5lolHbC7u5mfWA6HiBArv
UZ6XuXm3q2VY1puK5MxvGXK9HbWakNH3v+y/eSgYOEO+4CWXTclBDU6hKhII8/7qN6Duuz7tS6V1
y/+qpR548t0NGuBM0WQsEJEv/mBpD35ZxFA4FL0Q9VGmWoFg/woionBDUPAyNSvklvCV/PxC96Fc
7ImJDAZOQ1hkrA5UWjXK9WOzBaCvEKvhenKA0+6CbrYiX7lcqYEjMhV4TLhCPoMr+IQaQNFJfeMN
OGfC111gQBQFNBmXMV7Joj6KpaROBV3/ZU7our+TEVFAWQhpm6DCcQn1uxLcxc8ICXUKLQsUYwu/
8Y1D6NbtvC6QO1VaP6/+RVttlaWCULdiZ1iKMe0NPvcb/+Sezw8ceuTVy7EAwJEt61sIK0S/pO2d
rTy6CcJnX6UXK0qzvDoLUg8N8Tg0+l8T8qqFinnR+DsXCVIHOjI/r/NadkfzMzjvW8IJ1KW6hY0x
CYdwZqEAgcRJkPLq7GS2kIrkItXqKi2QOf+hGJnrQPPUYRLUByL6/Nk4VktW6mQ0N2UlKoT/TUGI
jjopuMPQS1PXVzzcKkEE612yWjVnbLxndlUZna9B2plN5Kp8Td00LqkNwlF5RmkweoYIrRIZUUXx
fyl2jfI41x2Q3TBRc584kPROZ1Bso78i7nzB3Mfymb/nZ9tW0QWYouP54EXH4zaAwsxy0vWXHouX
71JeMyBXrNMq0HXShUK+Ahyo+LMEK5AhEi5gJsl+SDHpBP+/0acAdlAI6UTI5IqD2DOdrbnJyFWI
xiMDf5HQi/nqOZycBZgY7dHXw9nVKD/vj3N4H42jQRH/sEg/Ao1HN+wr/VWtOa/j8ZC34eWDn7c1
VdLELHm6YNtjVH7HXKRPLPsxeTBdYjwKhtwCseGI4oVQEsipbZxgxn7P3BEAyW9N8gMByYwAtLUL
XsEwbwFD9aOyylZtIwO8OATo/0MutQ6QqV9/FwPB02WNIeIXp1DEoKX5FljQtRbyKF+nweHJ45am
9NHRowmd9iLV4QF2Xi7NACZg1Hih9EDYNiLxXE41Of+xG3HS8q+VTjOSjXF0sOWT4+JCoeTfqkqM
Pjlrzl4YaoPQmLbhfdj3sxZE99Oo+eUqT7xz9Khy7dJ2vjm97xh2vrv5VWEa5SDckFrYAHD5CfOa
jIWmnv+8o2os6wabwtuqJWZWncMBPO59ikCdMIo9Kd5MmmkALw0ovRcQEv54ZvengoTauLjjVOCV
OzFKpovuiiUF5tBMYXbKPF+WU5oUmQutvVt2Xm/W+0fUkCiT/M41t3bRu0MhChC4XlJKxJZEO2yN
JtO7Q6bQtf43mgNLoujYyJfxeawVnH/q1jyVdI43WkirUxfLMYiol403K3EEryQ0sxUZioQcjNFI
qYhhVV2JUt30Itsq6ibXSs7PFqaP4LJh51/5TzU2poFBYvepHREiPek4RDStzfisawojAWf9jTX7
HVQaFmFjnUBX8Jg0D59L8ZKUcRLJWfX+SAmMydcZINdEPKQwHSP4Q28Jd++LVCJhQ6/D/z3XC0WY
qIVmYiTr2HHxvhX6u6EpeYrx9cmtSrr0zVPoEFBMOW1+6Mc4Wmz0rePvb4GU03CekT6FTOaLqY3D
flR38JADRiarpvNCDE2p6rsPvVBWJMbabV3EqRHO/kRBybpIRuaDtZMzUVopRQt9DVig9eaYm96y
jtxrmHGlT5YVOah5xek8rhkpmLfOh+9TO7jG7jJOIVkH/fJrRJ3yE26Dx4VWz3PlO4iINbE+kwCh
/Ezm+XmF4Q6uVbfaJpJvwgraEo8ZJD05bL56L6qXusu8tBkoRTkC0d3FrhaqkXkEn/zIWp5TM1Wb
GIcOFaTBnCVtUpmbCouzh2Zc8nA1af3/FABw61L+CTsJUhOuPe+QJjxALaLEPvmeY2i6i4bO2kPX
sWR4WDoovvXraNkf+os1iNlpLxgi0/0dwNHL7joX5nJkaHSB+5s/p/gS1/cOPkJysJUivKtrtO5Z
cKBAhxiFa1L/u8F8mnaIfdBsoSTIT+NUPAAvZU95VyOjDzpHc+0sZd6511CCcVOfx0rNGYgVXTSH
HjBCCPpnCGDPyoWYdgd6ufrEDhZNOS46uBSB9FQwi6iY4hyxuJadv654hKRKMPEZ8WRaiQJsmETa
IDnjFooKo7r1CqLFlIqGpraYGnoWk7K6051kY5CwZ7zFUpoM4Ze+ysTKt2+FqEUga1iVufBjCw7N
8Ff0ZfGLBw6uRytHU75TKey5GIvoVVwAGwCw7Rytr7DoUZckWkLRH7HuPApyCoQS+IBxb2qhFIFu
oIq18crgYaeOcXk+EY9OlNYx99Jt/8O5ot2ozyzM1sYGA0nSHxVuZc+mv7ti8LeJTwMtuKnasISP
O4kD8r3Np8OIoSoWXZ/WDdQayDT4eza0mSWTsjPL8z9ohz65sC67P8H3nquUFgB4V45rhNAzsOeZ
yG7BSXhDOPnn+C1z0KiZp71jCzI95dsEhUeHgxyYGGgd0EP3o8wxk82QvFVe5DcOHbuGPrXsqkgN
2O69IWmcDNU+2iH9CY0pbUwp4jFDNgJdejhC3/QDrKY+bnDYeGy2lCPanK4nOHCxCjk7T8y83dIC
PMisAsL1/2yW1uZUhW5RNs1WWzPCb2jESfejApSRDDQDVabxcjq9tpN8JxtJn0C9DaTsjTeB7R4l
QmL9BFIKxtmWJThGJXu1JoINSrFF3WbTpWKGU8AxQh5zsKLTMfcBFbNZUw9w3HNqC0RKMoCLyQTe
35AaqfIBiFNhFhU2wN0ogdV0Jg99JKicLODpSLJI10E1t4OGSH5xN3obSnxnk4cQgU09cvpmUO7W
GABFIYtxKo7fUSlYGjgqhmPadS/RLS8uYcnwG+y9Qn2ni9OxK60T+8e+D1nVf4AMORZKS+hbue0h
Z7lkyyk/uR5VKWpDWGdBCIgDkgr9LHcETtJl+ySFW42+jzzzAVypRkA4SHe4MevtL8yzXu8gNvb+
Z4BWgemCwCWEXX7/GidUh2jxvpGFYLXrRfNqzbRhIRrMsa5Q7CIYy+YoDHcVwIC+PB+RA3ssXbmF
JHv1vpzpC48qQGPbCo5WtVnWhlZgS64kvLPHTogU+Q/rMxfCKIa8uqh1dBR0t5H9HsQVhUmQmRx6
fgkvOaJaWq8fsgpRObtQaN1kHh1JzQxyrzG8i1p0sg7OoBAE/RwHO/KlJeK2exzojtoPquU81ezB
874HIZn6ifrYsKDUTYj7e1qk0/lVwW0sC+m9i9DgezFs5m1I3wgkrodGxe9fPBc3TSPz8OWt73IO
oWjWSSbGsAs7M8oz6efPQclAFcor+solyRvgibkX/pVC+kjJ0q9ViufapeBJS8ouwUUittHBdSij
pHWzEZaqpuuUzrrZQkmgjtOGPxC+vCdJcltIxPTPs5/G0leX78z6xzrIw1/tV5S+8nRsDjhH5TzC
CBcCHhoGmw5T1NHoftSYNfW2kw3S0CSKAH8t7yiw3vvxW3KlJAoMCwqwwFQpjvQetwfi+skiNLmv
rhAXVWQQXzud6IGKFcDWWd3PDzuJJsR7PrB/22s6lYYnfTvNOZTKNegvQbdKwzHe2o4hcY25LY00
CiIbZJ9RKA5/ECd9HwLrI5WlL59wBqQYNUKL5/BqhM63DnEoTJDR2kG5gn4ie3bT+8S1Ne7oa3xc
jdy8wQxImjWA7XHJHKCcoTlzMaFiHyEGEQ76WSTTryIz+79HHItmTNaO1tE2qd4xGcwHHHZEcxq4
ry7IHYnvFegqGaNSSvcaYjYiqo2CkZcwTyLekQa8SBIUH4l0czvKmMksIFhTv3J/yOeQO8gEYUk4
K7/1ekvYWhKbYk/k7GuRHfY0quuwDA1VrJY8OTfAJihg8Ith3205NPnDzOwao9wgIu2rthkqSl7x
/Ijp8+AWP1o1XrLD0XTirOTGDN2zflI/iWzSlJhouephD17t8xzthPVgQ2VI4PrrjBAUmFRuqVIU
ILRh6JWkih8jtitkZqFJkr0wxuWPEpNF1KAQKO3vlOHcORVtqifYtzJT4dUgALTsSppHKo284gT3
cCl2ma1JXNr20a+6mPYnlaSf58mATK8t3VU/Tvg8uA1m97e+FAu8P1eHsYK4aAD54YjqOSpuFxmm
vSy8nRG3w2/7pWZKh2JO/7BgCMdDwdybp9x+HwXfG44dymNAghSOJ8VYxSLH80Vnkq+IRZUkrsBW
1qF+/QZ2PFGhyJCFzuW5py0oU6o1SRAfuXc+YEYGtQzDEhewG4eeC/e0ItRzOjEmnWB4xAYbCsJq
3yUEPOY0dZWO+jsXEdvbpU4pFA0yL4rPI6WMRaOImRLMZuzFtLgJ8JWY6Jhk8QYfoXYOJmsSHYJv
8UDeFuB2eDMpUQeqZjFuHND8nFDodhiC4UaBfCKxa8b3066se2g2ou0lgql9nxEJ02O8zAiIJu49
hot7IdO/oGBuB6k9GlrXtS71UtA6aaN5W2mvjiTw2fvNzVSTALLQv92UHh6p58nQs6bvCLv89GYh
+KzAn7UhcOEzE1VJ2fqVe4XFNlkV3MDv//wrmYB8hlrfi4Cpi11WjqfCj29lh/15xvcs4DxD0yCD
zXdF/7ZZXiVX9dWd9QzxjvFBDFc03XcR5ALHBMVi16UkW2QDU8xKfDZvMSpwXk5AQuAJ0vWq6ATx
kkvbMdihcrJmhcEleTDRGf9HIaA+Rwm7S+6jb2/W1icU7yy8Gwow3seQdiYx+xoVIb7+K6lzcAoM
36WfCh6ysU3ZELP2VuEgJ6ei7CAUGBFKkdl+gKkbLUx8Iomi0T8UGtccf89QbYkzU6b3GuGIENnR
vucESbsmPloTu1g1M/kTaY/qCdt1AZ9Rx8/UOQ0dbeI6pncG/6EPdxPHEsiO4EBAzznwT332TTGQ
4zhag4G9LySTB2MYkCAX6TP0tZf+avLPJQzLpaOHQndtJrtOdOBmDcBDhRDnknFLE03uGLpFc4bs
ojWibjrb+UJ5Vz0WhMBaEwCUhmNpJLaCNm5ZaxI1Kv4QtrdbcvgnrwIZ4IsfZWey+6Wn1XBB2PJ9
eR99nCSjf4tcKxDHs/ERfkP244/PZJCgK1Ugde7sH4EBgQWexPaaP84tjPn4pN3v/3TUFS1GMeLN
GjoOjtcPU9gBJ8KwH+FbnWlYgJr4uv3PWmbm2lHYzYoxuR5e52/24RsFF2uMxaoFkQcU1eT5KRRq
0SXBp/CgLo74/WlfapAwUq/m2wWNfiRHptm67F6hp7ChTQq5ayxGiXYfhnfQd9Sf8lSVhAt3CugJ
jZiMEG5gtUzQ23hT3KkrJLt43Zj5LT4+Hwn1fxQWuOvmhjoYMYfvJTIy0Jt+vBcv/nDT7V7D8ji4
pCMtdhRDOXEl0DEhDbQ+kzkNvu80OBD+z97ygOyrzAXGyZFVjQxrYQ+WhMANs0DhETqIxCbwN+I6
6TCPgcDTs0q3HOaIwNZhEz24sgg4CjFcTIyDGTBOkPpM+M2qXlb3nc4t3guORmd2n4E1WwsFRlMB
fEP1nf5rrtA1LeNYOmEvDx2GQESbpwr5FcT4rbxJpCVSwHSg+CKOEBqMiHicEL1TJQbymwBFEEbi
wsGxSWtldCLApc9u4GUMyNev7xg4LbKYb7McfPIjja9Hgx0OHxywzHY4n27aK57TLb4QSZNKOxXD
gcl4dyw5OWOLGyaTUZqnu2gj0NvdJHAMAoAbC0Z9uVdw1/aCVd9Slr5EK/IbgVkcA7oojMuRxJKL
3gbiSJ3DOUtR1mnzXZ73j/NdgH36BEVZNH53LdubOD/sEDA5Rz3dpY3Gmuq8IuENE4wPm+j3utUh
N9s3o8SNeKxoFDiwcdy9CF/Pfv1ddbBdMFiIkl66PwxwT9Vdyl6tu9SffCmK3nSTVfBYFEN/Lgq8
w/uvnySbESQv04ckee7Te0oC4Srjr1+B8Vv4AaNsr5l8jzIpTgpcQZvNkAiPGM5acCBWKTAkS9Ld
EMh2V4060N+jfiWRIVJoM3ATmBvxnWH6SN9K+B1aK58xXcx1FTHelsHe+h6SNlHHxv3kRQSxAvmE
bEXVmwualCSLruESATQ6tsBTOSkwcAcP+CwbnX3GQiHxTChkR7NhSf7aFP6QS7B4NKYra65EVB9f
+3zmOwykKn8FHb4FdY1RT734MkFHUwV/UIcsfxGVuo/WGuHkeaUb/fc3jpE2MDiCCFTW424uvPYW
P2T9wnvPLQroZrDADGN+f/S+GmabrIaEq5QfFGi/KzUisdcomwWFF0kp4WstQYxy18ENF0axH9Gr
iNlD/XqHSi8sopJ41Az8FrUHxeHPJiTElebH759KnCU4DjYWWnh+jUiKqNCRxbrYQIH5fOuYen7c
LTu2RWn/P0L3hzPe2M7rDf5Hacc/4FTpZBUxc30Sqbrv8bjh1rhupfAHBzxSEzPZKmMYdy3liqAM
ZA2LiPennqIMGGkqCkQ9PL+MYZKLXQLGSpGl0zriGsk5Ew5K5XV3fsaq6eq2lj/qBVCjUuCzYKLb
FKxD/C1xMH96w1z78LRiAjic12xeYN13W47PYQAp8BZocmSDEsT3dUCrbKJArc4fEIHs+b4FEi1a
MsDSzjyumvXiYrga+KVCePa2wDKaJY6l+5sqEj/W0hGaMUtNKG3AGmqXgt7uGQ8b8xobOyQIXV65
ysczbv1OPQQkQ9Wvdh6QNw2bBO6ulYIFb7up331QcN1EoME3T8fMmKHQznSeiZphJ7KjpRmwqm8Y
MJc2ioEnXaz0IvKt3Hgjw3lIGxsYpTe/T0mGZEIoJoYT0N/GkQbTSYV2SCrDLtBrfAQF+rGGgxj9
YvNaO4PdSJS+nkI1MSR07vbJ9y3GBWu/iUMoJklfMDIXmDGFMC3i5yw+bF8fvOscDkYo91/Yw57r
1BZ73CudqEhLjxBvM68jyxiMa6UdV+LA9iaWemPSxzyTYSuYlezuB4MZLZfYBk4JE/fDgQ35/If/
ASvV0j+IEjEIkQpxxncf8sa5vtwHwUmi1nA2Ov2jTdmyvl7aGu0M1StP0a2iu7ZYPHcxCgyhlMMw
ce90zapZMqcffXtB/nYnJ5c7+dMegvreqTi+dE6h5a4LzhebWRg0+azYUZKI9RyZxBqj4FJC3QBD
GE4ySRw/u8M9aelI0Fau/haoHD0DGHYuOQcFENgcCcCXcQK29GupIBt8RF2ESXiM5R04H1dp49v8
PiTlh7a355HVAtg192pOUH10RGiwcM5zXN/pQEec/XGgtTzCPoxlq8ybBjfh8UTSQxNin7/bW2Vw
ltLea7iEiuYXr3WCBf4W72pHyzA02WdagMEsNCgHzaoWA1Qx08sJrtoX6UjJpIBpSnQfxgMuOPAz
Esv7MGcrX5gm/pdqlJvoMPTHcU3ROgfuIaOMqagYSqkl8nqJULXayHPyT3g579UvLChcetiZwGKd
Zz8YRapl3+LaXM7yByE+QfH+mjU8oPjFBPW50nbGzNFVucN19ETkAyBs5rgA71yl34YfNfJf9nRL
Up7wuaqwQcg0Ie9wUknjuplUGh02wFZBYaIKF7v1hHflXvRuhz28Q5xz4IltYhycuQvW8mmjWWas
HQFfDAQcXGFdYyO6jXCAP+iguk3cKGAKhSsdkB2kMi7/cJD46+r8+fmH949kzbg3kqom1uj6H7R3
tEcv//0ga4kDZQgfbiCctEnRlqG8EhKcEhx99BVYUYcRUzKJsZmVpLAtSnb1v8QLTuMVwY791AtL
3k/xlv3+ZnqAPpoBAyyQfROBwm6KdAyiBsC0nDWu+E+EFDqimX/a92kU2vg/NHJSHufitFtbcCJW
6s+ilBJ0CFvadF/5uZCZEKBTMmdkZByWmatWdtpORbiv1Jqglavppyz+oZlNtMiVvit+9io+fjdp
kzwP6ExjhAXF54v4FDZBdaefQ6Jg6QRVWXscYoClI4DkBH5r7/9uQO4CPT+W2e3RpHlVOucCrHb7
6XyAPupTvPBtQ4dIyzphSErDaDR5rZsglu28hj3BWFfoX1/t77+ljT2ISYQQr56wxrAu5i+Qr/nl
JsEQd2p6l+3E3lQ7z92dKGvGO6cO8zMEzbgBwB0QcyhPeCTFFef3nOvaH9lUv20niz2jL6PmhMr9
rgfzSj6Yzp0vF1l7V0soMlaCzIk//+bj1QAAIINxMaZT4wupra7YePjyemjNQRmMMckvcLATt8hQ
NWderslR7SIuQxJfKMHz0vXhVtKRtOqCYZ79vqxX7Qm1oQ1FXkBhN0+sQADQqmT5ctkfOZnONoRp
bzDTJkx30hE3LUkrpYnk6rgdx+6KibHkNP/dk7us4t0rPLpTdGfa3oBUHbKt/wic/g9U27h2TdCl
noAImuN25anJh4BKiCyYBs8h3AHpSEcsooP6PQBsr0o5oeReS4k92mU8bGQaVtbJi2fU1vqCarpW
V2vuCwIvXDVbL87O1KZ8TQoXAaT3b/JoeqYWj9ylDbeUazexDNBE/WZxu6EY6x/E496NSICTwyCM
7Gg/QzFlcDoJRIv17r7T0HkGS6w2CrJJzwwq7lMxb7fOV6eiR4qIIab2Dr6gb/8zAPMFaBJXQZeN
Vqx+6vBBYXFun1ZhNOhMhjXGFEbJdM508Ko+KoWkSda0JhhEg1rdN2J/tqLCAAy1TXEiQLUMDsDS
JLFQeEp/i0q6dhloDRqWjebGVXPKTwXqe/LFaZz8VosZU1R/5Oa80fr3pSIQoxcqlFHcL+FQDqnA
GGDToU+9yYSNiuezAThvgbYONCrEPzOH0xS9H1KNrM0IoBUGSuovFcn9bGmyjDNYC1KC8+28pUIP
yzxGorYPvgkiTGp18/Rwhnq7t2nsQrbuPWabvyoBc6k/nZtOdhk5dSjT/uqggiUitril4HutfsmI
ImmtClWW0yvpYTEGYAXsMl81e+7dPdqhd8gM0GYrgLx1AE2+AbIwOGAsyQpwmYhvpv3SfGkHHo2a
OAi52Ba315iQvIACBQKcEGfiF6NrakceEl0RxoasMCfE701+OOpRiLEmb/bDwpLx1XHQ+6w7X2n4
lKhFjDDRkFsTOveeHb8rG8+Q5CvhHoSRHQaAtdyOTgMbM42io+b/tci1K0bre0IUw/X7bnImbpZS
bISxkfnmq0Yi/gnvDUrqVeFinNHdZha22B+Em+HF5/U5g2vtfqHmQUfO/UiKZhrJFAXr+WrzzSUx
w9nRnYA3lAHPP9QS4l6r98ZHDQr9M97/MFbqYlQ28A5kmeE9dOB1QfoSOS94QD1okLxfNFTx01Zm
OtxECM1muaUTbjBy+GJj44kgQ4efzu7YIYYxAH+HuEbOY+kQ/NowhwhEZojtQeedPtrYtYq0UAdp
gVMe9KWX6BuaWHmysvPvv4H0NqaG0pmMDQHDWUdmouCmoE+DLzyM2Zq5sGSWujOrRsUA2xUtEK68
P69zVvg2ZzUq+BBC/MgHlNCvaXmcYXRhs72dkaQFeBjEajAyzev/7ZjB/0MMXo52VsZgau+n1C86
20+t/zmFbspHRQMjmIwp0/Hk4Z1sqHHwk6cYYoOCUITZtNUg8UG+AmRyoVpc5bo7KyJvdWlRlQB7
1oMwDnC/cvZl5gxBufUiPsf4M3axitLP2ZW4RxSV6eBH6Ty474jL1kvW1AHf3x1yETOjPeJXzoB2
MV02GKF5nR4/+Gk0jmwraehvSxUjRw6f5sklzSzSj5sEHO2inmwNJYwXuBp3xtvKgW/nzvZ/W/Gh
Ii9v7Ak9s+uMInuUkn1QZRNum6BN/EdFvk+YfZoXcz9QJMVCYokgRFHKu5kh5oLVPdEkVOZbQzpb
zYo6cgrWB4sRTaVvj4q+pxfA4XnBdRZG0AJz/PYs5hcAn0dFbzmSKp4Bc78vczFK/s62ehdB5tiE
7z9yFYxhaEeVBdllRS+7QNrsnQI/FUlqdyn67eSUKQHUzd1CCpKGlYfqm/KJ6oSgY3CE2h3/RoA4
E3l1lHZxvJv3U/vaukdVVhrFljd3p2WAYZYd2SVKWfadLizXlObVgjkTziYvMxT9BCwpJGdQ85ir
vOPjfz3LKA+5Uqm/NTK4d0B93jRMp7zkKsB5qTGrNa64xmeB0iPaoOzrPjy1jREsV/4uGES8grfB
FUH5xu9HtwCFrdVIpVKdm87HCcz1lfg1OsDltJRG+X4x2noewLOYyQ+AyixjM8qOIVT7rWUC4qpQ
n+zs0jGGYnsKPxJjKdUEd2sGCHcszsnRBRxl7RCh4UEzWSZdpULn4f8p/Ll7wmuoONvGXDg3OEkM
HxG1YFoVaPHSYtC8ejP4NWGeZf8r3FPcsZpqvWhFmsIfXLoSWZ7tHv926oiuirj/A+D+z7vY2uRv
/LbhC7nhmzHIxNXhzKdykMEdLTww+fYfiwBJYAw0NqDNc9Pg/LV3VHy9F5flnaEkinDkvEBW7Fpb
XjOis83KUxl2fihaLDPXnrskmnFcNs43xHDpCmP4f+8T4t9EsaZCXAgSx2w265wjXMOe+/hxsJa0
3tvu/sc/UycqjFdTPuVx8MLEGdjiUOenD28ugYzOlnRoX6lk/VWtpqOymOyHZZ1ks8+QIsigd9QL
JwCMYGLAekj5xWiiMNfib/HAoRxuS8hCEF3PHbY5DHAJ9wezYnKrd07FNkCTrUa8jYaX6GxAqUtL
3rH36pAI9aAv5qaXovssGITsVctCv841Uol6Al8s0SJ47X9QCLMxSxSqsbVx+3Li2aGBy/qDkb6A
pwHDstgOQRWp3jEYKIm6hSyF50PRyLZXBW1vUr9UB8TfeCtBJgN2h/L1Cw9ZZTmLcWkEHRJbwmOv
kW5wxpoqWMX7LlShADnpd2QhsJb5ma5I8lXCzWia8QXuZF5cAQbAN/j+e5hb9vs7Vqe8NjC/1CtA
qu/uBabi7I+sF8+TlY92MY+iGffE1z1G3jKy8O3IQ2JPiUmbkEVdjO/VWQo+3GuUFaC4Q/pn3iqX
DxQT5f2+bEVV5Nzn7BcV09OBHyu/rZDszsnb/CPHjWYv2MiYUOis2HQ7wTm+nK9YMsef77PUFi9J
ywQmCDUaFCG6k/vJNaXT86pyQ8pZtmcmEZk1FWqP9RvKpUwcnLNPbtyjGNkTLff6N1tz6jAQKini
xQj6ztDqsL8reZq/FU3C3Fz4IhS1mti4ZDbsw4R3XQ8kwmYCzvs8+E1ShHCBmKuEJYtXZOg1Y0MH
bVwxp7Qk99zGkZmO9DkM3ScyUM/mHyWk5H3r8ibCr8SE4t+zXdGY7/IQxEnkvJEn5PhvKXSnyP8L
kulkCr1SG/6W3oaQTlcmdBx8+q8go+A/7Aw91PwkaB55BdswdXkZvg9hYB1V0FLitD+aMUdCP/vM
XUxn421Kf7LBaEwA/JiCwyl+vzFxK8u1jzyEQcF+f9QfnC+qmGIY+ub95yTlP6aUc0UfXvrDWmLj
FJTFoermxpCYCsrUp4vChO1DHJwggirA5ShB1fNEuYtdisWHW4iJVvAscBYu7vH5SXgtMmFB4UCg
tRCvnr4h9ian0h+cIG3XIEp2aSXS03+b+Aj7h05XjP+ukXz3Z+3IYSucNPNu3ydC8F1AmhPf87ZN
+3rv07kyyc7tflTfhJoWOcDdcCYNiTpZWOy9LJ5BMdyco0ymjHGJxbUcMUc2x3/okprYJjRRF+8K
leIKMprjA5dc0m5l4G+ZKXiWI4ilz2/hMI/DpGJUzT6qkxcfqzMyjf7pv6CQzJJOfS+mDaixYHXt
Q4AjU8d9vKv0+g0h8p0G8krmyTVKzEvZnGMi4B5iBiiSZ57fDslcbKV9j1z6BfKI+nFA4ayv37ff
0tleMylbjnydy4O/RzaiDLb0Vu4JD3OQBVzSj5SKsznJYj7pTrFZIGMXBEDnknW/POBJFdzgKF3G
67ypHnaHUUswjIkufkj+5B4M6+j1ZjSui3noarQFhClhkAdLx80qQd6bLhCgJf8P67geYXxakg0E
V3hXnLV3+o7WQ4UsMpP7tgLk6mOIcmImBYUH8d9nAFkvOmuPBFUJqsXtPf9Dkn6QBHHhwCN3+SzC
pALnKuLvRDDzyIcUKgf1os6fxu/Z0QlL0+UVtQvAE0G7dqMofGiScsi9w9vMrKGqYBjZnU6dIEcV
1cbjbdrPqMF5CkFaPmfon9H3kTfHJZTwB6NhhmyWFOoK/KlHxp6u1arKNtwaFnwFhojJd7PkjIwt
jqQKNFZqzi/LinI/3DR3BPybM4GF08In8CneyM1t1fgH2CVaHUUM2ygvQupamdvELzuOtcAh3Z3D
pIYzSD/+0GEGbx0XLNIUhaqLT3cE64jx4IbXlEhVI34Pu46yBSEw44b/YudvbHQnhNMeWjS0KyrT
Qr8FLxXY9qvSl1dw21ER3Q22Z0Wg1wrEf7Zolw3uLdOH6zjOFpx3R3HPlCpa0vTwlJ6Gn2WrAjmb
miWlXbjvSUwSB2gHVqKJrVedpQ9kHsCbuFi2VrZFWt2SetigeMX+zxGj2baJOln4HeHPDKxg2PMa
suq5OlijXXNdlx3PFwHv1TDhinT+AA+qeixpGIjuoR5HWE0jz36X5ofJGjoZQ+K1US/40e2aYi+9
6VtT+JTioRIqZegoxSmQfIuaGWqo8zL/Nz/vSk3JeGDGDZedWBpX0be8Q3rYt6BBpJF0F1ABu6Kw
UjQWjmqz9usfKhHqrwRSpijpFzsb/c7bfAatJpU2EAlDVjlZQQLekMqbHsHwBF87x+NZVh/INkxn
o7LnyCshN1e23zcAcXWYi4qGSvyxMBXFGNxcX1tlCQ7wKBWA0qzlW/FN0lGqZiZl6k5xjkUdATwx
3H2fRg6jFT6D6MLdfAHVxWNjFfoufxVcVTlFQcpyvB0JP4yNHwGuxvsKnN8/ZzEWo1aRAMZH40sV
Z6Cd7mB69UVE3SsicwQWoXy2vOC3ad6F26g8Lm4lFjRWsXnI4czutVBY3n7i+SaNj1a4NzhCEvmz
EgZG6xBb0LdNLL3iEGHoGa5gDpQUnVokhswo/wrbOu6Omdvz/KnZ546C9OJxxAu3gElLeFzkfSS2
SY5t3znLZQYnv5ow0QOYQcboBTwhRWNzFtl+JB45lsumpDVopT1LG9pKKNPaKyNlPaKTfXTj2RFj
4GWjivUROJjtUYp47d+QxouulxdteFdNf5SER58uzxoRaNosZian11C7lOEz4MvwXIv8V89Aokep
VYsZfVtrVij7g34EHdeT4Dl/jpwYpJwjRt+ebGM+oFBgZbEW/ddjXR/4OEvXWKXPx1ZRnFqANyve
tmPw0Qh6DVnGLmh2+EQO1EsLVBaE8jIcaR2G3+YCsacr7/ESHE390gIX8jgplOq1UfE7JmnSao5L
Viw0AQs47t8kJnXme0+jQpJTfFZ4/IGEJXGQIRGgQyHwVSdORTdZFQo7JQGcd2Vk6h2SJXr40/SB
OSNJ7e2GvYPxIZ/gYf/Zfil41rKkeH5ZtmU2CIVLBdvNU/77XZ/TEmX4JQXaU4tqLOggDHHyKECf
lvvdw2+blRBxxQd12G4b982fBrP5njzMdOI+lbfJWV13lJmtjL5uy2HNOIMKIfgdGrauChrAvf7F
xsxXfYEb9dqvldHRb1vaU0vNYsIs+RRKB0LmvSWdMLijazMPyKRA4P77WdO0mG9rp2V9J9N7fBAu
FpB+AOcneKMAEPj4uhCC0mRUdN8efK3XFbYKOkom96o+bNtwpp3ZjGNmVt8KbhEldI3pnrhkgkqh
oOq+9HKhVsF7xYTKaT93a3ytivSs3faiNRLUYl9rTsjbIAZaWsnVCYY6xmfh4JxaygqDYOc4Kk/D
xJWNWTFkNDti9DXyL32PGY7wm3Vxchy20Ib7ir5PvOE4TRy3IJkR3Kts26Y/M+pGd/inGrQz1HVZ
C0dsa59XOzrZI4C+cLsXksJcK9tfaOhEPx7PKRmV0Ed9trLOutQhYYShF8Iw7LVDYEOgIvBdMed9
QGkcGNCLIzSD6SXycT4CHGoejuABNA+arOGr/ZdKUAlCkE3RNFyFG44sUEV0EgqZiAoryWAAgzT5
ImK7LT9r75clhixUyOW4ecfq5K68ENsPG2klzQp54f9ws2HRFC78vQ5bFT/Fgo1j9L8qy4PgDIb/
2B0fqOFzX2hBAjrc4EvCnajEsRTNv5vRfnpVOCrjw2D4qhnfjxMMkfs3Ft/AHio2lRkMPVrnOu9M
AftWmKL4k2V/an+px3VILs8flvq0qxb/Q0rrYu2zm728/457au33Arhf6zGwBnbeObkBri4/Yw1x
71S4vbockzrBwwy1di6bmf7s58HY+VJsMpO+wK+RP3sWdUM913r+Aa0Z9CQzBjgQ3qnIn8QBJhGY
t8Q5kk9sOEgRa8srEt0FdaVC4Nvu1OTDmBD4L6iK99cKvSHXHV35q+DQ99kOZyP55I2B+JH+aJLq
nQCwiHrhdBWjZPqqWEWunShfpEm6ZJfX0A+OAj6lM7Djyapi0+MzloR7lIOxYeqQHs0zzolTW2DX
pRi6QDv/IStP7HUNau0Xxr5fE125qzfeIj/cQrfIWOEpXPNt5igdSoF40LgRKYo7SfZUPfVP5+8r
DVpBuChcXqprvSl43XpPE1Hu7VA9rJ+YxSJAzDaDRErU8yjeDeFho0sC84ruax96yVY1w75I4iY6
BjoqtUGTQTAsbnOGCG3lGZ35+FxnxgWBI1gjC7UvqG4WbzRpVBHmUQ3yzLKymus8mYOxibdqkPeg
icByws2IdsyDb5PCdft5uIOnzSeUoIoEWOgzNztCPbuEuxh0oRp/0xZBqDF3ie089rd6Z+x8Lg6L
gHZ5/P9971eK9LsLcSfjtFaUviRP7DR6gG2mRNb281GnHNQJagNRDPKEVsxLoxYQZIzxyHMRzQIR
KpnGSTvKOV6uh2aEFSnrrfr9uPe/a7rZtO1lDZJ7oqZepNpG2emSpaPLOopYhUmuk+3kg9zDSBih
DePjkyTmJzMTnaQy19sIc0DodkdzWFqYd6exIGbTposLdrVkw6DGiQbHZkHclIdbtuQ79boo/XIb
UHO889Db7zGcA7XW42yizidibNkEvIH/Hu7Q/5A9lEeEClRxHWPfP/+Kxf8RNIhA2p6BCTFJ/Z2C
2K8yF82ZA8TU00TeFBpgziBkYb4Q0fEJi3avQYNuyr9osl1RnJSdMBL/S6iOpI3cXmpyzeU9iObJ
vgfu4vSqDy5dsOo7m95TO3qghuJVQo+/LAUB3odua3Xx3d9j1pfQjWsOtDP1q7r8yuPMt0rgZEt/
lcuHOL/YcMZ4n2M2NkXIIbTMpztnUCXhc560Khn+12hhd6huDbu01NEng+IulA+dO+jvgyfQRDcS
he51eEV3EgkQKp6gwL5NOkOeW4+rrjpqKrBPe4J1AfrYNwVVOTr0GBKcBLyZmzPrT/7wfvD8UJe9
UX3SvVkYaf0LC9+IWHXcVm58Cpk+QT5lwNlfP1qGsEDdnmAnGRDBmCbVAC3xR4MPVtzH+OSAL4pV
JF92wH8Jf2ZF5TIG5ZiB3CcICJQpKreoEs8y1ZNC2EueyGayt2Z2sCZCvcWxOE17wCaLzMUtGNOJ
5unJPEIhxffFYACJuCeRUbHqe8bA7RnFdNF+GlH1Pypc+Cft8Be3QgiFeuIglwbRRdMFcxeaPUKt
xzp0hm4gywz6dLD7WBOsnxCYasttcTEkAnOug01naDLP64LPAORmMnwub2bYI7GxtK+zwgiArhzt
vTeahEyswF0wr3swxMosQuFp2lfc8eWjVyc9e84v8PKiR6fZTg4AIxY+PU5whcZTKw/WFEPTWqPM
+wzik3e7RXAzXQL/YnH6z9tvxZQkGgyVsaSctSe9bKkCxo3JPBYbKn/LzZ25gMHt9pI6gvGvntzT
e3dCpJvAplpYC3WU/uNHH5FqicwMg99vpBVKW1wznWopMZCB3ubB4ArdMrfXfWcGxPt7/dRIV1FB
N1FXFPXZbJLt1mX8R/wKCRMBvDjnVI380fQZlS0x5/58k3hXUcRmjLWx7oTByAMcxLcPp4OCv6kZ
2TFzT2TDAlCfaVQGZybf1s2PvVG1KL+HATz+htKLJECq7uXpSlYmfzf9tiJU33498AuXZcRTfBdW
OkRwlP4hUq2V3iNJPb1bOIJ5HguKMpTM707wcbkBiOzsU+bLcJE2hymWEH9PVwMYIicC+X5X3STQ
1WsdZMgT3REAujKBukpwngt8OsumKPM/MRM3deIiQyRKVXfY5VFLAnIP+g6R70bwna/7xvV/X5p1
IuQexPlKpSZMHd4H2asHASSaSq532Kmna/pdL7W0hkrX3AdlnVEoEOZGAO+C5vznAlzpd/Vro+v9
17zxKgaRVZl8RCaht0pYSRzGaMMj9l/wn2YBt8atmbqIokp1mTva2GnZGq/eToviHRFmLwHoO9th
Jl+kSoFKZr1FoslIhcZX75b5J31Z54w16mvepHMIyGyLt9Hw+WWnVYSmAsNdlxJNVVE9T/ii8Sqg
j0Vs1TF0CYeVQgA7Zw5Tp6frwlsmwmnQ+wwT+GjOSDJNQ5JrmzawMRWx+YKOWLzHop4pDnZtzh6w
qytvz9Sby6YJzMdra+UX6bvI5EhcGtNwkROo3xVNzjO/bDksTJ9zdwIvz1wzRycOm8lVXmXUDOH7
BEUQpbrivSe2s4w0nG1t5w8NtWGebJJ7tVnn4tDol2iquWY/OUhrLxvpBKXURAV4IsX9il8m6SpW
UajoYesq8BXF13GXz0qMguNFoHO9PJmHVXIrX84Ee1aP4gUm03RYYM9BxeQb08uFx32I+X/ZTJRm
RuBV5NnEJ4kSeb/8XNH0zYolxofKeWGAK+bwuWP7hY1rySEUsoeZv0i39HuFK79XarHUQYvcmDX8
WP7L+iDrSXmHN/ExrNsvMC3tuZYJILZUgmM4uFN60WL2Qi2kOYuIFejXybto6lLgl27jG1Jcpi26
4lAxl+R05ocXb9rvfOzYji+Zr6d+W/d6PHDvUtOkoU9c3OCm2LQmQHks/2bhpg20w+gv4YAq68fb
ANC86XM9QB28R3NuH6S2nylSp+5N6tLm5/yT7CK+ensT255cEYQSIGJE6AiJGcmK9+0S2kgrZOXm
RS/t8eh7hHo51mDbuhuSSkD7M3qAhISiGG4Hv7BqsHLm5OhfRG83mwNJcneQGDGOgEALQg/yQRP3
qj5CzbgM1BTusfwvzo2Rszz6SwJulP2eab+I3aPvKwyyyn5FpFWVIvkjn7d6Sy1Ymg+1yGFsXFuw
nr/QKVQV6pbtPe75dSvUIrKcV88zX/HWx8SaPgiNmJWSQbEFOasEII2/lpa0ItLmaKRNh9hOulHu
rsAAvC6u5014tqxWFK4P/8q2YKffN3XSA+ynzbKQfYZAl7NQT0KndFCuK5/3vx5TKKyH4aqpJo9b
bj+Gw07XOMvc4DOLqrhPIz/ldDGgfJ/a2522Ofy6NVfau+mg1JU/EOp2zehIbSBvWhMUsSiIgt5N
YHPuAC1W2wQSaDOaegqSReqqKiQvYcl7SUJalRatKJa+aNfcZXvhs7LFMPFlpCqLmd9yW401sj0Q
2lRbAWwvhIHn041+7pPjjzEzKBZT5vJQ4k180iVwkNoje+CC/fF3Whk28NKppYncWtrLjDYkM+7a
K0J0twl2aEeTp0hwAAHOxOkSBQ0lDJoy+9NsfXNjxDbWe327W70RknGpCaMAw0/TgaiQaq/ExJ6M
6MO2f3QXZlzGqooKFIlIlJkJFtdPL0OVN9KZ6ekkZ9T0nmhTp48TWf/cfVvZGh9yCwhnRY07IDjt
NPQ0Lca6S2KOUNrOWWF2xYZHoNcc3dmzNeYs4VAVeMiT+s/+Mt9arTyr9JaXTYV7HNDe3lOXKyx5
7D06v8Vu7GEjXn378Ezoer61dmamfYR2IYpUEmoXg40wGQIUx53MMOih1R6z1IXFwUQMhwkGJOW6
2fUB+vaIcqUwmlD+bnWb4WmNgoTzIbZZdnhTGbb/tOpngGrPAxqqh0ceL6niP0rPXJ7trQB6HDtY
IJ0Tl3mWeoqtqo1QrzrkYU9B1S5d41uvISjk1UIYcDk18fQFfQqp4VSohtaeBwuPweujJzEA3BuW
p+TUim9LB1Enpvy7Jl1pt+5ZaTbIbL9hNNPKOd7WQeN1B2LUud7VN/Hl7vDGUUniJHWrn2e5tXQi
+mMoln2xcanCVkLefr4Wc0TBEcaOppmYkbvkyQhQPA8t6B2DP5rXckERraJmC9nQ9Du0Odh7FKxy
4tkCHtT9IueOVmy+N7SGMPA6K/H1u4GotSTFrr24/CCXT7cOmI1X8S8s+YVQBI7285fqJA8vEHfm
JW0/B3bmYGdqfdAyBNAQdklxT0rQBYsozYydQhkPTbfv9hmC1FjO4SKeAiAA6SHJGNQtaKI2+3xy
Ph8TjGDRUp+1MAKmp4Y86GoXKxhvAP5RfPxz+4Poj5bHIWqpNvuD1S5TBrEaZRTjI5rApH8uC4Uv
fN2Vl13x8p5owYfvhuweFHxlX0qPyuwgjcFJVTv2pNMw3r+nL5HtVWI4FCIQFWQapqRVW8lsDxQ+
18NZeCopGslnSCZKZzzBlftfrFw+qxmiirLxEwGk2hK0HLp3JMIem0sNZEe14DtvMCahZAn3xnlq
ew5iT2LU8mIgOIJYBVOaxRzlnTnOkpU4WrXVpDPb7kXke6FffHwkLzIkxnJBmTYsVn+sJWCQfJGB
H7u0xGClGblm27NX7+XYl4ZvRTKhJOPG0gKDjSqlV/0FyHOKyFbhssFMVxxNRuy6DdDxWCRKxXcl
RSYFOK0k4bOXVV7r3KUfsM7YE9vHDZXftSUi2ojpoeon8MBPT+fG/Oi2kQXv4h3zqk+Sx2F6wc4Z
rCcpMcVnfZApDrdgb+oxBlaPps4lPsNRX7sFh0VugJjN95URcctI7j92yLEaWM0zAYmqSyaYTfGL
/j+7rWkA7Brp4+8pCWDNg3yJBH6Qdq4TgzO1J2XfqJJv06bCL/P9O+gm6rPekW1MMwr9ADEfqD+V
ysu58Co9paGdvdEZgkypoS5gciO9He20bTBPGY2dH+YYNCWJQx+ChGtGGy9Wm2pKnY61UQ0slRFA
J2PTaaBzE7iPayzAwHnVTiIoJvEvoJ4ILFFYYJqe1nlXEAHtBYOAwJM/PbVxFptZqx0Q6Ce6glE2
qwLJnagFuSirqWfu1e6o2gwnIJbT0n1MXF7CG29SUGuW+ENkfUPVkBAEGfhk+fVgPgd+VdvOoOaO
RAooaPe9ONT+7v8VBjomuqVH6p0hbXDJA8kSi9Tk5nQuYSM2UkyncDBwnWjM3/HYSMC+emt15T8M
tkqJgib6b1+9DcUHQ5lAW/yXZ1di1YYQCarRBj3dH3cnrmU4wtbPE7waM+98/QFb+pXW/2mKud1h
nhE/OfgxBxZEGNg5fXjR68h7cP6Vg9f+2rXrRuTmLL074U95tpn50o8q2hbJv8WCuQVFAMu/bOhP
KrQw0renl5xTWCUxVNzeEP/IKX7mHdjSR3OgShcsKzZ/EAUM05pOvmKTFdSzTXduuCFIAQrSEmCm
V/kqfy8C9XSoDIzqY9foCdh6lHQp+Fyvce7Zr1YH7LAyijMhXMX9Dz1oosHp3bJn9Ps7EIcacDRa
2eHOPL1CitMEOSBKWiVvPlqwtQg/187LVb6Md0TvlH+uswKUzgLnY9swQLwtgjkgTY/En0kmQ7eE
SFZ/bRTg9C9JWN6kSBut6/WkBQfCBShWM6/I0TT/2JJJ6XsEHIB9yZQAIkXV8oWSbKCztHfZ34Kh
fF+D5yrh70Ctp0R5Lqu281IAB7Oatvit4Zwng1dda30fdBj+NprL28b5Brc989zFCscJpj8EADQk
HqZ2dOYFP3mLnO0+DQMkopWbH8ZZzqzIHmpW95aTdkVFXoCpUh0SH82KYUANNc0mvaoW/J1bEcfB
dFGQPlOMhJjV/uxQpGfgIKNhUus3qsQrWI5knnVQjeLCJFPPXviQSJoNH6Wr0cnzjqR7TTK8azj+
grYjwY+TKVp9q8rY+pBtDE265CPYBx4OEpkv4iiG77wKwJYTa3aSeWxp4zj850O1tKhgOkshDoIy
VrHhx8Amw+0Pr3rui4TfvhA6KSOxKZ3Em3Srs4NayRRtK+qM9CjgfNwr3r66UqqBd7GsJyLzJ8c+
aS8OniVvXGnWCQfKNSxOtSmmwX5l7Rs8OnUPSS024r0y90JngIYQ0i5Tx6FaPs9jdg3M1iUfz0Qc
ulpCxs73SegRR963STpSomI+AqwAm7hYCNxYyHpkZZwvZoWztamnpoEp1TCrEFqoyZqeCEkvEk+h
/jk9s2V1O75R/l+gnm8kqqQCbS4FRpOs5QFpQf6x+lg13hjR3vvP7BUKM5RM5CUFeBUrFFNxTLf3
SIJmkgRtP9hq7fiZG8g6kQeWdIIef2pHsiai24n3eVvSyg6Pu/IfrF5nlrnEswQPQkctxBsPFMhJ
4Q8tiKdedI40sKg+QL/O0GMM/o0IwtdV1EGVLEROdq0TQNqBsvyJsKnlYx6gXHS4Id1o7aBSiZx+
iNSBEkZuMa7LoBW7MTo7Q+6bvhcWlsdZgmYG+QuAxZdPsE2SFCM/z/oetjfWGMMl5oB/RSYRExIe
FQhslz6BkFF5v2tvRJ3wEEE8tFGfnY76OqVClyQX9rgPIapOkMr+GJJ28ktIR0wgj3vWYRBdfg8/
p4/wXjUInoxkBktld3aM3/FEUF5f3QOd7hkF+eXAQ+T0qrqxx/iwlfoamHctt9xrjDW8i9IIjVxq
2W5dK2ozWQ7dVf2HlK44AN6wZxUrYL+ApQv8PgHTkcSOtxwCgG+DF8jc9j/mAKpK3BAtYit5xe3a
inz/a/8rjn3xoioe5LUd1cUhHQaARohGSSOdlGo/Z0foRaxFSTtH2Du90ETRtJuTBwCS3B8P8A2u
x2ukVeKu+nnBWKFpOtQtIN2bOWyJ8X1qKLcE4OJj+p6jTW4TX3DJE5fNgBydrOj7aey/Nm/Ek1X+
HnjWoBUvy1Bt8XW1AYwK1pLoolV4+z9uA74lNBBxvh9R96loTy44n9A73VTY00iM0Mb4UWUhK1nB
/Nw6YtFaMqb/KoLALqDZmkN/0l3lEgGHEEYd8EK13h8cT+gWoe4KlMfwbqBfsnvC5V3ac/1Nnz3q
gSZ1eQdK4/6sa9q4xqMIIipsLaVTI7+ivpUBm0xyxbp+0D05rQLj/4Nuq0dQEH/Y8CZB7OKeg5bX
esEjP1mgDXsZ3YV89YapOddvLvi/kDqKVbeVVdEiFIrqoxGqdK9ds9kU0ZWWYw1Ko3LWL548oaH1
Yb3Sq4snMnynmK+6tCFyUn8RkXjb0e7Wo5vJ07F/QRlzs56wt6GHEtat9VpmD2jLwOY5ONRjkhn8
AJk9bBrjq3YF8aBYt3fCkfYRzP3wIT44Nc53AQZBvaVMivpyGg75C1aTiUuKw4OUCvCNwBJiXhj5
PRFxVUpBuSxSC+nhL9ch3CNB8UGsnMnTz1GamFEKJFdSCRCdI2cDXfgXZBHxxpZyBbsGTKdBV9C8
1niShHC9BJyHfgh972kDgvmz2tUTt9SyG4E2DzsFETGwRQKFC3THspALXk6+1fXmlAU/pJLeCNT0
Az0STKNy3AY6E0YucFznulb2MMt4rRKyPfGysZDnHiYpOVJQLvByzg07YBDUtlYjny4aVcUABftQ
tdCmGwIdR6OxbhOKesEQv1v1T+mzmhf5jZ90SiuE7M1xkR/KbCquVrp0OqWseEOfXhmcUNLmHwcX
IJ6oT7fp5Y8qwTigPPLLwp9QOKd0fmLdLCHLGBX8fjT0012knSRiWUpRS6pLlE6u7HfVB0upKN5k
L0vFyYLbTESd1xXFu/UtnvSevxtTxXANh1LO3nj8n8Q/OZ3d9HbyYOcQdoDDgcoPr7ZnuDP++dFQ
JiBL4aNRrOiPG96YuS0luWF/Xi/0BsodXfJz0mw3ZY5lTBLKQVLwDAlfi9kdMd72AeQFRGd+Ol2P
fpNhFK0snFnYqkr5xKy9QYM5929umPpsQij+wcBctb208X9mQlMD4A0MyuVe9kxykmS2L7+9EA6a
LRKB+EhuVHR9LIje5WrkHK/FqOtcYSfrdKodh04VmJsIERGNE/tSd7ZVnev+FehziSifL3U7nh3X
IUQoBzk4y61KWebU4PNG63V65Qx1h7vfKpEEgbzp2BFVbykqlkWR+aDR0plStTrQgsPv+u5JPQzA
6JEc08rHsnm0R0JX5JsT3a1fzHUiPLkTsCtJzc3S/5hIK74nWuoomTW/biQItDze9wKCQ1p4s3nF
DEVKW6Agel2Gy9vFSrroiYmmvrL54/zV6Xkkmb6UX99uRfScpTaaDvzqAn4CZrtJsdNuPxkeBOzE
p3kIeHSBB0/AnwAeSedLV+87ElUHNSD34fZTt0VJ42UXUExK+pt/rVvwyNfwVSS4BG+LPrmiJCZe
Pk2rhEwwkN2ufVJcMAvkog+4L0nfiXmif7GKGQnFf3Row2TR4fhlvYLLtKfDf46hDNACngPS3DIv
qCWr0YiZAd8SLWcMWJeGYNCdeDtACLiZeS9KOSyvT0MhEue5tOk/39H7CfqqNFgAcDt4wSNoH9FZ
2ITUMVgCoOPbA7GqeM6TDIhGN6vdKdaYx8xmNJiKEC4z1k0SSN3vjHeib5TYOpLosytdH0zYMWUn
ozdgnVqvtdp291xnkdeETquajYbDPHjZ0wPFAX5IkPgfw79kzSMkuejpeBbifELepAv7U4CazXkG
aVZ0SAPSFjgF/Oa7Cnaqr5dCC232vzCMFQaTkDkZ/6FuStzmc11FSl222zGM//x7Rl3tVgU844o0
gb0gOADRyAEAoN2MZloWdUlgoKlYOAjyzvtEZXrK0MIK3pb+KHCztCsux3+fQT1TBb3drF9BaDAa
BpXvfjQunLnBJJl8TJSGpRuKNQcGp2Ef70dbAMlNyLsRce1TOaxqpx7phT7ZKTJ5lKZYXjsTlM9V
k2rjALL8ughAhJe0eCFPUj6fN+9qt6XIhP8XASSY045qdJuKEJ+GSqX4jkNtHwhoLoxWjukTtpHO
nnInbBx6eq2/Iew0HaKZJ91pUD+4ngavcp9JqW0xoDWjKf+rQpDQiB7fGCrvKJguEkNEmeDvhpEl
zpwMh9Q38tzMHLTVf+wCQKML0JrglnVeyj8zE6XODLmBKLJpuqO5mZTXUyFzYI1kLmCIJ5X13CYx
SKZSroGQTsYcR5HO0NotM21n2vbZmkBpXxt5B83iof0unyCoS1LCr8caGyWuXucOvWTxOjNArJ3s
shrmN/lulzmAwXMrpA1Nw6F5jxy6UT+zIEafA3yzKiqn7e98h/0ZtVSsD5lvB7LedXIsbrylFR4H
qvFuq0EqfOAZcqqq2aqP/pTT/zSO/QphBd8LrfeAXPCZlFaJJd5Q/IgT1rYPNiMzm76KFPKQfJ6N
vOGtk5IxoPJQKXlnaXp+C1bO9Otfm98VGAWcxM4GKd9KDAboZe3oyPgqiBI4AkaehSVZzQ178Q3P
jF1mTZ4sMhiAjhKPqrIyAL+C65HB3B2zEZVltrupmTSZYlg47js46q3+0H9TpKQ6nrkEcvdkMnwH
M51Q6FicCRdVO1aM7hTo65YSci0SPLIDC+z2XzBdH+I77LstmSSa+H9DtBWpAWRCbBA7+kHkV0Cd
lAseEJQdN8y3/Cp7lKt/mmm560QLm9t9Bw8dpKZdni+Q4W1gXzkKqMBD1Io/QlLWnrxlwAobIuF9
fzMk8JTlEyCXJAZDU2uoIhY85vSKWd1MEbp3eei+uf1gTzPhppTkqqvOvV964Hj2fRg93eAPCwWH
gvwYuzQP1VrOwwXnPNUs+1g9+EPjMepVfePkzeFsYXEVZMwI3ggC62p94BW8gYYSOVkaf/3nIRMt
Rg7GCu0Iwa0Gu3MNEuiy/sw9wY6vmA0HMsWLAUC+cGdt5ehj1CW/gN/8ScUjNIBspE1Yse4myehf
EEz6IFKLynFVMp3TiCZ4tsRKbr3fR3+vRem/Yk1F1xN05ZDOVoCfp9kllwwm7BAZNBVM6SbG57oL
Aru5EA9akno0Cs01Aat4w1O6uyZ5J0JLGkZ8Nxavdur/dp3+nKAAa2Wa/qCuYRj0QLxebNOl70eI
P8UTMINvSqlD6Fim2aBNncoQAKTsgJyGzum6u3C8ODlycMoYDdJbU18ea4F5dr5RfGheC8+Pb21+
cIBx6L/f42x5rfS06rvcKU9qr0OhJGVeKq3Mc6TS6z3ajcSYEy0x6RHYDdPiAYCWDl6povHncYw4
8jvqHm2NEhzRfB5SCHd7eMaTG20v28HHlJ0jLbLXbQMPhZ2EyY6H0RIWxpt8wrqbjZB0Io3m0tzc
lQ7yW3RF8agiBFRYbphf7gE7BGrG/rkjjlcM17q1oHIRDM7Ww7KAP3hA6iUQP4AAEO+jBKZ6JILP
3GCSsWcVP1Zc8ZlyNpfmXomHX3tQkn7UkVOrCLcgDyP9IOnFGOFc5xwvQsG4aHWEPzC8jKxuG8Ai
qoNStmemY52xpe38RGuFCz5g6oXefNThFlzNMX2Bd4tlKmpFQZTNUc0afl27/r7pBB2GXWr99frD
0ntzWfwUYdl8MSoNdE0TH9xg/gQtJVbC5LxcbFy/jep51RCYK1dCpfXNF6c5dT94n5gsajj8dm/O
z2BNWkTPMUvq+6tvUq5VIxymi2iY1DPqn1GvqLGOXatE9GRI2Rn9Dn0LrnpkgAVrBWes1aULjlkV
TAtf4L7wwyjmtwQwvKQxuK7cR/Ts/T0yhvs7DcSQynHb27PtiRaFzCHxHeypBiuQceWIsIeaydmf
gDB/bSKC0+xd0sUhBp0U2xeb9lm+0VI3C05hefTwz6Enxl4TVG0NZzhmdXh6V7fhP0PRhIJ4fIId
Zj0Fys3Md71hJCjFpCfatLByAyFh43uqjlz0AXYXpgYpgtVM8y7yaOVod6UAIbIL/4pC676OsF2h
mXtROOc5HW+pGRpTDZOQyd/SmtXUnyD1Ipg902DfLw+vXr395W4EZId3EzLMzgLxQWRJhAduEHxa
U2rbKmU/B8W5R+WX5Ary3/nhyyUnwUZaRhbeE58QpYvJyFpEStwr372dLXZ/VuSquHwendXldRdg
FnqSF7Z/xlZoJqs86kB9kk3wFkozpek6e9lIFJsEpmqx4ulO5TRjRn8DP9RK43UyWQ59MEWo/DoT
qDSLzijjYE60CzwF9sCJRsIHJg9oyPyiUWUMfvxeFSCSB5XGaMqpuu5/mCLEDnywECCX6e00mkIz
gZU9wM5No0KHLnvLWE7QAeMriowsqMIdC2uY6RTORz4L2jprirGNAmiLS4/6Q6yE5VnOk29vcxIq
RIz8ofAQynIRenoaBBYpk1wKBo7tBIp8QLc0yb8WPJ2XdAhW2Te7QVFvzioun6CVk+BYo/d1NH2W
B9x0NmpvAJ+ufT+QH412nae9m3cOuS/vpFVe/fwyU5/c90nq5RZaxMkXEw9DqX0OvtO8ZAwrbudf
wHYIvfb+0JI8KTWaJ1efcJeDsP7o4QrZx+GlXci/VCXMqgQ/VsDQmMaE583zK75CwowJ6WrrPmc4
LIA3pN3MadfYeNfVZDFdU2vDC1nNwavw18OEvw+wXJTUGQ+TUF4IoX2g7DKBeUlpN/JzPNBgUpKY
SUB57fJWi+qHVf9pzAS8JdjVKvsxNZwyyBslydFXpKdK3StFSI5bNGTTvFmOhVwEqV6cDjne/Ccx
8Z5mfP0wdB1UXBsynJ9BWyyhmbbz16AOePjTxZmVp0D9j9wGEBOBxQBD72dD5G5Ys+UxXznmlSwC
IQYIBKojx88FXasrh7MSS3vDPlm914sblmA/5FTf43SsX/O0dvkMLwql96eHHvwCBBn6yYYtz0kL
kLZE1vfR6gjCPJjjAO8f6eGhNgQdZ11Ss3nNfAp0o9J8+KW1MwEugqo44fhIhprs5XiX+zZu84Zc
49xx5PVIaXrtBQ1TK8ss3ZHNA/vqHWpDD3uw56xuDraEXSKZ3yPNzGRlVJmLPflWaL46xdZC2gwl
BJDBTNug6fCeWhFwN931oQPfl/eUAPfzZvkw4qZgNLxcsza7BIHio4xGhf6Yo6H64oo6WkSJ6j9e
nN1hAAxYVKWeMSjEn7dFNXozKzM+YzWKXO1rubmyH5xRTbGLdWQEVkyut4p9mjyAaMGExa/2dXmz
OtvHw1AAIErFKhlfRLTD25uXwg/pFTaHHFtUJo8Ns1tLP82f/xlLnB01aFjk6eMoV1flThHxN/FH
VchZyP+YMXOBkPp9Y5eFRVK6NI00ctEauA1FQYC3TP2a71rquApTt5JcG5NrURG5YWpym47fPEA6
aq1IQIo+kcz0FKQrCsRiYAvlZTmk9Vdh3xrsHoW4jkUjZmygScdqKI2NwqVa/T6jqtJf8CNHnC4v
2zrudCNsJWUQH9AZEXWPnj/lrGjwGuKHzv1zFntFS1y8jyeU9C1EnG803tvZTAznk4ldrGgaetXW
xZx4Ac3bhZ6fPbBFuzWzhvu3iKMX1rtnrPRLRZE0Kzp8iA2BBsuGiVuwvM4N4mwXK/Yn7DF04pah
OWE+ehlm4ovx2szjiasclrz+3NnjJAknw6LVdlXv0yfEH3fu2AlpzpHtQPDS3zpnvN/l1LdRrpsZ
fV3fi7PfiGS5udgJ5YFyXz/5ZwUh7TtwbU0LDKbeS0csZiEL1xUMdpg9diL2IiJvyIHwVD/GzISw
EmQ2UR+6Ty6ANOY2gpwwTHkiLQXfj9VIt8Yi4iw/zpNLRMn2ewKcLP70JJ8oCT8kbyBhUYpCqy43
CMG2B01oYZZXiNtyCQM6CQFWQAz4OJMeT9gaYH2N3a0euXyZMbHAYYTzuvsGs3Gn6RUY/5+bzYZ6
NNka6HAOgpjXttCVNsVFYzSFYpEVw63PfLoIFG38pfDSm32AHVCr7uFuVLXcJ9cMhl5E+Uen5/pw
qQFs7ypoCub5BCLnwGS3tmPMIxgdN64RHfg+hbg6IQc2sjxktLpgsoqEI7BVXEX5wSeRUP6Zxekp
PoZWYmRoR4n3m4OVsCuTQwvHrzFIzHt850H44Dshx/vBsvUxLspEQ6M0mGMQfDZJRa2DgSRN2m4g
E5BTUwHTMuYeTkghlUAi7oHsN2yg+KZD5o0g4fYrAgyGOoAdW+7gbM21ZB+FT0Jy6IV5Vmy/cPRE
f4m1tkTQgLDFzbFf8lG4sh5KWt1COgn/eeD7iuIYBykEPBuXAdOrvgjI+hXOBDSC0O836CHvng8u
pWlfAIxqinW0KTeSiCmxvj6MOhERxWFlYdPML5w9z43z2gQvVjo2iGORW6inuqbdDemnuTPJfQrp
f8SDUzd0f+k+xghq3mb0t0lYwjBCnxNCTpKYzQw4shudPGRUM4pRd6d5enphGvxeswEhaEZGSE/5
RBb4gEMCUIMAMPsiWbO61n10xGiPwP2p0pOO6b75ZXBSP3k1lN2okbavgXEXWxILlqu2C5i2pZw8
Tz0avwF/qdgF1dhJsd5EoIU63tFYSXpxyMCBb+1RFy8vwAziD8tM63yRZ+xPMc2BdO12m1oEeWKo
HYFQQk+7s0Mehj3sQ/4tDjIk0lVOAVrTMQP2xd8HjSufmstO5ZRmilyiciUUd+CPcxJPmucJiB0/
OAe7Gd+9pnB3LXwQ5j57lTrcVI5Sqqaw9BkifUVAKuFViqFBKOtKgUvTiokaV4289OfrnLSGpoHm
5TVnuX4QMoLEyjNDjOQ3fQNP5dGPkC0K5t7KC1sZblnCAyoSZnVeCg5Aj6WxVwp2zIvsdAObX7ng
kDkw6FeGsJmJ1BURH+lYCHC7jlkkBWwIVfpfgvdBLRbMxxLF6XIWw0PW/fr/k3fkdADrgn2G+N8S
Keozdady3FOK6toFbx3fpsgExT4YdijiGPbngDXBs5/ah/gAZHrir5nyVMf8NoUDLkqzRcqpNZz+
XOtHHGmE4n2yFxqfDH+zZ4WXm7Bzqu8lKe5xT3Twfr2xOz4Z+/sFkbK+8XLIpmFb0Gx3J/g9GLxs
HOlKxAv7b7JB4mI6aej/hRPav/ugsWlGmbWyj55JbkudX6bshOxlWJiIwToxzJh6InJRfSlkMnYz
VFB99bPkDBKejbg/ghuk8m4OBJ8xKjdy64mRYvTuwQbSUO1bSlp1Lba3kVZbdgLDu1AgsKMerHxp
OOPCysNVfvlN71matmlv26B5amavQBfUVN6kY79JZwqSYqQdFd0ctqbpr8lI9JOAL+9C47gKPhAJ
UrZhVojVF3n1eFgToQrsGvRPezJkv/Wqj50/vfFp2faUXxLDfbcIOiJhO2c3TlhPs/6C34cWW8v/
gXDRh+vvUieuOejceSDpD1puPWuSJnyTPR1pYbhipUV1Q3JZo7DPKxOSRVzMKkFJSmppoXgVQjbm
N7J21ID/5XSemagCuKOe/GWdnHhBXgJxQ1oje+M4g8iw9sY587rOazxNdDxTvemAF2WnIPIZTVPZ
EcMlVfDHY8ExqCRsqToKDNhTR1YSoo2Y2m52R/MRr1hScJv+NI/eFY7bj4m6JZwFXnV9ep3AgLCS
Aq3YOi+aRFOescalqzsfMpz6bPs+CTiJPCDIiXPPGP40GIYmw4nxzBiaZlEXlyocYXXFBAscn+WF
Vs2WVxfBVkJ5zBUK/AiCsSG2ROA21M3STtjb5F2Z2XjLdRDHJDIkXrbFnY95JGiP9zyzEA6qKZe6
lrGh6gsHLjWUZaVVok2LRFmvHLpkGGK/ucyVHl2WG8pmQR3F0bIan8w8BBp5H0EZJ10IsZCnTkrV
xy8H5JKHkWnSTj14fPZpoTRiAZF4oiqFtuGrsWuEL761mCvfmkmG7rauugLqBZrgGKNbr69eEVCN
dds2794S35Lrci7EuPlOuopcAucHCgqLjgxqSHzyuApa1xveWUHsBY2+AhFSj2T+j1Zv57nbT7ig
1TVlOW9NKmVxL6FVzCnSEameEyMv7goETRkSpKOkwmuxb1YLnb7momO+s8t7mUOjTWOJQ9jZ02v1
KvHOEoA6MlCy1kPVGzca4ZUCZ30Niep029XDUZx3YVxK6zLqTYhtQ7mFU1rZHSEs/O8E4TsbU+C1
cZxB4Vh7ReWv96MWhsLK43TWAL1tLIrXzbkCw56wnlMUiLY+sf30xXmLybZywHeoxw/F/E0Wl+7/
1XWqJuVnoJ7qP0hGzvOhdcBd/AyPwDRqil0Zjv84sP52EDUGtAiTxRyERmHC1XdO8Rv50AY2cYCD
7EE5Sivzi8DJs1lmcdjTz0PJpvKLWViYxCqnJg7c6tCZ2B0oyGlgx69ItlD07hyvfRC7EZ48WOxW
z+OdcXTtcYhlQRw2/MnjqrO+FepRghYCgS1veO8bgjjkQ51j1KfoPbdcvh0gkmNm4WABLss0xzKc
2I4L11aDjOhG4D8Cz/BLN5GKkwStQCZ6a4BwodXEJKPJivVYKY5HWv8qsxM6FpRc3GYIg4uPYaol
4awwzr+pP0zbmM+0CPntYQOs2AbagUgVK6Cd2hRH9zOU2QFOAN03MWqxqdsdhufkW6KFkDO+fjUg
7/Detkg/yk10h3+CPb4aKveB6MhocDjy5TusWz4W2tiRkyvvWRzeMjglAqeRfSR3X70WHUeXJgab
8o4VN7omn1kTNL/fJWzeVWN7slfXaUzD82v8dE/fJosRwSjfN3cD9Se+FIu/BKoJ2IucOOUhkMh/
I05DgJIg6IQ8TvRnaplFdLQg8l6bVb1VND2oIeiOoCvPnC/k1gAl3jnpys4ZqLFD9+YnOIEeOk6E
dGfwUx6LIhQLVLFzxQYmaeQ4HU7GLrKeE6MkyjXjwAw8xRXCF64iz/+uSXwS6eYEjzpbJZtRiVwk
xdD3rWO35TWLAxbwdO1WP6lyIE6UFIXMizX0fwmo/6zq7WyuZtFBpMlKpDxRVUH0ODy7xwpSiMt9
b3J8RxYj9F39qRql0L+UzvmTRvQc87BRya+qOgZS6yMRnFX10ImbyHZ4uWxH0QrkJJzUACLZZTXS
yo2ItY9Lu6w+8wVtv1+L+mD9iIJom/NaYkMuE7dQ3J1Bmtsl+JVFOsHmGaMpA8RvtQ3rEHcojVFg
UckojH1ezmD4SKGCc3jmkuBP1D0Dika4lJFYdzUlXLNHHSErFW3P6eT65uBcxx4QOjEgkenRZGWW
cej+w/K+U+bbFfMTwsPRSks/6PF3cY/JNwpHTgowqcKTq7skz4TlSI5m84+/pV2QThgDMgDvWtWj
fpd9M2GOpWRtj25CoVRP9WKE1aHndcE4ypqZSr1LtWD90rdP11duZt1a0ZPgd5DCIrhQ2cF9anHt
v9IdouE2kdalha6iE3ZJKr1MI+//1bhSVazwddFw//1bxK9MAllMpFovxaQcAXtOPFk3T8pBRct4
lV2KpXjNQUWdiqe2p9JZlGurTFErz+CKeEAvYTKONZu674GNjSrtPQjOyK1CPKE0VX1D0v0KW+7R
DHKKIHdhx1f8tyDhRenyQut3zvrX0DNKCKFG/fhXaPaasJSRjkMO1GRJuD13MukBqa6rH2uLctEt
AWXxbEkWrDeeWtvV64FC00Q5cg5WGeoGBhMOIUyo54aN49tVMe9v8bA5NcNgDERE++KBVxEK8WU3
pEL9iROATPhri9/P6ZUcK0ZfoJxl+WPhWAg7srxab0MO389kYMNrmaA1PmmS8bjdDyPF5PzAXxT5
CBiOvxUXySevSXXEI6qx4v1+yy4VwsNG9H4C0oeHTJIcXRr6cC2rpnQfCx6wcpLax4pGfyKC8HM6
yoAnRwIgxyme8/hk/nXCDXomV+6dLlrXhLCBSLSMtftS6HhJ9UYkKgUbLny/xg/sGCnu/sNhG2jp
1EQwnCKrieTyi0QBztaPt3L30nqzMzgjL+Tg1mhckoQAiDUIaBtHo9YBreBGw1WwI/wRestR8ERs
GateIhHvrcwhm+aj+ZPYX9l1wQPGGv+1rYaBp8Ekxxb/tMgK0Yd/cDpp9lTd5M2AnctcmbTs5V0M
KE0TDrsBq6M4eBXcbmQKfj6SOwJOtOFObmmrQmO63IDHBD5P9KcQDBB3REo6fgK7yOGVnMdrkBJB
cEahjhu+4fTkJuwgQPeIHn1dcFWoFGJ3xGFxf/xP16ozUumy86GnpmZixIh4TZFj5yNLr993cCkB
t30qpky6gW5fWke/QDWW18W1TqZoGUBQK7vKhhq8jTyaQ8F9U+nvTubuFErZXQbYPD3Ms/7Dws5p
522nMQv08WMNKj093ja+LK87NWMkeVMy87NUD2Iw3ULcxYLSE/li/qphVwGtYVW6nXES10dcGcuN
QQMhxKri/2NcriPJ0KGPVYnXu09Hi/FHBSemgEEYcK7Q7WTkGESeYfu8GQmfou4xay4JndlhrDLe
rOkn1b/ZVbEvKkpfdTA7ivbqdpqpW+V6pT1C7QQkCl+swz5w/dR1IhTLSk87UTHHcCn1VDV2ygRH
5Fw/PJsr6PVNc8JzAIY2F42GQGwxMCa/NfT+lIW2jc6xP1IvZBvjC+KCbDiHnv2PSvt8cGLVuPDA
og1sVcLF8YMvLUweb2NQyP0F4gEsTTtJBK+4Wj7NPEzIkjtK7SP2oT0SrEuutfALqeiE1amU5+QW
DhLKZisLpnwlQ/E/ENqcVKCuDYRxh7WdPMDrqVvRobfKT6jPPmN9ANOjFtKEUx6hCfqwdSwSRbdB
6DpDzxjIvxzspx3GBx0tJixG0kl5571/S4y64dI89zDwh4npeLGZMRCMEq20mM17BgiN9iG3/Zil
QXOMnivmHmfSyHerpnyZZNIR6jlulclZTlChREkxKCRKMvLZHXub7Wxl7ctTMH1/XMeLY/V31uKL
PRkwN54A1HFyaZqEKOttUXLAyZpjLIJ8zOzbzPeA9dUbuXfNpcAS8pD0fH7gMibiUtfRjwPIc4zN
VAFcy7mXc46bNPV1g5dgiNePPpAAjfBjnzn3vOxvTKtCw4CnZ2vVh8PYsmghu6Z25N0OcL3sBLTQ
oKFWTv74JgFnOaxxI6/Wq7VFLEVwRTb8vE0pPwyDuigSwu4YPBGWuj1XtF8ckeZMZk4CFQ32T38e
aGCvJXve+MrHnIooiVZIU8nXKDRuGvY/nL4V3DTyX/3rsobcX6Rgm1E0MQDGc50nYybaAwRbt7vK
OLGGmagA/Gnj2ygu/ZFmpRoOxNOq/sMDN0wbePUJdmdipDpOKGCIOvVWPJbm+td1uc1e1b3tzkOg
ECw119cr92Fv5dvA2onnPc6iQaTtux946T2purt2WI2b0ruKjcrUhRF+70tpJNWo/w0vutFkVrW6
b74vl/mIQqSiU4fo5OQJmtvK86leQXT5lfxy8X1PetldchHp41kywXvPWSqVzvDgdrLa6L3pZzOV
edvpllaLEsn9khsEp35iNd7SFkH9Y7kqznjCr9Q9v2gUXhcFzV/zOHYtJGvfyuX8BbTM3jxHIzhV
GsIcPhwWV8UwnJM+IhOqRsZADfUY/a4C1YMpZ9NT39/YOS5xW8TAPxnj89TMYOf6qjAmTPQEaaXu
/kCgw2b8nqrW5OqyCRXsNCHn3Y+Kf+2gd9SnFs3e90COHcEgTKU+NXBno+BQaKhiaWVslc0+EHgR
k6kcDHqgRGgKYC73uWMrDtKsevxlr5LgtXEck+cJwXPW8Z4A7FMvkWzKCSdNZcktkCu7BDTBuoAP
lmnoHos1xNs2kv5mA/JS6iaqq1weGWUaXXa6NoH1PAGcO+PfkapbNarnMwVbmX2Zw34aZXxiVy/u
BM4yi84gycKFwcrYu76tML92OURwQdRSHgy2P3gIN9G97YDn3kvHl+f7gu2CTlM6kPrSDGJ5WNt3
PIPru+gWL73mfrEmHagI4n0tEwv2eeXfajilwMlVgpo+TXlNY84sNCjlhicfXwg5PXRs1sg3lSYh
ntXh1gF4fIFRUsUuoGTobYb94jwEXVgRzGFkmyq67YpSPJSsCJSRNj9Qb5MBVSe1EfAbB7GaaUN3
WlYcpeAbjPcVq2WNKXYQ+01G/x1tslbL8ce900TDxpNPUdU/V+8NcHPUxIaD28glgdN7IDxnqh/H
TmgMLf9wACiWjgjitOmPLxy+c56bVOryVfyPkhI5al6vP6OyN/xeiOVJUoMk+H7bJCZXnyWVpv9L
NUcKrKbcitPiBhCIB/ib+dmcoH0kixMJpcD2rHSOVcGH1Axedc1dRNm3h4sUaHA0RXTpmwf3mwCP
kqNbNwLdyKQ47eBpu7iQZwJMtXMZyh1l6pMFm4arttRGuP1LUq5KEJiGzSNvxSVQiYjQLAR7NsV0
UoGGeOPi4d++Owlxa+vr5oaH7aekoUcr4t8VP4HmGcXmibK3X6GmRSC8s8ev8flDm0ZPEU8PY9sT
98QoKPxoWPUZBC/Mw7Kps93AlxbBXHi/5YG22NWS7o5bMuRtWP8v20qw8LXlzbB22WVFjAlsKY1y
E9TDG48Zu1qax7e57bHIHWnx8nlubEn0UVgG/IprJdPzRn2AgvL57yGca2Jjd2g1KnWJHYOy9RAR
Csa3QaQALwcDT5M04MEWvkYQEYEpKpN7MdAonqMbLRUpgu5uvaw0KT+vkCZcfPgaTjtrTr3eqzfy
YAKQEMmIBjq+Xmrx9jAPHONnPezzG67s9TIqvJ10+VIrJnWxoyOUVsqD7+naw/LNw0qVCIEju3Mb
wtENi0EAsQmommbqfMLTVYeojRCDvFUreIuAUf7T2z8Azde1pb4t9fV6EZDfY7BKTU2lgVUSN5z5
FIi3EvGM6sjroiUrzikAjJTzm6ya7o1oCA3+RProf5qyukA9MUAnd6OTrsDxh6GfHUvD9sr+vlk2
V3TeATXYkDsTaVp0Ivu+Mrs+oiAldCTXE0k+zCxBZ3a0tH7MP1EcqkuZqB2WJ6LkcvWRpRig/pxF
NokzhiRJX9vpAcKfiJngEizUGv4FFlEVBMgg28bKGhVI9v/gfXQH+j7frUJ10p/SHKFPPUXJT/82
74lKAmTEjKOCevGl8Qw1pR93/Jz3e1miSTHFK/slS4TU25AUGJd3ysuKqYwaLWJbrsSwfh7a+FiI
6ikGqTLonSIIzJKIfAyHVpa3exIOUVUKhK0o1wpg6zMurOqF2GP13rfc0krbE9RdRM29l7yZ5yy/
kOJhlGLRHYYQPlCy51GoTv8obmkFk5g3mM3M/ortUWl8tapld2MAWtbB3WWErwd30+i2yACpliq9
1ph7+njKesJ0v0jPgVY3VpsRvGSL2A+r/fsIr5jdEP0d7BHdO6rXU46m9INR9jn85FhF2t59XjmV
9rhfOets28I+WgM198q+JiFKi5RTOoGR9qrpMfXBXXkqvrLtDglfHC1fmxFBzU55lCyTYVJA11RH
ORx462hIHOHFEPFBxECsu+gY4PJOq+rKCBJ0NLfzpCxg7D0O/woaigix6kiUSOfERQRrbLVYPBVw
0mmoLuy/LwW30H1vejTCNe+kj9+koMGv7ULB+PBn+wDFocNE6yJ5ufNdVuWNVkKsLFuFSdQIeh6+
2bndtuHfpJaf4Ae4gWgkF4HigzJqZMOxJBU0mynx2aJZrJwZz65X0hLsJmZsBT71LEJVk5OScKPV
+fmnQxbnf2b5jVaigZezvkWKMLrDejtC4zie71kFPD2igzXtMb7XVuuct8DYIcyaSZAyEBEflUMD
zdxqqk2ybgCYPFg57oSUXztBAgNZH2emQXvQj2iLQdZ2HRDAvNMNyI94DXaf3FNLGmQTG+bGME7H
JEANiRU8Y8HBtV8B2S0fxxd4sp14X7cfuVE3gugj6hSFDJVnkiI61PM4VxOt1L09Z89Z6vma20Bx
NwwKaPxtirAqn2at1C8sCYr/4HXB7C0rRg2E7wcAWX4olzoJqYRV4Ab593DfFkFR5NSiRNTgzNx0
4VFZz9FNMwdvOwDxxjHIKcsBUGP9poD3a6Vr6pWhvjtTK2inF8ahiSF9meB7XtomGCXXG/Y11T91
Qul0xCqmjOAW1j8Nnw6kEQq642HGO8oTCXNGEZdbUEFIpsTvh4ypDwh6J2X3mRMn2F4PwuJ1Yys8
yfmN8I4dmuyZG+P0AqI1+8cwNybaZ7adjl2FFGbwDz3lO3Iv9KLY9NeBLc/1biBlDvtVWJEYm2DH
+qyRoU8cjMFvuGAAvcwma7PNqBBdw9sn365j8laKQybPDm3wlM6Qmvw7jxpCO5IB3Ytie0Bx1u2n
GB48CXenXSRGtZf/A4U491TDT3ikMhXaX9G0yVbNomjMNjGp5OBSnz3iQaglaY35k9gAMy14qWXv
grawCbQnFmg+IjwthkbX4ZYb7eVeOjUdX2WpoQCB6bYqTzNzgkUZCvpfXto02pm9F7PR0fQa4aBG
lY0P+uZpLQrHOjAdlPlgmJdplGH0V5eE8jN9sACrzjvj8sUUNQ4Tmt94m2h+ebIPOpDINHJaI89s
n/EdVCdE27+t0Ei7eftl+WFXqeyGme/wlq0eUXUL7BoFIicZ9PTsibkospRaxRkrGwd6M9kRJsc0
ZZRZMvC5mYzjVnlCKvnvIyGQFHu2OL3iPaweie3tM/AvOFRSI1oUaNeU/A9ylbR4w2KS7KBQPGFC
ls0IqP/Ej34uHwoqla5Uo1PyGQCXHfqrIUusvslINz8k9zHItt369nNuY9lrHCpvci5ewnnj5JYP
/xZJf6MsC2I3AxSXJk5RztDVPmbS2XzfrAMltRYqEIpLZ27jfew50bhqtuROxrCUoNuKeEisYzUI
UzyTBHS760KC4ATtxCJNd19h/LNntkQ9Hhp5HGVixiI+MZA3nJut76ck+cV5fg21lzkPzTh+WESY
lK0IiajAKILlCbGkUhE/hRUtBI4GI+QYB+EAIJx1jIsOurUbd2c+nY7dczIGqrRAJwtiGl762RAV
Pmgp21Nob313bce3/JqwiIEdN7vL5nI4Rn83rVeFYBB9wtnSp5QNyQteH/sGtVWEpxaqQDyz+6an
6WkvCuRfdNB8gtq+asYAQ13JpFD6las7D2cecCm5E9ye8NPioVYvC2GcEQaWgtzEbnIdABF+cDl8
mK6sD16TdFbl1FOvOa8mBH9oi8ntfw0tH9x4N7Mp7fXm30rOY+xQSdOAE5BJGJuPtLYpb6zhrxqd
TfmfAbTZvHTWp2GtkDKwZurNZXt0KQj5wY2spc4MCej17GiGxXlGrOsV750izi6ZZuyJbD0qaAh8
BZFRC81zZu/lFpz6plLyTMVPGkiWpsiIGShBRaVL3m0A8eOyfcILp2PIhoHTv/Wt8XrsA+U6rmIO
4ztOlXMBqcnNbUh/jSx2OY6m3lFzrQXTMRbJFjum9M4Exi7r357auvPk9sXXVz7QEESbfQEgtHFK
4jaLe746E1zMIJKMq9pOLFTZhKRHCkW+RO+KQ/nLSBIffVekNDrrRUST0PA5ejDEYxKqqREc6vDR
9M3A7My/NiKN5pnc0cH/qEs8NA0vX/XQu+zt/GqLSTmRmIQIH6gSLtw5DD9IFfbPfKqgVyW8doPE
VrqJxLmzk/fMNN8lPL7O7NDaKGBQWdPm52t4w19OkhH+KWAPBjRksLbouFB+7lDe2LQKaMVOCfY5
AoIEFPzXr7puuhBwfOpU7+8P4uX2gi1T7KLub8N2jIBJpg9Q4ZXgmkl+1andYg2aZUNFr3affHb8
rP79n6AS9Q5VqmsDENvH3sL9D9UcUoGrnm3x5ja06FX91aPNp07Czvd4ma5ISBjxBfSK3l2cZd+E
ZGe4Cf3cj1k9ic+6bhakofTLvyLsGJIBLmBURpT1S3dAqO7auvfS2WXXSLaCjR6+pRyA5u23lut9
ohw08QpcsjNSInUfGVRsuWxCIZQ2QhuhtnLFGurwxHbP+pbWgXzY3xxkC7rqmFCAYOupKdi6XQXl
Sfnl9fiYOKLGyRh7AtHSrtIjpI1X1oXjGeiYM76CZcx6LAl0nIQlDkjLTAmE2DEinaOkKq//pjeK
sjKiMa8Y0ikp4OF1CpeXlZH031TzuYAXX+uCWUcV3OJRGPr5yNdTCTEdPwWDAg0WgiZwwSIk3slO
Prb9ThSpp8vA12zfvGeQ/Bao5LuGTcKSHGnlmHJr+gcKPOJfv0BYrj0JRMMuQ0s246MJUPF9bx4r
YjDIIA0S8hT1mYQVn78XnW3CB9fTQQiexL30LU9htu7QURL0CFyRPK1CTZOBZ6ei+c+dK7UtOKBw
jx5SXvzNhpa39/WWe3YJfk0ovjEbR0yYg9txHh+49Lpm2PVaFZ6E50iyo5ZoWoVxHanwRe+z39y5
e9l2CWagSrejuWXx7KirVSm3zckhCKtajvPg1ym4wTZZ4bSvlof30MWbpzdS8dl/HGUblS3NsI/m
RDuOCNw6a+8fAtvubWQa9ZjfX0U9kqMmWYj+fbQu7Q7HB0UGpZX5Ej6LkC86LHn5KzhxAgR3tmum
YiDqlE11xF9zNhpe4FO7Ueg/s6sTX7VIWdhZhLpX+svuiBiVLxQeEvGDQPVr83E1eIuxLxtHK5SM
Uje/kX2QZYXiC5ovhcg/4yF0UObI5zuVvmgrT/Gf4Mmjy8KFtSWlxa5JLFahixAvewZf73q8UTkB
GC17ItA/60WzBodAamPwe5+14ADX0W4Z72vY57JGN9qM+Ig3c9UV5Lu0oeeaCK/1LUYCx2QKeXvs
8fAdo+H9U5D8MxIiVCNCzKEbtO6NulqiX4A54Gv7ki/t3AITTicWBO/RtHGQhnYeXgencLdLRjAR
4QP2ceGz8b9ApXiY8Q05ApjExOGqIpQM1hfbNWs7MwKOgHCpeugMPgCp15jQa0L88ym0+dFK+p7n
7qNOOeLbEEXAsYcAyrBhA3CWJ6gC+zQQPYRhtofHoAfodWoshrxc6Y4aJDbW0ShaHUxdfgPddbTp
0+eD0yD7eVBHHKsJgmNUvCXSFfFDprdYofNfkL9SjXPCoLTFW6B5WuNVxKfXnpWqbBtEUA3lV4Y6
kbCT3gVDXSiauCvQKN2iL4BSYBWR1t8oqwlStik6CDbI2YSP6epSNQGVk/PWhSsAKZCnxhTmovB7
BE79g9tybOqQPYrCUI/DsyN9Uy1QizeKf5d+lnEMAbUUb+AyIWl19A/YTys4VT7+O+XFDUaOYMfS
AFwsCjGpNbr34Wrtff8tgNpvzrqPtQOQvtebLsU8pVw2Nb8YwD7U+9gz4FgdgQFvj6s4mdMBdc7+
4dM9b/FWX3JPZXKsA/DXuE4Jdl9wwwoVjyLmifSJqJDXhfj/Ve76/gKJKBVDefwe/RLmu4sh3E6J
2tz3z5Mf9jrXhoRZsN5GZ9QdVfSE4JQH4qf4oSM6TFZM8IndSALp8JuZnYj9fq5ic0pWCfOmT3oY
UdoDiA8mJzPFhmc6kUzHdPQglqdT5buMP/onL+z8KO2nL3vxYp2NEhrt3jz/oK9ODBg5fo7srq0G
utAMcEhQEUcDO9s/RPKiYcNrrR/MlFr1eLaO4V4APP5Kt7KuQmIywSWc+FVGGnPEzcqZU8PwL+6o
fKs5/XLbOFRk8jbkjF8RBmFwjY2xaQKcBhAozzJLMibb826ndTdl4Cor/5A+epsKuomjmz7PpT6J
rDJiEfj+SCczqsKPSzD3JZplx851meqEe/vcb29FwybuRQ4HTvWtHOmLcv0lX4JgiI9zk9XNsVsu
mIiq5SHLkNGUbB3+VQN32Tn9UTL0EztqfU1f45O4vv0s5U6OCXREncxVdK9FnNkqVLlPehGVVhyi
GQFB2rUMCNuna0sirfRR+N2lPQwAogp6HBM4nWuG9nEQX/YyYSFkPNFhi1HxSsC+tyz2u0pPdBqW
Tz3BcYUYcJiIMvCFORSGhRwhs7OtMwvC9nlPG9QHX+/o4IuxTXE0SWm5gyFE7rm3qaENfB5sdoL6
BQluLUGcU66dDLVR5F9vLxNww+gcv7ugJRGA4oQiVpVw2XoIvb+fJ6Vi0rCqLjMiMM8IHOE4whTJ
QkdfnFUX02rBt6AzcnoR/vxbRCMEqQ3owOVkT+q8INx5sFAH5v+re24Aqsuh8vcbN56kFB0DkDI0
4Xw+IGJJUDa9civQ6QWgu3oRfYwejLvBH6iYhHZ79jQ/G0uyzNwIdm9iWZxpnblUdkT7cpsRR9qW
dJbVvQTxijCkVxo23TuHyszP+nr2vr9TvkHu0jZvBnZTzdjpmebpANUlZGYdhRIMW203+5TwUCfo
NZM7lc0FbdPOGc/M2Hovg2fW3A2H+1mp//NCuV1Y5rb7VXefzsNqAtfEvcp73VGs5ZEaGcCLzEPE
JYiCwpeB/mgoM6Fc5Xcsi6ebl+Zf77+bgTUdJLsulEVSwTxV2OfodxbO826a1JNtm/uC5qNkSCi1
sqwQzFfYmLz4aWhhxx9FHGu9MbeVcxP4GCxhMojedPm44L7XiKgaW30NKzP7TiNjW0cJeGC+sz2E
gY6kz8bdg3y9b18o/dpBjbftgnV1+bejZgk68KtGl+kYckyLzdzkOwvM9QQiPc3CeWPdJgEPadq3
TE1gv1VKjPyVUO5QKkSXkMOL7q74yNkIJsWDYztK5fc0EEX/TmdoAQLyKzJgKSWYKHpraymW7Wi9
jB2HCEftuMRsO3iMtBKFv8b6wo1wOnbKuWR19JQ+mPi5agQiKl8WQZHNly0nMGbAVxhXhql91f5p
XQ9+n6VNpkqTpmWY7iJAnqTUSwg5rgp0rCL6AEqJOHRVr3IUfQQ8EVc74PnaiKXqxoERO0OH+NIo
pyP2+iXk+dP+FqMct2rqG01kPQKYbhSpZgv/MfW5bV5bEsvdtU1V2NsPzARGSBIuiFuQIj+k3LXl
jOOWSOSl8GbrxawpLvvup+0z4sz6cQtoM3xkF2aPYeHVaT5/ctmCF5xt1aBKlkcQl/A7bGWoFM+y
IMkkiwe0NBLgnBgoxkYOhRyRmFbb7xJMMEqlMUie8ppvOUfJ5UCpZqQcHOrNRiErYYLJqSOou8Kg
i4jpFK3AP6MTzhMv864KJP3jEA5CZWzt8u5BIkO2sc9UPlWxpAlDe+E1uRUu71PLvtBwYtHQcSXX
Dc6LqJ9X1QBtwd8GERin0AKYSDFWSOwFrWAnze5ZehLuzK+3O3ECuqh6OzpPMgRAWAqlVZL/MdX4
5wRxba3kEvaHY3F+hBZzbZ3lGqiyr0MuIllSV9mURRSqL/ByfO5YlqABAqJsAU978qpcDDEt4XIZ
ots/37oBGmtLaaYrOLFtsffFmQW3NrNWKCbl15XecWab3I6dpR9IDJZCK4s28tPCCcc1Or8mciB4
92A3GS45fgL1TWuQ3j2xQ+wt+b9D1p3jK0oeEqMMqvh3uRaSaO3z+iSZwonzdr2KdGNkZfvhLBm1
tn1NoFXiukF5l7vAi4XtkKvsMvLOn2ZfvJu+IGw6Y9uAjPr5jSelhE3DUl8AGmTAdKuK0TDTyHQA
wAj8pfOq6OhKNrnVL4n5Njpwg7pCsVVYoUtR30l5rgWnLPaOk3m1f1qny922pBzpHWQK0CkJOaKA
+Khmfl1fh9CRhV6OW37DpL1/P8Mzitl5ZVlsh8kILxD5f3nlWlKCtCeNNGoxcb/IBabYcETt8fOL
zmR5aSyaviPvZdo8JtI18yncjqrzWrmVRbShsMxYFQ9yarWLTQtkrjHnn8hislHBwEz6QUsrnM2f
HjOC4/p7IZvHCjSSTHmPWXVDMNcMD90DSKYfyUdFdDvVCzJcXs5y2fxxwZPNgVjPxivbGiuewQZb
C/AR8nDu1KVKABrfCtkkaTeu4q8MhhnyBHooLSvLGy2WMMjJ6AHiudg46jVJG5OX5aaUvMotJuQ0
w96jQ27dc3BV5riD13tFMHzrb/fS5VLgu8s43VbEGYFo5Oy9pARBdMiKHjeKacxeJR0lXzOvIHLU
lEFxdb1YMNZnAkHrAOjQt3CWTWSNneBScRRlyEBSMFs9bwcCxjT5yrFmVif1iiojE8VCGQqIIBDz
nYWTX5EL+brreAjHlC6PbBR6qP6ZWkWzXxAfpbM2FRtCOlrjSQf91EEY2ZNyEkuueoqL5dTccLV0
sfVJhM0YzOhzRErTWpEE/LNahHJy3FAXsa/Oq0J8JgJXY6l1ycgK1sTXrHx2FZjCEt/Br20/LAi1
KbajfmP5oNbSr+UphTBCJLCgX2pA8rYVDr1BSoWo7V/uphZkAJTUURsv9Z+/oDFCA2N0nnraqhNP
FV2sDKFW19PgF/J6jiZQAs2GdmqPjuR6RthZsTeSrbjNaDaOB8IljKN8SJUXiua7VO2inPhWsXiZ
olGwm1flV1WKtTMsMRwevoiAPFVJyNO3hjxkbK0PIyWxt2R5hgPoZK+mXmdbLCPBDocxL+rAKCPu
aOD/aCXHfIQln9N1lTNzbm8Pr5DiP74ka0Yi9WORScN7zLXyh84m9RTuSXpRPRMiCgtVfjmtHEvp
JUtCOXxEwiAOJpytpzHwISjESUuYwTZboSEljFkMcqqYUNLLmbetjo9fNmlRGYKApKE2257tm9q0
srvV1S6g0kbvhWaF9S9Dv6VyBW4PyfrZjFuOD6azmFyfaB5/C69S6yUtt/NuoQMvBWMJoEGzP8PZ
jJxGjOhuMRiWMs8+o0zhwMHaFKHtPuSpLgBNgZswDNI1AzQQIS8jZ+Rqp2e817QYYPeKwXIbfFFO
3q3S44+NR47OipHoY1Ch+hYhU7MdflEgsC3VMDpnzFUYt+3Nfel8z0iXx2S7KPw/43Q2lVz3WsFr
VamRw5GYYajZ81RxVCWsokMYwSYspobxYh9h0sgC27VI8z1TaG2LGcu5TLtYpJ9VbCjOmcKBZzYX
ETv/inNkiYiWSl6QGeI2i5WV3uQmxG5YvhwbzHFAlE+L+rDnRYVYSqUZzIfNVN50U3PrU6ETT1hT
0BOVBmuwguN+31llm7Qy0KzwAPeDBGZZWx3bVZYPZyOCIb38noP29OqgRTpu1XKo7fUyPfkgWymT
sRYLab+6YKv6jur8RiUqAfMAwSfAsh9OQoNux5V7fWr7A3EKlWo87Yp6uZNlZeOyVYG8mKYnqWPN
um2chnyHlHa5Pz5Md7PJG5nmJ3ffyUcRjIB0DLIAfvtJ+1gvn1URgYyjRpcL8+hPhCGHw4hC2zlb
debquX3KpjGKuIGuSh+dbd4k46jOIYadPkYzukxelt9qwpX5l1nRtSMh/zHB39b0f141M0blwpJ9
Am8dA8hfXFaUukOwTMyI4e9JWSdzT4tjIbClZITelCFeDfUSglMaAuiliLknSfSLXKzcpq0kvNY3
vsFuDlVUsveUP0tOJXZ8A9l/ubVvbUBrVdZfLyy4GnQ+FNzcKfgMR0fbt3jl1M54f0gRwYz3YC2L
cYqWl6DP0KQxJP6t83AyWk/qRkmr4W5ecHdvWGqrSbweo43i6K9JKhKlXRyLJjDsq4Vvo5Wi8lBd
Y/UHCe3PkEvDc//AY017dVGe9uFYNVqMXyx32+YE8yUXQNzSD803NRQIL5ItSMwrgwfrBvVlcmNV
3RQCGJOv1ZVYx+nJW+vMWRRm0AH4AopkUBIYGMAxpO8aIoXwitnwwItLX7/vpTUL27b0x7V2gUEP
SzwwiJqfUvgYP0zM35S8Pippws2KljB09XoDT9kSdov9Q5x9ujpgcTLankkG8gi6LsDPnu13rDr1
iHuwLaeTWA28W4w7g7AAdLqnmqIt+/tHd09h1RabhwVnk5wzwt7uH3HTfOtGzjZAvKSRmut82ofv
LjrdJNj61uhcM9RO9rPdJg1x2UHgY1du0tALTubzXjd39+6saY6LWKpiKUsX8hbMmpvKczUcJIfp
WtT7J1rjEZOnGAKQztpTPFg7dkWHjkyHiRPsPFlV5w+61ygvHZBAmdb/OQIrWo1sAXPbWLad37/Q
yWu6FkemqMo1MsAsrMkCkXabYTO8o4lp0Zeb3L6iENja1+6K3NfLv0Hp4ciOkw4gKCTmZ2VLeUZr
+RblgoslJ04WMJaw5g9xv/FzQOWxgfH4P71uBDKmf8HVTp4x8ILxucL0+w2pHEmyN4Zrcdb2BlYw
3yJKL49b8y0Hth+za7ZpZNMBJzuMXrvvJoEfucW9cN4741jfAhNbHHS82nlZBuF8PqP6bqpJc5ES
HfG7MyEhJY1U73UpSmG0gxZumZTvyRlRVsXJx9VRQQWAgEJnjqcHTQslWtvT5kJmbkETTufOfBxm
vfZmgQ85v1Ki9newoaEyfx/hBaHTdJnq80BBqE8NMGq47BmazyWssq8IFVuJe4eD1jFPgilBNFjv
7Wlhzlnd4GshCdTysKqhDEU6sEDsoeZUyH83xfW6xhdHlRey5dbvnQi1T9FZsNjl+YjQimREhbLd
BPXWyXJ8IPogBV7y1s/GGLsYaETDEfWlg0GqaZK0mZslp3a9ZMg+0Iw8UUcNwdv26PkeDEnpkrNx
tnN4cVREXAoz/6b3HtS5T/xjd3rrF+tR072xLk7PJ0c6sIw00lA4QMSzf7kLsJDf0vE5ZivbF+cK
3+uTug9Lwb2aqjdU5LFb5KVgP0RQetv97mKy++hXfoCUtD1EkCHQ8P4pf6fuUL8DWp/1VppI6TIz
D1fZBs0IMbl7LnVDUryZfeEqpSRDLIA2VinE1a84M13chNPUc5Bew6Z4UH2iErD1pzP8X+FjlFB4
7nwO/GKFoXhw6VnoO8NKo8X3l/OR87XsZwKy81JIq+UzcnVWUDqd1zv4gdEvu7ivxTj8laRE+l56
0xaF7LGZM6rka8EyjZidsIjKUBZDvZg0SQL07qk5N2XayAUgGEqce4EkRXZOPTAiOAoHYAIFMyT+
wkR8UKOR7gx2W1piPJmI/v8qmv1O1IsyLo6KrqnBAP9f71RmNKyAQ7ohMT3vFyjNKFWQre7GZAPD
ce05yvU+rwbWHx9otqEdCGZitA/2vfk3/tJACNsemK3VpKYRwVriLMn8Gmwds+dkePDybytITIsn
0HxU+inowVdlkCMPNsUnjTfG66hjzZsLarN+T+UPZgrd23EC4F4+HOorN9qxMOAy4gLJJpMH3jdZ
+0Nr0B/4xVtmgxEofYCdPlqn0GgTVSbaWigLUR2UwEgxphoEc+Jk8wbHsSUJE2SueV8gaDJ8I6yM
kfx5dAt4l43nUexFLJneyrT3AE5B2DG0yNQiqUBmVFSv7SK7InXGaXpt0bbbdtKeprNKjanvPHx9
5qM7i3pyW4yTkvVwVhSIrnjn4/wT2RhDUk1Tz8s5A/4N3Rdn4DQoknXOOZKsrHAcc+KbBRZNWUzL
miPRn0XnT9GVHmwz3zDGkS8N7YUkB8RWYN38dimY22W/+IRDR1BaAkDAOA75R5/T52O7rgvGSE2Y
ZSi6PO/7YOpWBpQmeu+st8HRoc0EL0ovFLGPMxQuavHjvBuNbzqdqdzUDX6w1Yj5WWZqPoTikTKv
YvQPqFbMRJlP+PelMVfyGWpP+zBpDFD4EjQ+WCS4GsqQ/FnECot76KUOY2tusuboo1O88iA7NrVK
zNPZ0Y9TQ7pwTnCohcWXNNpFf0LyoDbh9TMExI/5w72Bt8jDi4F9jiyiRIA6vy7S95BUgVrMCbY1
hnFibNI3r228qV8yv3Vwo1YpFT4PS4nSKSIXM1ca6zvUfsHX9dTclXaFKrfwOyox3htdvRsvjiF+
y1WrDS2GzKXbz58iTaCcdgKwqu1XJ2FpXWotH2RdHzw45eqStO+7h6fK56kx0Z/Jy28EujbsiI73
xhoLJdFGMRm8OIMfoU+S3dH7RP2BVrZWUn5BIIylAchuvGsrX/HIZIkRSriky8W+HdkZAx6HAh/F
303J4NShr3kOL1Prz78RNIrxYiQ1v6ANoeXHzr3FnV965mASzjm9RlA9ifkVuQyjvG3nQuQljsvJ
ITBsaaTmEqw+B0TFKRlOwz/kz8gfDj9QL51Vi/c8/w48Mk0NVWfbr/EBrt8nIK2Uv5P/wwuIPsQB
JzK2pIxJbiMEj6pNCJJuZV6Zdq8apyoiNRTBAUi/w5h8kuSEXPQe9+HcFYw1CCSIKow7I1pxB6lv
r+CT3jyXEmXSqpS3USFRTOQNnH2hvQPXwDU4IbZ2S/ps3eKpO1XXX7zM2g3MpW8XWJ/SffJ5VKTW
N7GnXMM1ANJePfPoW2+a0e0KqFKttdMcM7P0J2coK5t4/Mf1y1Rdmua+XSShyc/Ij04rP8OKgs0T
VgFvfCocbQ5MihxI0zSBN+XsJYSXz2bfIhTsRxzQ+wjWD/LqP57w1CUEhdGE+D7a6w9QpA2zuuAu
pCoK5YmjtsZcEq8WT/7StGN7ILtywm7Xv7rnkRcXJD/9O5YPNfofigvQwFay/wPwhrUNeE2J/KWg
N+MEJEDD/MuficqJRD4VTRSJQQhBfqV1oT82uUnb4dUCJBsQj0oy/OIdZaL7vfkg5YGFzZ3pmqX0
YMTUp2D3OQ7d6kgrhLc4Ps15oLIBAKQjFzFIMFYjjmbtfCX0T+/77H24C72TlQ3uZkCFiKAHg0GN
K9W1Cy37suRQs6g2p1p2n8cYtiLEgIOUpqUSJaE9oEwW87OYTG/Ti5nELR5cLyaCS9pNlXzoUoc/
th8/V3d+cIrQmmYr8aayCpNgbsmLV0E4tqyMhbRyGVe7OLchONjiIWmzFREB3aWZc1YoFqATbXEL
a73nCIrn08E8QJ7e29Zmx2INhtY5vIGTS3hTmSY4XI5Ptv1kat0U4NIYd/khT1RTh0/4c0RcdpTd
7FKSGVbazEchEBJTE7Ec+gc93KC2Tou6NiVorCT35HIY31v3a6HxHDaEkSZPHW3nA92EQnufUHXM
DYNqH5FatSMEmM5xQpqKR7FLM8sPO+zRdRMm+o41P/+44wiOUoniIxWZYjGmHnWJsD10h3YmBaaO
eQk5wqmoaQoarWeiqnwUkFNOk7ZAqcI4lDqahE35/3OvuAVZ55G/b8BAn1indigti8TgOcdWNapG
IiVjeVrZySoVXqaQdCXp9Ju5GzpAL7mso2vrSg/XPSqxDQAOQ0SNQUn0GH1edR4k9I2TROyK4zMQ
ghDpFgzH4Dao1JO40ApW8zHAgsyBXJWgxZbRVLgzngnsr1Lm0KOvGFG0N5dCHWfwOblDMfsJR4Gt
3vOc2dJH6tqCA2rIqrguaZF5lQ8lzd9rAexAxyQqs2s17LMDJUowBRz5bJNrZCTZJyt7K7mDzruU
iJhuojYjnnwrEKhi930l8lrASDFvIZMnzvb3FBuLugQa/yASsT2TL5aCSndjI8Tji3Etoo3Vy8IP
vvoHdEXih8i/BBUVggg+CcKMvijlHp+8pAgZzDAoNzjXQ4iQYLX+RUGBYkTco497gNHG6cD844QO
egG0LISQcxEN4NatroAteJot2+rh8OU1ALT4Hu8bvSL5CPzQUnKtPX+oNpIXqzfjnrYjZ0BusciN
Qy6BIGhIPCPUcarnWQO+YXZZTweG6YCP26ubRMXzs6aOBjYpGbODHIM+CpJ8cAOEUVdXNOJLmThL
3seKmg/YsqSwiYTT5RWgCGOi2IXn4/7BRI2ubj/XWfnroAM9VtLYgkGN9wuhLMIVU+DoJ/JgJ5MM
9lmX6lAZd3ehx/d0n1zmtYn7yi6tgGdY1GSSjx3eFED0xkuj4heLdA7Yol26Jgzj2yrTR79Bf9hp
rZbRdporp6psrv3ONJO0xGmAd5c7sy1SjFf163kdXj0DNStv/wsMQGF/wOuxiY2uinlgT07L7pvJ
BxXcaWT9N1YKujt//DTbNgQmmdBXetdKSNT8dQ3bTIlySmuEfZPxM1Io95XQgnsjdQhhqxhB4KEw
QqlPMzJ8W4oGHZtEQJX7Hzm5OwCsVwHyWmXGmsTm9OGhJUcdeKyC9sMsn1jdF98GD6kHAhB3Hqwa
ylAAQFDOOaLziWTFJ4EXql/K/Pb+70VYN5R8cbEgcv5VQdxf7/Y6YD7+gHntVJe8ry1EURkMTjgX
BgHq7sh8VP2cE4OlDl1iNtS8yDb9e4b9N8oYZ8JYx2PRoiv+Ggi89P3KQydX+vUgNODv0bDNoja8
0HTRcqR8aNAdXKSREXDrjgZ4vFkYntxe+GnLnUX33RGK3NbIMp69YXe/sGR+IoZgNOKdqTGmAUfN
KsnqkI9g2Uff3LUKXLbiOSY56NqdpimK2kQfqq4Xe3NsxONIgNEokUbs91lzVBk3/rGHngH2HbxR
bE1D+gLrJcyfHJY0O5Csv3hER9/Be9szirOXwRl5Xu15tTb7wPadgz4YMGH4oj4CN3nERi972YYJ
E2pErB2/UUKzvRLqjJF9y1HZ/+GxmnsOffGr08/F2Pe8fQf4t04a9YnP49+SL62ZUoQJkuTsl/11
IdxbfR0yPvEWvTRmz5gsqy35GWAJcHu9CeoUygllS9sBsMcQE/O9nDX8nRp3uAMLHuO2DbP8oCy6
3pjCRRIrdMMzt3mCw4w3YUqJTHcIQMWnHzF9Da3GVEr3veA+3QeJi4xWHyv7er0CXmFnzL6azTsT
d1g7RF46w4iK9FcwapexXPmdgAivCH+bTdF7MWrmdENm4mTojB9LZW3aC9GI1Pfuu+CZVc5U4fV0
V7BLjK+0cHTOrL4QXo3bEMugTgJGbRoBXnHcgGisc6RttY7q803OMnemZJsrFyLeG/jpjlhN2dz/
cku2a3AWseTcY/65B4rwIg8YUyvpNweJZ1YnoLvRLIK9PMRnvBe3A2gYeoV9ZGRlmSOQepP9vGUf
8Nl+oh785TsaLPbnIb65spLOw5/mJ9dCM8F98qjVk47hOhvuUvaasGxA/Z/rIZ3EPd+DajqJ71fk
dvmNMwDzlbcYvBj9qCn4nsdLo75oD9dtzrfJNHUgvvCRMRejGv2awJDre1n87S41bCfgWu+5he1J
/7BaEg+/ct1oDqbzEgxPq9Dd7B6jDDQJRqYZovn0Abeq+0kMMoJPwXpHZfDIy7yUKs1UqoxZ3gYd
rpcJcfP9HmQEWJIE18l7CbN4gX1fu3V7GQeD5R9yOINVe/J0XDCBw1YHAfgWXmC8NK4kzpsp+a4c
FdMnUZTPX78ZOzCu0fzYAhAm2Kl0vX8a9nwpxDr2bSjzJwaGkyPfptBFdLCowjhvN8N7C9S/YFIZ
O8O/uwT+9N0GcVyh5kl8uQMxyqGnboM/hQWGqY2jD9AREkLOFjVwJAdegvnVa2k8TMXRcOVE3xV/
pYj30Rihyk4Y24bkkYT5aaVacCpKKBNOHD5F6boNE7pvBKIIqa4M6wJIKJXOZx7EtAuMADVt9S6R
4owbODil/H+ouxVRs2yObiwgV1wgfqR4/OXaErafMhXAX21g6LcSsxipyt8cLZqiitAJOZOYaZS1
NOeEzZWFsA8AyjP/lJv3UO/0Q+y4q204uI4YC+PoEjqeBhwpTgluXKnVmjbyS61atrF6XtbaU3Gi
gLICmomum+VmP+UlNRpHYAXKjkVqlQ7Fkkn+TYC8f8xaDSLCXSbS48KdUnSx5HxKswKSy9YpFq/K
cTFBtwEkOwW5DhCn6EDw1Rcc8YjHWDcgnI7dmeNhFH7gX7dwMror8XDwVsYT6pfJ196Prvp60/u1
fwRnScnKN09rIRMiIQT3/pR3I7fP3y2m/2vBxYRAGnSM8tkPXPqXmC1E+Fubsnpe86zaREXx33a5
qH/FtmmYJF7INlCKFC/OCAoJpkddlQc7ta1xZmAf0OlDMlQHqqIeS3NKIMkfGqxZcb5xOlxhd5cl
9Y9rkoXTu0tPNT323yQ98TdAETcgaag3Cv8XkjUFy4oZghs22q/LnpySGabdnyqe2P/SWbF8ejHb
uHEZ90xn/HS3QENrYRMv0U4Zcpj9WuFxNJVaU5PXDlN3WU6zcxJgGdhuCS15gyvqg+MSvy/vSv3r
ISrpgTo7RHSGjV6xIl18ZVkfYjmUoH+4RBJZdMBL8A4iZ3hhMp6EwNq0HwP98wW4/d9iS2+vEXz4
DXHTAsnmFQPLaE7JJtP4PdKgqFl61YYwnuPeHtZzrGffiNNARXwZvAk717ZD8VmqIAN6SgXubCnx
p7T1xmMCAMmX1ef3iIlEZveMT49JuVQ2SUfVOLBe0HN3P461IH+WL1PSCau3UaKVz1+J4zakAwCk
vzmZfShHhcvqMXjPmAi8IG+LFMcLU8hJh8EPCTHbDqoO9xP8pv315BTHgVSnfT1o4M9Lt0fby94O
5c+8DWQHOIYGS1tNFbTz+MKHw34IZFx1wTFyKKUd5QtwGXp5WXUY5wHWTXBRPFRXcdITlLFfYlGz
l2OCfTIjHMpmf3+8+NG5+MpZ0Eczq4iCmuCtudXlmoXydOxZWl1FRD5ncnlik08rcgaEM7Y7256A
ItAB/KQ0XLQC3VJv2204iuRC8I63cJ3Tg1JwDgLcjtSNSsc3hjMcraMFGZhJOvWZnJaKLX3GYcA9
7lWn5yxhC8qcyO/fz6919/JF2XV3pPtzdRcpRSzcrCQruOh+fnBmZebIndk/c1TqwMI8nFlzuPDM
Mj/e7ZbitVEL82es1YNjiFWDKgbWVhyvsbGsSOtqtrgDfTZW2h68ENaeZQXLaqJy9WhUjg5AzcVC
iQ8qbnBOKx2eH9IVonQT+SegJnCAC3UZd98I8jyzFQYKseHsnHXlfCzHGIkNzfk1izKxbzmRCj0k
fQ8j0pbsdQOm2Rx0QQLVIBj9a2Hpx9vpfzG/xCoTkROWiovQCIs6yCwmdpZDhDllzw4ZyQeb5CYK
aiLqqJuECTvG3Reu3Aa96mdo7V9gRUPOkiY7hqC2Kc7wHl2peKhGbwCKlccx9qvKQaNRTekauDwO
OEDFLHXuEJ9g3j7y9Ezr2dWFelevrmWlr8noAud/uN4LLWNc2wCbRjQoI6JMQ7KNfc6wPtwUGz9Y
1o7cGNWCiaMVzFZ2GkDQ9TKXTL/iHhRgEkmoW+u57cTtpact2y8V7HmE5WtajymAOa8RL6+YrUKx
a/LpUDOJQSErafuq4VkmLTtN/TTzAKlRdXd7Gw0XdT3kYMTWldXoSUT3r+aSJkmJDN4AGqd5NiBJ
q9X82k2Cn2tmSMg4InEa2J8/EOKHHRb0Jg3wk2t/JqKFZspHXPzSlI254RSSs89vDzXrUM0RQUNp
GYu7yFDVZL6zrfw7bu967kDRj4mbrbAuROig3D6El/vtUxuumAGGI+coMlzL1NPeFl1XAaV5+JkH
AFXilfJJRjSZWRz9vPZ85X3u4om0VufA/0h8gqxReMC27AebfnLFf5qvHo6dtJlE63eWPX/0JRru
z/pxvKFA0yw1D42GSdmsk6GHfFgHBR3a8m9j3SWYkAUCQvZhr3h1QClcmfxL52E02sMg+75tsa28
Mmq7KUe2aqZt8jVcosTRMzv3FHicEfg3GrTmj94aAPxgKIR4PF/nqmyniYbZmCeGvc/CPuuEtvcx
co0F9alMbDDxgFJiL/Ip81RCpXAhSAchl3zV4zNRiGH1kg3AvJdR0UG/nNFel9cNtz5UYg1ownHj
LizmsqAbmksnSL51bNxBef5GE1qxHgBo6zX4/3l3AUc3PdY+v/0PE0eRlH+NuP7x7d6Id6yxJhsn
tEyhlnQA3ngED8/h1VVEEwfYSBrFeZEzJyFMgNpucf0ouGdu9iGQaiNe1cAmNI/8S2u1OiGB2LfG
7pXZas/pbkawhOTPEXS5KkUXNQUci3Fo6u8krxNJmnRHfnnzNOj8hRdmHqwPKDrqlKNxuNsR4yol
KpGbGdi+rTd34DdVY5Ex7PUqmTVv60ZLoAnO/eYjk+cwZBHHnNNxX7Q60ZtBKoWMiKg8DaFnHoqH
i8FCpTkzmIs/q8z9TVD56cxk5XMOiHPyQVHG/MQTd+VwM/Ju63tgP3bfv2vgwJ4JnwUET91fpWZY
guiUwj/ZT4xYCniTzYz1yPZ78CZtFKh+V56BBiK8sGBafKhIMCEWA4VBmN2SBWhN4BEALaxU85gs
rutAt60J83HghEuCkBA3Dg7bxGqFIfRgI2s1i3Vn2P3zx97jcPaOeViXCEm1B1WokznCzpHdY6cx
Gbpbu4sDkLaJ3uG+s/UZWGh4Mr0r45SN8aGGvcCp9NriHD49SDkflbgcIrhn6OJhu7TE00/imxKk
3ioPwpBlwJI3ucljvK0OHRXHOoAO8iwBmBVTRiZdzTIP0HkA9WUVYJXY6Q3/DYBKSSPznkg2s+TW
jZIOp9ZXGkOC+3erf+ngdqHr6jvRsNzVxHdSZW19nWuW9BQzxC7E3caBAA1Z8qNE9G4gtht6Vope
a+ZhvT5TojzLym5giqzqfy4dYaTl5iTq/lMvNzQZb6AaL4vXXNh4b3i/efex8szPe1LvIeC6IsW8
N6GpSFYa/jORMZSKAKc/dWKALPB5N0dJo+epqsxdL24IGzhLdttvfRXXJFeHqjRdMaDugWKd9jQ2
JcHTvQXMXmKamGrPT5UxRCWUAQZL1l2uOKXApKtfJ1CJqxzf64uFNMTyEk0zIHHs0Ck8D6wZzwl0
sQ0NngJF7bX03lpPLO4wIL4VeE471gyk9o/bOLt91GFoQm5DlZVleuG9hHxi1x8szB54P4chuKri
O3Xro9T4el2JeKKBqP6/7Zq2Fw9zzWNOJi2Fg2LXDTgHE2PiL/CN6mK68POnNUxfzVARt19tRKwS
KgPlP1FFgu4/yzyr4hEOUd2fSI0UXG7NQRSF+qu6zJVqoEdLCzrs5pob0q1ie2+UTehFr3reMtAt
VpBH7r2SEhorasuMSO7vCfVClJrbE0rA4xDyO5VEoBZ0g7xwfg2aM82FA87PmCDLzHkvytNskWFF
HxX0jFmY3V2bC7pszVcVBfpyOL8h3/EQbTgdVkLYmER7f0WUWROPvTv056JR8jFuJSYOfanGNTPk
CFAgTibKlLF4yvPd+Y/Yqcx4mYfyuVtAuTOqqIuw+xnGLDkqdtsramdsXqtQ+NpxMxjrjQwio+UG
3mqBJjnz3nKaPoq2s7Vg+JM8jf76ZC/80y/I8GU3d1WYzzkIvf62+4XEghsiGN0tL2dO6h2K7d/+
p1AwZMnop3xNVD6SDArDC6CxU5ktSkqRUZJqe83aVyR1yhAKW/YaCUmR/nOq2WDhSIpGiuk51tji
x1PxsOTsgfKQc5K2e5aTjiELNpkXHhTRsYIIqSWbSDodv1JJSLGbTKsW2XJQfi5rYId/sMSz6duf
GYDRxCTSFB7uICpqj10Q1S2dmdDehcyb8WsZXTZZDfoOpWLE/wChK0hdGKCWnIB1PpbdtdkJLZMa
5XXl7+mRUAB4WJreUsg928b+RJOwTqCgbDziKorfuT+vhKoSMvQgM6sDzClgCjl4O54nOVNVR7Cc
+FqTzEmGL/PoFddiuvxt+gR0tg/WDtMX4724U/a9uDX820ZZn7qf8kcDtY2+T7FsUUpAMc4rBqcx
Ji5Ar5QEQPepqxl7ErPkT32F72x5+US1R9VKDbg0paH4OB6i2NRzQpThJsa1JTs1o51pksbYRRUB
L97M5vbEcAGNQH8ItcMymibi1ODoRoeu2k14AbguUbRzi/MUF33Ln0JRKZhRlwoAYHx2N0j8zrz0
6+O8fMf+F+WjhBnJLy6m2ZLLs3zca9JK3A2SSkuccTV2KQDK6m8d+9aR/xJ5ZRRQbSDiQwKZp0lq
KByxIx27FTxjYPfMnbmvJ6ajOh9a//PwY8Ss4YT6CxjTP4OyQOHSYizKChIAubHKYC+qrvmA6hP/
XkSskVEkIj4qyGVL5zERiw55rRBEGT/hC30UU77aVBDycTfjg8J5OudvGHI+dCOjKup0ZyVU5jAv
gQoiJdN9pf2Lj60XkqaFOGgrg1kYGntVNaNqReBjSDFqGB+Xqq4MYavxzoj2ZjeUzJhOL4L2Ti43
idQ410tqA9NOLOBI+/87Wbxi6BT2fa4Ltuq44cw6ItLNuvLnmKwdOwjDc1U5Nxq7D2Gz8bbvNDDe
57Kf8n3cmC5AMSDYckQsRhtUOrBDLvex3E9DoYyjidA417u7b9itVVmoDdtjJeZ/7ymQG2gPpAHy
RbvUCxp/HMK8DDCA5BognMXYi26wVRCSZ88bL6rr8D+WgrTyXENI03uUkNkRikHf4fUcTs/TzJzW
JXJVyMT1V9ZXVXQVIA9an5LaGc/nYW92fJCbNoLmABipPpLZ2531StFp+Ed0T1VvHdjZ7Cdpn6eD
oakVBpO/KDG+6PrCWSl0jVycPmapej9GhWZAHxCH+u02FAlhU8vOosACTNdOUhO+N0fG+Kzw9+GW
1LDhs3sYmVALmohKdprUg+9oSIAq2kzexHnVlYeIZRSOZX3v1MwDGwV40zCQVKvhFEEHFoNRZuGD
3aIYMCE6r83PFPqYoou3zHDwH5V7nF5silZC8DWgr5Q+bzXcuSlJI9HPh4dMA2LtZzP2o0yPhWQY
RjXAYKty9ZDJwAUwSlxpYTqicdnx/CuKfFDb1bqvmOAHRo16l9HKhGyK9NBJ8TzIqkm/mDO038/X
/tDRMsYfWlEDJg5x7tnpZy6FeP7faHvBPqUwSLLQ5GIgEoy/tEP6x+ydIsQ1HryqW2Rb9q4RrqvH
ffg3AudS2WBXauCIzFqT7tJYcyIMDPylRN06nVcxClg7DVkmEZFQhjStJXaD1sjIj8WVYG0oM53S
riQYP/g82e7xB3ZOGKhRFiSxDz4DxJDPBq73GIe5Af0wPlyTVzfSqQOeed5KcTj1K8yEG31NuImZ
MoTS3NGKWheHM4mJlPE9mX8qeRU3FY4elrBTtrtqyXX3osP+4aWuO+rDQKMd+VOFySuGKRjzhWhP
FfXwYK6g8mG5a/rarMuP9EsvPcS8bDsKK1isLvZBFNZoSZV4fkINbRBzRz+3HE1aomgp45HMwa4U
fOixRvWlT1ANDqjW4d1MPPzRAlKx9jBKoKBIJEtYJ/vxu1IM5lX8txhz+yUdcEuzXfcnH0vYAzTW
oWiQu1WCWyPK3uwNrJdDqFXxyoXVPB5Zdk786lZZiphmH1VweofR6gmaTlAhVKbZaeYHwaALB4qW
U4dTBZ4WDpb5/0h4st1Shx56++lZWQQwPnvXGXDoQwWXMufhnjSIvyg5B3iPYSpkXADzBcqaPvKO
soUCBEaLj+ap/lPh49iWzJ9YePZk4wpbM0p+rmFXW/SAD5xoEj+ixdaSo+dkmfwznvbb3p7gU43K
xK5C0Yqjyk8Pj7Z4DVFIpowdJ4cpfoqUeaXI9jyaCnk9GHT5SN6Ht5WyRNQ65+V1ZchPIibHZpN5
skCUKfNg9VtG7BnTOKUbGD1Q9TCc845+35ko9cVuuIPCCo8C6uo7VeRC1+xFhT2fQ7bKsasjmrPn
BN9IVnr/DOGXYntX0w1eMPm/6RXmUkIiNRn/b25jb1huU/PZznU5hWJya9PWE98ZxVv5X/nswPs3
98PdQzswsHYaObxCJiVZCZVipoHCGybbbZo8ZTUh1zBPSuFCMoxrYI4v9GtnYoYkHgq4vZo0GKAN
M1bcRRZrbh/uBuEz9GuEJDcQbVPHt3ei2jtpftLotqEOnUT0qedp8hgZKEB3F8iP88WzqQdXCd62
iHSyjsSVwyWjCmNAeRUouOkz34r+mx/dCWcvhtQ3CTwtw8kVa4ddZiURg0ic3qhmlD4ZpCoTssYe
POMrs2HtVoc5taeMS57KnBJx/qDXJ2SetclKmsrfKLHItdquFeJaH7tVES06OjQuUsDKDRxI7tIb
5I4vyzvi8casm1ql26EZ0/1XeTWe3BocLmLj1Wmf0Apf7R+/QT/3hq5yRkQYALSbYbzfeTyMdyDU
6YF1IoT1LPTWdTZPuugOljzZZcYERHYnqtWd4LhfwvxyHUGLxzfeJcO7N6Cm7Ug3Nb3zl2ZnTChp
6B8GnXY+yOEbn1O/L1r9n7A4vhtJWQAI+6QpaEjtMp2xaClLvCE2mDxy2aY83qEmW345b21KmFcd
G3nidUj4f4hlyW+3beJQcMD58o8LpK8+luymch6kfHAP44Vl6d7tSAwyc84JmvENVrUNP8bH5oJD
Q+lYCRTYcUHuNA8IccXsaibV3N63DFVjDPQgrq0hrwij85TFHvJjOwn2rBsu4rjSajCqoTL3xQfl
jV5ZB9ncEgp1Q+hdGgw5mekpAYhqCUgSUeLtJn/+IW6SGoIKWdgxJk17tkLDhzM5uk+HPhabf1pT
ahOx3wDUYpjjcSWKQXUXp9Gj/VwH9Yl+GZOIGbFnSJX27omJZGuswW2lRMzl8gJwg3jp2KfviUg1
fg5vnpFtFh31DHy6GjEXA9jWTsJpMy9BZaiskwSr2OB/CrF9n/jxJwt/6a6bUfJkufMBnZrkjHL3
yKUa3o4UbZCsD1ynmFonrXQvH3c+gaWSKHKahtD654PykG9ygg351ULbi/pA/nIzD7LGxs19CEMp
V0Tvn4gE778sk0DD1Cii8bG5JQ+OEAsApUaF0NFWZiXEMq8WJ/Vt6T4k5bQRKRfTlSNojvc9rd3/
hMG9VLNkz6GbndQp0wMp5y1knUqB07yDka2VW3DYcbKGQ7iEC044RKPnObXtT/Pjk1hRTwLCF4MG
Sx9o94jjiZik/KqmIWiCHS4ZGn1NmfhmiQYIrSTTmdjBUddGQXZEPRL6cL4CCq9EvwVJCKy35eQ+
Ai4SGuXCWBNpo4ClfMmG+Cl/zmHzSrDH0mpglAN6ziUZxC5gS2ixdZJ3dASr8P0kCU/IsMMJ3vyU
ZAcXN40WhLSiURAh2vLiNGyKVaUfxKFsvmNS8jpFVFBu+rPWqMREKmsRQOJFhW4bnbieCPvTrYB3
uGXmAYR6yJE8F5YcxMzrT3Q7dOuSeNhS8z/Co+do9mq+CbpSxLVpsZQcrLYYGJNrieGkpIUjZK+F
8xqAVHNwoIUDGrCb5eC56sj2t8ILCLmWRdgMdBdFaaztfagDFVF2MOZuRoT7nNtsKW8L137LTtb+
L8tXBgt8JkHnQCQkMuXh17tqlaAh9R11VCY7pJ2888eBmBq0sW1uKz0v7kTyh8B6j/osqcJvSRIv
KcjGtZHBb+I4yy6iiw2gSDkYciZX0dd5EtdLqO/tnbZ4ymsRa4OPWYe+RshMupqfMdqYmkzn/xKu
WVCbf5jxojQxsE3Qv5vVkrx8cEaotJwG1rwg+uklgVBO9oAJZna6tkQ2Oi4vptrx5rBBHSAF4rWp
p1mzUrP4UU0GVfwiZjVz9j+U70Ffck/DGUJ51fNulsxV1T9Ior/4hQACzhCwFBn18t4M0NsMkp0u
xdVeXi/wSN8cN6xiCOcp+/d7rEFkufLP1aLRa/lO65oCZ3Z1RO69mjWWxac4zVoyD2dsudj0KV9b
0lhTdsfbiUrtvmVz0syhwrBkCBQ1FnkwYOP/dJqbrOPLlMZHy3DqpmW05jIemxWO638i6aa30P2q
SIVQBZUzjnPradKT/WqrMeJhyFgk7O7Pe1Xr/M2toh3SGMVRXxsnBjpk+WIr6yHlKkgaIOKZLFb0
wVEzxOmERAhTJQKEkJeI0IzWiSk/t+OZS5h6Ss4UAEgeLFQChIcol66OmVbRWLgMXl8aVE9FBZeY
+8JBAFo/v5PSr+xKAX2YKkNmce4/U/7adKxKxDeSDrh779C5W5OVR8mdwnN1XdiDJnt3BQeTImz5
EU+OTq/xOyEVggC27pBKpKnlbilpWBUoS3s6ULm6qIaN829NJtDRWHZBGsAwoIzFgP4jHViYvpBg
ZPSotafIwMYbh6NkgBe+yuzwfcXKwKrGbCaPiXkjUOEo+9zWD7zz4oUWUUFbErdpjmxHev8PeJb7
3J5I5RQspQMQSCQn2UJ/0QBo3K/rd4mtuU58UIE4zA7/Zlp2gncwXONiQj2j78etjkpMALieM2ky
j7DToGuSEhmBuNsCiZD7C649RVKlul2PsxP6P2hImLnv+QmLl9szglLt5hlztHCZMkYvFvkewaYY
/2xJ+mzZZSSlEQT1mL8Shu/zu7OVfbBfU9sCALuF8bEmNJ2eLbpSKSnqqMCZIZpgbV8aZqtr9QIk
1RDQhZP7pZrh9b0hnmTNGq3iKPpbhhiPb/fimyMD22H6ZP/JOf/NUIoXRzAsQzUT7Hb2Z6JLpH00
g8sDlVWpIUkWPQA4wHb5AbWpxC807ti2VotPMvqPGAet0/TUvpbQrxv+laELE+UzUngBEm5JteKu
0arOfT8Smao26uULCEKiBV/54bTMDa+y5q8DBYblQOv2idjJrOyL4ZedvNoC36NGEXVHDnzQ+JsQ
ALaRfNn7+pBPiERo68rtovjjGaf/S6SqZJsQ84mMSzvXhIYggojAv5cmPWnj4nMmkwUkP/sIoDpW
ufC4TSmf9tqkufAlVvGYYWMCnt0pLJfh2L6YEXqiMtBWQYg0oU5QwFD+jKWXd57t09OE92k4ORI/
l5gY5IG74VLEt/Phlgesi24k9aBr5uc2xGIbR4P0nlavjYkCAo0Owv9EKAcLaIumTXfk7Fs0SRQ6
LfKvPugoPyncF8aCSmv77HIMXZ1YSxfjKmpMimNU+UjUzNVczeD1NxrFIssrG6vtoMbp+nN+JcB+
ls8CW9/EMht90C5BTom28xqRZUbW5xbqSH2yj8PwhcJ1zyhXotzp83HwSvuiw7xHt3P/pixutez1
f0Y/1Nqu1k9A+HRH4c11rAE47FNnisc8L+FHBvv4hYHmX8thNnpxamg5/FUucSPejlMOiaV9nAWK
jhOJwZSBpnzSgtDONQv6YCWCDczIeotrHRu3hQ7kZbRToNhOkUdgLhSQlpREArwnZkiWiPShfd+n
ALy7QrXcZbf8dN698OXA11Jh1XHHol/tWzaByAaBQvHEq2Zzkn8MtA46ndtoX7+YsCdSQBogeNQ1
+9vRt2WVvBbBoRjYp+5ioEmZoMgJBqlL0/p7UlG6zThlTetoR1mKutqVoSm+2b9LaGyZDOB3+Yrb
8F9GfafzWHxc+TtZA/Msj0VVqQ2/Ds0xEOtgkPeP/MTBmU3tD/uvFfKbCSHf6+uVe4kLGQy1BxaM
M+rC/xVJCSrzZ7URd5YpovA89PeJ1ple9sRlxKt09aLEIT5NGzAB7BMqtK0o8+ijCjE5Am9VEJlG
PWL7ChSX2a7NyD3TiLqcMXrMacFR0R/qslkcU0Va0lJNr/z4zcIt375O4+VtjCNYmzSc2CkhEB4Z
U9x787bh5MgDN8hJSC4z4AEQPzZE7LHCQ1tmDA1JGistR5E1nciS4DwipRlAqniPz/neTaBouDqL
7cgh98CdgQBm/OALXjJTcZOavt++Tvp9cEivN3yujQNGMvqBR6RElyc/lJZ6HJUXIa1kIWPoyAI0
BwnwQcIMpIC/K3rmr6Cpu14wGxj5H7HT1ZkzVCPD4Qe75bmpEIPbNjwkMMnrG17ZrsEIc0xXare4
ODvzpTZHeBin6W13cuRL6g2f/ldIG2SHSSQK6l8DYh6J+KdH90p5AoWp932/u9/qIcJ7R4OH8zOF
+2aqZx63dwCXJvlKHz1aceSKCGSC5mwb8NsMSBTX95qPG40GpRAdZuXxH34qKX4wtvTx5B7FA4hd
yWqaI2cAhRBAPlhUdBfCDXxliq4+YHn3VAAXnIfES3zPUDo6tUk7G05yPpf1rxyrYLaf0PZ3PtzG
JePvchZ0+mbW7ZKnWsVpvos9HeiFjSuwhrMVTzgwfYLud69uJjfJeaRbMQtKByutT07hPSomL7uE
YgUuqCM73mbQmn1ivGChamIjbAoL1aNgc1Faa5u81kSiKx6xkxJPtMXwwPCWi+JevWyPyVaonMKG
brGzyITaihijSMHyxh1lwrRYrxdr8sCLlsfWfBS+bnlP5t+q7EgEIR17/Kdh60YxREBsov5qEQgk
ZdMwCu0BJgTi5kfTldONr0tbrZhBcYHydJLde8xipJhLnCZ/kHrZy//BaKrcf2qg7UyB4YFK1mFH
ub93PhQsZkp5n0MxoWzwWpAelB30zAq+yI9Xk9IJO4vK0SngPHpz3mp9YNHbB2hsHgedJELlNUEs
whyU17+W6F4xEGFFx0ryn58tH8BqVEgcy3GoZq4jsLf6CqwVJ0Tn6RvjATQC0YKVaWmHkkgxvqkd
eIy4scY30b20ADLiqGfIZdw78CWPwYju+ZstXW343mmXBR62vm/NcVuAC5lWavEIxEBG0JUq0vdJ
kBrnQ7B1UO1zLuvSMe1ibvlXrG33WDr1tH0FtGw8hN6Kc6avCn1gUuT7aBvuo8bmI7+/dCpqg3+C
1nyZAbr1s/oNLN8tRHu46BoghIJOvg+hIkMx+s5n+zeoeW5AU95iAOyoKfQ+hGq7wU6cjA0mtd/9
6BbOfsGjzG/70AXO4OEOCHXr5uLX/GYJcUVcHSy0s/A0u5iHlLN+TkhlI/+jskdURxXknUcCSwfk
bcSvE9k2tX7EyC82W4Lr9AMJzRtR85LGZLgqjNSksZ60EYtlLNNZYYb08Wbo+w+ptHdzmwijPPyz
m+PjXue39d20obln/shLRK0mHpp6teVQDjxJh1Z0+8cnog/4txBuUQbmvEMdqrjq+cYNnKYF+OJO
ayggj7DG6QpTiKFvqF+JuFZPh3FPvxU6DrWMJ4uEugvSiVW/FMumBy52ActbIctef1hez4mb6NFB
nU6AqunFSQ2/7GOQc+EVIbD0mC9Z7eo5sYX7pL5Q+bAx4bDfEKz7CUeuoRDiJXWo9OWC8I8/0CZl
lNO/hyr/30GP6cX4Xn9WQsURGhqjRHlDWDqdQo33Vq4Ee0av58AHjl+vjyNsKlItDaLB/ImEokLk
AwchyV8corEaThGRk+A4BqyKAequrLy07FcAmGXd91RNWk3T/mQ6K1yy3CHSm4exWe+1gCzAwepY
MoZWZUbLcPznzMZPIFmpJRKcMS4ZTyijrEEsE6ioaKmabQSdQOOu1BfEUCJo5xnpifVc9AVOPzFa
3YyKC64Timd5iHI3tqS0qbr+OKNzHabWvDrf2xcqvxLf8CglY0oHZFiPEMEZGh1NgiS4StlsywgZ
GyohqTL8PvysLBY3jW01dHHVNWvAXpijxTyUMiNS7ypNSz/rU3xAvFGnzhO3xys0F8ktj/OOCg1Y
SjnH/gkAW+wb3yKz6iuslI4c2Php3R5EX22xcXYhwKro2EH8/2BI1WlszkYhd+zmY1LJv99ziHEV
CUewUIr6IoNGQWbK7LHjNl7bzPUayxD7UKJ8crphqda5h1jp5+qnQOrN6pLKkmJ1S6Z5Ep837597
XSJoW4USlHl1S5+NSVjBJ/XlbB7ijo+rHTJOg52xkwsO19mdWExMgxc40qFzquR8O8m7YkenWErn
mvs3TkRrm+MDguaq6VdXvNp0uLk/hHZLytMMWnRhdihPFtk7sSh+47+d4m7cWxvtKBtNpQlyZVxl
+06SGb+VIL12bSu5GQFUFkGAtaJsJ2Ho8WCMEWtXKYuj8YLiLDh+qSOFwiRn7xYMrBrBEk64lqxj
C8wvAh1whSEEZJgHL0Sk4Dz39IAU420b+fPnBpWJ7PPM8TRT7YNn42KtHtEzOi8PRWK1rbMZGSSq
+SZnPxAAET0JxeJcIcCHIfQz2OYvBkqIhv46WBTTU8M1nDhUqZKdZdT4YKfV90+COk7HQ0A1buv1
RidPP6c0R2ujbXhxtbHfgGlsGydUeYv9hfXjIXjt+1GPWRIn2nOLLtUvm6JsH4ati6JmcuNJXq7B
v7Bonyt9ToQRagt+5FNPL/wkwKAH8OMqILIUaPL0xgdenhJy/nMYXihfDIhORNj5FlcdwcoQTyvL
e3Zp5gFk5n+4kGvpkOoyt9Rs+2B7m+hYcp/Us+baRpVTXReqJ6843uYnE+FzmIp/+J1It/EPex3Z
G4E7EIO7PEDReuVXNnnlGxPHmsA8hgywxhyjxpNFhb9I9xGWk3T+qisPTxZGpTXqBCZfXJ7kluQ4
JuU2+4VczmxX/2Wbx4XmpU7Nlz6LNlnfYCbLAg5aOaa102WNUNBbu2oxKDbcZ3CFHAnXPL/iUDEX
hYgQLuinHiW4pmtQnka1HBa9OvzvrzNpPdmgMtr4a5Plq6XqsDK534WI03Qs4aSBtZCVJ52nvNbv
0m++sp65+vhOQCMyIbc+aMVYkwmDTwUSXOY/ro/xRH2N4n1xMNZ+K8ms0jbdJ954/gCQxnqThZy1
RFZ0tCCi7VmfPQWBZCVKyERqjDl0zVGdA++TjFKb98RCXCjGoC32id6YFgLHxO0sBr3IW1eHwodh
HC8witVOGT9V1LGFJZy46u8JgaH/2WTxCTwpfGoC69x0Uz8mLaNNvUS8iV2KJ40c0OvTF6K+vVI7
b1igrELqPia06qJdgxYbbwGyaACJuybfHUWHvkKXxDuuXOFLd4EimyJZCSs4D4DXT2i0j/btNcAy
Bjy2jGLhdpQM9ArRxr4D4biOCjnfVN/klyUmGQ6z3hbuEQ3DEWhEkCQO0AhW1O+UGjuj2vksMr2w
5MPG/54IrRl+5eVSOC8l+m1MUFYXRNnh8VnZckvY1O9oxwqGlf9WX34d0hb7o5xT37fbOZ8fzrQc
LTGwZuSybYU/SxMsnv3Y5my7bacFOfHk/shHJQTimhGI2TDL4nxFeqRdnMRoFKcMI1W8y9fptSwz
EMqapI4ks7Gaswg9JWvKPC0HwnIG2Vcu0bpFOWfKKJ1D7d04K1geh1fTq/gyRlOhLelgwB354qIm
hXkWnIEw6I7WgyZSWTmY9MLs0E09T3FcyfM0SQAeBkA+DhlvzJRiHHWBMFcAfiucBN5qZVrpvhPU
tYrFVS76HjXH7W0Q44uOLzix1gBn9mfrSizOPOobXCbHNwIYnMOr/8h/ilRdrQGpzKvIcVKqJpQ9
n/pqViYdDdlVJKZ3P6k9R8lvGSzZbe7TrtVfnBdCEZueGn66BzyedGHk8o4alJI+NpH+JXCTmd3k
vm9gXYDABrpxTfBNbj/tflRlf88Pws5eeVz3MM/skQ9Gs3VciYmETHsGXT45dxssWJfrSIayihY/
jGe+H1yJ1a/Ar5grIJux/ndAMaO/zqLoq6jcWlbvD8d9gwPxtlHiGXHc62uhRbm142Rwp2BylHYL
txt+0RlR86yxv7q6DRihYbRH75JQjBJOXw2DQrC6BIeZ4Oa+Z944gw8M/EOwGujkEsYN9/vbEWdn
0ljykKqRQKixXlGlk9KjgwIAhBO5YUfCKWKonVpY7O8UYKOWz1aVDI75Sv459GmKfubsLb1k35VJ
jykneBrEBIkIxIhRjCuZJA7+YC3eusDNkHmX6nxYyHQuB7F+dZKJDDrIcXuURxSTH/Jy5+IPXl/7
hPXlaEkjwCjYxP0Lze+0BBZ/ZuEGCDL387L5sRX03Sbc+xo12k1iavbNBJBsqV+fb4Y/5xtjl8vU
/lnPCR4MRb6HxnSrYUi7raGVnXYATExdZnMaXYr9veaa78rEaqzwN3fc/YAJK4HpPjmVDtz+3qb5
nG3e+5QspF55dXlyR0b/MPYeLfWcyt/K5JaVxhxKtxl3IRM29vDOfUOzYjVx9PHu5qWNU/JTcLtp
pv1l22bcLU2fSV0i6eHXx6nk6Y5ZaQxkq8GypMUf6C7TeFYyJL4Jyg6EUrRyp6FOAzrii3c0IofI
DTQzPctGpBhE7rIPGZxHIPr15wf2ANli8LBsFNuE+1Jxd/AnPg8lBonyKJfW62Oz1GRiKyx7j14I
uCu2UuxJHmjSTilvdUYWC5sKx8vrX6Cs/IbymLCTCCWfOGFajAtKSa4BrgyZVAXoklKi6DHQPie5
KgM7zpvL+I0k+M2GOpy+aOU3YU2LXu10zDjych2Kt+uQLm4vOZeqU9mCUyKdXN1c5InfSOm8LQRD
Xtk5AJKHwHZMl7K21VLgvVlNVEOnEp/n/e0+9372YVLqZ+YkQvQHC020Bnw3bgWUaypJzTV1tUtw
1dbqjyWgj57mamWvw1RpHLlUSTDe31D129hfDL+cRUMrPTRYWEnC9Iu8gh95/afqYPfGmuMy2vAL
nJzYU8pB39XhuH1AXDpNdLDvgyB/oKp9pY85Ms4rcUDHha4Tkh6VXR08TgWMZdmYyuR6E0b2z4D6
J6J/o32eEjlCYJT6cTi0R1EuZcVF+oI3Jtk/mSGJlH/29bPzErkntFuVN7Bis2t8RiZkzFSaRatW
i7sdq9OWG5wrKPKhu16isePqsN2pIFPDsIQvu/gQMpDaC6em6A5iHWkCMPVhcBX5c0zSHHtfGdo7
8PhD1Fuu5PTNyzy1Dk+zsNzebTugeLxyUstnbkB+eYy/pbj/jvcPdyhOx5vAAwgf1FKgwHB5Ouo4
ZEMBnA7YFgbUpl/niJQSCPCulAiHp+pApjrn3ZK8nxl2qcBObUt3QMksoy/Vh7EpxBC7I4ve7E0D
cwht4hWSw42l8lNxZ/+Ctg+qoYmApWiv5sDFt1KDI1Y6m0gcMsNgcTXE/RVRdUkoNkG6dTCJd2OZ
eTk6189nDQx/4gzqAUKgNU30yQDe5zYmz6s00a7pVCsNOBEN9F34wSPQ8ySnjBLF6/PsLFJTn5QR
6kwGPI47+QgBIN+X9ewAiEc3rk5YGAlCrS6koJ3Czok1mMn55eM6O4TMhi6yenwUN+ggWgVFTStD
Vz1RdszrqCu60mIZlnArMqQRU/dX0BOYr4BV4Yhvs0rpVSb3jSgCJp5Pxe+ZkNGPlcLvNUgAywLJ
u1fINVS4NrbGazMC5iQUAMQQSN/UEcZ/jPLVKMnoP3gE6ihSjEuRBEmMYEpcZi5NSyqErlrpt9U7
0RrvcTkVzT59pndOsWOm54P5BsgIxMMcy2SG9Jc3zw0pe5BZ8U/Z5cxiQja8TQJsYthNOwASj4AG
UQ3WyUwWtAnCKWRScPyoZMWFMCXZqVjWHxJtczd2sVkqgO42TZSAXHiIm/oMVWvmPhf1qhSkG0a5
wu+D9PJCo9MmxfoQcW+D4gij2TylXJ+DKzXtDgV2zRyjN35ZHAe9dS2yBFNGWysVFYkGloQLkApa
0jdPaWJoxsJB07lMtDo25V6RB9mL1mTDU7WOok2EIuao+MLjakyosYW5NyhmMNS1tQO4tq0ubtgl
puHLIjmoGdC6MvoiKMSCc5kB4mgqvkEwRrgHTY0J/d81fC8oOkEOfCMBb5ozGaFqz/vfoonp6zN/
ZQvcrH/K1scT4q3vvN8GyfzM+8Pk1EYe2AA1UwV7Ko5eOA2jo/QopItpmkoZi9y2lViva1IZnC9c
nYoMhUFfrdZ/8eHzEi2Vynv1zjpl0pdLalxbej/Mu98o+rOgluvO//PAbJ5AG5MrOUwaBA5SkvaJ
cV9NpZ1Ld1wM5xtYBXoz70CyDm6YM4x1B2hSdoBPkrRr8dIrdtroDBm45tj8ZDHV8fknEyotkaFJ
pXzNrMOJulITfQzPTF0dXdWHpZpLK8iqMUCq+aw8DdR6TYvyBIpO45uLNq4Is2oPzk5OdjcF77tU
FtxUsA2iK64MY5/HHxOBmiSWcCmtw4WWjClN1Zb3u4sRZDjF0wfpzAESX6PLEWWLONggyXvUiHPn
C7YJ3JCTcPeKTqIDjSd397ZXfN1nfHTST735LHlG0hNZJKZF7oj0Wb9gfX/H1YJgLgz7QJoL+ZcI
1960wn+CSo2DNSgD2K2AKmVKM4IUP15wL7kNFajTy6/SMBK2EMs/BRErpBsDN/shX/oZ4JBV3Z6+
t3kOeLCiOpiRhOl8roKzmCCcc2B+XxQFSuShabm1a9resUR5l9gdwYW2JVnMG1dySy3swKYYOVof
5LC5DlPB/zytqpAqNmKDZvvIRTl4y/xs20j4eyzZYMSCqyVyyqEaiKiAVX5WHqVICoj2tVF4HgU7
3TU23/AjY5GfJ1IROxw0Sn+yuEr3WdGsFb8zrIToS57RmxZkSY/ok3gV06L7988og4i2e458GI0F
QbswrZUVF3Evc8on5HtoWiSlzU2z8eZf7K+PNkYDu3K8r78SAftNysl6VdvY8vLqBsCiXhtkB/9T
yCGBqg3Kz3hE/7CQJ3s8rDqjyIabn9XRmfj/B8D/ra90jRUr+UxsiIdGUnR5TASPSxbPSdE0gd8O
o3XrymcDJ89+MpMqPWLYyUlJzIkhfzJ+i3NbBUPstIHymM0CJMaIZ14Qecr0wOEbEdcqB8xSC5Rw
qGEpiveJK10wn/v78BBPPYeA6Lw3SFlcVB0d+dAux4h0SJUdhNuFA/5cN849gU6P0cSjqpTtULZr
RTYtIYbGMsRCVfzFFcF1vQVf5rm76z/fh+YDZawc7PPM+zzfI70dksyybaqwHf4f+p4MP6fd4izX
vP871+8VNXxuacotyMKHJqrHAU2PpxtWNorSWdVDMpawEKvlwYTjdfSkoVVTWop8qs8ipFy6avxr
v+Ug8WRpLg4QcIuLNmH2jR1/52kzy53KfAgdRNlds+UISXv3QD9BwLaXurV7vodww+L3Q5GOXCoX
JfsHZZdjFKFATgrxT3o7QudEFQOAI+k2+4UcTD+F8yuc+LSvnSzpJjlKc6wT7YCXByfqHBuNv7E4
TQtQ3O8m/cX3INEdAaqgSYTpyQDe+/hfjYVQUP6SIAgvzdWXYqfYo0sF/NTeu0WeSh4aelpiSmaY
a/D1TA35rmHnXK3EzJ85OwcQBsRx3F/f/D3JbZ2wjKGJ9mx+8wquxSYpMwATVv0rC6Bwj/eytNEB
oJdVbdKNdpyv4mxP3m8xZH1x0OVCe4V7d4gxvEvFvYPNTxKeo1hiGROqRS5FaXTBtZRN7MhvFbft
XBrM1S2WNgGWczhbXOORxRzHegmyzBUwFkpKU406PlnJL0F8ZuGnwKHbdqB2+M0zBE5fTPbZ/Gc+
0Qdm3uPvXQDOH/qNtzcCBTDHhhEbywtUyPMSEPOP/ZT+KCk0CjgJbDUWMLGIcOMCbr5l+1POHtXu
9LRaXpp8E9JycEg6f5N/gwwKNy8yA/tZC5xL8Be6ysuK1GtB3oL+WVKfQn3TMrx1VTiW856XyPOi
AV33+0lgTo6yeHBbBHMfpiRjal8JJ5qsdqZucKok/6IJStt/K+osaCY8UvC8VSckh0t7c3Ffk2at
EZ9Y5quxcE06YmSRXeIOlqRBobLOKeJwmrEToTaiGL6xwN0evFDUNtmRwKrWI5rmu7fVcxFt3hs6
j5BpSK3099F9UlcpmPl2Zqt40B7LlnGYtQuuo0ZTj3USWJ4SemEQBStl+xyqMYXXUhvAU69YcKzb
KEAmw7sm3mvT6UutBX/NJ9iK6qSgDFX6hFLekD3Xi3TCd/iPyo30lsojMs8ZHmlAr+RGo5LdjkUf
BCOG5wHjsUxZs29j0QMN8BZtQxTLmkHywoTWmUQVdz1OedDTsMYvkNpQZEgsFagwXJAaEW1u7y2K
q+LhIXGtCoPYit3JmPE9Ui8PitmsEV2zHicnSOXDpAv1nmhbNORHrbheiQ5oz5dPbfZ1fZATXIsf
tbGCDllF4WKWnFIClmi5hWwTFZqIkXfaLzCsg8n8K6RUEttY3TD+noSGeZwuCP2NmZoVrAmPX0vB
m4OyJi0Z6+Q+Chz09gb7jtBULKZ3UTMcVPx4ibJw6Ln2WWS18JX7y/fkllxke4XtPTW2hffPfMNB
p74Is17sfzRLhi53EiHxVpDNSS3oe0BNcWiKIuhmZpMDDckDiWpCWLpZX9QDufR/yAFyiuuawhXS
VkRZb9OOih695uoa/lzM4PlTrYm7+GOQgBcyi68mu8TpXJpd/LNAu/VxWu478LYXFW+S9XArDVOG
nvfe5Ry/oio4EeWnnr12ElMM0tiEzySofl45wLewgmXsU+H4O1Cv6/vMQAS3iIjYULH75IAHUEaH
1vLxSqfkibolszLovuIIObT/AZh5U306+iyp8azToyHpOp9tu1HXM7TMgdVuq6p7enBNAusjHqL6
YJvf+aaO85YTMCLOiSeMc+jhgnI+q7ofbHJgZ2AcaxyneWtUJoi/FeEIt6bC6dwzbDUHW00tnVHJ
Rrvd9ZkbmwpKoUjpz5Yik0bJR8zqqsmi1aK53Z+JNVu6I2Wf41wrkArblff4wfKOE6B8vrDm1hIQ
wIszpBGN91zSnYbHkwNJ2UbQqLKZDL+eBphR6OnYoA/9RPmXEVLCQRTbeW1VJbXNbgqYB+rbu/V9
3IyinGTeQEh54SpgdfSA8JaIN8yu7Iq5EPJO9yu1J99TzBse3c9wgXX62tiZckIG6v/qRCcnMr3s
5eP82TScI6sihMg7A1iji1ImMsmzBlJN6wJrhHgHJtz0+eKN0LGGsu8efTUBnb9OFqjkD6QtLg0C
ANvUbachwrKp3KpMPK3dwRjlOONRHVrHiu0CEnfZGwY40j3C6mpBIdF6niNd1ouwpWu4SqfjsfQo
XO7tYUO4sMs45kOlZRHfwkuYUV1PdlPReyTJ3lT0UjKTwJw9pVB1teUgyH6wBKnzUbQtmfDC138J
wqUyOgbuIY0p5wAqJIGrNfvgIJNHhZ6gS4gAl+pr4QJQ+V3PO+X1t0VYPkWpfZfv21JuDljH2k+F
fxYge9LUy4FtZrCtesiDDW8s6FaWODIQ9fjiSelm+XaTs2Jeooj6wZZn+G7vvozk0qh3K9Qk0h+g
7TO6P5DHamaAzWonUuZ0C31TTrcebzd4kujtcSZpFa7GmwNMxEJckOKKwMNWNQhQ1aT6MJHeg4Gk
szLjOdB4eSMFMoxouZQkM40yIX2HxsEhKtTQyL6PbwCCuZzfwfU69uqv4FH7EGyutTjEKJUT2qym
9oqBdvcNfuhsqxsaZrhFWrIh2YVfyvYcUyTN90oR9rM/eFlvmM3nu5mHecHoFJrcgpAAUud+sSun
TVGdJZ2iMUbcuU2umIAA9myj77DpkJfDKjQUZ7rE7KsuuIdalIZ7uDFlCxwE4bVxd/hFb63lv+UW
i8MYAY2kYGTfVTxo4PeaRF3AtIdvPoVgIF2eEiMfjrljdbhHsxapHVK7aMwe04+yGj1ni8gWG687
vfDCqg3ezMziCEVTlLY8sG7IPdxIWWf05y7Vrs2lEFyZTAik2xTJJhw/IViAVwtQQApx8IsTdWQj
ewv5sTiIsQW1xARSg9ze4nIjUUeUzsAc8dl1vkkHP/sfzO9qn5Uqq7FP42Vjhxhh2CNEFiNfibOE
eaZ//42i/XtspRje8bIE63RSA3RTVqGd1pWvac4cZOSs1hQObJXAh9Y9AFbFesWV+1Y/fPQZOJtC
45fsKN0RV8KkRXuQCVEJHiiK4eHedDqUZ6i/QqRrnKwJTdorKy6KC1ciryWWZRaTw4tRvWCGPJJP
QfIIwHMg2UMem+CyMKXf/q3v7ZSpmtgx5ZzMvG2CSfJRDJXT4l+c1qhKtlczgYit4AkcuEGJIN36
QZ7HYiH6ZNq8Bl8jnm2o7rFiCmLmz7liewB3dGyL1dOU3200lwxjtaL6SfXER+tFpopOUQOJjeX4
H5nSMJSujxH4EqgwV60n1FSHW4wRoso88s3GrvHIKpWU2NUpVbKFXEpny10zSwSSo2zDmlwhFRXr
Ic/k/VHc2CaYMS4k8LK8Ctt/vCYJw957xTm/pZRtSn75FE74sMuX8VhuftqhLTBWmEj0lqrLlEbj
6WK1CYG12NBCB1bXEr/t7hIcE76Z6mOuvq/s3aAUjHbGc19FnzAWch/6/EXlIE8nkIqR7a8FaKTI
9WpZNLIIpqaTm42na72v8bjNOra8Vn5KgMwa+rf+eoV0CGnwH3wY9v4yV4JrSBUzQRBfv6B0JIQ6
jZGZ9MTBSazD+onl4APXP1m0hFxIGt+BdtBr7qFaMsb47xqqJPrI9kDG8ubbcQ3gIvBkZCEFeEVC
+LX7o0dEXg3aADRQ/fvnUOpRw6yWsfYymBqR8J1PHETKLF7s09AjElK9sr2lQkCUlg5VK8MPYeVl
uOJQJ0gjOcREKzfrwx+rpneImpBimPs5XN1eCVzQ4OmoFTXDwziqova3ShewCWqAUYsSd8mClu+w
EQqhgJPA5ykIQB4QD7tBdjdlvjFty+jBUrhGd8uEALoLn6GOoPR4f6UUcmnwafXx1OSRQE82yVpp
UQf9sdyb8bnuL2MnxfquHyVtf+JtuwsypnRZWoUM4SmKiT04f0Bt9UOEx9QkxS64hpPj4oyadOsh
F4rWT7FFZ3NyYRXMMNm5loEPxrrq+MGzyeOCw1QsFwp82Xm/fiHRSD4/N+cZBo6Ts4e5M0o/J+wc
bi0CQu398jnyuL9WHZEREVWoXn7zxXZKouknreqqsC6TpuOj5JuZErYrERpDZF8zUnMcFvdlmKBA
on/YnV6Nx8q3Mzma750ZSTDaSnzLZ7Vqk0Ykbl7jyVAKeNEC6LS+UGggw5mzT5ccYbpCRLq03v6c
QA+HetmxvFO6N0+Ii3j0cfB+afpZLccaxZI/VvZc/MR1yWOkDnCs2WY3qv+NeNXRFwyLrFP6E3Dl
eDubz8LUkxQDDn5OLKStPzxhurR99XpNE84FGi1I3edrvrF+wcAytyd3YSSBHXNyDUYwFWy2j8pd
qgvUj/mu/A4wCsnWOMm1wWhhYIMvWPZDyvkMJM7cxXydR2hr9xD9EoWFn1RXiWVdFKSVgCxSG7KA
NhquMsBPn24awI7SrRZOtTfk4bQcWCG4IKBdnB6gKhquaOmlRm5WoompMG2Un7ZsxQ9w3fqKrvR/
FjSTOKXhqqOXFM17tHk8HwYqGVzG7EWolt2mmdpv7KF9FzSsoTpnbwzHLN/7nxUHRz1Dk9slaevy
OOOA4tYH2BetOaCyGfmSW6bN28cp3rwiiIsKrDDXbNOIqj++7hdq3eo5201wpngaen8tnM/n79yP
YuqFR06mefdX2oCpUMXjsN0aKUPxB17SQejioAcsQELCWsRri/mYr41m/mEvOxuNtsCQ28X1Bq3T
CplcLL2qO8CehC3QfOOshqfBREVVTbrTMxT5CGme0gbdzP20dvfXUA+30dbhcAcHV0eeeastnozq
jE5qBVKytXmBeEdxiUg4pYvt8scSa+WOV7ZNJE5dKqN3yALdnEFnc2pSYSoI9Il+M2VZ7t6A20qA
kYQz4kfzUfieSm3Hk+C7wyJnPc37GMXfS1XE/qbDH8YdfHiM1SXH0Y0MZ6OhqbIM7YEbkIBQY0Yz
20Q450CWRUuHvnczCrgB+ldthlcCYu4U7fWxgViXWIX+QCk+w26x/1LF3UHfp+wAqU2odw+LffHI
vAEQX4mQeRUZKUL2tA9UJUDkf4gdoMM+hFRidmyBHZ3BWctzaszeNKIkLmDYq0m6CPTdQtduY4XN
GeYfOeDnA5dzchcqJvHOKNk18jqyghBqM3ma34t1hrC8WYhfrmWZ29vukR84SqWrMWO7V46X7bsW
yEqEHDnCVqFTJRlxCzrNDWL/Jd21zRZsL98miyug532gkE8XvzQsVZV8BnlDVobJ8TxZ7RcpafzH
eP3X1+YvXUPZC4GgTUD9hHMyljlPiNptMkFANPbWqFiu75SbBe/o+I7YjB3CjT4sPh065mkUkYdx
dpdu/zXL/5K46bZGOmAbe8I91r4qgDlnD1aAugFEHhWf0moaMYA1183xnKWhCTAPvsE44bTgggHx
DhxdaknuShrl5LBDURwg1MO2yz5VdYXUengdNSs1cIP8cbKstsJtaPdtb5VT08IKvfS7pmJ4kJEv
PtOW2eky2IMbPMbeHnss//O+1jCI63eT0GNr0InU5/Wd2JsGQT03HTwtmeLMFi1lZAJfbBeAn10e
OaWx0AznDpze80TUSLg/92MfSC00YobJspo3aLMX+r/Xn6S/qEoOW+CkIZNUIqC1Ua1zl+6HJsP5
svOnJ7/ccdUTNMkadwDwZxbx33EkdjiDAEqdGCokx+R1oUKSCHB/CyI/8TTaEEZ7hmn8VmrLqGNb
/K0F66ptsgqALzvVdhrRsGOLMs7L9fKtZpSDyYcxjApH3zkOEGaUciZnZnLL534cbaUSFmHEMwi+
1fLsPJ1hokjYJxakxXImyTNeB0zAGUIzIgkLTlYTTSPfHHqyqz+x4XiwT4vlqnbcrj+qYRSt/l5s
K0PkQ9mhuwNzvZFUF4EhafroGYm8J6I9p5wuiYdjn0xRKA/8WZxsMrYsNVmKdk68HjALA4GnQJ7v
q+TRwBqkdGZ4+Ql2wGfnl+MaTSU6L0JD5d411vlfjJBRN1ebu+Kt+RO2fiRv9HxboPl5pXkrHC/3
k/lqocw8Vc1ChENXC8pxXMSEatkgMBn3EBksRrrg8WoNlE715iBHUNGek2lewwYVrkEb3c9272YQ
DlziPJ2aQQLZu9AZ4mXhFazlvrjwQZjOQYrGr810HTjYbEi2V2xSPedCIs9VTj+lW+O/nceGVe3g
oPazZIKZF91dKqb1PZg2Po5FuZzgrIY82GABbYhlA7kqi/yGSA/jIp5Jq4BWVXlkE8Yhs1i13PXU
j0Bc2mz1beU4zH4kg/ybe4Z78KQVFvlInKSQV0Vjoblv7qGmkfTSFy21xmC7OuYySNYFbVYwec0d
GaLJsKMXKQOwLsEQZx3K9ayT3FuesUPUMbVVJn2DCSrqYGArrepSEnFboVAL0zxvFN7pxVWunC/j
1KbpogoWqpSue0UMO/OnhKPT4QR+E5aYK9FvffQcboJ5ep4fCbGd2z6KwZx/fLk9brncp6vQHaE/
NVoiQDx4UnX2pAPvPatBOiOU7/lvOhnTZf1BT+Jifrozj73PJRL7PrtIgNYESoXL4nOG6l07aVen
hpKKj243jezCUd5MUipoMb335hQosQooQZEcYhhYtz/3DSUvLG6xgyBDQK6NVnrJLiYtHOox2Otc
6SZWI32JamsrWbB9yWeuc+u8Cp5tGWIZClOHBVzSbqmOc5sq7ajQ3aiW91JGtZA8r47NGqPOw7xk
n36IUqS/dm/vfYKvUITpUWdB3W+14BwB6R9Zmv8pV0v5sgdrUs2u9UPZpsKD/HdnlpJpAZ52S6mA
SVOqrI+O4jcTYUQjqRb2i3V7tfPphqQQ+v1OE9N66hkXoc12VwaySkRIZ7zbkMGoOnakfvEctd6Y
giSqLJ4poUFg4CzBvR0UmW4PE9K6ZdaZW3pY2RVejDAqiz+Rg0n9tCqk/730it/xuwONgOZ/cwou
jMlbYQG4bfKBpmk+I0aJnmOKhcHEiBEAzKFJKAteXPmwxZuiu6X229mWSag+xjJlTUD0rKmX5aaU
N9rTmrcnaauIU/WAxwlAVGQFRz9oFJcJAFoDlxoCDmNM3fB6vvsN6W7CqUQbky/XBhm+Eqm9dSbf
ZYek7XzLuRzc6ZkXFb0ZhWbg50xzreSJkJRkxj8754D/CnL0id2PccDJ7Lgt/2b0IGDAlNDcOFvD
IG+K2gklBcyXAVE1WVQj3AeEoCkMJZtLpEpd8exzj2cNhxZ/L1HievSN6k6kqHo8DP6ax7xlIvj4
ZmSJngkFjRE5F3uP8naJ/vngzCS3Ulcm/ZBtISk0ST2GlOxHhcCq37hQxGg0R5M0qRDoLz41HuFN
Tv0BgV3g39UwsMxhAln9OqpYfCPkWQbYRO+JW2/jytTjsIy9Jjt1mSkS6g6TvccOSx7RY+jqISxu
mlEfCBNtreryZPYd1j0ijK9P6USY3gGO8A/zSQYLLsPIeHTz9vE4HBQVF+K2d1gs8ix0pCGe4NPK
4BkWymuj1zzu2wQ2OfgGbs+H8Par5kOCMdGatkfCH2NTnfhO8U1kmpOTdMYKNrjOkdOhRHbzWSQZ
7ofZE411e1O3EpNj9PpkYArv2B/o7iE3VkIgCvSkHvtE0d3hi5H7LCyEn9fez9TTn8/3gBV0rHb2
to9bsDh1TI42NlYhx2tF2fyDNrJyKAf6BE5Pq1GWAAes/pZ1j8a1Ax9DSwUzCBSR1A4XvuQhH4Jh
jT3FL1LYwv/h6goTCZlBPBizJzaQiBngSsrHOjp21TVpuMlnpDVC3tP7ScPI+LN/4w/Cs4m9j1jt
tDKxlUxfsFrw14gejfRgQPiian9cBFgmq3xEk4QQc79CEsFWqyACC0vkkYN0RyVI5ZwcgqepjLaM
B0x3xBKpaqB3DfydRDpg/+0XxfEAfKoEhGtFnLyPYRUqeZLI02HnjwzbgmBYO/rNJ4K+C6Is+CB8
OTXpHNpm6DVAgUYXv9qqQpgVus0EebaAB94Och34+T3+/hIwqVu9zMuLBmXmop9Ex0tpT1BuGYGL
qcsaRaa/nPpxEQ+ZCu5yvqdstQtQteuPWUhXbwLAZXVAFNHUJ8pcbFPfTlWj/7XJgdTmB/3Q6X2A
A4n0bSGTSKOzldPIHgBV9muv3fNIRZmZMbJac1ZEHzFVRn4BJcsMlQmFgM4Bj70InsM5Jgrh11Lp
QTi48Z7f7tnxbSWmljn+6AlPYvjQ8gD3QWi5nEcuCKwDh5+/HOnd2XQfXbJiq10tFkKvNs2o919i
uY0NaupwKQOteaT4EklWjH543cgfsKruGIVX8FpRtYLx4jBjG60ygleMYFz8Lhc5r37pZigJTiwF
uBUd67vou3OYE4pqrk85n7eZOdMh4G6pK58W5ZaAswZYorwOfFfFoclkHPOs0iJDn3lati60knQL
3f9yY3m53DUPIUWjtJMqZj6/L9J5L2xXbw/QRkf7VeHpZ5qOebcc/bBPRZB8PrDhT65zFe1jPo/T
0NuYOS/8EltZFpBngM9xt0fkSERNUEYKxpzuesLg+kDxHGjQFB4EsDEYuaR3NLxTY9do4ig+5C4b
1jWpWyNTMDdXMSQQqCShTY3gy3uQGuej1sHi7E0pqx0jGTz3YFswGyUMApc31f0r0wpmqbDWILrp
146jekxbEoIOZixZ//sKxdmjQPdjMOc8B6BeY2jz6XbjNZ3GIi7fibv0fSbcPWwa1EFobB3v26A4
2qdcMdY3mJilEjJWv/+TlTAz6O+W3FedKon/07R5Eqq5TcnWVjsTxwBHlT/SZcZnlSFYxl12mJEZ
WClu5yOT8pAyr6HRAgDLOIbsAxZoxZAHdjcuqIERdbOqKz9sGeBGkj8y8PmHNCLMkMrCiwuwXOY9
0GuMayr2Reej8dE1uUhayYC0y+kYVPBuAwgFKFEnr1Ap65iLTWoOKFMFnYQ8ZUPom8I8/dcEB5+c
aDVfpIuSh73pEMLzQjjCuCbh3TUq1rdj5s1tQWSFN7Um3qHWJXEPpKJixoQGJeYfx9+BitsmjsFs
aLuFHfc4WPLSC6H6+Q6N1M4BY0kPZWUtrtlPzjdR9frj9qMW1tawA1JQCv9R2NovNG5FSJkU5QeJ
S+0uxhyCgfW6dtKlrwcQFCHGSxJHrVtMm3Mcy1sWtsghk0W0eSuWSal6Ma4GMfqVHupIz/u7iNBW
4QVS0RBRdDy4h+80T1u7cUfKDBVTKn8BcQDkbQ+eUoGO1JZMUveXXH5g8BWKAQvYgMvFkLXRO1as
HktM6upRu+C1ZzCGi8HgiLk4Yu52vOwiPXqJTO4KB1IeQt07hdeeFnxhXL3FXARjVRL9N64VM4q8
/p3OAY4cx51TXix8HYM8PD0z4ugz2ghqEDWZojIMTt+cV+3AvRQpVp5gsUkqe8hlHzVZ2/PIfLmp
uPX9oOjTemzgxiOFrdiStsYzKPGK62dKC4lODdmOMkb4ok/qCiDmQ42N5u8GZ8zL5igw9/voqlcC
OOpaMIMsNO0Ob+vay+iIgjyWGmRk0i42NaUmVgcuzrxubctZ9fVGIYoR3wNfATPOscyIIcS2qkiX
T/sPBoL76Gjc2Qi40JWAg07/rmAomacoJNPwuiDYKxpgn1uvQjc8kiRjM7HZGOBIN4BEYQcPSlwV
i/GS3LeOi+vxy6ta466uUBJlE/D9qeTl9fyj7ad+afccQeO5J/AFMVbDybqUZuTc317Z+sdLIlPY
TDXVUhu2bwYjLEMYhtv2AMUoic3gVAWyMFnY/uOgTQ0x3B6/1F4k0t9AMunr1rPKwVBe52NQEJms
MH1Q4UQJBc3l9AFGCO1iXms/ouCBFX2uUC9g7jd4/2WOGsahKMcpn90/LV8j3jue6tkyP76jHroV
Reo6zE2dylNYVMq3e8GoW2ABiakZaeQ7biYtWoAXRuWvAneljtU0l3na+jPpOI5tVPHEIzWJvHHN
2GxjhTAyUgLLM5XX/pJy14C2JCloMSUpn29Z92J4BqkGF7nJz2j2gCgI46VcYLROk1HaHD77P95x
a7QU+GmNiSjYD+y5iST4kqpYrCKYyLHm7b28dOxph14NmPnMxQEE7aFWe+xBxerVSjcGOZ/qDXMW
ZgztjjR9EwaZorgo/CGY/hRnsDN5I8vOi/xxzZimtVsdU49j0Lqke+v+P75kIvPP/BVcz9NtC0rd
MzUUTHsL4+XUwGSjDpKkjuPTFrpbt5TEB5h/agSmnTGBwZEr9xNQ5SetGdBPW16MqKfzuSNtwsUz
wS/GjRRUnFNEeJ31pplBD47BGh1nHzWteHys1MrgzQ/1IkGa2VWK/tn15TeAzLloWnkGQrWeSsit
K8Dg68i5KB8sKaRfGj2SZEnFT04yFhuWETUBwOi0h1ui/7x1EPbzctaQC/5ySAzoi6HwQTMMG4YI
Ni/F9vE9N01hCjQqNMSmSek1FZKMQledRnT3BvcEs1to0/IVtedqerUsJJkS2vXqvIKHQACKOwYd
Sr7nrMy64ZHFbP6wD3Cpth04tkr/bGAVVxiM9+HkFf6OBZTLXgOMKWBY4AnKsM983uZx0giu7cdC
ZrXc1IEbb38K0tWxfzIDi9TM26u/gfm6bcrYeZrxX3BqbbfodVqxPiGb5MGCu3UjE/+hJ/lLisl5
BqQPVV+ENxRCz0LMyFDY7UveMoVCBWUaCkRiuE5kGPjWW5Gxf76Tc83XAt1Ni4JHLUaNGrf5sQrb
uH9WrjDMG6+pVtE5cuARApsW6yRXOvG5eqfw1w1u+brExLdZ6QTB1VnSCBbKJkuRIlBxx/UqjkfK
Les1/KrM6acUM7NDMInsGL8U+wC6Bg93Lyj7JDS7OlaniSyCRprM06tULUSXJzNUtItbym5dvCFY
tYvVcgSKRUU2TKt9gfO9F/f0n1T8pXh68xXGwqDEA1Wwkt01I0r6/o1ZR94oGurVhaIX5jxosAsl
o1hsxZCYAfmtEfHySUvT5aUICMWKHR+q2OJ5xVR7bHYI+bM9S3BB51a2m7qKMuQQxptJS/wlI330
v06OopJXO+zH5hsPl5ZGZinNbrbo4dfkAa+eHovJJyqI9Gc5e+pcZs5klcQeDsr8cX7aaPo1Pp3V
6SNdAM+06huZPQOxOWDwrtq5azqSbLuK4L9R1QAZfuPaU87/3QiBJPnnFv7FG1r2LQF03+93ZUq4
f/dmh+SQaraZvdZ78Ls5Ilm1veo5bf7CFJD04VYPzFYy5Dz7yWj3OAzCCzyb/e34daAppEgimtqg
/Its97rAJ7YjpRAJUEPlXw8XfLbbHM4zmIKDFkR3vSX3ZY2BLBsxHpo7g4QGFB4vllCtGz3AGyRZ
8EssUsfH/C8H+N3Rllnepoc+f6tKYFb+EP6TUc76rOo+5t5iF6FN8qSw2ZcXXdqf5QF9P3MXYdIv
PAXq6DFiNHNgTxqho+nK5UAnicD5b/ApunutrD452oG3krbfnJ6QqsvMYwGft6eQ83RQtzd+W5Kl
VbyYGylhbJ8z9xvwVi7htoJ/4cL9YVg3WvtrO1z5EnirDdfetNGIRMTAPLVCZ6cm/9obG3Htuyh4
tMK3MY9TbC057fCFAi50MChKWIduqRS64o3+FxMnpQUfC5T4RQHWxSBAst36zBIGPRjXO8hpnCag
61uIjdgFCAUDVognO0Qa5MMxQbCuadMyoOwRwQjualqH3eYuIR5MJ4Y7zNjR3nHIDSKE5l/9edOI
aNKI6LPhs8tJvhABKkpb3qWevFjNOs1aa6IjUouYKC0Rsqy7NfIqvj0B5xcVQ/EdUMP9lI9JbUo/
X6xNnHBLzKpq1dNDVo0BEuJij4VlVNB5UiL5Szrjm6ZDfcm7HhDE06XQBsirtAM4F6ZkHNXkVA3r
71+IkMLBxmx6edaOPZ+vTizO1+dv4CQrzdHZDSyDHTm4irUjg/MxctpOMuVIpA39PTzfp1ct9KzY
1tPDMcPZyaDi4Gxa10NFYsvIfu/6Wp+mvgThe3NTWKwCeT2LLtQ0Dn0kpVFZXM+lmwAyQAYw8lPA
6nHhdTHzrUUpDtVwsalST8l1JOHNMT/4cjDRURWmOj1icLHYay/tIyTV87VYb0qrMvdqQlUevsr1
K2MhoBmqy9PqUZzWd4qO1suRO8nPHwZWUF/emVnEdhkfHw8rJWZMH/XtW5gy4RRJx1fIv4kc20cv
NPMsIF3DKSjR5JPisqdD7N0rMZJzRISrx4PSM1kKEiRsnr1iVriE89/Km6WNTcRvzPZTKBthCPjd
gFymWbTsXKKQvb53n+JK1999KIDJcyDNaG91518/W6xzSHXOS78pU9KsLvWsP4RSvKkECL7BDpf1
PziuOjTI4FSimtyhB6Lq2fRpAAPyglniaoMxEkD1aL6LAE1kCYhY7l/vBL7OCylne0CKelNc6h+h
otWh8qwOww+nPmvq1QwxB4tQXonVWNb87iRb1nTxR5KrXGp+aO2Hw58QzK91dVmfeWIEBEas3JH2
H00Nor2roaQcSWXrC050muWISBSh03CA2hNz/jJ93pSY5X+tHAWE3IGKB4lrIdlJjY1VRfU9yc2X
wTbeptnE9Nfeu/zH5DKvKESL4m8GpNhYaRE+LW3fl5XD7GVaPbIolrvlBANnQ8p9F7MKEPMjfarz
btsKdE+OpgMtWTIkVS1ZqJkUVHUSKxqTX4yxn3nV5u+YgzhSmTE7A7HIa5csnb34Iesr2jIDLxuY
uyOFh9IkG6li4p54satKHPkBpNg3aUG4gobFrDQ2LaD3QEcQnxvMrsDsfm3UDXkjJuMXslTmi6No
o0M2J3OtSQJNhSmWFHB1NPQJuKggFxsWtmWhQ1ByyTth9ohylX7f9SjtLjtN52D7+/9AnrM7H+k3
MvuZ/HZEcBMwrVsAUz0BB5UEQzFD2nSsftTrNGvYjIDQHlKqjARMl4rxUy2G1caBGN7dV3R5eLIO
88RICw5qOiEcI09JhkTfSuvhszkka4fEjQHjrITjxL/T7DY8349w+O/JuuAi8K87NrLfL6NheRlt
EUWvk5wtcodtRKu3FiEBYM4nwX0WrspA7zN+s8rlnkxi2MkKLapc4txtolHN4g9D5T6lguO5zoKe
p8GVS5wFivwVdvwJF8HsnLI/nAd1uAslMZ8OqhkSbo4uIs4cCLPT1TK9JGMOlldReQuoMROhU5Dm
ROLCHsfN44/ufWCzJxe0vMGrO5xmuN1AQuGb6LPfFbhhYCKz+9zLInlBAAF0hPNvN/CIb7VJhycn
6T+SjSMrHMDcrgN7TCEACpylmPjK1dB8xdCZNQbMuMH2z/q+Eu/YeGREPQD56JZ4PrR6A/kiE9wn
aH14s3ayDuN92wKp+RartBiMaN268J+R7zrsfplUh5dcH24269lt1SGxPkf2FsxtEmDS3HwG1sJ3
z/OWgYJ6V739rPZljC14ztykXCKeG9lDnjVsgvKJN4ANMeG31soc2Fdvqg1dBjD7ORlGoM7fG5f3
+u3ReCmGxg5s0XlIXfBMPaMgnmosoufRcdtElGYnG6b0ysN3436/3XHYSV3MCHMpz6+AWIgKJciM
3bKDHy2pw42T/EDYNvkLI3Q+q5QhI2aAsAmyVodI4QF3P7SWKx9O/KZWxBgbXvkBvwtWNMNXlNwL
RrriGPUMbhAD/kD4JRrLejZzAlfX8GEd6sWmkBNwoPcQMt7A+HBXaN3IkgWWvgVqTWeX94whSBuG
0amMgxZIlm7tmExVB+nvqscANQVSSsIbOWPFU+FhStK1Cd5vDm3xa/BWpjZWRAnpUx9Kuzup8Z0M
0nGyTNISv3Lq8giA2IZ5Tu4c95ExIcEOQQeKkXm6dev7gh37xDIvwHQUFt9oZ4oEQP3A5m7h7qyb
g/lpUJP4Py47Fn0scI71no8RFvxUPPp0KYQbOkR5UO5Uu2X6RHZ6FFCO2ang1h06SsYKzpIUW4h9
KMxvhzQwgflVMZrXFiw6XhkGuBHYqn5CglLHpCgm4Nk/UvjtsXl4T21pUxmWQgKlrlQHHWwFAaZT
pSqhdxka0ot/uR983IEOJrOx6FPSxP636cvIRMgbPtcBQ8CoSL1Y8kkQnlnKNcG3pOCqZgjpo8I3
h9Ft1RTdtWbPAswy/qaOzx5MI/e1w9G42ndmV5R/xw6V8N1oW4boQoh4d1cClqVsUqWZUj3gnuu3
RRs7L7l5HNl8z+LeshT92jEYRcLJQEdbspISTVDoJsXe02HNfNMjo6WGjBgcWut8+uOz/3XvFLwL
mxn2ctiVYnAGIO8MtnD3zuZysp5CoPOMJkzVQ0fY8SedwsI98sIS1kX1r3/z9UYgQg+7E5lbB5Ps
ZSl9GbwDV3yD02AbN4/RqCpMXkDzdqsx9h5bSAU2IMbcVsUpk89D6Sm+kdIS50tvIHnRs66H4P2e
Wzvl6kxJeVCkDMrH32N3MaKeIgyDjKEyd3UWxQxdukXW2VL4cm0e3BlzHIbpkaxDTVcpkdj8DP6W
vEkN/YjLpdwvXS+ZP86s2sjsKOTRvh78YJQuUj58TtYyQCqbERg0MgC+o/UJs0v5DRCa8jbUb6t1
oFp7D9SPQYdDUZysCuhjwMHgjD18vLRNVJbFAWBL4FftTQbF6mPNsmLj4l9xhE430flGGi85L2n9
oAFI7dnG/2Otl/SSGs8VoRVvt7xiwyesZcPGYhv0Sh+8zmunI4JJsmrEGlijHMaLsdyZPtxHvfUO
bCxWVawBzQLYInByW+e6qRbe16RcunAlE5W7M2BwbzV5cg4duursS2lqso0JLGvQSQUEGeV2yKgu
tGyZUDSFIklPlI+s6hX4q1TTYqt1qkG7DXFI9kml2UkkfJ74KngzXjadIoxYt4Ilpr5e4eT+QmhH
i6zrKnu/m1HnKMzFjdDzqu4ZoNMV9qLqBepoNxjh81ZBMkZC4Czn/JrqMJDPktEn4lBZ52SOgMN1
kqRaUYfbMRf64tci3daM9hwGKJl4UWWMTon536X88cO6IbFR4r1O5p1eBeY5BiawKkiHA/BWVDl6
q+fgwzjTxJt4mB0qrS/j2TbDM4TY3X4ZUXBaINM3YIHfLSWDmy54C/qpMB4JrnMBCcDK5q4uWwwa
NI0ucmDl14xq+AHY0Dqh/O+lycHruQfZ3xaNh4u29hEABfUuxpN68qE7SzSKYe2LBgx/ubr/mcVB
P1fj8onfs9BgIxYDwkTE4mYAGmFpBsI1Mz8nOHl0Dqdk8uiTzfG5rFZltZc3QNVfJVXCkuXPe3BB
p4R3Ze2cMYaE7Js5+UFPz5vXsDVezTL7S5VpJJ9wnm2uzHdrjxiyBeomd1ctOE9jUARxNjmRiLRx
v3lFla8538GAtTPA9NqkKhshhMHYASEkk7iE/6rwI7gzKdq8Euxzhr6QSiv/MaGDaoWzyOedTfpr
niD34S3ZS0u+1jwSpFnaW/xon+NXuudszVlHRccmM7DL7HEt6BKwK6hsuSxTzZsOKUet9JD8jtn+
W49doVk3wxzVz4v7Aw0u7GPFe5YjGzkePKB9V+f/BILSsseNggGBj8LR1PYwRaV/nzJ9ikvuLguf
dwu7DG2NwPB3mzE5+O5fHJ/KIDdPFZJv4nxFFpiABoJJtlbiSv7RDrkaqakaIUDjm2/HFIyIdoeS
7c+J0SoD1p1QLjZ+IGEGCfZZ0xsdZneR/0jGicydC4qY5iUiumAPmTTXA9p0/RScXF2qtyUSDipg
+RWIfbQxXfJjQ7GSxcoFb1XX4vg1hWTVGZC9PMqut8vwpaqObLbHwcIcLVtHUOI1BcX5xSEj1TLw
ddTCxaEob6YOQRA8QGHr1/7U5GWEsAiE/Oe5bTND2O9QohaO7PKdVfR6UydoQxIYx2PghCxMa6Gv
iPg+rRWfXjOa+OACzEXnQ70wIiG7PiCOzfE8Y8CSrkNvSPOpnO7FnPy3RkDTXx5uBLHayWOOBarn
6nY5yPlDMJ3APzvmIogcb0e+vesCStKeEyHw8t6a089JM+EJ/NjCE9pwCpUsUINkwralnwkeqTdo
3RTftuXoI66OXb0lJMm3wSiQA9GuoRpbfKYX+RPXY0pXQy4mehLY+6FFaT3RfdylETB9Hm98nTnr
mJE50z11BBf7Kg+JhiLIdZYyJJEDgqv3NE4zVNd723sCo5N3hVaN1OUu4RWy1IfYqr7339mGtSD7
k+p0PNrznSXZih7uGXfAVLUup+NE5A12hnySMY1uYqyWrUgfddIsxKXE4VxlD5NPN357KJ3k9rPn
WRn3wHLqhE+S4mTq5ZF8vt2vDyByCal/3FWtaLJqqh3H4Y6wjxjEYs8fwRGFRIsJU/bOvmTsTUPZ
6tDunbn8GXsuTvK2OW722kshClkwkKQkP+HQiwe1vImImPAfcUxJo7vdlvKoB63E1UQXMhFeCsXE
etaorIkcdmH8JQqWnCunlm//QMvA4v9ZIt+pA8c1gl38AdZqNvoVCRdhxgvSCB6P4H3Hl180OvMX
DrAqgYecPf0G6YivTXBkxmNm6t+pSEQ3Ki+2YuiXuSFNZI0EggAGBUFBiFMypHbTqocSxhMvpjQU
myxkFSchRE50T25NgF+rEkkMQgN1+xprJCPs6FanetsHY4TmFK/JHxvVAiYdEu9J7TkTogFcfY48
6oKxMjmZj7dq39H1+4LrRYirC2HeJNOxnC8E9pmYhZ5NPdFaSTBZMkUyxA0JT/QxI4GX9T7HMLK0
nZTYJga5kjW7UAOSJ9U/qkXy6v0GWN+yIJVpY5cZNn7VbsQJ+4Yy07k19MAscFl3d5O9XwLdowhw
SDQfmIhGAr69igZNZzv21a6s7WSOdEl+gZj7U8zhANCyKn9b3Wonwabks0iWfV9eoX8aUWgAiyJF
ZNfZBWsJMlKLSSHwYaHTF4imbv8F+285gmooC6kMdboBQu0DhMv4vDiftem6LL8BPMdWbbsTyMJW
T1uB2+Y46/XyDeSiyAyCozZbB6EPEny1MM355VB0Z9ownhjhd9ncGvzvyH04PGdikXqjZad0C2dg
nLkI8DLspSzu8oyf7Jq+0MGEQ2G/qgPtBnvP2dLS6y9EhhiZzm20SM9GezRhgUDrgTb52kBffMne
x7fu3tDAGtvdEGdAUop9Xe3OziWVn1VZspcThWf502kH9Kkzohx/qLJUnyrYoY5z5w5vq/VlTRMe
vMxd13+EYj+BEialUP1dKtIHnXcft75tPXzXCKpmj+5CJr4l9S92oJnL9VQuO97P67GYvQrR2+ag
NT/bs/lvH5d907/hzX/rKi3iMulhzaA5YMjHh1oH0Ah88AiGf3bs5IMTVZhqVyeq+Hvy4MU88jcB
b3GQLAG/HR1VFAXUrjKmIzN7LxrPd/9fG9zssMgNY0vTDBjShOCgIYyh2aMBzWonZPnP+WOVapG9
Wz12XshulM6XOHZ1Cqav3glbuGq8mJP1dL9MLsQ+tCReU/q3/ksXk0hRbm2XNC/XrL7MN8X/zHPm
ZuQPY5kOxPt5/vOOAWaKL1f3QshPkYBh/1zgbglub377RbefPEu1tUuQWeSqSAKL+rqZOOGqqzRd
SMF8E+hlHnpUg2ALldZ5gZANfG5CYA7m0o+AxmLdzm/clsb9lazhcg9u63ZpOGN37cxu5VWpZ+/J
qSZZnTQnEjhBWjqgQ1fOasXf9Uh96u9N63gDgJ56QQ3qzzgkEWgYqrh3SZ9Ovqh1R+ONGCfcu+X2
p7BHDUu99PMeRmnFYWZ3opPzuqTp2tnfHAXl7zWd8slWH6yNC+UqDFnATOscLsyJQ008wfedvIjM
QhY0rkUh3ThDjRELobhTuA9PGBYSFs2lWjyxx//9F6q5X2D2x+0nAlohjweiLguzf5vuqO85t5Hp
TeqfvXwr84BokBQ7opAlpiWogUf45Sy/bhwdJwwouL2Tv0eIixbFCvNRUG/ek74voHPpncnUPKNj
QQyA8mOY6Rmlxy9PsticZ5QfthC+IY2liKM6dqVE+K3AunvZDG+3XNM6yH0ZFgaa2s2TCSlkxIbt
n9P/lyjwCJkFvPkUwkuMbNt6OWTZfPgpIfKud7Ulh9Tc0AR5KNk+W5Zb3vg5a0qxF90baH5nB1k7
/xN0LObIzXS97JFqjVkQRzc3RHFSF907xhVqNwma75SmyrngYlKxMy/m/2N3rG5go+r4Dfx22vk7
s3S5BwTxMEf4zVqERN4ghSd+2HqOXCNi7G8TzrrK8a9f74zzC+kXxQcmWxZFyC6+W2z0IJPiAtp7
2Zr0ZctELI8f8VTbu6HjFzLWLGdJC2/YFUQ8oWtIaYMZA1BgH/KLeKI1hz3fDYktdPJQam92xvnt
nPSA4fa8O811LmUeqd9mc2Jmvk/JkN8wUFshA8oxuszSTpp7T/bmi1By++sR0oy9SY0ftq8oibNQ
4nyQm8GjvADszvTey/TJFBl+qrLzRcCVg0312rge2delwNnlHvaS5vXBU3f54tgzXeJ5pDesGwmW
Ht0Amff5ctL10DBrj19jxiSO4bBEemHMixFJB94gBw4ccJ2CO2K89T3qYDAM8QyVwqI8IpKopn/n
XIs5vU78puB8on/QB7B8dQ4sY8W//RSt+qVlWboMSvRQRIJTpi/iUOzc73kqZ7PcTPpnrdAKmLue
O8eCtaKv4jBU4zZxqoPZrT+3ZgyjWd+qkrtwQgWRTxqxkd2m9mEDRQYJPDIqb3y6mRS7LHZwqXTR
rZRkgSil9EPbt92ffGgG65o+bshpQ4nVcO6f1oXpxI87X5N2cge4EtX16+sHsvB6UEUQRbSQfNG8
Rt0dVeF8q7xx5Sr7ua18HtxAjzWmZD3SvJZ7BWw75Ihdx0WA5Q7wBUYFxsARPKFWL1XPJ0nKwLna
tnFKd7QEQv8PQQq9EbHT1b4DZ6BxPgBsSG+8FP/+65xWoHX4+KSnYMHXN8wy9WyO5tmJZAIR3/Cu
C37NtydOU406gDUrsi9cVy1FlUSlxRBZiZVi0DRHpknlD9jMY+aomGwv5YUyK/13YyxuXZFRtBm7
odu+mw+60QG4HpGCxptC6PrQUDVXWZKlbQNGhOqej1SajvW1FOiNYrwT0ZAVLKpfTZVj93AAfeJ3
8tgpNZoPBJCwMa96tm27bhlsvjXe0KvpShZYYufQXkk7RWGVZSgbqurTrZMkmqE/R4V2hkJs5Sxi
Yw+GNmpNN1L5guInyIOZ8w3132lwvss4nNAdoPBSpHkhK1Y8rKd/0/EW8zwFx/0hLrqNYGB+KTVi
vMTNs5vriZYEjhj6l0OXeROc1v1y/bikHz2GT1olUKnbGN5aVB0AVavzdrfcPgMkIPWOSyyUnNEw
H5wOlxc5JanR5S2taS1caTiKZr4Kh2ZDYYI2uB/zcKD5mZ+BX6OEvCmJ+HEFmuWbUlaLKbmV6S7E
KxPiLPpqHRiQNrMR6SdIEi/EFlsESJtL6YYnkneT80u4VY+aPxuH0BhxdpOJE0uXk660Yj6lcyw7
UIKfVtbBkWLwIB2NUTyMEze8NIhjxdpHBMeodtuxYskT+LXAooi/7EyLI9DvUH58zSi8XATDnpGG
XJyU6JjiuuBC1k0q7hBuP3vcmWCXPpADazfNK8xcrgKDa42vAz5IDM1yXKAsMTx9LI2PzEwNfBva
rdcI/F57PWzyG+L5u+yaqXSMU8S0RbpuD8RFXOvc9I48NCiPk5fSfIhnPhw/AN3/IlsXJgN2TpwG
pTRQ03SNVEBqZu6BKzX+9RiIumL/7rEIxNn8HHCBR+YtGehI36kdU6xg6MbC33JnY4ftVihhmIzd
UzsB+oaImkGs7DXpAaRDNyyzTL+Y20mOeq+MJ4hAEFbRLstXPK3BHbe0PMvLKAPpG8KZoaNM1bfE
zUXS8aXZ3Tu4FD8GmyFyvBpreHqcYiJNe2jUAX8zlgFVmP1m0ii4Q48/6Oq1drQXdhpYhNxj9A8J
NOg6H4Dx6VOkR8mMy/MOG6QpS1zVVdG+TMMclftyO0gVGXSVfNPhzF9ossiEiwr+Y0IkkP0wipsG
5ORPFqN97xYxNvUPUjnrpGUrJLzgy8OZ4dVV1drdrEAflY7qtA0qFgPT2GS0mbUngQzhe3uKRity
i+tUD1sZyUcoSlshqxfRk5Gdqw1tbuCOeSSIaVMiGSbUYIG5YuxBGweDaqRgvNjscz/IuhaoZHBH
3NS6CdE+IoP80tcuqyH6gSVxWnH1pcBe9NEa7dbeC3SH7gmUM/k4xTeAZIZ7gOKjP6M6wj/n3H3y
us3Kzv1izwLK5W1F8U7YV4tWrcTGW7Dp0/FsIRbi+uvSLyp0TD7g/Uh5MGBUFDFz9g63O2AgCY5R
au/qtX7D0ZynPMRSQVZmIqOnL4K0Bz+gKUPUuCWuaa4HSLELeTilQSnrn4Fm+DBDZOAQ5Bt+Ivks
M4d1F+ukxtZ0eHyXxAWXyd8qJ2iP9u07NvMh3GcECNMREhgm5IrYN1Fr9fhDngFijdDdXOZVH+vm
rCJEM0TXDBJ7nc8Wsw373ze8tq2AgSWn0YUYnRvRWq2fx+G074Px+MuzDIRViAuOzU7AftRSvMD9
m8IJA10TMsD9OXFBH1pLQ8yRE6zBPUVyJQxuMnvuRH/5rPx0KVYqVcGOfEb4/UjVYAkjatkALJwZ
rvaPOfxz6kNXEq7q0tqDadfSvvIiL1gPp4Oo75ANen5f061T1TGNtJgQzOhLDZ12zdgjL/6/kisx
F1Uvd5Us8Bpf8SbV6j2J1vYEq+Km0f1XMsxG3oSvEJs3eZI8br84sui4hqJdafho6nwzBMjEw3r4
jI+PJEdRhLf9QDLrJCF+dRQqseu6fVFqSiuPDcZC2ChUuqY+HMfQyb1R0Vx5E3NCS1VKHP7rLRrR
A9ciN/yhgPykCDNwBHI5TQqyy/edcqP8zdrvdeTa7Bn/DSX1dOIuX0VpwF3Xrn2aqPzt4XIeTb/m
OQsqiI4U9dSjiOPUcniS/n0UiEVY3xPzgCtJdMVC0iWGeYqymmfIwSJFsO5qJ/GmKEERhBVdP/yN
sqYd942GvAyBdW/ro7JN5M+FoK8HPMzmwLf1X1RAzCrOxPnDT1WuAOTeBVrU8LlAQkNeWjbAS7UZ
lU1sUm2h2EXCR++NhRAjnMMCgVQmPXTjwk/wOxMC/0NqFhoiGRtgK2jsIy93R447svCIjwUX2NJD
GF09rqKZrvUG9VoW6FQmmDtaxFwyzAVLVi5NSqAPAuJY9jMJqwr7tZsWFZClT7PksGWPvD4PJKb8
dprodB3R9dCyHp04o3Maz9WAvGRvtHKb6wfHxYPULDlNnQ9X/M/ZTuuiMqBxxJIfOvsQXBGL5Y3l
W3Uh6nbYyTb2DB2YLbdcf3Wn+QLnj9Twu/wIqQL94v4eyOjIaJjJLqX2vJVIqoC+OpXWDw0/JFy2
AXXDXIU+6yVQzL6YQIrSSw6ZLnSI+Km7TB5D1cR4fthbUGkV8KS+4jyWXC3oQLZZjl2ywWfuwEYI
L+zsx6GTpRPL63HtuZJ2JUBKCFV2BBYF3lQDnCT0Rz5keUcvPN5yVJcuSdb7cMF2zDsKZWcNHJXx
METV26pNvjz/tonQvuctE/FpC8DKHdLsfjjCYHbyiw5kCABS2NHnQqXJrjFFDQuhBeTEsv/t2Qlb
a9GBFGW4R5FRnUZCqirEw8eI/DxVRzia/RpZN+d+HJzarj6u0d49agKgi9p/XtKeJQFGITjhTtx2
I0sQBK3hklZ4u4/kQBCrNEFkHwrJXaO0wDvXPS7mkjNWPWVO6SPTtdazibEwMxnwgQVhts3vBG7y
XLKtZ/+b4LAo+cvkSqr6DGzMYInJgL7CEvqkc3CQuUYM2RATxX/M3kD0ZTkYq1DOUqelyrkCHelo
oC7e2snSXITLwAROR/UtVxvvIjMMr7D+El8ZoQraUnScIaYTuU+Yh1CoKJJl4K+iPMDLGrDyeRvw
HXzfVK9YnanFshREqGGClv11U663b+nettXAv9pYCyNrLjXhORBdPZ0cUa9cnqx+/Jhtccmms8dA
ziXw7w2sTSpQUwKjqueLeNkYA0bIbzUC8S9Si7M/O3I9kTZhajzVcSGO95G+pFhSTYnnibkpcEj6
1k8vbvgTgIkC3TgAD6Eq4xACroTTBLHLY+9r74peDD9XRt8mdgHE9DAWDJOZYnBQnrRb/ETjKuBr
AqqRfFtb0UH4dZWYojIOCSVBEFqZYmnRWQ83RU/VWHLG99PEVnSitogW46niTrXA5NPUuxC+5qVt
sjfz5njqFOiifshT1kT+xIsxYip22bMns7Z1+WLyyzxuLQW42v4uVaJkhyq50/60EQraU7rq8zGS
5rDL2DgZx8lmBWLfnxZSFaA7N8YP8Ls6tQQpbXGTHSa38mEjQi/+SzVafH5s3JMJGdhHLB4j0wqN
C9KviuJCD4juY7lMfUbLwjldw56aKh34fROROYIXKrrbAVqjHyEAtzl/JwnwAUBstw85VQzOuXwq
8tkN6MEiuVWo7+GJcb4e156R+v/WqJk5/iYxSS1L2cT4ka37iyodI5c2iWX4KbeeXjWIU87DmAKn
UapgTeAkYSGlZ4BBKPus3XhHjjQFT+PaSROm6EUA0wGx5beuyzFHqLHkHPR+8Sl6yyoQ8iwa06BA
+7UcamxeOViQRJFgR+HQk6PKsIdnHaYlwQlRYeYzPiCNnFjQx1UEiu7SMpsszTrAODP+HE0z7B5L
bR85NUJwNc8n+2kf9fOYlf64qCqlrXGGDjxKtxahDoXSh3+kdbm7Q11MC1L7GmEX/sI74V6Q1P4t
EJF8NZBXdN1dkd1QZtJD2iyxWjO2vYSODhHNnBrHGe+jeOu63IBffhliMT9HQM4p5n5FcxNI3S0R
GXfqbZt05Qj3VNpHD4GVZNGi8CvKpMFEFMFpY7DAqTX/Gcb8P6GWZsIzvrPbwRZOXQ+Y/jPd2zo7
J0owE85jT5/qzcGj9eeHO0Kd6q4mZJg1autFVr1Z7De/AAgbz2YPJLIpfqvvMW/S+t2Hg2osp9/A
QcJ2LxdUvekSedZ8ZpWRkWx0DyzTKGUjf91ag/qXitERydvex82Sd0UxZ1pceGwU5Qrkc0cEWTKe
nE3osSn/FlhO6UucMKRzs9GxjATnSZP7UEVcr5Tor0lsiikCz9GE7CMVRRvH/0iM81G3eZoS66OC
LcnjiY7zGqc4Z/DnE4Gg3OmyPqX3uuCFvNqBrs3q878RS8QmXM/5FD0l9A3cTuhqMUSZUo20lx/F
bommb8D+YIL3mw7RdTvcEV5XzQ9kWC5f+p86JKKo9c2etswceeecwgbk2khNA5I6PhIFnfsY0j4D
0alPRNJVYF9y6p+OkXkECOUrMplV+iLx7MEtIEPNgpVu1eZqZ3kAl5O7GYtM55GG45cXJwn74h4d
ilDZ3vVt2leyJl07AJRMbMsKDronBE5QLUnk1SrYLh2HBUwvapYZBYeB8yQ3dXmG96gbFkzf/KAr
xk3u3hevFFCInGkgngFl9jgtblw/oPpnnBBnYQfXL3uVQ7r+R6dgHIDHXW/2uPR9SvpwlpO8hEgs
F0Ugy5GYf9J9cuAv3ba8ro/YfUyFDj96QTGDIIlp/3kB1Y0p8X0Y6mHdbBjbq9VAJgjmRkvVkdc0
QNZX/PTaOxPmbT1tWDadNxKfOCB1EXvzSkR34H7ajuifQr+/pHnh5lXq3avW+YCUGOtZ4P+995C7
uIJ1CEU2ByMy2NVAgu7+MN/79FcyR5kzZ/S9kAdzusFYLxyWGUjoxQm1qY192wxptnnuW4aTGpXu
wQyQzMTbBw1tB7MNnUJxARpxcWFOsB666LnwUyCEYZ17ARvv1DJ+aZ9pZi5UCDt8PDj6lnopcqvP
/eAEIPwIMeH8c5OvKaCTx39hNaH3ctaMrsI4jqHC8fz19XbuRfHL4ysXZ8kusFc0P3DK45c3PeKT
k5IqNXb4Bqh0jxKeOqr+TzJBagL4M2J+V8tJ60625egfq7YV+at3efunGgO6s36FLTqM39q31uTk
1Bj4QyiHyUKw2zBI5wWszIW+tcJ5NaX/l7wgxtycevuBUV/jDmuRuamVwIPk20wB+uQYMV5t3xkU
k9PXH2JY2mlpQq9d4o/RdMn+hCljtn5jKteENiB3OfL9g9fQViUqNa5zqxxUGgvi5/isEcg7aQiY
X6eQvh9HmueIKes8mW3TNg14FhjlikG8dRC9cYgdAeWjT+QhAedRUXhcBQF+Rj4+TFmrGIbSjEPM
qqzi83Ackp0wTN7WuCzA9M9Ztc/m1kRfufQUlFOVFqCYzWu3PGeR6czRanxZyj02g+SLHQbThMvp
K7O58Lp008Sn/24GMBb7QzYL6PUye9bBncfRE6LkR/EHYFu56ytFHEhO5Frx+AIRNObolEuOranN
N3QqGaqPFStbdP4qtZaPjY9bGakPSY7pkjdl5gNN8Yp1ph6TtIzZ0gTanmG0zUFCeQZ9AXWRyIHG
M+Po/FlFZw6a45aXac6ehTDhco+QA2AjgmyrnOHL1XjN43NiKHycIoXeWBCyQpxAGVwy4DFhWM9r
8EtjSdd6Ov7kEp56WQRXY/C4SoXHGVDo8mrpogpghb9mg5hkuca+hrs6orGfVvpFle1sjYu782Yr
D7v1QlWHXvq22BT4amt3fl1n2XTlyleAaIu4GKKyxwGt+yRKn1pUbYKvRVJxYzodjZptuzIFzCsr
TIcvqitZDOjtKxfeHtuog/1lpVI9658tOjjaQnCGTsjLFke7q0DP29pMAjgy7ozO5pIFVMPaYtjw
xT5qonkxaFY1VtFR5JoaW0uNvGAlIYNFRn1rMWW/TYURLFCCnap62EqV1Smkw6JYkqcYeN0hl2Fw
ehd5b50eMkpHEVwHSlCxCApSwcfAuycGyh0QTzbKWUd8l1CYJscGoPu0aeFMTbUSRwRCyUiSomx3
D7Ro4++CeXfPk4bcXtD1uBlMac2R+s+2JO6t0j3qQwdY8MXs6kXAXUQqbwdrEbG26RvDXyuEhnbc
omkKhHVspHRw520lGWXGt1Tl5J/gfJ1gt6wbsJedW2vjcDWqczCP4YYImgbTq/Pb2Q4MmASrlwYj
6cyF9nMYvkNMFPwufGqXGbOr/8lG6Q8h5njrDtfRstKZ8zME7i3eO7me4/duHWsY6/pR9r/Aci6n
tmrL8QAFYwfWjGM6/3Ahd+XZff58Ub8UwQgmRWZGP2U1gP5qKcb1r45RrTXQl7gBum1dNHaDXrxR
FZhEHw4hM/YISF57M3XhdKHV+V/Z/B+LVNb4iKv+SXirtg12aH5EVMRhorn9JnCNRsKfeuDU8qXi
KRih/kO3UpFByNAZ5FwONQbxs4KKlDva6OIgqxysbb3PQC/qPHc8AK7VlVJE2Nni3jFB0KvrhsKP
aXNHqNUJeMpR17Vdk8n5MHr++EjWhneJ1w+htDiqi4Rv8vg7RE7H1Q+4lTpgA33DLH9uXKbPydHA
KTFS8LWjmrNg3FDhMzsVtT3YAZDRdV0y3KuXep3Tz5KxgUixyOUEDOwT2fFyzCb3HEj8Q/ZP13NR
32iK222E9cJm1Hirq8IEFjSARd4NRirfj+a0Xmc/LPJxkVeysXPLQPcRUJys7E08Dqiim/9qKG52
JJ8Pvtdj9EYPYyAvC6JiVzJaD/XELBoYSZNnIyWriDotvjvFtXI5eXn6j7yJGYO6DZv/VRih/MZM
rhC/fa+v6Lgcdn8MFF5wEMiBnF2QMCfrawk1SJupndJl8G0r2d6RX7cZKznAXO7ZtFveo7xvv58y
GK3C3GgUEWJi3pL/ob7t/lP+qJ5kbV1/QBPnpNkVwFQFfcDBvGHT7bdyAa49YdvB57BDRKS5RAfj
xNRRGtVFjrRsWu+FSOYkRfsg7BVowkp+DoGFTyNCg0C1mKJl5wQ5Q6LaJDClgncbDnYvDlHzFfGO
pGMFEbOBinIk5KfIA6zgPcOhBoW0cWjzoMPNqqWVdrTDRYJZ9kq+yBf7Yk95Xki6zuxTIDBGuCHf
OVdupstd8XSgNoBUm8NaGYaGCueiez4SpQLMtzxP+RoifISCvaBh91zXyV6aFq651i+qDO+ermSq
OkiR5OjV5wcnqXTs58LKY7qHF44CP9k5PR8eqX6J8kkKOcLc4kxc0AXZtjDD3UpXC1T62aD5hBfS
c8CtHhB6lTxTAiEfhyZvBAQ+ZLoBK7OL89be8WoTxX1OeVKevUr4HXCwFxRJcuxv/6vsaZo6M4xF
DPrPzDXeg9pjCGbTQvVIsLt5Y7SfXupD29Z8Rp8EhBxULaBwcGaoTj6a2wGbTbotw6cu7KXJ7KKh
9mooipTultGPdcoHB7xfkg7BL8HKokNm1enYDfd5OqnRBuN5VpXq8Y83Hy71egrAytWeSbIt9OX2
cZNUCm2fremWE6yc5A05JEiDJBaCiwR0hZ+0ugnxfhdmUHEanM9I2aWNbryvkp3WEVC6ZaK6n9m3
NkLl7/DE6X5JYSC1tfoReN0avmciY/6Vgy3PaEZQJu0UkCFx3kklsfLPbCYdIN5DOkWTWBRJc7DG
YXXkVg0m3BPNV4VBBr63nPsbR5XsANXlWiuCCOmZZRPHZ8z97HR7VRskcrZifTUBow42CMABWmw5
9uvbyUdmkvIj3Z3N4g/WnwbJu5HU1yJ+xOKALf84Oqib/PHK+ElYzed7rxjeV4fbgu5/6dTcRcG+
DprqH4Sh2fyCJ2cszBI74Dfe7i3t71SCusXtDq9tOZ7qYZFQEPErqgMdlnbbbExrqTXo6D4dgqG0
5c7kvGDdLHDKxDUMbbhFcKhntoPRoybPsKcIc8okAqiJ61SQy3+Q6nOpEbT/KcYKPt/Oo8K8uc03
seCSNlhc7n1ftRI1ph00LCtg0iRHftjboy5cLioKRUmvqemR7PR1vXkOmcB/AfXAZ3N5tCDdd6jW
rufMNk1fHHQvIpKgM6yoxv89Ytnc2twzwX5MNnNuxoSrbdpQGs6pCzIm3IWM7YE310mrXAWm645L
eKHFyp3kgLXItrB8ng83UL5+YYZGJJUFHHfvHWTwvChdKCZWC8OigIlAEBfg9EpmE7BZam/6GrvV
vj28dveYKDtzQAOt9HB4UxWgoOCuPIuHSzgQJGUmoAVUsNVhl/g6n2S8RhxKM/ix5vXZfMmdw22a
woUcfqJgjHgxvz9wBdrjN9cW68kL9z0NVvkOBkjBaUylrh9S5EzNmoJ9DGINVgStiRuILIRC/L3a
/yMwYPUbkHyciC0MNzoMVjP/0dnpXue8ZrpvstSHekj7G4wM2RBEf0p5Xk708rFYF4+vd36BW+cs
Nj2WGbEi5N6oTOK8hE/zycHftZ1zZpr37zXqJLOpa9iL9soyL2X62rW6OVr2QDOO1r4UhBlSWq26
+Hnhb9+AXKxaDNsibGNR3uI7lW4+UTzDlmF4SngwOfGiEB3q/dzU3DxVC839ioY/oI9QLpiW1Iut
U5eFi3xeqC6ETi6nEitc9pz2s9NLWiY5Mu8nl0JCmFs4RzT/tfYJ6qGO25lMqIzRBsak3crKctJI
ht8I296aADrjy9ntzPH/+haPOenl05QvHvXQvVFqA2SDrQOOqzUEGcnDejG5mfcZ6Xbqh1lg9Oei
0EXvAvvycVPqOW2jOu/UQlK2jNC7OGSqIB1djLAaBIQqzrD37VBR1n4RJYqFUr7KahhoLDr3NryM
290DkUKukdt3rY64Ff58TqgD1euZHxnpEptmbunxenL6TANQeshvD1XQgJHyoSwwuTwi47a7Zv1m
WCzyrsV/sHo65vFsu2Ilorl2AfVywgX/7Y6uVwicF4MdljuTui+CKLBTsU3SgAuas96MH0Uyrtwy
goYTqr5I5os2WAVcX9hpYHi9VJhgXF9N5ogC0M6FpDrkSP9UQ3AjCxIAVlLU6n4BH9h6/0FluGoD
q0QJyo8leZTAVKZ25pJKkndFOkZ/F17ml0czUcDFe3SJDuj1/Jyue1RArWwhKgHK96tFlCfD6F3R
VBnrSrym9aAroEs/9hdsZNz+d3FG2Lep5wEOxeWOwlkNcCeDDzJ10Kvp1IAShqjYjg5hWAUEFUcd
g2LICIJ8OxHRvg+Dkk/hqubLnY0rr4nGV8nLGZ2NpwHL/qyddpzQ4IbxL1lUwPrxejqadKhUvs8R
XlcVfEXoN3OiEDuFHufwe0AAd/jf6hxe+V3Ar9VjYSXIYix+xLJr74V9CRPKS/Q54dPz8KundHGi
iOF09lBwrYfev9CRBmDbar8BF8bbw2fSHbeDmeEoKhZlts4RfBKe+iSpjI4OQ3XHMahea7G1SyN4
S75cebdthAbkMKJhs63pwFpHGUM2uxK7wU87XkSuvgiLq0PqLdbq0Pgh+a9QSFFzsSbmFedsaU+7
qvQavAKaO0c5+Y5+9LAt+yOckSszzsmIyvNR86iVxSpnfiN9lMQF8hMNBL/Eer0TUC1wxqn6CIuU
+ebi+1GXxjNno+h3xuBDBjPnheWZN8s+GQF78TYwwHK9lCUAX/LJQBFjsJjL1idhAOmSqdWvXvbF
80ikazjN90BLDyza5qacK7XgeW5HvUYwS+qqbeuFI/HqOON3sAujpXdgt4qx7QGw/KFt4zuCGhtc
5cna8M2fLeUikg5knju3aEAA5JtnoTCydm3UWhTHvdFgqCHmUvUV6mTmSoLQmuvJbbZ2SEsCJbTa
J13C2W9d8HvUTsg2pQcEl4trxSTk5OhoSFprjRxZQuvNh8PNgkxIxmSctwchYDZPb+vv+lcOh3nR
HY3RXNv/CKCzZJHtf02bec7ZgwjSb7RdTY5H0h9piy9aMlw+5A6jNRyrIn/FtsJlZa6xivc1/vbh
wa83B3eezi2hgr2Qzsg60N4DsKj6C7qw84R6qM9TDZK2w6pEDtS9orqSFVhf+u5ujL+hU48eb1Vk
eC2EtZrzoMawIC3wQFZVeiy2g/xwQI3V9zngvzQlfW/2kIChM4oyLtQ1QUxN+DY49zwgySBcm//O
6B0S+/2J4kqXrwwgfJ/ifud+kaE5S4GcfzzXwRvoyKGHcIViMhgLLSpVu4z95x+froNX3ojUtNPx
0l8sUFkxalSf+D2Fv0QqmnSdtkeNRliWeYBbiFUpMFsM1nFoX7r4x+wuYGkVx82Ml6s1x2ttUAmv
enkTzLyae5Uo83gtfWZ6d21H2Ehzb7PaLYjbC3IkDDf3Oj9cD8aCphP/JG77SFcak3Tuy2vSE2EV
yFE0uPfNzGGb4ZtbjAd5QPY43yaITKewvMxVpyA4OzeQH5wM9mXrDy+fK5tHcwURuwtzN5CKzRUq
4Y0KWZWhDfQgDbs5o2/iKzU3U0x/vmZDeVB1hFcK7K5e7Wpa7JbdgurUXex1ihSGvZbqBSTKWz25
4zbLGJ8MCdccfk/2AMETdwmF/Gh43nZGyErLcf/d+6u0ZXWUp22ZVnPwCBu4tZ2+iLx2FsQ3aWTb
yjOTOV6CZuFcaSJlIdsPcQQGwuyxc77ogqG5HO4OYp3ETs8C+95JnQjOeYsC9pDB2SwIrwvl+LVz
nT3IgytFdvWp1XAiJZWuyZ6mcEc8bQr/zQFjW7M6Ow9OzGE96syvMRuzPRhAy0tbZKwc1DcwLOJd
98aRFmC3rw7Epqnr8zzynhcMjZGCIftpL1S7e+8ocwz2pUwQqQ646FJUHtGWRTj94hsRwtsd6Sgq
FmYhhlEbT4Hx5y6LfovJSV1dlvELK3RPmgmM14U940I4zRFLvlYx6FQTgkrfZ0J9DlWqfegzHH5d
OHUE8CCaZlAzjFxvqit8aWUJtgz3BV1qgJiwLz1t1PjiQ0Agzj8MFbkSLxgca+BD2VOVa/jVl1/v
M9EwLnklwzYal/a7c6Lj4T18f/Nok1vLrkDUVKyIBFUdOIMtucRIm9z/dBP3j1o5ZWYt/uLfMQxQ
RStns8d93D7chiY1b99hbiGwWrDjsV32AMwkcsM8syorhQciGhtwp3SVsDDjFrYVqkEcuFCddAK/
AyeV00I6mB+ShZWybeJATJXPSQZXyDBjo1YRo0a4GoDGweul7qFgjOcuYgUQZwWXk4mJOWWHnYEG
SUOc5j58DwMMLZNiyRW2PdcLqvMeEOFej/UHAieZVkHKbNpBTI6+8/tAyGN2roK5Lut9TrvBZFUm
CGvjym+w+al/6kLCm6Cin9IyI0cbciEERicZonBySTF9EYRnkORwBmJsyBJ6SoShzxY3ILV7KiHK
B4RVGzQSjFpHc5Wi60Z3levPeVtmTO8iTPAw+V4l/uo017rxz6fa3U+3FRQso/cjCajQL3u2K21I
+wvmQWh4k1R/wCG03x0Tk0NZ3ooVjD6K2xsdAWaJD22KeGZJTSpX5A4sLA1vpIVHRyUr5DGOMpd5
+HsfSgzXASkFexFLmjl6zUWON7gBGGYXCG4TKHa3Gpu1qiCjieS7P2dyRhaRgOZRt6Lbn9Hyv2Pm
N7IwFxYiVDuZpw9egvV3QPvjCen6KNpCpX9rJyRDxYWbEbcsaSDP7ZMM0gkG92aDpNJs3eijS/Z0
YlMI5xIPVpkc/WDT8g3KcbMJJcNjNZ7Z+e36FNysnnKEXi1d4+H8BN3ZVqhmWLI8TTJ9TsprTclK
qQ6gSjwjBf/xnIKJEo3NjdEbFCmzIxvYbtl8c5muWzycQnUwU3elkNTz1lMif/QOOhXon+gn6wZB
8tm+Is4bE/6JOx0cA8/u/HClF0dqTrSZfrwgPVcVdJKolzbsq8hFDdnfXyIwUfyzmH2rd9oHxj5R
tmnWdGT1c7JJScHgAsrSJv9ju0afRSbgVPGCgGyuYefTCJuQPJa8fWGkEbGjHQrI6oGc1AiBil2b
PzKNaQuyCIK2eb621qOvY1xl0xbBNUmtpQ2Zv5WmXx170wJIXaj7qpZma2NsOKS1bE4LlxSqP4a0
7js7QH0s/TWzofID6p5y1VH0Oz7D2vjlKDl390uuINmxBAy2WWHdAtI/zUwt54/m8LuYs+9evWWL
TH7o1brCvboykA1zOc9NhecSa9e6psOGeJ2nYIX4jgJOZQU+s7iqo+CGuctp+PoINVuTjh7dNcRD
cibzk1ZWuXzzZHnKZFB0aB7qibS/heLoG2YSAG6LtZ8wlu4Wj1Sf8OJ448GuVNdbNeA6Vt/UsfCw
LLWK2C7pxfPRLTshbo+VQX0jz32Yx5OcUDWGbEiYyIpMpNqmPgZzRcF4eiBiQ9c7goNHz13lRJPe
TYrQ+us4TkYcvOul1s6lOVCQc54ElhFlrI2wkzisSZ8i5tn6T7fg7XkmF8I3YgtCdDbG3VIpiH50
r4sannDoErlRwYbA7Pf8GcufSl8fLrDzuIHLXtMlI/IF8NR2Lqj5Nz+f6fou/YTXTBExA+QGh/QX
9qObvUueYf7LpBrjIfzdb/pmXXS0U27eGDAH9XC+An7sCUhR5QBmfaXKg3Cw0NE1mimcnmSqKJoN
pPOcoqCopbYkJ9AgHLC+Kr3Pv/AST8JnDxbK3tKHnUNjQhF96ZXhKMxgUNbfki3JatzB5m6+NOdb
QhWSHFyalQsz2BN5Q4xM81zDmcwn3bU6pUsRy+4ub90sqCQdbyknherN63rzLkSSPEOLWlyZFl+y
Vr8cB3PcT8dm4Ld0UiWZRH2wKy75Q4M2AmoyXDcaHTODE1bLV5sAnq/TxIrtd9Ob+5eiu9Jk0uaf
e+3M3+k+DCKsFOo8qbzKJ3LZnSiMaKs2hVG3TVSO/Q+rj6CRlBhPNUHlDtBd5m8q+pDR2LfzIWHO
xgMhVz1Mg/9OurrGnntyA4joVr+epwlw3lcBij6hoJn4CquFhcY/U9kx5XbACk29nz7vahH5mHrv
PQgvxpe5QKXWh18IaaZnlzCYxZZ63nWry1Mr1pGrSivfwq1bt7Bt5HNrJFwlnUYCzGpTrprnStF1
mgtJuyd0KaeGElNnUwNtVHj+hh+zyVHMVJgD18uUDbiBo0nPrbMrTUrAnE2hdtctWULyqDBmubsB
zDVicVlxwDTqm9bHfG6JU04oeekiYv/ACiEQqzPX33JFyyP+5NaWlwYXK7t689AnRZMVL2Dmax65
Kv+0CxwRN2v/5PLWTkVg2rXOnYPJHi0jCbSj+cLfLG/jqFmOy5oWjHmn/DP9/y449eqnGDL8Oed2
jRzhe7xadaV0rGNlDnZJbEN1ZoWkyqQhPUt8xcvtJvwQqEA7F6mlpeIE+jkvN5tJOq7JhF6OBtJk
DmMvsO2j4VNND6UYMaM0Yu34eRfKpCrfGZquQCSnSnR7zC0W8Ccx1A2kv5BXSFkTn1giTDFkWo3p
kbjKYFwfSfEMRUBOVcJGtfqIjx24TfZ3IggzLMzBQi3/7jCdc4fkowyml6hoih2M2wpUDOgDrJRO
01GcvL0F0w+PTSZfwQDoA4r/dmB3jXi/dhGz9SXIzFCVQKx3iul01Ro8HR6jmeLsRpZ8zHyyJZJE
mHgilWtBdBZoUlmatbt36d182+B5go5melpOXu60ehjj/ivdHMrQ52JGmJmxrwiwkSYOxSnYFC0F
YgLKVJll60lt+gUHbjFWCuWYEPibOWnG3JEoOI7RIGf/4ryKqUNZR7iNg92ELeQ91P2nJX5zbOzi
kdTEQTMyFgu07hqJd+692ro0A0F6IpEzcCQGM/YG3wdhExt8ub3dMKc0QFHlWv/HlwitMDnwO/YL
VtMppGol3ro728g0VZSu0yqVAuXY3GtDyYQJ04wfrAjgrwljo8vGnf4/qJ1A5Up2+2Gk20fbDLe2
lOIbv6bZO6OOx/qFLmYAgoSzxNI97xe1VFhUxr/WvZZSIQqxkpsbJ6J3PmoJUG2M4Pgo6fTKhUdw
IABlvBRrE3qhVpjRjNoDpFXAPfyfJsB0KYJl6CjjxFrdn9ivRvXxznVw3Jm2xnbyUZVJxU1Jy1ig
1NdHIQS+lMQCMlykLBiFrCs3+mAU8IZ8DqDf4MAHQihydy8eMXFciJxT12HHtm4lFBw97+7dad21
76vF5oGFigThNtZjS0qOTug3H96fbmTSJp0E7ckfL0eMiUf1vb62YFyDrqjoay2z2hf4iQ8m8qDZ
Hn/2voMi/Zuv1ujukbqLOKb6fhkfOM0WH1VKOB8wpyJtbjUUdoET2qnX05GGVhE7EoM8CPlaxYVo
s+eEh8FMUAc5HC8NjXKMv6NoXULdy8wc3Qt7heOd1ZQBNuWLyemMZB/JApoajN1OBPq9CLE/UYxx
l3VJiv5YKkaQVyTYlFgxsvFH/XiKn76zirHIGxb+w1Kp23KWMYf5v+P4LQQrOf6L7mj/Ufo9S9TN
O+hTeC44AmOzdcQ39kAljcPsXw1mZT/AYJMNHJyxOkJSDdRMRHT+THt+xl0+XwvaP9idqZfE4HGX
90VnXeTsb7Un1RHSpanDYw3jXAEyEbhYCsmOpn2tCEohOBBWTp6TX+wR053t550eC2iOZvEQ5mkZ
a02fWjloQZr3cVnPXuaszu/rfOfVfl4h/2U998lH0P4aX9R2C416+dtD4Ka7C0xZHs2NI2SiRR4Y
kMJLnbDBZU/nvkf1kj77kMiFn2bxvj6qvQFCNlpD0AQn6Ur6a/i86RRe2PB+arCtix/fYcPS9d7k
c4cOre2nLKr07K1bv1o7/w4p5ZH+vNNGX7F2bWd11DSTCT+ZdJDnRXKaHqh/cAROf8f/99eLggN6
Ynyc7jf1GkO4Gqnemr4PqS5wNqDfUbtfqF/TSJp4sQzPC/qk5D7X3//TztUj0Ns2XCTXvFdit7P3
ftiy/QA7xY6K+BBbgHJNRCkAtjKy1t7aHQZ7d8dang6u2Y0KwgQrnk3lGneXKkx8k5omqXyVWoam
t1x04J3fUOsuHoZkYPBXF0OCH0P0+/LdDqAoni0temJzsYIafYbxBmDfgzGc4Y1uJt18jTN6zmIO
Y/1HE9efWBZacmeiOFW8OFhprc8mOdkd/+baZL9MIRACuTnf98BWdToBQG4qOxjB5l8Wx77mcMix
9dwvY3oZ6Zwm26/ZNp5Q/xoonUhJ/m/q6e1lmTdbAZoWtdN6Gm5vNMAQMkbCbKMQjqyGFljpGkHv
r4C6gbtYJEfuhLOZ/2mKt7Jdm2FMudKjxnkbhqclAnf0x89Mlf94stqKeMj4LhMpOFbiX4RsEW0J
BWtggfOD9f0vufA/jfxcGjaMdABZ0t6v8ieDWXrj13ywvQWbSHmufEJkgpcSY2zuWgtyLylMAqws
ZP1weWfUm7QWbkvemP8qFwXVGcdgzHkEeAoJcucjJ2FpN3YWwXgeHuHpx2RaDlwL2YLY/+fh1+UN
dYPvDy4U1wCDxGXwJGlcrlP81rotPydqGc+ngFEJN2LRrzwoPL+T74sp6tmD5QfE7aKrT9hFu8Wu
gXBKmLckFos/MNilDH/0ejoETfyxDV4D9iosiQqduXmG8aEPu5fKmudQfQNCMfZusU7+a/F+rUiF
TWNuB1Rfdnn8beTYmTLdCOcF2ce5vlHoyGpEzc8HaLnJoWa2n6OZHTg6oMNiB/us3QxIfrVDSXGo
ox/9/mo6ebZjSbt+uYwVzZX8bvgznh+qqv6G/E31f75cC3SDciz5I9G6I6WlbwIZJHmk3iO0Mrwe
1NYlz4rNwzQZjWZL1pFUom6cO9CMV6XUMx8W646ZAIjnDPHrn9wq+8fHxPS1NnGOCznghcYZRbji
su7HHoHzEnTRY0Z7r7ooQho9QoCWQM7JUMsQi6QbapvWvv82tWxRmC2cFhfVtBh/6cyhUEyMs6IF
TQkdxUuhT44qLp2Vh2CjPSq8B67TeJZVPccISPb6qWL3ZqATNPcITaB3CnLmhhOhAO+NgEH55qsi
dojGmk6HyMD/BpYZ0V/FR0hSxna1xs4lSqC9lmuUgcWq/E36KIOeUVNZP8BKhGCcjON6o+Y/YnXo
9bSE4OpqjOM58FpDKtLLWD+FGVhrbtG/axjVZzX2sLBhrBe53NXcWLU1tuWuWDPOCWKhe7DWiUbT
4ETQhQ3LhOMjeJ68fdmpldmYJRJvyZl1IpSdLDB9UtlEDDZjF+mhvRgmDtixNpxhq2BwoUyljRve
5EXkUyAyHodzbJiUCfK5AJB/1QKdYvMxeqB90uHPs5Z5dM85GCDDi48YgVeuVnGzx5HqeOLaJF3p
fGUYliGbwZgdbqdn2BCwTuD0MVQ9fZ6I5K0cxml5gjQoOWNJia4v9jm7E9o4T2ETtTOZImL8rQ/v
XxjBk0NDEN8qfzIzhq8MDZrQZTGA/Oo5dR5AE3VBqBZQwe4DASD0ypGzCXkfAbZxB7wlon/paEIq
eM8zKaeAh77sTWHBiffNh1vD6KePOfpi6GmfvbJwePcfgCx6HbJ0aQAuB6Day+97YyUHBJ3jmxXZ
n3xt21ZIzVTb2XAJTl8NfsJY+smeUF5Lj6Cy2qpE1vbeuiaFqc6UG+BH9778mkNJGvRJX9jawKbF
/zzz4iWYL0WI0aaDfrfM+1QDzkqE9fKlTys1OzbhIYbI3EWcThuqXJN1fOkrYMKk2vUKq8U5gr3l
N4B9hpM1uSZ2Ggemn5s40m0lM1KNbSCyAWmpmhgh9SzRalOdOOhUEkf/qpnGYGIqxvppSbqkkZdJ
nvDPsdgqyEZ+Dnq0gL+PFo8odtwtvqhyf0UXSwelw+TRxIr0OM50asma/D/YupyLrvJVBsOOfAmP
yKXKsdLUYCWkNxYl9ZGRhEQK0TOuBZ3VcdEoWH6wK2mdjNWdIyjC9dY9YjQs2F0ky5nSpwgtogut
KNR2bwYve2U0F7NtHrJMy1v07lHbuk2tefn1RPb5grSBmr4Mjk11G6RkEqZ5slFaYqJflt0bUTi2
W87jsmwzhFmbiCbr9pe1yZR9/35jGtVgqSB1kUTrRfnTekmhtL4+LYeuVNZqI8kwdlAh7SUgTMq6
eklC8Spiq/cbJ04XDyFcqOB6fnojn55XdRlpY/jKy/YtPnPC0B7i8Brl7WIPPpqhuCP+xPmDGLgZ
krBjkyR+yxzzc3VbdwQ1gL7ZLSD8I4FXS8yw4+EJohtvOe+JfncKTgYm1yarR2QZPMabNXw1VrgE
WipeXpYgTWe2HKvruluZ/5207nEmgUUnoQWCqir7SPARkKwggR3QwjBPiiOuPJgNBx8z/mdNvTDX
u2Vn7N398lov6wJP6M8ubjZADDzn7CcrfC6IEMqmZnpOHOw6+5TluELm1hR5TZeHmzVVFaIjTFsH
pKlyGMJnFPh8w/8krpZEoDDUgKozJucjg/cvkIi3gaYjQHB/x5PC5Wp7MXzoxoSc0hHoRlmnQbUF
am8UYq+TJiT6O7qQk1BNsL2sMC4cLIK3nLfXeLXULLg96A6bZVvA3i6jv0exoPYptkj+J3R8WB+y
Re4tBNfmKNLp9h7Dp2DW5bOCTkHzPqnPcN9DO0npMZtR/BPKnV9z4Te1elROB3fsnlbAudkdHoUI
Aj7Z+6v8FdE1aBgGiJFDydvLjhTMywnniwOTOtr/F7GKi/XYE+BFOyTf4J6D9/v0aJHrr8R5K25W
0BXgI/Kqusi4znk/hnO3AyJWZyNGkQ+GgsN/CCAI9+sr7A7i9K2dYc9zO1JX+51DCw9Dfy8kUQpH
dSNa7Qs6yrcuXyP7QbMwB3Ch78eKxOPqBjlyKu7/ir3tIsYh6afKW0bRRTv7aLLlh9o2eKYYuqm9
aUqF4dRqsIxQJv7R6kLwd0U1f6PfKP9ctq8Q0D+p1S6+Ni5o+T7OG03aNxs2w0rI7Y0RJAhF8Ltl
sAUromP2T43/vpXjuJWrnJoplBWjlr3AG6NENLT/d1Nx/qrXkkm0xnXRJAK2DTNIpRn2dXJdahlF
b0wGmumWwhpVAzrFdsp4/Wjx+lH7Q9yHUXYRnDATLq7xvpKkLzxwLU5B+TAkNclDq9zkJg99FGMJ
HP3ZHK86HeouKT2BqWBUKOp8q4RG3lol1egQMqGGNaJQ61R9fJunjZ2KPW1g0DWAG0CT2YuOfFAK
VFsL38Bh5UGnxMgCRGyaKHfE0SkZeYJMKnwjFWp/J8Zz4kk0J2IPxoW6Lxvq/CEfex4KOmatsRs5
a1LhJXxCkgzE6f14ZtdhefjpX6x4UYPpbrYOTaYIgc+KdFW000jVlhrHfnbmxDWoOG5FQu7EacKv
ffOm5/fWsApIgycixvfmUbv8XeEvqzF8aWp62L5A6yInZ7pCqS2u5F9/88KZKnqLgzbnVfX8NcpF
p2rcbQcGhOAZJyx09rXCMEW1aTg8qAs8djp4+b50KiyGS3L46IW5oRdc89ymD1PS6h9Zs/0iHG3I
+zPZx1Lpxz43asFySrMAccAAIcrWKtWYUciVr+ML2MlM6HeuBHyiwmIai5M8m5pWWaKHa7Tf44JI
iB+mjldUNVVgNKW9E1kOmIqv1htqpNBsxIlQooo+WTy2IVA9MSU9WnYFEBIA6q2sgpvEq/P2sjDE
JxJIxh5D6UoZFGdqyCwr+jW4sSGC+vrr/80DnpRVUptArDCXlNnqRW1996QJKQRj4fQaQ9Mbs7Xc
ldZhNoFmgaWZKT0YRnWPYfLRp5SXiaZyuMnLzD0qYK4B8tMwUgqUeg/fWY/eHP3AJyrQ1Dh9ngb2
mtVkwyrW60V7oESwKftkBxXTNXx5YcTjLHTpBt2yDNMsPkeJz5AkbdwCYzLtmGxX9fwgLUVabujU
e4aHrtzmJv1voUR99kJuhEZrck1qVC9K5fFlDTyebz2GApmmK/nX2ISvq3xBr7BjYkedahKNxcy3
DiaFms1brNqZuzL5HamUYUozw/mfVhdZ1LgCb5FFK3rVkprXJnRRRm2Abd4Z1VfGjL1o/AzrELwx
gyt6CfNYOEV9tDyvSOaJZJrHUJQSPtKYUA6oL3cHesJeeiuw1kxHvwdz10mI48WFxVUTIEKRU2sr
PTjzVnwosPCmB2K+lBceQT22ZCycBk3hUrca+GzysRoBFsp0Rw1udt3LUKJT7uoXKk5yZ+TnLO17
olxXNYQ3imV9D2uVTg2kIaGnOybJuQF/EHxMddugANwfSLDUplRH/5JF9OKyRuV00TVr0PTvLd1X
8UHt0sy1dNwy0Zunf8O88PDvuIXis88LoeB2ih+2zyITUipIYnUS0xfbVf8Fs2Tyi26S9R+zZbpV
xe5r4/LwfE0joo5o51tQ//FZNXvkoh0zsPc+uDKa2XihCQlnZ3HaKlMWBdwKXk5g1eU4tMOaqQ96
Fxs9jPzpblvh5D+S2lPo59UhVvZMSy5/BbM5VEGrrVYLOkHfOifqboLkPkTSrgesbBcK7pJ/KkQl
mBXXg5csf55bxsA2kOrSoCyEfUeUlYtYYuohcsRR9XImiDvESkjT2e7fvW/4wM1+CuTlYCT1Olcx
+G3JAhE/8RIDe29Nvuc68Bo2YuOXlF+lVZXq22PXxfTFk0ujBlXGqOYSwFWvhPs+XlYr5ZK6Eq3L
RA5y6j53rDrRC+ToIge7N/IlRb8TnnQvROc0h3R1t5n+niXEYCj4nj4znrgLbideRhf/yYoxJUX6
KzQBc/InjsKAP9x/6CMdsID8zRghdScE/4jo2qmHeHA0ArUC/E7RxsxDbsGCoSNqJ4+qXSdU2Slm
a1TlNuXH4ymFp5SDwLr6w1ZjfgC7aE5lGOGJ/CLT+HnNjQPqbDwmi8iqrlEzIWsXmO9DBckl8uTq
XxXfSKJ9yzMkI2+q8PBC+SEm8a/y8QfsMPMt2p6MKZmJaRPHykCNALppmnvvpbJH5lI3aXf1noUr
c6f8BcVoumUWeltGGHv0PdySnHnmvJS08oboDPAf+JEtMh3hgri7IOJVyuqrT17L8K8EGurD4ocQ
YseaCZtr1PX+4xwbvp4oY+ai1uK70ZcWn/sOBm0vMYtjvL4VQGiJrGVibKRF+AnzbwLQCqaL2mR3
xx6Z+Y8J51G7Fqnk/cdhcSJLgBtQoS/vPeBKnkj2I/ELTGy76JdJiLqbQ37KrACZCHoJxYrvOgsM
thGpltpvSXPzymXMxG7QwEteqmemGAh+MX9FuRrLw5/ocNtr0vjBxPnyvchBjFplOEZLA3ASw6zU
zlw1HJVBoTV+DYNU5vkIoemCwoxdzb1adEIG9HIJ8QTn3R5LEh5YEbiX0c/lqBsOW1d8MUpIWNAh
WnWEcte0tDWCrI+NY0zXzljP1BN+B7rtcD6ESIBjV3kiEml0r79P4LnmxrayFZKFoS3g/HFtlFOR
drG+Z70KAuEsu3plq9HUmO6zOKOwTOXZh1guTN7p0TLlUjEvmpVmP5fnxgy0bxNg5hBIZ9LaYwze
ob7a+m3pcN1l1ldD3tmHEuyVwwDiSvmPkKw44cl3av/j02NI4fECm4YUT/nmnTGL9mZsl/M5y00H
GpP6DOGj93Yep++gzXyPUBfD01B++5eB/onH9ZX06QqLp2jh/hGIBrnZg0XBk77fLFpf9NJqfHug
VEFY0Srb8gCC0HH7pQD1/nat37qtsWOhe7+f8gANHx0O132gewzqlmHCr48p5gQvzDwdFpdp4oif
PAZzPmkdea4mKWXDsCiKlplK0ms93O3Wwheohc8JHIFsw3cRt8kiWjMNPM4vgJYnHJUJoxfiTB7V
li7vNsEpepCsnmDk7M9t46lGNUmg7bg+7DOnuxUi394VgiJCYVcbJ+wQpvv0FTiwkioVTlvp+EoR
is1FrlfaeqJvWhimyfWcYX6agZ2PyeUYUUbahpFy/YZJiphcrG9r6CbLwM4qid+Yn3nBKl9rJJHh
Uv+WqzURx1E9H7DCu+hVUZGG7V0MOU6ZE4i0No0ULAzyRPTO+6XSSVimEvUeOWN7OZtJqyKNQmxh
gPQO/3JcKb0BCT3xbqt2cGSdq+BeHWNTDeq/NyHxwImzn//8ah7hru2af0YF4URnimE5bXVFKjey
44zZ/lTI7Dg6rnjlREXf1A+uqyZP88uccymhZ1DNgSBcjeDR1Kxs044lSz09oFUiybTB8pyYEAKo
SgpNOz78fgDad4iMT7lDX8/Z00adL4vWId1AKEMIqtkMBVM1zenywPQG2QebjS7S4gP1PiVi749z
0snv7Z1mdy2w+5PuBIASzcDeyVt5Q38qtHIkiq3+pvQ3civ7iTABOmA60u9kvm4Z3iMACQkKOjLB
wNm7+mgcvxpo48tfkVXt1klBzoAXiftgCrU+YVKsDQLrV7F1JliFdil0SpKhM8tDK+cjhPpJ/zoL
M7izs2QWWpr5FRN/zFNg0+Qkg84N6/Iw2NXQPd62Kt3d0Wvm1p1JtNX65KuiiGNx3flSkz5CjtWo
oZ55hpPCrLeuo8GCkmmRVpbp1pfCSUS1X6GqkWl8uO4/YSPTPCrOpIEMxWMIDlXBsR5nwO7dG90w
LJ+u0wdVPacPZgdkZjNJWn18ctCFLvxGB2j+Z7vQc9Gdq83zpoJrsalgY9SF2+Om7tv7zPC5eVoP
ohjX5ou1oR1tBgy/MtsGWdUL4vb4fsooPbmB44E7T7dYEM4TLFdiib43PlJprExeI4IA+OuzC8dC
QwNIfFq8egGwzFSnGH65LOGLWSWiWapQer+mbXFBmuqJcLUkUxHJJLhejUSjs6XZeov2Yc/9fvbV
9M1XnJIab3Cm3Gnx9twnutK7ljaDxfgpGc9wwhFPx7V3tqWW0mM5+JSdjscHSA5kUBAf+wWE4Rd+
Sos1mkCX3enU2Ke4o7XxjPCMu30zRlMoVJOg8f55HZfVk/CZkGtHZJmITpkn+XXFwoFGSwDWxTOW
2aeZTIZ1+Mw3BxUUOGD3hQlJeA3nvJ2M5mGsDqCXWAAsvxd9voJGyYcsUuAnsLkUALF7/s66l9uD
YVFbJQ1MSBigqRTv8iOmvsmJtMrcWG+bzIgyHvP4yvSaX1GdLTHoCWIEQ3v0n7DFrcR6VI+S/EBl
feCsBrON52Uch6VRQnonuxdLzprKYPOK7Dgj1RZ3lrVcbJyTF1oWyxwHQtuPg1Bs8Z4imXZim6a5
t5/DEhvL4FzVyvQQLDjmqKjnuW0NKr0rQOtphNZAfi1E7jXkgOd4iHXojw4vl2XT7cgK4sLBqjVR
oVMHXHrKcGsh00X0AQzgihKd7QVmttStf/IMR74yaH3im4vzzthJzxoPi1GIUchkuGN+WPpiQ9Qx
peheKy8SBzjSJ0Vk0n4NsmEKc2TuyGlPXLhFuFwkOhzB/84HkAKBiCuBeAWwhGjbVNFniXdPYw3V
D8e2/40J8a7Ebhm+7CeJXI8Nr2QV5BSu9T5UTbwrwMBTRYMEhvfD4MW8pm26mdPftOSkOxiSfa39
yg/u5MUtkslJEFdQY7xHVmxZxvymQjgdI2rwYxOtoX4wgcU4j/AvM/cfn1XKvFvZZb7xDgrdwnX+
kBP2BrKkBNmdHiDrqkQdmW00BIo+GAhfVtJiu2tNrgxuygJIqi2ORzUiKTH+SfVRdJqEbIRw8ger
cd7Zhq213K0vCf3RrE0pQdlpIRTamxJUyfhPCCGUT/12SGtf9iTBL/LXrYHsQvpH9tqSD5qoNQ7x
Y9VQ50LYRYsSbbVP4kzz7Yc8/l5g9mS6AUB+KypsRAZ50mOFKWtedwsjFBB/EgJB18yMsfq4vNo2
S2n0ldM5U3Ov4rB6dsFL0c/88UK66j+41mfrWpbzRtBGRZX2J3WKkxgU21JNBle4VBHs90OFq7PU
6K56tp5a2hrvPUMf3N+7to4zn8JDBzVLIpUt0tGA8u/0kjJZ14GKWT1PenRIOJYcvaxD9AefteA2
oslQSIYX7KuGFvIz9wAsiYPpS9BX/cTN7vawRlMw+9TN17W/dbVx8HrxaP3k+cEGv3UPyjO/qW60
RdQ4GxPUwgsLhB+PWmqeNgI3I/QP5y2LWHEnyuaG6H4mOruHaYNED/Wrwl097XXq9A7b7tvcyyH7
riQAdE/6AfHCCnkZ6Ie9EaQ1/wpbS+wy+PH5dhquZWmFKyWH03e6oOQwHn+kVjfgmtKzw/bO1evj
UYsrLw4YvSI3/MgovjM0gptRqFEOQxtynFbSrynSVSGxxsLqeOtaoMPrApujSUh1PpvwNqvfQB8q
HZiXeMonkajywmgp5B0m81t4qKahxryae6E0NEe9FmJN2kblxX4eAC452XbD1yJj+JvtcLh0tM9K
Jwlc3OOWatHjTHHzfZn5ld2l5ZX7y6mtR30+xju9FABq9m+03IlWAF8wimbbuwXJFGk1ZA1Wfi8J
qrJec87yVCTxBhCQBnpl2tVH48pfmLBrsjrtmNXBYh3p2hJFXTyUknaC2u25bLzEoWex2p6BUcrl
HdPmCWUl7k8b4k2RexM1Pqr17PK+pSqMV90d/Gpd/5uAHWQzkAVtw4ONQnTaHfgpW66bxQL8EGFM
kGY4ATt1+HFy2+NfK73hHOkO7dzxgYdp2SQAgy8jZopO0DLJlnNddaxUeB9mZarPhTc6CSo8RfXs
juR3ZWJiO0XOv3rKUhYudTCdTE/i1jmKkaC6N9l5niiCbB4ly2GjKD3tUafkpwgsN2k9+i6SHFGB
bqdVEmq6V+FdtsGXHGtEpHHj14Cyn5VZq5vzeb/NMZCAzCEa8gGioIi2kYPHUCUSMY7xWg6MioEK
gAucfyZcQDxKR1Ygi21UcePGkWA/kTz1tW/Ph0Zuj5u8fkafaD7YC9N+YrMHRDKHRhMCDrBmtVmp
NjONTdtGrQwsqX9O0lIosxbTpN4GIHC9OJ2v9jrq747L1Seiz99CR6Mh3Xx7zdpg5fGQZyoFcXGA
oGNX8oWMzxeQIKuB7I5lQyEBbRltcRfXuufTA58Xv7EVrSGIeaTu2dHUl21PwM951o4slfWb4OjN
I1bQoAKVHftz+cCTpZck2VR+0dbsikZdSoPPOwgXkPdoxmwWJEAqY4bmQGWb8Z+msZII+uJfcPGY
vrN4GOev92YwvvYfjB6Syxpxv2HSUS8zEUagEqlDC/Vbv7eT8w0BEEpPTEY/BgeAo5m3nqBD6hJI
3teCY5otTpScmY/Bj9sb/98bzOtSSPrpsGWLlqG1/iU7lFYxmhkoKBMT6Zb9Y9uJKo4mZSk3tfCY
5b+0xRvbqsXsLyi3uJ35kGNn20RBH/sJk2DWmCB5QMZtjJgwCgzfQkwyTmrBfkGT/VkjBgsddwv3
HsGGtrQntgHAEY3VjF2Op4DyTDh52LybjyzTvnTD1PNrCt/IwMFGzcKOIq0jzlaVy7j0L1jjGFGG
00+oaHGF8dScSZt5rmIHQTI+DuIg6pdEQpOptWyVHRJfRp3R8iuOeXPGfvWwqjGwjrqtV1qenoA6
Bav2Pg1R5a7N/3NfpBAYTCd9BAha/KgkqBWTXlJKZFMOsTdwuBg+MOZC6xlbOs9iTkGaErsFc8Ud
B27gwReehI/B9fTnOdur6ZPf9u7M0nzhuS+S2tZSs5Rr9lLa8jNk74fTnDW9MsM7/LaCpASopH8R
t2fw1SDggeUlbFIa3KDD1Sr+LZhAhDEObepTs4RdQHkFQib2Gb0sXS34gQ8MdAWOebOMYy246Ddc
SPpfbj9VvOkVLYRDzSYtaqO+b/V2qwbFSerVt9Wcj0iLEpEuZNelfZEqyQ1RUGNuxlg3g6mw3NLR
hSGIxT5OWDcwYWM49wDzMnHapfqSk2ldaI7jhQnuOkO21obDGiKTAAu8y39RdKt/gQr7zqZ9pQRw
32xbBTxgCZB5WtI+BQAsMktO7r/Lh9tW4Zlpd1JdT5TS+fh/6nkpRh29TaUIFujZ7Ol/LjZOmcv2
tDH6sgoNrXPFVqL4Vyo5aTk4n9YBTofyPCkxFYwODxfKTNcIKr6DrpiChELGSJARVU6KFxrYUeBn
mgiHEmM8Z+aauvqaZZwf21ZZc1btMQM0Zhh26DmlJGJb7Y1dmbn0q27+ZTcxDzC/MUGK860Cjsnv
4UsIxtxaaR2ue5ipBqtfoq3HMZyLvZkqynmgQInZe1RW+qykJemktuY4frJ8zB+qa5TslPYQtjO4
ZwdDajCr7p/5vZWJsn59nBCqCCoPKG5DcLoi0XxQqowKI0cS27/70LlFd1ey//fQwV63tVfFV1TD
NPppkoz9buV4a8TLDTIK6B/okH+VHcETRK7CuJ/1q24Vc9In+dXng3Y3FeRwL8OGi3RlKaeFYAbE
iomUFoZrAlhYGaaMZ8Zp2c9MvSVG5zmcCRY/bu3iAcCHNKmlczdj+Nca+YJPrGMNsfoUxeE84252
OcHbRzeG+YKH2zeRe1Jdv2Rr7xU+xbOJY3eOqF8NVnifb9tHOH8FEAP7XgfajbADBZzYQhmXIHeZ
od8rxNYRMKWi1DbwYRXGyPaO+vQ73XGfTjDZYKIg5/IeZFN+7jcdFEE5qfkWyM8I6MQy8eEp6Dok
WyRYc49n+h0fE3toCLUapFufRCewIfTZhy4ReM5SXZyjDndK6V9FWJuov0yEjWKAbfsof2Z58gbq
WsQJLOlPxR4GFKNeM41uuBIE9pvW/SOvKkj9UxRD32ZLJCCahgI1xtrGEUYKXtD0hwLrJ0CzDkeh
S6Jp+ViNFpwjQ0KOKYWqHgYlKLn9xWlKoF/BfgySCqTptqNU69ShX9zmbTzvKauPlXQ8DKxHmxH6
0SZsHxXUEm0TbEt8vZt7xgfvThzPIrUHbCmFpqUaRP/x2zYaWF/DZthBMAavp4uAw4fbm/tpzMpk
E8acvrkkA7Xw3EFDXejewpke48EDnD7PN/tHtd2F6IQFKSjPcuO9auMbP4T+p4lC+8I+mDfSIMVU
2Qy25eZ9NnK2bW2f/BuajKRiyE9uWK8I6s1lMdM+Wfh0ZqMogvlgPechsGQjCcsf7CLswvHNfZbd
fuXf31M+TdpVgNJSVLvGP+c/hMHkOxXC+wzXU+R1cgeXLFWqGup+6oNdNLF5ejrmENdMGqGeqRrM
4vSSZ8LRiQyEAhCS92MHwqLOGc7tA0ECynhrPAyhN8WQNO75pE29vZ2s5e0tcq93P+YTywf/1NUC
esLJWLaSdZqAG5B7c3nlTvSlGIRBoYnvMTpVxYqGr6NsnY0qlwdFh4VuUd0ZGRnJl3FITRXMdZSR
5KRtd/rCaFflRZfRboEs0YstXZByaJAuR5/7k1caPKiaaY1wb1hptHTHr/Up6BVLIqBpnn2WwvO3
U2OdwYT8dIznT4RF81LOmpIUiSPsHare8czv4S3Ruok+DUXaU9s06c4082vg+zIzcydi9fd9Wy0L
ZaNhYNOMRkcCUZDS0u5KVEVpeqWDM8fnk7/s20naOfafjZMAk0C0a7ngAVEU0eY0z3UyEVjRNQt0
z/UWNzoBczT3n7W1FPkwbhQ+zi3xSC1GDiM7RRsSCYGo9XztaYWQIjYnxM4uwm9ulxPOLO7plXyH
FHGJCMICUbQhL3z9rw8Y7e+To/HHTf4jEdXgxJnn+TGvNzALfDYXIIPSOgHwtBXTFV97S7uoIWlC
ua9dqrOxS8y8AeMkfVpY24kavaYFqDiL5eTC2LsrAYY64Kv08l2vsAY2N6xq7oedlcxaGBHF/qB2
nePBLE1z2Ji4RngewqHKlkls7W8gFrbpJKAGKQGCCwfs5ZBQAdUI6Wiee49Ex8JC+YCLYRAGcKhD
f3dskeZqqPVor6Ro6W7Yj229vYUqUG+8SvpojcN9ZL1T0SX6u5Y9AMio8CtZfo1E8Q5eUWblLbJR
aJWt74jA2dVHiyuiQqWucMNU1xQqu/L4bUzvDyVOIMsIFB3M+KFZkuFGVy7WV98kwzQMjGtlHiKp
uCEpktCmnhOFF5ETSOFxpMZvaTa6i8BtIHkbxhcOPZk7RmMp6N6TJghadz5eK0mA4yzDudTSsCF3
7inJ7ONLVKysCRQh41fDuU9VKCAZreVlsTBh1TaqZ4VN+2QB/Z3SKehVjDHaodNBVAlI3R3dR7sm
6OBe/TdJc9jPGjM83XSGJ5rv6zwPfK4H6NpjG0TIFk38QQtY/hr5k7PccEKGxWaKSsqI8os4/TtL
HTDeyiC61/II++TNftmY+NKv5baOKPMs5HvyrYG542+62KgDtnC4bh/pVqP4HFBK5xT1VfA0fZoF
HudsIsS8aE4UwCjoKvaVlAZXfyZaZR4LAOdusE5ulbRidG8G+0NUnLVpr2rf+EIXyYlsdepBzq78
Djpw4CLczssl7lgzy45ufqxw6My+6lwYfpz3mpRPzn+eRv3nJ+rMwl2mMCXXFt0byCzapMPkTSZK
0BLaCo4P3Q6s1Saqx8On4ue5BBO0xIbDgtc73rO8LQaeVfTqcyzU6IIKR7zVEF4iU9YibDitHrwZ
KvO8SqeTujhxUBa2Bdw2wYT+RPwfKLt6+/KSDAT+QjSP3BFvp8s4wY8VHdfGiB5WYDD1S457eqAp
MtLUQ8wvbqPyQLn/bGrp5cdtK/fYdZ1PTLVHThy/o+3byGVj/KgcQ28C46PTOOWyhWmgTGfLUf+/
+5bj5dSnv6YfPKQ2nkJmWHDhgTDM3twiLfRktyB5boMkJ2aA5BgYLSnrt42gXiBAohIdBSouUEFd
x7EtrTbS9UKqfhcEgizGEf0/GWcsGs5rFZ4xS3cRlVleYrVBtgpYgd+IPWSd23K2K03noVYfIuA2
RgAA8wyGpbVd6N4OZuhqhhM8a00f8LBhOx4pIV+4HiSNw33yd5Ye+HXUWf0OUPSSF7VPg7Y/3JAQ
+Rx1L9Og7A2I0LoDCwRPwob0C9VhXkRPAMHB+StXM4TLzEq9v6gF1N8yY6px9RZ0prU29TUGlrLP
85MK1uTOIBuQ2Tq4vuceTXtTxtJP33HqVdBNO0kyb5cbV5xtrjCJIfL++Np12mYzRmMlHFQ9jsuG
Zj5aF5KlxkRHSrZWNtBN3J96N6IbVFbZmHPY6Vz6K6PfY0dIm+HpV0CcXKv04UQ++v2ztpgK+dvh
sSLQxdH/UflK2nltOKItOe/9Pa0vZ0Sl+nnyr6SWskKOhKLQvnuB6qzRtDzy4W40o9SyKa/A0BYs
KIw6SC54rTxmYwe2WcSyNi8qAbGsZEgOBuD0f566ooB3gpnrjdtrFYvFJyAqij7V+6zfUEWOz16d
F9sEQTwGpKK2nouiSsI4MovBqf2uHI3juYDWH9GRqN29S204k05o5ttDSL70fz9/QwFb99o/NjRq
WPJdPsE7FMDXWrEvyZdX7A7a2ikXMCa/ivfT30Q+KsTsFWJ76MPpJrRqELlBz8NODmhU+jof1An7
hbpwQ4YvFdTewSTcwcmu+R14V4ckm094beTjgfOxQ/SgcTPq77uBhqLxX62Jwkzfh59U5wxp9eYD
0KkbS6m7LjdDWwkbkTL5fXH9rSMR2QWqaUsX9cyB09dn3Xu4PUjrikxvHSOGGnDE8tJ6NGqExqYR
n9ViuooWmoSvoOAyzwiNpp/0zjkIzEjxYY6ZAXuygjNB8q0d+14679VHyxAmERP67APGvj3v4Xu8
bmTqI3yR9zfxcusv1qHlx5TcpYfpC7muRsmlykHMwzx3QWnhG9JuKhLoq/yeB4frPLDCOcX+1PJC
qZClqU8nWAs7H/JJH4nu10dxqBlSk6K+EpIxvIWrW72Xf5Kil7Mlhzr5Bf33EVf2mw3+ySwPKo7G
Lfc01HtF8u4o7On4fGkphyo9x+6xe6Klsm63gyMaBzUThWdiQHQaT1bpnx3vS5bLC1fl9MW1c+MJ
j2STpJR7SZ0EN9U0F1ESdONO6aKIsRiVYX+B0HYb/iW5NHk8+1CZhjfVWaqQaH5kSO0qtqHpgFwi
PqLHX8JSQtYhYlHbnfxQaMn8VZ0z53O8oNKFy051ep0BMQXC2frPelFJXi+j9pgU6ufZtDa246kH
ZlIA152L2gibmRta0AbMNk4yk9/YfneTfxw5AUVwyr0sj6b3U+EJXFcKiPwv0dOmgDThhBseOTbD
hiqlT2HLaOLK7P2nRNEDoJ4nB4kCF0PoYhRs3xM/OtIo8Ab6hCkkSHT/PAmL+UTdDEsybKEJNxjd
hNwQeUbcpl05XKpjGSw95w2XiPcUvT+BYb2ZMMJfrwbJVpjdQsrmzz7F1rzoqVEe2jxgl3tPpQUp
qHdpz2vrenDOE0+JF4TD0nSaLNeQNVCf/QbRvbGvC/QsNXsD1zDbyB8Q1j7JRVTA5Nou0jvrp2HZ
hWknqmuvkSWT7s9HO7EAcKQRQ1yGQub93y3q8AE0iDVcYr1QUk90E7k4rvsiBrIJrTXGW/TC5ybS
X5t9m4vgFdC8tJrJy2/SpQh3VeWOiKSZNpZNt9AeJ8i0QnKLODbQCE9F9QC+qO9U0QIw8q3rU9H8
ftD2liVCyZldC7moUu5/YdeEZ7oxE0rVmuG7JA8LOAs20a/kqGhEQcxpmHLUwYcVR5gzWqA9sZ/L
sbFwe8pyk66qShoggwMt/PFJdgq5ZfbLqSQvRl0Hf4xI+2DhwJih1xExy7jkH4hNIXDs3PLkmJOT
TvtPBBnkz4IkZhYhmJM8SnffmcGI6sclUMjUect3GnrzRRvgBt8SsR1L11VHRdI6GlK/jHkIHt1o
drqb2Ae/cUt0WXCdZAxfkNWRb1dNmI6S1NZPvKZ4RoQ28jJEVLO/W4cnJaE+fgqlw2+YvbtgYaWT
tdSomWFou5MTImxLavLjXIbkBU0Q9eVYLmalXQoi0YlTeL2Zj3rhhFt45mHzuWQxD22BTJyAXefl
5GE4XglG8fhQDdhQG0eHn8z6qtDPrblJ5XU0T52J296yVzwR8VYon0rQ/5f6WbO1ojNSarXm+e9H
C4Lv0e99c3c/oXwpm9nMMdMQ7DFNa/uvNlM+1MjSa9Br5nBBAso1hyq53QOEpDHemoehSPaWz0qS
XHVDR8uOUkXJUg0y1KVm9S/yDNFRdxYSUxnm+C7IJkXZM33ka/l1nEo+Msu75b6UzX6Y5MKckr+8
5bCUnay23MwSNv7E1UT9ZIdsA7GsxL4To35uoytgQKEx8gTMzEYKC7eErx6ooj8T+rm+anK4TPPT
M84YGuiCmxvpOS6Ua19SmhleFMiDJ4+eOtBBb82SBbWEea7GFyqvR4+HgBQQ1h7G0sAeFhlzDqfr
GLJ6Z2AaOXGLhwCG2vr6z/C5MwR9d3gkicdPGqbncvlEDrFnF2IrJ/NIg4qsSxoa6DQgsWUizF2J
MCDIkr/u9EdmtpN5hIU3/VegjuLh7ALdovcP2q4m8nd4qJvDF9DHFWa1p/Rt8li5apXmtXEKHL4q
ntsQJnH3aS7IJyMndTPePh26tUko75ky7kSRKyexLUCozeG3zTkuXNrMNbHOKVHWCdVTJ/zEBF8c
UzKnGSTdOW3XxBHt/+Fj0Abg5/S5yiLnNRcapJ0qlpxwPHmBAXH3AHmRugCkL0rCWznFsR3ifjKV
PpymAvImV5iU9FqYpeTzB81gfSTzBNYOQIFf25+gyiYhE7P1WOtIc6w7LKj1NERCogLHTTqaf9tS
F3awMmekRjEr9dF4MQAf6mu/0cTwdWXsCOJsV8ILJzjbomCNslZ8cnRoFN5NIVY6S/XxXmxktoVw
CeshNBvHBX6LbOKLEhnvbp7AM9TZq0Gw6LehNI3ufk6IonG2GmE+V++jRbG6nAjUUzU8rdRTmX3g
TFgKfBHUqbfIrsg42F+FyJUj1Zisqgu+msHs86bqBr9zYcDn0H3SUkHVdJn8tukm4BS4HpYD7Oco
hya03VmHWgnxpIYEiuDW81HdIt1cKuLXd2AYMb92HotOHG519Z5PT869xKOPBvxesKP6Xyg/ueee
pX/nJ/wcUQ32OKymfklhCNG5Hs3v0VwexTcrUFnxFj3ZBKBroqwxWIWILXpmtthfFIbM12oK0Tip
u5VAfuN66cLotRJ0g3gF1UOXfH9oeWSBxJ1YrTAAOg7C8ERnh5rDBjaDCSjmevCGVlmWbdophdgn
MZvIk4JLEfxaP31lG3nbq1Yf0o6K4jZu3zwAHM3IFt0MpzxaE2UFxeJg+5MUbaBXysAAtG3lnhsE
/GxvRydtR6tAZCS0cDPErcR8RZLedauTW/yvj4tlY8Bfrht1rfAEafx+sxvELr7JZgwCa8ePlhvQ
mUjc2syBDb43rUQ9biS73gV80VFA/5RpbwcnWDyrexJ85GAiQ1D0jJvGW1l+BqoP2VWlJCzoBY4l
RRn0zXoYnMjb716vEwCPJ6d2x8ufWY39k3X8fw3DVeOZkvaHdRdTAJ0d0MFFxgauFusUiuGtprAd
FC5Ush+x1ZvMIUTApkavb8V09yQThhJZZfdRyh+VC0+oQmzJplkg3kTTYH7bYUDRl0OCmpgvl0ns
mvE60l4DHETuEAzrI2o5EGmi0KK2+3d6Bau5CZrv0BmNiaWL2Y+2QxQeeOR9e4rqGMk+RWGeTdbO
0Zgl6CtU2FJ2t9ePu496pVWE+gh4/5AIEeNpa1WcQhF3lH9Q+Y8gSWbuUEmEfZfgPqXkenk516JZ
9dsbDy01leUtA70l8FdfZbPWbph2o+++vOmTM55+BiP00z4fNEVtW9VbeqDqpuRkz59VBJ8Y1Uq7
0CoVMO4CpY6bNLUez1kAy3qHs92tveFsNCzPolBO7tDx/XKbrSz71LL3nsqo2diHmsbUUBYJLnSV
KNKyJH5rK0o6xNmgnk0w6cA7Ko8Q0XKNan7ZgeGJyCSXUFWI1W84Q4/HCR87D9UrJ22tc0FAWtuC
TQ0xjM+CkczaJPP2xSTqYrYjRLl5smzZkPG6kpJFBs1NNxD1KBrer1DBxKXFE6uxAsSo3phxNM/b
tc7fLszh7GZ/noAVD8jJcXV4Z4qt/ISdInnn9kI2eRVVw7LV9FigJFqVNgH3hp7tb5HWsoDP6AbF
z0p11nbyCLkzhbCv79o0jkq00mOqGNlp8Pu9vwVn5RJD5YPTIw+ph6xlHS14ZxuRsSy5ywOdT+49
ufSHiukn2t8eqokZtchLU0ctTh4FIz2Zqbh0xi9jUQsv9613kGzCU7kpSraA/EqBpRq3znNA4TbW
tVj/0FLcuC7TbzcOIIbj42KIQs0M88pWlckVZVHqOPE17dPKeYhjNcfCYwRQ8ro6y2XB7KlG+hq2
xm4BwL76S48QJp7j/25+AZj24fQX3MBJqZV5dRQtyf/RLNKGULLfW46Oc/ctW4M8ewfSS9sAbrYf
dQPYdBYbUuQtCqpyDAE8IjWq/QAcEne/UpuM6gkgBsZknPQcqjjN/+gMTEE87+IjE6+nrIh5iNY6
5AxpdHhFNgzBp9qZxhx5cmXQTPMvtos5BjLehulgvdJ2rB9abxx4FDywevh6IbPBhyvR3jqt4Wgp
FfJwJpjKP6iidvKyBAClC4m/PifptVWGThACgAWOwWiXqvjCz2K8xmSQ9N1vRH9svzLzfURQ1mzN
RK7X4nCNQzDOi+D2kTzzEB9RO+XJQu7E99Lyhi9kndr6HCFSAOGZZpuT6oS9DY6la0Orx8XGnrYh
2QpjIBcPWzOM2fAP1ofyiYWl8GD6DXCZDQmlOiKbAnp0PnpoSxF4Sixwc6y0GbJpdQ7uWzdJYDzZ
N758r8O25fDpomWnJxOJtRVPXcAB54zydteqttwkZYLAxbiq3o2ZnnZekWOwB3LIFbyxnd+DBEeF
tc7YUZDAVUyYNSgdA11eM4+GeMlUzZ82yp6lAGAfyICyVu1UHeJjnNGVk5gskhWXxHLCqLkSPHb7
8Bo8/hKaxztMZkSIpDIpqEPBNtjL5g7gZT0yj9iVh5J0toYACpDTbKEyH4J81B9lSCBGzJEsA1v8
9EMFPKs3TtIwa/hUN1i9B+xVUII0LVLULSybSSD52teYH635wp7i6gIhJDbwArqrMHtRSq1jaS74
ZrtoHZJGCtHlk2v2/EIHDRkX+FP8/U8si7DVYZHYe/8BlRWcvQMTqksuMRMSi3fwit618aOs4t7s
+ZjbhDgp/EXU108x9BM5jpdkmKMx80I7Jnr8Cm7qBFggEuvzutfB7nNEcfxpyKXSgjJKk+veBMDi
Snv3TW1SHJ5nwvgij/daGTTPS9fZge3mh5Pzk3Uo4kkFvL0UzGeOVfb0jPe2QmFRAfbePz/cc0OT
cEycsA5gBmDVeKMGoyz4AKDoQmc7oNkp3m7iYssLpMU0JSPxRbDVwlk48mhfWVuMyizfiPjG24b7
CEVyUTsmb+manPue49tUoob4cxBgvmrEpajrvmE1UOxsq8k+b2caywEDmBqiNlJBuCiKZBf067kX
csfqiU3dHMKuEUUQV9QrkDRDeyelQZqG3kfMRax6hh+AbbNA2IidMB02vCD2X4QOc2wCbFPKMVJY
AZtPrWVM5LnN2iEhA3BQJwOEysov+WOd3y2Sl6i/Z7BYz9dplRKMTsiBunu0sTSUeMath6J7mQ7z
ACwa8QGtX2hwMaqBcNhY5ZZMgXUdkwAxpbXYi6/KlTzq6vMsXavtmEdlCz5EY08TG39btuT0ZJts
i+PiKwy1f196ciryymkRngCa19UZFNebnQLSj01k8xV3JXwbPW0aYeV4dfhBTCed2yia6I3HBKIn
rdZg92cyZQST8XEmyKHkn1JPj9ZN0dEcMUXxp4DBPbenLmQvMB+HvsAfx1C3CC3SmY09KCBTygfg
KL1TUYQvnDlo1WreaWYzrnKSJ1cYc9eJSkUNaTXWpeB2oD7BH4FCiVRMgQv5wDKur9NEKkXb7SQ3
NRYnOtdorTv9mUKNzgpbXOkeVWy17gqsyvLVZwQGvLqUE51g2b/yFu/ehbPShhNnhNvuysaM3vPQ
qGADPw+CumjjYwAJEwP9fp5QnsEfe/Abjo8V3NUczeRR4sdT3P21g5yeSDeZmv60zMwin+bhJWy6
hGxgZu31nLP/+dZhaamYrwLI+EdpUxWesA+VTelASZepiDnuW9ellz0mT4PGeBNC0ust8liB9zbR
3LIoTj6sjwYtQgYm9PY6IXdTFc4PoA673n1MSFLwePLOE3CH8qCSTw4LQwxVNTZZag+dgKux6SpN
YM1fx7LYztP8vSaDnlvUM5k3Ioj34iZ1z1Lqo1KcvJnny+LY9pInYd/jTiOjmy+W8aPOOGO3RlcK
U6t2XhfOl1dQ5ZD4WLUSfKHSUAjVBiZxEVmClhK4GET8bg/Pv3VscQdE8td4CUx7Zpm0FoSDfQzW
1SdqIVtIaFtNESzwZGx193F9zwlv4P2OejFM/GfMMqDgRlx8Lyp28o1dMTSg+35skaii5ErzlpJ6
6proS/GKbTn+Y2R4en1zI2jkO+Iu5D/o5qBPi0LJC0Dzokx7kYUmKG5sMwIfGGy44dheI+LtRe9V
uMJM/JHOsvScDpOqkzMuTmLWnugR6RwH2QpCXwaK3603p+PCbta1xc/09OO1hyHa/DpqVS5JRQ6Y
iTi55IYKC9TbVd1LOdWxUjs0kGXDJjjR3oYwh+AyD/p97zwwWgmXyC9QZPMzAwVq/Ocz3Thlaw1J
DViIpyPlFuUTh5X4Lzioq5+Oci9/H1eRR8aipGWBs8A0WumWS159Dpq7x3AGt1A1mSeadrS6O+B+
nCfx/Kaw/RBoaHScegjLRydfgsUbH8IbsPiua86G3J3n8pARpnNStS9ZwY25kRei/Uh+lDkwVxY7
9Dg/ciBDvDf8sifW9F8jobcgPX4yn514LvX0IaP5nxK6VtSpH5Fw0d1atbw9DKHsQKj0dA8ybTRs
nKdn31nwy9E1xHx97/Vnjdyyidb1PSoBueykjT0+MKugvCDNP1Lc7t1CmJIIVJK+IT/El/yQzNqu
egmaKkcRSqMdYGtrcsRiMPHFTHR2bJB9nDUSHZFmEVmAlDTldFsoC4R994ZV5iZWfxmkDLH0Cc+7
w1Iug0r5ioLbt0KEAs5xq+74PcEuZVd4wnh1ywaFRQydhWFO8PWJFcbM3jkJ5K3XzhQQfqXpRhff
5YNxOWk6iJAt/3zAq04ZrvPQ933w+CL3TXC5o3Ms9WSmO6iWZ9wutHJQuVx+gf8Q7dQkfWDGMkIe
/AoxiwufBMQAJjzdmqTOeYwetuYOb6UvD6E/IN01Bqy3OmzI+mTdiJHoVmcyzzzHzU3RPjCsaOqk
B4nwZFUJWQqaGJSQLrYniKpuj+NEWXQqHOJynEV0b4UO4q8ygAkIvikyTvtDqGjqcKeDJkPOB+Pm
E8WkzwWnXN1g1tXUJvPjBTq4x/UCE3e5yNk6NgjJDW5QBcKeodpKs7TFRJYeGf5IPz1R4nPggypA
j7FQbW6YfVI4bZk0O3BAVEHPUriLJ2U+gFO+vfqJuCwd3KzMW5MJWS13K6XI2z6XtPgo6/TjvYRg
bzHYUUgmLGN1E/hFtwIybjDuepee3/Oy5onlC9hJQDKNGErIINRLEkHF1MOJLFkRdwVZKml6wgt2
aS95rfjsvee4jtuuyIfUqUrZlKfigDhh9/Z9aYPq6JByz5ERNNk7fk1n+0+iGhyL7BlCGMjcdha2
Eqhm4g+mzicj6Q33/+MayUcwpu9Jlf1r6VnADHo+p8ZhVlpf7y2sCdU9O1zO3Co2P0ZmlYolzTr0
6X7rfPpsoE6BbZhMWRBRJT4N5RCZPkG9dVk66ap4hocKfIhGvjLGi+HcoK+44HcStKi7nohIBLff
Xgf+Tlix6W8S/gqMFTBCb7ltITObs0wKKous1bg8NsU/xZ7WXvjWSotVNmyccWNhwcZyA3Y9rf5h
GDqLJCjCIH5zf3Yr+oazNyJqQttdr+aH8Vy2DoeezCl+X38pjjT7sDJ/MzpSsGTCY+0pkF9/zwWX
eAHzPLN8XHTt4DPnA8igp7nPzI2EfJ8nqzh0pAjr7TUpF2NZivEY4EZ8t2mkeDMRCL4bkEVK365S
F9LAU18LR97SLIJntpc2WuIxI8n0nT4I9USGwm/qCkXwMXfEKgX/PO/Jqh4imwaFbE3R11kEdIZV
AcMiGvMfLCfEpWsgVro3YUxl1r+TzKVP/hQT4OpbJht9z9KHjrHCUvMsSv3I+cmITlk4NeTScJjf
MsB7xvrn7fVLF3oShOFSaWObDbUHnc6XvTHPb3ATfi5iEoHbs2RWinsHxDQMgkbA7GthcIr+LTg2
nncf7q4TUkQsRwlMkcqkA7VeU0UWfxaF+QZ7ghbV9SE/wmMD4Za6cI7rbeojqJ8Ux+X5NHvRIYMH
0Q0NWOdZuC9i1aJqvZhO/D+nyfmIdSmxjPAid+NCiWFT/8AiSa8pZ5DX9gAmGq9hjlfHYZTGnSDg
/IGgC8sfiQY00bBP+V7wUs0yrcjWP2DOJ8uUQw2g6CqodhQe90TZPw5Ksv5uf8r0PtL+w79hLoBz
KOsdAgINx0MTt/HNz9Nu18UGePvRDu7fqBpxG0wDWKXLdsEYSZtzgkUoR+vvzYZPzsi15cSZnuqq
LnXBvqnGBhfsL7oeq/twwbwTX6INBepu5FfwCty8jHBFWj8z3YV9vrC3RUmB61nWAzwz/nVMH1Qp
eS2cKUPMs48DzO7c1a0MOkL8F7XbQbBrkdE9kJl1n1enEsRsYFeMWgEBPAwIsUTheb+BVfY0jLdg
/gS9DkRWAU+G9HhPFxWk1rYjcBHgkeyalxsuBBPzlpC7WpKiM8y1fw9hIv3iB5zowMPbBbzJX3Y4
acprGdsyO4L8hdm5bDyIYc++2pqk0toTQkNEQvX9BzaZJtkUT2Z9F9Iasp4EnG2yJMJof+GMHV+h
jK6jp6R3MAbIBGa7gfmiGUFIxvavULH1lWhS/v3imTGjUjEZ0T8YTrbousLV+5t2K54961zIJ9CA
b72AaKAptz+dpCHsOkU0XH7KlJcE9C4ivt1rhoFkNureaa1CvNg1ZP5B+DCNL5pmZA+w6RlCALWl
QiWnEPCq3sXXs8QMgVKcGE/YablzcJrZrCo65Ob55pLLgS5373w0kolHRaLvx36sjuvcE6SS1Qeg
MH5PSkPmks7uz14x6AWcjX2fbop+BvQ2oUJ5oL0/ffDf7wed8yr7KzC+PYtRrua8zDq742K5wIJC
LEykWvUsl56qVYORP/okaDLSXPm4uRQKitDru7vV+Jv+d/nJLJbuLwRky8s7aRVbidU445HUn9Fj
fuP8lPyI4Unnvb+EPAWFNTqTaeebXvfoYhZN1DM0DDJUTfNBMtHTDuc12anVoawzSAmviUfw8Vje
OENkdL4BRAIZM5n04Ad88oOYLOAenJLernMiYPWW3SsWNoDycRtc1dAY8cwpZN3PqP7t3sFm9Td7
WEZGBgdMDJM3Q59A6MXX/fuU9hUUNlISVgCCDF8tt4H5PUXTmyo60b1CYDwkMOlOPE6IHOLw3Af6
kMBhIxnu1L3Ty4IVhqNoy3dOi2fdWNs1HGSeDHr3aSyUEjenioPFrmzeTlDHleovErbQ4hp3k/rP
WzpB8YtQwgBnWqWIirJ603pTXCPJIDPLL9K8ykjF3l/WUAEcp6IFH6gQdy9SVn6fVedoiwnztGiv
NXVc+yk9y7nc9mFWeTEtX+Cf+pEuekhyODR1xFuyIjflRA0e/k98Y+pUMK48diGVIcKRzZdFZdQr
2ZsMh5TltVrKLxPaVvCFynS6mcwKsc8ro1jo3yL1PY1aWN6Zkc2xTePd4R3Ks0BpVL7eBesTGxDk
JZ+GPBUi7CNSEJD2bwL0VQZnH9DlO2o5UAR1k5ZdcKV44ZJAEsep9nOJapoBdGLFKdR2DnYh9KGI
XZ5Zx8mAgJ/IeaNFv/fui0m5LR+AEyhaGQjz6Ivf3RxJUmybvyURREcw29hxIq7uc9UO05U7zbm3
C3VG6s5u94D34000Y+fc0i8IrzcD2piP5c0mhuKqCtzDQaYp2JLx1CH2iMsS1rkyVui1ZH2WYjes
vQaS4mRHCdfOYIvqDSrV95YxU1/zPTn2cRzxeMp/e6Hv4AC+5zriDBvFIPvkynYwgzGK0a4Bx6zj
0BbWwaGFFeu21rjZPmymBbgVJ1nJrJE+kxKG/FckGkmCwPybeQIzahi46fMEtGsculZQsBAN+xUS
T++x6rmOVg49tmlfvhTGFnt+oEfeqLKM3oS1gnV0hwi6sioi1MU65WUnD7PrDVeEjxiVaFn9QDEe
K9IO2vwA9kUnTpJU328Y9L9S6VD4HRFLqUY4QAlep1lupXxYwg5QKk2v0A/SjgEWNnESR6a3Auv9
j0wVJDWYABRMHs9iZSFfhVPLf40sheqI5ktMJta3Md/1L845FC76Jaodq/Nme6hh3v0METDW22XW
DocQcZleq5FL/bcbR6PDpfKRz6TkJuQ2CRovftwhxQs1QiDPy2zbM1XQavZQNsk0XZoe2Zo/TyBP
FGCQUGpcWBdLyMX34qb7tuWHuyj/qMcHFekMi9TGI1+A5/vWlLGKw3oWWFa6qyqdW3PXVwi/gKZw
KhadycBPQ4ilS5zHnBwWPQUG+y5ATSUXxg/3AiqUi7SHBTUrIAMY5f68YxPpVW+bKGdLf42TqpbY
eWSTxWnndrNjSRLboCv4ldgvsMbJ5OFmOu0EQxHRq9vm3Q3K7VTfFZJITLrfkJT7n/Jx2OJmM9Y9
F75O75bX7BvikyzGaZWFzxfeP/nk67tF15UpoyxTq5fRULUlx7TkCTX/t4FnFpDO0tWGlzI9YFli
q8mhuhfmXpH5pADRxqvk0e91ukbaGYy9cPEqZ5kJgdkWttTBmk0e2Z0WpuqTV+13fhtTFen2r1nD
SbN56//AkOfLiGyFH8zRQpP87rK0s2lbc1zsfZzzH22Qvi8bLG0/eYAxtRnI65wLpRg4H5NM17KC
01ETEqN5wAsma4yFgW2HJqtRCWSUA3Zig5BKSxgdgT8voSD130kcGJ9pIBEJGTotWkL7Cs2OB+n3
yMg1w+/jp2jW9X3koFxs4c+hlJeH0NQrUJbfKi8CtUb5W8mA2PEEpp4TBV8woG07uDD6pUTRRZNe
5DddiMgpVqfec8CVXu2oYxVEnNHne/A4+Kd/T6rZtx1OE4aEuj3do6aKsgzAOso5W7XfhDiCFjHB
zG1W6uQo7yZ5YDlUUGcae8Cr71UvHWA/dAyTfIZAjNEuJcmHOzyHe88WChreNqyRhpW7EZRqUyyW
5BT6l6/XrYXtxEGVGXP1LohREhXr+4J4p00EUOYbgG/a38lUWXYI/HlHXd2FfILFOtx0l+Ta4+b3
WtEcy52yjfR0uhHvbaEJ9HTV9gQ27GELyEXpBfoorpVvF9xqPmCajND6Fxv5Efd6NHDqsswzldTG
scmJHvzbPEvRb1E+WZF8zIEm2JTPPtWBJhdRSeSPl1BFMeKDT7WsDMrDltRi8r4DaBUjptwn1x1j
KOu16vl0Fs4Us20Lm8qDhAZk3ci2zMusYAPejwL8G26DLQ26S+f55peNxwPdLvrcvaFpM3mB8ybJ
OBAnGbOb4wOMPE3Y2i2VAIM8VOKacJE0rYQWvC190udXurtGfKmUV+flKk8fyitPcl1cNIPCzxIn
f9n1R/Vasu7/E61B3Jpfc6OtSwMaxHiz/O+GDpQicpPytCa4DZQbxQid8YrLimtrD7vPEGqnT246
eiPDf26UJuOaUOE9WoZWqdXj6qJmVGT2mjdqEpnPqSL1VV0nCYeVzk0qDLB2H/TVYwxsOBzijadt
ks6ceWd6Fy5IyhA/N0Ncoz/g4wCM6hpC9y3ohgpmtqAARv+sab8muQNmkQa5XPtwAgHsVmrKdP+v
gPBKlf9A597u/WM9dBkRtwA0htpnTfFKYb7LxDqAyrvY3L736e+u5Ogfaai/RNJPVSkVNvNRQ2nD
a5uWcLlrVbWSczs+F3Z0SsoQiqKpFkmWc3mqtcf5yxnwLTRH/gZaXHOenxqjzcRac93S2k6mOVSV
sO/DJ0WjUoSCUJRgvsbkvufO51tk9UvqheB8DKhLzgmSJoLz6b8OaRgjf8S8I/Wb1c2bl8UDeGBU
e69IeSzsNCJyqhQVyPaUWHhcbtRU51zLvfyiDYudHNB9kE3FfUNJJmg9qd7uGV8BR+IMGKQ8MPvs
TTQSRmslcDkEl2F2QaYvWVWF0/7vo1XMeNhTGdTBbFiuB0XRHAd4L64RB1OIpz0kXmuaW7D5beny
Bpu0SSUN7/JkfmcNoq+Ox8eT4YWGFlliI9nG2Bgb66hQTPJpgExr3cZuJsGu6X5B4CRfNqnzPS1r
EbP3JC631ye0buOwG585mI/x5P9Dd6zuWY8VkWnUxOoLzFqSYCPIWjZbwzaKwq6pCvhVVb5Qvkib
mscFbkZYPcP2+1Kk8pog+64hKzSmorTcX8VHXxip8DS/mdt9cE/R4Gosba2WseQ1+B43MgPv2sQn
o5U9lL4KqHLPul5jrrgtxIov0J5RRWS2jBbjgQjO7tOJbx3ZXmxeXZu7HZWKkJNET8h8Rp0NlQOM
Px4XNNHiDELH0tNVp9ZZQodPqLbVlXRRxbaqEIofY3tkmGFRu9gyOYaRqjN9ufsKgdgt7w58CFMG
asYYC7pFaPEQmZvTq8/zd7RFORvuKytC5lz2TxheYRfKCzgqp8VMQv076EOr5GPDw13QhjdicImZ
AfameML7fF1hU6ZeMW81fuYAPYsQIlNzgeZWBpItRI5AhTJz2RkrnCKwWakk1StS1ZhmyajNgaLg
pSbSL5otRiDggyr0b9+v+Kn/Db3BQbyidD1FfJUK5mNHVvsvT1UvIOncYJafZnzEDpCOaPBPJDCQ
xr9OuRkZIHPjrFusmqMVRhVMBzFQQBgN0jopvD/1IBJ80MqOb6o+KK9Cbk9r7WVauEJh6C9TnMBk
1HdmCWjA70AZvqwM5Rwevp0GU5xDH16WFzCKzgqz8rQ7UbfrIH3fzOKcnfl7HEpn2qSaVApgbba4
6NaG4EgUQkLKuY0GUZJQ+Q/5t4Xyzv0GS0/u4S38QhU0LUj2kkXWJE3P4OHA1MqiLMCEjanS/bmI
eNV0ByUGYb8i7XjkCH7ymLrsvochKConeZqeQ3C6eVE68qd7AOVN53g649T3JR+MG4zP3bF7vui6
h9UQ1aqbqtcLAlQnl9YzWd3yPSWGV4fdP8dGG8RPOulpNCwa6jxoyAlbg3R5PsEbLHVRl5eRcTQf
FoJPCxx8Ougr1g1fPQFPs7PwS/cJEzxuWiCX2QTDpmNwB2Zz73DiWBokOvUUSCR2JkknA7+Wbvlz
EcckO4COQdD4q+c+6Wav7OzxBurl0xLwZ0BRNK6NZezOvyeruHPnNDCB7hmmw/vSv9ohOz5SwlTl
itmUw4VgfV2XHS5Af0SiNVLuZnXD0Su0LRdYSOtqTaGuNIuD7CbNb637P/Qij1tviAIxhwirbT4h
rKpbItdOhS3byZxeE1Cr3oWz+S6XczeytTnEzyjvHDhorGbRkRsrSGsOEpX2SLCOHtdDEpKA9yig
zkN+UYV8HbX4gZXQFCadbvFLUkerIDPhwW70wN1gn3Y0DT0tqsEwsVuqvaEukpYG82+UcY4ApnD3
s1hhNdpOK3yrKrMjCB+v4eHpleZGWOnq6hShf75dYEwcNWWv23j4q7maxw4DZ5X9VFs4UwwW7qkb
gRrzjv7HRK8kweWsmDsZSC53UU+WFb04DaOjENMo/pqzLnuUUfFopSQLRQ+TDKdJ1LqDR+HAMiwG
uKZPbKsE4qtybg/DttILcZFrKQDhtZAFTxHgoPCpllVsdDLc3Pgrm0f9EOJmZbF+PyQo2HlU6W/K
1UMpnNySzKfYHlVPqpajZ1V+fiNY+MW4H6g0Nk84W6vkUANZ3i0WUG1tkksZpCXWlRfkiWLZtMg7
Eh7QyIQE2aA3qVXSvWkgEJp/IZGj4J9EM+UU72+CupuPg22sDCvyT2W946ndCnk7x71uplKt/DWg
KP9NZAzRSoxoIWMvPYL8f0pURFTDFJxD/KH+mscqgcSe/fg2KVj7rCTYgfqjU7CHvDY1Df1/gqHd
og3lvdegCENKnyj/KsLKmX9uICOb9fwBI7cONEEkCg/zg06VzTfcmJqtxgrNuXFk4SoUO5tXlCVT
6ifBTqsC+2JCwrIs2LPPMPRXH7zd/3Y49/hN2LWk9oZxrxylvL220ULGrvZ9RDHGVhoFIMd4lmCV
A1zYKf7bSGq499trqIXgiQqI6icZyjuwc2pLSglPSQO5c5+6Gsyjy+W83L6QyaRiy3o3UJv/nsRN
Zk/zi65z0LY5JHLhcbNXfSoGb2wsqrDWhot4fNQWzhK8Gk0JnL3l6opYxetrtcSuWESodSubnJmp
d4RXaxBH4KMNzMafAgp3XgYmgnqW7QitCsyQQcQZwMp/VJa9NRPEbWmcjn+q8vTBOLstpZK7d6z3
ucjT34u3p3sNEoC2irw4AvwVYfU3anbBiqEOFl4ng22W7sKlSVEuvv7ZxKEk4wWKmiiPhUoWvvqo
PTttgwbl94kXflqsMNNZ4bLgAXlV+YDnJdS1YsUlACtgaEFHNGOzEMdEPFvdGPBQTmoLlUZvXQHC
N1129LztDNQGjnSZNYYE6B0TfMcNrTTnOMz3i+tjXDz08LRjm3YmEfsGS3H/9/A4bVTiYTlIyVVx
5g8dGJ1jjeEVwJ09l5L3kUo2Qn+eWXE0xJhdD2ni2Lp5J9P5t0Igi4nMe3AOIIkpZ71i7cLwjHwc
kfgVcQ8m7FiIechbfE9fBRUknuFnW7uu4cHaFgpc4f8JlcGYglpf775KG8CrZrkTkZZ+3R4lS0j8
XHmdPeOemMqRdj7cb2BxOiJt0qsDd2TiHZsGLnW8S4YvNkOf2fDQpesC+bL4yt9wbP2CYPakalf3
642lGt7NYsdTILfReCpCVvSElLdIJEae1iLIH95+MCZKQDq4nvKZ1zPfyxRf4/OiN7ca8uivJ/Hx
+kZdEHi+w26fnghWJoojV6TXa/txD1AUjob6iFKIiZigtCT9tI2QozBUicEbYQ6wjThticB8YgNa
JR74jxCrbHexfOP4hvaw56nptZ/fVorbdwgEAXOP4jCQYdfscqDhZqDJQwYBTqlm4NKyNo9wlqsz
HqapfD58CDM9DFHYSEl4uyNeNT/6tYtbzUgmmynKUhJ2ZaWmrf3wbtXXEaNE7lW/qISkUW/9MiN+
9eFNoZMU4C3pbVdWpzkvFkeZtd00y7F6H5e7eYpGw+u/guvENJd4DVbbcMnGIuNCgdRYA2kYIj9y
3BrnwoJ0Li9FCASo+qhm4kUQgPMp9Lk98PlpYEDHW8WeLsZLfkKS5NXizgngeKkvUfC6Cs2crwUg
yAbq3b38o0MEGyIBa80ZKoE6Cd88Qqfit3EomSJkmsKiKqUufxClhw91bVRSUnsZPySiwjlPIdk+
I3STZbE/dm/m8ytZYXVi2HgECwANebd0Crh9mnRKYMRyO+EzzT+x2HwNMzXeOPPpeB3tGbGwYNWB
PDOcW8qdzzniLrRUBQX2vU6dQQ5nxvqyhAn51+Uh0hXrrMPmOzhVOFLBZdJScmZqR6q+oUBBr8VM
XR8sONM/8/gyw12N+EAJU5VZH56t8zzMM+3emFseXLqtzO74R96B+zokZigph17QS9MONAvBfHO0
W9Wpc0lSqlm3mW7wDA5xcCWfcSpaeSRCa7PSKNtfN+99+jdydrjoRnrujaa1/QGr9NKwf9y2QiQs
hg+Mj+FgvBE4Jkj9bvC/JBMkPWb2PdMmZbRxzA1Q5vH4APIbk72rcguIFvgAHxSEN3TAgrW6d4Xq
DiH80X90hl+EbRVeuEyKX0ntj/7aeziFovXba7eCamp8sEoGvbfObNGfkgbyXkgEjrSyVP+iN6MO
hJ5P7ttB0FyziyfQEKvdNJTZT8v6q1avYwpQ4SaYQJKi53thnsTcSApeX7cfQg27Puj3LY3CgQB4
IkK0HPOcfIPFLGPauraCVWaoo1viL0W6xD95pbyCiFCybsjmUOdbtO+C784NuLWI8oUQ+JmPzA35
GuN884nV6yKcl/iATXTN5DX6CgGHp9RU8UmVrxbVIU329UxnkHtqA2KUZV4GSjnqp0iJE5pVet8V
jdq2Ud+se6PAwxUj1IqSpdxfYCIQffRZ+LFj/Op12h1qwDsoyhLV1thV/uRXOHqdw0Af5/hGifVt
H/WDrf+D4ffMm5TkoQF3nXdBlIQDz53WF69RlT1CQsYYdXPi/x8jYyxJdSMcFikFaglFCew5dKn1
0LDNIAtcSPV1i8tccJcQMHYECs9jEOTCSYb2AkEq6iRI7oTuY24+14al+NXB6plKtzZO6WWaSSMS
nTA5M3Uv1QCtqbimmuU6n5vKAYfDnIk9BohIqg8RTdnvPLnzDjRpqRy9q0cWYrpmhASyG9vLpaJL
4uK2w/j5MVIpSF5qIpmi00cpHpsmGJhRGyd69YjRRqVYctxNq/KQFbTQTbJHqZtm3nGlbiEPydKP
RizG9CU5TWYCAq3UlsNF/eVedXsR9b5R2TAWACy2XoNEsgKzysslhe7an0xQ3PDX+/xQn9Ui9bvR
ab+i8LsNdxWWUxF0EqY+ACVCwT9qJYjziZNsotXhBU50sn9oVc5oFS6BKFvT1LmeeP+JAwJR2gXI
flVZ1QYfQtztHsiX084XbbCBtdg/dsUs4u8U3C4NZivsSRDpqILwZrvGZ8tr/yo12rIuZQ77zTWS
tp1OPZdK4GST99mMvLJMEVfH6K5f3VCmaLIKqv6IVjHCju53wYVmFDJ7Slib6NyfVJJNOhsibfOd
tPAj6+Ek8AnbE+LuZVKgqZiDJItMXd2At4J69xDhidSAwHUFBbiIN35x22ikUdutDCI6f1iZfVkD
Rm9HjOB9UqSKnnjR+faYrAqhinokyl0HupygF1yvqb4W4N3tBYeRW2vliKGBtz/tUM6GTM7sxUQE
CIy4NcMddscfC2TOqCPsMuUBlu0sBkeXHq6bVMqFYxZuVxd88CJu+yot1ZJsrK8r+3bW82NJOblK
P9ek72dKmrGNL3yCjjqc77YStssYPBnt1YRoL3tlYJOrz1i6enqxDxhIxdGltxLFrEyDsDMAQoDn
CJ+8il3zCsK7xQI4kxUN397IL91Xxnrj1iPgiKVZoA8wEPk65f2dE0AxDSLLq4S86K1ASYW8PD1A
MoH5zoBlQqasz7Dbc8OE77r9K0ohcRlfY54+/C3jmPTEMaMicYaVJaLMp7CYalnF2hAV4LI7/3/K
L1n1JEXeUwqHVbnOOgmHo6F9Ogk8gFuKHei+RqbT5wkKUYETaI2sT8sLNLBENXka/Xkfbqx7FSLe
fJCTrLi9xWOibCfuhER3K+aa7imyvhRyStAyWhgQ/wjv8wfP2be04hVMjEvf6UmgkjiAWIDl75qe
6DnhLABMwoErtN75q19BXetAX8/Wm+FU8ANwgnyYWR9oGT4QXaXpZDK6sIWwuQnrOfi9w4FLMNJx
cwTiDXF1newblPTM9+r9lvT4iEpHAENi9PBFVHDUtXPgxRxsPOYTwwNiJQQVf90gAYMe4phePl7I
IftVdwvJ2OabB3ShhylYP4Mb8+8J3bvQq8g57e4DnXqmo2F1Od5JNlYwZxlWZ5U45Ivm5wPFkM7p
XZduN5Y5MbReEcWkW/1OGhP60TAz8jheZk3/ca1oaQnJDhhhkGIsEwgHgkDnXCe0KDYlfp5IWifo
Hf+WnBb9gyxiTtDwabAb4fnIJh1EvECyifTYem3pCkzIHe/DCkxfbAtSu7BsRkxBr/ZlR9g8oguw
YRQeKELYcXQtX4iAN4YWH+0MQfrcIVlag2n/xAaY8B1/TSR+CtclVsLwU0rON1+oVcF7bAUGEPwM
lqB+VjxK5yqlD9ZOMeqGpiVrQ/A4nnSU4A0VBNozHF5w2a3krQQyiDvHS5AjMybpokaglCFU4TEV
0ZH/5SVlxyHxSj5BMnA1xkEeoPBr8HjWLQuFxoTQwMe8j8EzdPSEzuibC3VPEqCspztiOY4A8m6I
81rFrACFKXCyXjLvFsFcYi6ApB5hAqsVfVErf4srhp1QFr1tHnFEzQeq2SDS5PcAg6fFHSAQRHBb
830aQeAywy/JpdU2fWdiSyf6+aHTqUGQkcv5hvZ1Zttx4Z5n/aoyu3cmbuUp0aoBVX3kgw98Uvwu
Dm2aapozBT4BmHyzX5HivlFdZvwMcL0DVtUXaBjj3bN4W34IGtmmbpF30Rvk64zIMfdFZZ5W4N6O
/i02Jg74+WhwxxSabF6i6r8enpaxdsNYYtzxJd/JluFtws6iM/i9XFI2S1rP3xNl/RjCNhN1Mmo1
BC5ppUMZuz65wMdF9LZ+DZNg1zIG4RXfKehr+YBhcwfa2jcWT1gzdy0kjV2Zs4jqzoODto+VX6BT
i1bjI0x4A9F7bR/yW7mXiU1td1OgiMhM0oFYACntBmHrPyCsL46kDbTtYK8u3oy5wrgN8iYXZfvb
pF3fi+JoDDtdloNYtJvHIKqefzTVttTIBWAXITZMzl2azAxp1MrKM17TwO1YYQhBJvkBxRGTGjGq
2gUbDDxkOpaMZlA77sbUh3AAuV2e9B6qkja6danNfZk5znrchKWLodxEWrbWZJsvv/xmFI3x/gJF
GEsnZqc5gLOJJnMaRlNZ6cvJDA0wuyCMuK83a2GKJ/leUZXauJUZUrJGIQrAc2475sjMnGC9i+jQ
bWWxSjdSA4Hyl3/13OOh/ngxAOdsAxmavMKsLHn/Fck8rjQTX0SdCOPynT5hc80+bqu3sgdnW47U
Apgk3ED32okmvdX+UXFEv6euDNb0WMCm8BOaPXmZiz2vfe70v3N+YpLX0ysvGCfNROJUW8HR6Lke
uz3Lpd2p/g2ivgV6qpPocIjmgdv2Pi72AN16VaI5hleXgVsyJK6EeUbhnnnbCDP/h8/4ZMH4cQjz
RQwUThyVxhrrJnRW2nWN1Dunn0R4hdzGYIX8QbCscH0lOAJHw58MY6T9jaOjjzwFCwV/pF0EED8y
mfqllsGLEZw/81SoyAxmeKOgvc9XIBzj+ByqpS2Yaf/0MTwJgwYOnmUv/jDGXmQAu7riO3oMTkd3
NLB0VwdTO5fIsfaBWlyMcDJxYWAoEkRZdJf/12nJyoyuFa+6mjF5wl6SONIpOfHaPL19p1r2A7k5
Pjes3CpSjHxkPHwmxYf/6BdLqCscufuWNNe53YkRGLsOKNAUElU/wxtpqapVkLBRh+//FvIZAqBy
qNeqTFn/VeelrbQGF7iAbLq5eSvOaANHpk/z3Afh+ssTMnfjFoEVYxUbvbSRiTSi9B1tu8eg/1//
QtkA1XdkeWyi6Ys30mY2DDhArd4mIp7EToZhw4tmEO/PdJUwacYyHdCkJ5aIg9HQ5PbxJmbTWEfY
X/Na0z5mA0tI9+skYAYVAesfRPIVSaFe2SJYsOnbi1qxQisbb9pjoUs6MmoR8YwvlQaJ/mplZ1bK
LovNLvCXi+3IJKGWXZ9xL9kEadd2PTkfFg4yx2UGNPM2H39pW8khWKQ4D4T6N0w7u8TEfTf6SEkN
swuXN5UFba0S0EjrQ7aezB7bMJj4JAmmqTv87WnvhniaaagmyIk50IYBcyFn5qh3E4a2CV0NWqSj
fbo1ZE6emXHMIcFOa8stcpLzJH3wGp6RdMFPqzTfNmc+45V7YL3pj3Nu/s3/IlXNpMD3yOGNCkbC
2zokAbTXS8374Zj8Q5Zpmjy8Hzi5LGlscNMbAoLO6RihprpLY7SRmp90ZzV4WnXFxmC/cWdSoUBk
13fdNGDGfJZ4xouDJC81mQNi0S1OXiV3yECWpchpTADTlVP0CNlwgri//rwM6FBXnd9zXjNRubcr
IpkqpIPOT0ck/HJU65POKpHwUPD7/KP98jcVonsCG5hvWd+SP5gl8yIJoH1/fJycZ2Rkl+F7QcUI
dv5AL0GMTu99iMD1tkSR8xtLwsz8swQSoyNduyR5TiAXb5T5wiZjyfHrH6J6rkCfzqGOZ5agxy7L
OStKLr5AyyI8vJpMj7CUeBGn6JE8MS9ivdKAncvYJ3Ybn0otPAMalhRg9jhy6aLaAIGt48WENW6S
dhuW69lgYeRTzj+ZwYVBbGGVwIoYR0vnDzuQ4iIbGtVWlbnt6V9kq2dhoFpTzrt6mTyQx6pQBGoE
ckWifnjOziqQ6BCwIk1GLe2AQiphEhLAegjNwq1lE9rSfHzHrMizkL98CEEmabqCAmzs+0+/jySc
A/jaaeQkkZFZbE/R/JeNdTDIvBRXx2WPKzl7+TwAumO544ZBa0aaNOP0yQsihaFmtXZKJz4vUpTN
tB001AXvUt1Vnh2raYnkDSb5JBKbC9Oj+T8g3N714VBip20Z8TbMPNUt5HFTuG2ncwHSIMfo1leM
GaiFFtaiGGjlMhvcB0j3RRjpdigJbIi14pvH5Q8XEHnu029EQu7YCdf2lNMskAaO6KISFZgx1olm
lM0qC6SrX5QMQE7V6MxFyVxEJa8OQBaQaFbmiYgvLm7bw2S1cMHADvogPtUm9zseGL/oNWQoTUuc
kPeKm0vcz0Bekp3IFFbV5MMT1ZTTrNEnUijpopTI920+bf8rJZHuRa+P3dtcVQ/xKGsJ149/QIOx
JIpR06sIAH7PlfMm3QrIPyh93IoekTzweG6xWRqfBV+AvsEwas3MFWGk0zTkCZS8RB5t3V9R6Q3F
rM81PRHyHZHlSGbQ5uyD1lAA3eixP+IQWLO1VeJWyM5eJH1WBzdQB9gAdWNFiNIk3b1DocWAeMSb
LlpzRGIqfz4yzAe4JtIY+yA/xmbsDzEo5UcVZ94ghyC65x9mV4igAu8g5JcWyeFKzHtEWtm3Hlay
/vnflF9CqGhcow4mUMs1U7uZ7oOtT3QCKrAtJN2EeJ8BRN25AbD34cOaYYoO6ym+XuSJHtVg04UF
cc+RlnqS2O5Ue2ikZmxxbcPSbYsC7si7ZrdCeChteh+sWsEYPvrfTGoYETmF2L5abMoSIyTyCQlR
gtS9J+Pzr2LjxaIsWgkCFunPrvljQ3FJR7n+fTgaFPvzWB6hCdwxN267QPTuhpWATCn5b7fS6oLp
oxyTALM0YyaKns3ahKjO+26tSU/L8so5UmCbuHhlrfXYFsEFyfP3267QH3dCSeiKdwBBBEm5KXag
TRb5meAQyVqrVceJXoG3W1pjaxjM3162W0R2PRxMCV5h5M1KjH81vLt0gdTDeqCBjk/2dvAFuFgY
X3g/sXkEXODLRyfWbh1XE7B3LiXWeZD26RSTzQv8VCiTZtQEiqzXdDAH+PYc0RXMaFtvEe0ZNvq6
dUfnkKnSZAcj07q+57GUzqxxsCpe+b0W46G+ezS2EdYuTCkho5BjMC6Ja2TYsQI9YVV1SklodC8P
dHR7Tx1KVt23H+IAEu+6TGvDpmi9le4Bv5zfKFQshr1eDOFzF3Mvf3jGULo3GMe3MtNuZBQnPIU3
PQDN9JMjnVPmiO9T67HRShJ9EKCGLwD1PE9j/IH2DU8FdSBrrBJmjO+bpMQP3N47uoGKI9dMcBX8
POeMfnFzCpt3iAcmcemcgBCGGQiH/rT2VF9C0PJCjPbIczWDDH6svpn35TlEK78LSKxc8DckbQ6M
ExiRS1+ojBKBhjJWp/NXdySXDjFAUi1k5j/S6CMkqUPb4yKGsNEloXF1UkbkjU8cenw23dxurbkT
bl9LBbHQ+YLupnlm8efxEnsJ7Tr47HPZ5gX685WITYtaXPOmznT7Lg2ahOHbv9fT8/N/plRv4kUM
fKenZ03yvMg5WESXSBl7IAikRavBbHlLsu5NNo3Qlv87bXtxc4er+t+wzShOthL5AJcOhd70JNDa
0mN9Z2fTUihXNsH2S/da3GAT2KgbZenCHwd+cLfHpD9CM0n5DpQlLMrAph7Xmj/KUX4GqddHtosl
gNd3yFgC4OKzvhcfMhFfB/vUQzsFcHrCSsE0mKXoJ/y7McwAgyc7ij4TpSJ+dNVnu66/nu8Hg5fn
/UQndNM3f4Jnb7k4eVBsqvXTfPx6Aib24olz7uiJ30jyzotvdANlL8gCOz0FWI8dNvD3Gnabigqd
LN4qg63pEkIbXjQCDSlNmjet9W6t1xalDE97A+G3kL3eN06DIM3mYPYLK8hQK1ufgcC8L+CQETXq
pcEuvSOyXQCxAuGQwy/XEAZbIymFCp7foQPlyqO/jvIQnZRxViGL35krdix2nnuYUKxxW2sNX9zx
kASJK3XTV8n10GDRSbXpqRLLkkenPX2PMIRTE7nvuBSz5zOgpsDYEmqmib1hF2bubAwTnQwAAfxE
trb7fuo6KySECkAof9SAv3sL1fv+yVYLsMItGiaTCqeqGlZBfcikdUsCsqjUboYcpAXmDhPhiz5j
R3FRll5f323jvPiRI1jmZXyYyA+crgsO+WjLw+hA2owKACwbuL8g3D1j6c7nyZJYZ0hmT85gUh6K
EoAa7LGWxUL+vojX4gILBJdj0adGGcODJDQX6WgrNDX2YLl2695chUUszZLMtK2nRHPs3L6wEdZW
QQ96JT+svulc+sbn2sDZ38F+QfQj7kQcJqwHbn6m+zD/S3L+wUb8vD1PpEldGALiB/mAvLhZVg4u
rk178qSj09fF1MbETnMERgTPjZRCujx6enNBxtx9KkDKd2JFL+zSlmrR8+TT7IwxgmlpXNwWDobS
h/PbDKAhzy7F+SAIQkdvm7Ned/aflyMY1haMgGkiOAlpO697n0kKGTPHxeb9lxClOJ3Wo69hfUCg
CQeldNsVZ4skdEIufcZGitOorsoBdU3LHwBTRUeKWagh/1OCqK6PDiQVKSfwP/H0LWmclIstPljw
Go+FpHVx+eE1ocZVR8KPBCyb8FwDyPuR1cHNzq5XiqAAzCGu4fd6oBKw0OyhZA407pjW0PrZrADc
uxGSJIVpQQdbSgDiXmty9QERcQKyyWBJTPlc4zQyGEof1RT1A39QuU8DyYDWyVRCZJHuDCKlbSKB
DcPOcf3ydUWrrJfDWMOhpoPa2AruegLNFYCbOcJh3AwqyTjSM4gxj33YTVrHFop2Xe9a5D+AZOWa
+zc7ycmRdFe93o08wcn7aXkGW0POWSkkSevaviTOPwtHMhZTVZdM184OwCfjyikcOJkRso3pdSDL
pI7o0xlDryEhnLdwKpt0xBEW45J6f+4Faz3YSkengG70jrdQd1vhP6ysUKd9D6ZDze7U8l96b9cK
uc0+Zvmfa6YGPzlic7eN0wxyQk5+YfWC49EmPJ0yeK6cVPV4tPl7fCKWiP8irr+KEoi6kIOzGa8Y
tu2ah9LgQb+4iebxr7fWsxFLop2aeo9D28nMT+CTF/yBnMh5cvBkD/XqbhvNNK5LW9VGNIX2CWsf
JiUWH5oVAXagq+zQZUWt7XsMgFqgOLrZotX4jUAoSKv1mIk6e/dlvIinQEhwrOKt9i0SBbN70J8i
tuttChwP61D1WG1tWDHjwHgPyvkm3xClaafnEFG/YOO71SXImqXpLjXS2k63xHDoB6FqeQCfCuhv
eRnvuAKlLYyE84c+EpYYKq2uAOQBZ61FLIh1SCvyhKUy19vpYgJqo69KJAM004BM9yod/SJuL0EL
8PA2WbY11u7uWB9E8YxGJTKLl3j6heTwO489jUja4TJOc2oK8J16x7OENFBNpQ8/GEpaK6bCoBeV
YV3hwOsYsZjhUp/YHjZyS2G027v12MX4RWkLSSpLydOG8vmmHi+DoSxB7hsmWSogwVV+ql0pU76/
saJOind8UJs5jHkDKbLyTHlrdGJMeYTRl+A6CwDscNrk5w3g/aWMPJ68AJPJifDy/6xInYjxuUqz
6qlkaFDwNGbA1ExaZZLdirIo7W2QAV2GID7GBBmSLExnQslzy6uU1OxiqmX4r6NoOb3JiPlcMAvh
PB5vs4ethBw90m0+EazN7vPtK+DlptTNNKhEfVOtQUnanOrh+j7jvnxs9Gdh+dFS0w9g1Ory5B+k
o5ZMo1rupP9Pi7LeAR2Z/ftIMKwlqJO1ZQ30leodfcoOj/FnGF0zdykvZSouGQe/53Plz9HV4ZVs
ijvYhuZ3JcyNW+0usbWSyHv8MaKqfesZmFjoD1T06BB377x6L7ySMLrIDXrXGGKpShUv/fRRB51o
E63JkVOEUGyAcZ6w4UCgBvg7Hkd3FzWhlzntMoqaXA7ChNBVrJbWQ+94preFND1n2OHR79oucVhc
xvRquDWsYC/2ki5WiNdR8KVZcGCU1oQ7l1KwCDRudZI5nLq0NL2BBXztJz0CR9D6pj8PH4v21ZgZ
WcZEeYUOxO+Ry2/hLP6Wuiqdzs45z6oR+52NzC0EbzPrrIX1BhzLEoXjw6J9eKbvLzQlnEtBzVCK
s5J3MTcJSxsFg1iclBxVcoKsf08Z3UELrKHzwvVHgkuPx0EuCDoAzBd1aj2bfi/ArT5emuLmTL+m
RPpK6NbIGds8pPgv1V8vusv3MWtxLaLu8Rs9XCqhTA/f7kRFrFRL3GyAkSBGX7u4g/1A7sQZutLC
w2fyAwixEbP/jsNVq1uUxLNXNAslTconJ9N15QS7zuSngJHL0Wk+s7b2rLjiWl+IhIjfmUyKVLsi
GlOGOU6wGSJMRNcRuMpwEJQoDzG/B8GbqcuDKPYuF3AxZRfoQ/JFAYBf62rp65VJQvLss1vwPUh3
a1WsbHfbhu8Mc2esClylIgs+chX1zDtmEqsxA332E6FTlnILqhhrpLBCuDJppo1YzHTHFJgb5e/Q
R0sTmCxUSD3ZrIn7l9U048yCtVhNRc1PMcI7Bc9jjETLF5iCx23y9cYS5J7gnBgBGGm1mbCEWsLo
HhORMFF+HTavMysw37ekvSiFdAbGTbp+YQ0QEMW+DqzM/r1BHf9qIZItJB5v3HR8lXlhaR2Atfyp
BjDdL3mHslj2c35DS5R7rcFzYvXkUt2ioPwohVuwcbiRIXKgrRmhue+A0A0o5d8tL8SGlNIojeDF
Z1lMidD8Hbdzsujhb2lLnmCl88SjBj4aq7svsD9VRjAxBmeI9z78Y9shtx9x9O1NcpzNeN6bs/wW
avVAvNcW8ZpD1T2+mFUxUPAuvkVpzp7UfhKSovlDEVohNj0EegJfiRcH6xyN+x/W7a1hluCqxpjT
SdPfOuDOcjrqckebVvqm7ZBfH2dds1taCig4eXcOVQVL3b2OjttzwHjt6c9p3sTpFh4w8RuPHBJr
eT2i7yvhTBugNWsPWXzswowxSll16O4NxGrYCJ22OAoggVUSwiSKRWb4R4LOM7r+WoE2gvPRKro6
lfvNyfnNnCLQU3UGpI9eRfnrhBScQDZnCzKy+gEJNMhPN0TYvB48DF8yYw5oJKaH/tbpmxD8/FmJ
ayN8ewVxJP3ETIjQARrxWoswmGSQ0hwBhn21+TEEo3RWL8e+sT8pSwagkn3NXvat3nhoWTNvrxBe
Iwz1hkucBFiTV4AyuiHCt1t2cNiAhJdCO6d0YgfkyT48BlKlDvPz2KlCGU7ixt7OucgyUgiJiZjV
Yh9NIP1k8c4dSthYqWVoC5WORrGwnXXyAXpqmAGsQ72kBRDLPRfkOPj3wsyX4jcbwhuWXK9bfEwU
6HfaSN4s386SBw6AZcGdnNuQpKSAhV/I0XDlLeqLxbldoM9K0ZVt5JCnnvw47iLDfRuUR0tAFNpX
AMDCkEE0zMyCrx/VyR5oJultuCw2zeMIouPU0aKkjcQ2YDVKE4SpDTPaQcfW5zflZmekEH8JiqDF
jKp75K/vV4HbVdrJJRBIMJeMyCRI6yOkrfGqLFYTpyoGNmNj3pnqmu8AM69cDtlQvM7BYCI2CsxS
mH2darqWT2dKoE0Yl9dECo1/dOAlmP1MlVVD+4WxSY8kTL5NkcSgvnK8QZOyBOxctqw+gfK/0Oj8
4+n8ESggaITgGb1q87TPqAlUIT3xxaQzV2y6Skjhc975p+dlYfrh5Gzrp0zE1TkJVUAMVV26bqgd
un4HapFKpopICimzNua2scUk9NQ3FqAu5Nb4Ywf49FanBAoqq2IkCQ9xOqVYVp8Z2Diie41ar6WN
BzOOd8QMCFwjZnbve3dsRr+hK0LRw8OLbGGDI49tcEdHbLPhS70fLnoagrCb46xC48n35woHgj9s
XHuwFXZHKppzBH4XfWtWq2PBArn9rGKZ5YGkwiwtSjVIadZJ5izsF1nQe75kNPdrpLm4Q2Wbf9WP
lpOExVDJs7hp2yC22WyPSVexlSk0+YWSukrwgnF9cY5P770XWwPgKcHHCL2jif6N7H+4vjvyfEAT
+KOKqmF23QW6Vgden6JGDnox+qWim8vwY2qEAuysE1VAm9gEsRtUC+PRRnplhEaTyHC/OTr9lRid
AA/V9RkarzWlSnIydp9XZ5D3ogfbmvm+Sw/gX61GBElp8rwm9jtW3AweEv/kRJzVNXFyzYY27OX0
W+F0zIu9ZnvS8fEL0BLQ1/zTkCiFa0K6heVinAuZwKx+4ng1lrRgIngaxR07ujWxqwO5N4Ndimyj
6VNg/mt8nZGiyPecMy+QGq33GFsq3bH05eWNMIQvyUhwk0y32oYpzqmMf73N/jff91w/WSeEXJJz
Ro+MNxhxnp3Jbnx97AUBW49UlpiCF0/cWDyXNtNl64f92cf9YwWtruPkwyP+TIWaR0YHQgrzOD1q
4bAiRdIhAfOWx5WHNokn11IiZf2MB+HmSmry0BszsLVMxWnlKtayn0dqTouLCQhpLOzPpERqeAjk
Buji0eq1QYq+3ylx9VnCY8nBdWtet6neaA7gmqAPhtABTFqUI4Ysm6YO6PNzTcx4X7/8wkQsNcIC
JzHxa6uuTwHjDuhhrEsi7/LDLv3jNXUm/MX2BQac88LhfU0FMsRQ1RWYvA938xN2as5qn5zmJCRp
KPKTlTEpkWl/oOcD1h3J+SqUaqTaa04JdXiNkd80DrIKMZsNVmyaXFwqJdnZIZHaHk/XELGJfFu0
Xb/8kOhiNbcOT4JBz3uVFse6pGG7oTFRiD732prwOMhwIMOVzHd5Nk+4pZV8QR0WAnkP24npLe7z
28bIZvO8l0VOD3ijpepq8g1mg/DuYYGeKjHybmRqp7VDkEtV0QFNjfgsyt63XNCsQuj4mj/dbJyD
Fx+o3TuQA5NtbEn9t5ujLpdVOdwLzmC6/it4Sl5fwhyT8Q5OUM+uTzHKb3jl2KL3F57LGsX/b9cd
yq9kJPRbHFAj+NiDtti2o2vJdrUTjE2PKVelcONaE2PjFWYQ8g63uQAxAEufpGCTXj31oVRH9LhS
NmP5/U5R4sQRdBMpyVFqMgMQNewB5R9TmDCRLrmDbzw6210cKz7UIaBRr46l2OqnQVGJJ2pHxRii
X9UN+4t7wh6nTPk2QDHMiMOZTX4nuYBHnV03+eFXsgWBO8Ads2FW6m/Ewj1J4sl8Cklg5rAXN8b0
ysxX7D84KHr1UWoXl0m2leoWn/rClqR7tAyImSufoc3f5yTJEH13zQ3KNI1+STS9rmfTOWCh2UvA
xEEEzLnxklkJwKiGu47eahh5/z1qIQhi1NKjn1HLP28OKb1S48BGmdsiDqUJ1py4JhIdGUxMPsrW
Y6XF6mJHjnocBByGM6q7QZtAfQpjhsFu20Jj3cQSjJWtpN46OhgGQObzYazCO2eyqh9dENFtHk7i
6EcR2mqMLqj83C/J/cQU81pZ0eCTtm92WkEx1Dnr46KST0xDVSEyQFDT7FBOQrGg8OpcHqQeRFYe
dLZWos+wKYib18UuknKHQZrCQ3nQ3PfcsxgmU7Yuf94m3YBOFti2IqYp5BPt0VJlu6FjhX+DqKu2
bPnpHjAFgXVmCeOiwUClDUN+c7zYoT8V8QlWoowY8GWfa75rli4ClXqwCfjjvv/ZFW+2IDUMFyI1
jAZm8ttNWxBotId4vMMfzyjLfF4avVKxtP9GqqTyUBvm9PQyE+7zphbjinTacU3533qDbFV1GUxi
hlAud3B/7ObtdWvuFABh54yzV7RtOyDgIL+1Ut0QvXSDd9mInmSlSEpReHIU4FsqFjpAsNUW7xSu
6l5PSFH8xIA9/I/NCTgE9l5/GOlXggzMVLmn5xpMS3ZdBC+YGyuqdbDLbCfuuSGnuI0GAW49vva/
A93LI3SwJvbniGRkeegzSNdZO8Zy50bi3X5TuXXP9cOl3PcOdqtrg8Xz9FwqN1oQPExGkHxPzu2e
jDMTFBt1mo7Qtp3bGMO74gynVe1WS4lQm0dyld32ANkpFlCxaOLGL7lgqAnUTPeDKGTFbYCS5vgQ
q9bS8LQXl2dqlrvckfzSGMT1uW8s2qCgVW9HL3jZctuv4/GVUwbqttTH0t9ob1KY9+1xHek7aIyQ
FjHrqkQW2DZn5/MxNAT4hUquqP7tAcpJWEsiecbM4kH4kZ8K1VpUvUuav336Sk1H8OZLYAADEMwb
Ymo/pi3OvVcSe6kA3nosQq9jiLkuo3euwmXzLTtchJ+ZDhTYYatbsaYyZgf1A4/1i898mpnvYodr
FnyIlIdjfLHilKOK9lGj2haP4s81sjSmWyhOhDHgQdSi4OeQR50cxutbiKpPUkCtDvEgRQ9xkBhq
4JXqZ6OdyCddNZup7cTcQBrRwZoPuF3dmUrhjRsl5ASLf5QqFUE82DWmLCmA6Ucyr+FE8qduNchp
9ToH1Ol4YyPhXdMFe+HKlUVMjaCbN4dLnFFKPfQmyFOc/LzMpmAt7SwGBwN62lkOQSy823ORuoQP
jCXdU9urph2SOPv1zwywenbmslYYPa0zerp7SrFkuLUnn5xJ2IYxSUzvtgmlAoCDfPNDdDuTnCrz
3Kxmmu9p1s4yMn0rYdKzXW1pLjK1fPSRQh1NJevC6QdxFL4oM9DTn+vfeNRRSSYzU62j1miNMg0J
7Jdt2dTyO0P1izV8G3yA/wXGBS4qWUyPBvE2gUTUY/4VOaIZErq4zhzaStTWTw6lEJ4YueVg3gOJ
mWRlWQciwod6MQ/1DB51N1IsHtGekrZkqxnhaHIxm/c0pmfAMx38+bR79W50nfXGtINM8BE9km7d
g8KkT52slUVbxERWXdRc0LmzGqsY4H+4eKLvO9Qh9z1Y3rphq2apyNWcsarxY4U5eKPG1/freAlp
D5vJXnTfzlCXQSNzGHRkB/j+Zol14WLRRoYGDgIpXjGuQ+x2myUbWsscRJy37QSfNAZVOIwYs1VD
YOn55CPrjmbb1dLD4934wV5BaP9RuKkXtAyqHlSIRJfAat21unhaHlzbDCw4T46DDqoiPDzW/QZ+
yQajz7IHZO3du10Fqb4P6oE6NWEUXcdJjpnNTqUgAzql09mFw7bhlCGQSL0z/Z2OfwHP242oJJJl
VI3sTlBDNk2MrMXQZbsw20/QQw7doh490+am1lcJNNWwzrZKbokcN0M+2WTGZ3FwTdlTl9VcaZa0
IDWdZclaxuQaeYZhbZybJoknkhDSBGky6013yMN77YTplJXnnDSAjyAnHxPcU3IqCH8u72nH7ksZ
Ih59aeC9OFSVoeuLW/TMN124/ncbah3t48VvBGuqObo6Frh/pDcbkHJjE6khyQnfN1fdGH2oLyOr
c6ZLFV+BpNQkfnO6p0cNrZRQOXFrpecL88P/lhWbRFHzoTWM0mv18NmRM/5ZUuMtNHqq7OwNt7h3
lozusL3GZu0bIbABtnVSMCP99S1B2r+wAKAuevCfc5T+ClxK13GtKM/Sn3ueurVSqbIM8gqJUsaJ
XkOYDgiFDCZ1HDzrzVpfbThz2THiDJc9xUxhhRBmxkQSftq7piwEHlM/t2sEHIUWjWiXOUUdoqll
Gem9p51XJBCDCbFFuQHpbezHgCC72/wO4aCR9P6Ph9qhvIvFevmpji30X4u5gPvjfZIJCBMba73a
DMAiMClgDZMzFEbFVRAk+7lmzXLHyn5UAdVq4iJmQ42M8o7/lUWk8Hr6MkIynekwPG6GZm8pRK7A
o7GELMBpKamUEkFoHxyvyiA/qafLZnZ4WcIWr+xtYMP3qXfBlCZ10Mnv52x0oHMbOS9+WrbmyZU3
UZkPEqD3FL57sNrlLykfuOT83T2PrqaLGj1BIbXutztqHJf+TsAJwdNb7wGNaAuO9KfIp/V+Y2j7
jxaAkPqaM4/DioX+n65GezN+uhqCWy420Q7Xq6dw5lNzo6rEQUJSynFKF6wCXMCKZL8xsf1VtPYd
p1X71CUWMFHT8JbeWE/1krv4o/ACR7N2RY7ZqB0Ircmzv11p43frUy0S3vuZ67WStCvTwrRfB8hy
OOYKwmWZz1dd83bn+Rv0LjeJ6kmINk2yHgH7Yh92xL8tIIWqWVLmNC59dPBvyeb7Etnbdp3Y1Rug
81SJcGsvlC09/5PiLSgSiSGOaTIj+51wf2tZfsrELW0sMJDBlB4wM/56/RDF3U/uaiylcK4sN1FR
RVgJq/e/NJ7dU58jlcELhY80yOTLQUBV9qaYxJiO6v44J1q/0hmLKKTn6hGZzhwZeLgMdA/mIRR9
UCQsp6YmuMjIzbGRVDLOkdpIlMuUDGNx2PBxePtsKXuvCYewyhCPgS0udbZ4pUg+jkYvlj82hVOB
nvxBX1Rw9K+mKNnckApO7CznfPqqwFevTpvE+xfmGh4UW2CMsddvqu7F6BUMxcysamGcK8rf18LG
TBltjM79PzpSRY98EvO0y/FVBGXPedsmr0lrnX46woI3i1ZH1cDiU89VAt8PF5HdPhpQrUOL2V8a
UiRxM12LHwq+z3lGpVFpn5GZOvGZuZL8CVC1B76DvsXOsiy+ovMPQH/AXaJOaPIT8w3E5U75OYf+
I5EcWh5TqAESdmirxa/KTkj9cw0OF3aVH1x4fKRIfdRfx82+cJYlYrPYuPcun9BCyEbl63CTL30Q
5MCcX1LKJ+difoz48zeKWDmgI2M8/7Mw8d8CJRjkY0UKiQsCoNc5a+FfABItz2XE+T/BWK//PjVb
jjlfHXp+EQfpBCfxZO790KLCMwnVPkCNjh2JrcFLRte9h+W6hGHm828VOsJ675VCohSgLgV09Di1
xgguqNAYfJcAmdzNSaRe8PjwsoQCrTSkRX1uzK2xweKx0OoAApMt/b3yaIzK0Hc6oO9epT6MCyXf
PJhanuwEcpprkvgq7vTG2MYL5XnQq9A/cAVBrymKlf3Cmm3gOqCmZOwDb+SI1zV0tiSY2UHXOsXn
AzBoU6ksOtzE3hV8IxVf3ItrhBTVH63CvPpmI9FRubU/CDhL9Srlaz75UIyAWQnt5c4FYIdyeKd+
VfveOfGTqM4E2JbHfLssYd9ajZpnVbcXh8P+43Ubl1JvCvrKIKVE6eTxO9JbqA5d4I4Dqj/OzpWM
JMbvr+zrQZzmtLmwwYabIQxfmio/39GzSHUnhhZsrCks/8f8fuNTNKQOCIXhxL5jFDGzV7Or/Dhi
sJtN4cgCcmzce1Y0lEkRDgwwT0nuUEUeZE6OUz2l43+AX+z3NHVQqrZ90N8cx7yzDUXPbKy0TvIk
JwJgA1ZWmuMdy0D9IUTWG5Kx2iTxrIWbQ2/HoNeBaUxQY1aFERLeTiFB+AeVv49COUPSnJZ80PE2
uRDjzFnNo2MjJ0bJPNriPgvtn+16nSFO7LGm0LkFD94cZPaEntcNmwI1laruiotcfQy3Aeh0ylnJ
zc15Iw/JTax+ahCOQik1KK22Eirzff2ZfE/PsmGl404MbiU/BDX84NHO04/kij2Ht5nKMK4dxnfj
7Nfx4uMUXGv3HzyCjnZLxjITM0RPLhDekH1L5tVSmql8bLywG60RbaILzaJ55ihhOXR1Nf7I7WiU
2FqbuVDBFWbSpsS9WN5Eb02rFTIxLbIIPMYxbmP1IESFqNa/Ap15K7I1164qtpkSmdFbRbFuaEw+
3NRTKL0nUwSRJlRD8Fhto/91M5fCY1lAG/e94NCx408qu5rHa1NrRmv4cuBP2aBfL3c1ho0/YSLC
mvODtUkFNjEy1qyQsGE3hs21eXOFyqiXv393w2LqX1wRO8jnQya+MDUNnIcwwbH11UgyJw+Nojyn
7aVnRyFmXroUvSM3dtUX2wUy4bn5z9/ds96DrRXNVMzprNVHNCvZYv4nsB/xmrX2wfF7EbE7UQSZ
koe1BpkiTjLwqMy+OlOBw+R7szT/76Eq4V4GyljfiLjZrY/5ooNChlQFQNLffuBhkKlIR0ARzGnV
/ZyBoEQ5O0V0LEurefKEqSGR5d4BPlBk9iquxZOh5vDpEl8gn09/SH7ks0/52+uQGDOWDbDhrh3Q
ga88LvuAjcJ4FEK46uhn79LhbjSO6s9ktonzBd/CHAPRPTT20u0FhNrjLmM44xMOuYwL7YDkwK0H
rwA7eDNbOHda7iy7r/bmo8lV9ruT9IJI0YxCiwWbnqQxrP1lJIVgIJGxQ077sMYmNgsuH8TXCr+y
5yH53HEFk2d/8Oowk8MTbPMxMp6NTyh0ewB3pEPb0Ftrxo7V1EbnXn0OwhzEsnq9aJ+xBefTD6sZ
6He9lBcCock2YAhuO4+CIixzv8InOdxlnZKWXEj/MNEQERf6O3EK8yaKosJifH60Gj5MG/JZ0XET
5LorykcL/cWzhQP1FL48Wk21NsbdmzxMzpteqRatLXr46VjulfFeMp0lzAl9Io/Z47EK4JNzxyhc
KNC7E9f8X/lHR4dlM3tpB8YsffcT5+p51piSmVpI2EsL2fDgxYS9bEfGD4fVsBadnp8SfifE0bVV
9qtpzGNVLEpWTAfEHISG00wB4juGM+i1upv4wPejr9XYYTMbP+DdaHsnyqz55dYth50OQ6IcMyOH
GmTuaG/m3WujjXODoJSikC+eU7JqGIBJ74tJuDBig+ih1J9R7fOy6OV/yfvBrr+VKV1SDeGj8JDJ
HT/IwGiCPuQbMp4AcKGLlvskdy0GYV3wiBHau7NSJDkaTqBKU19uIa8ugdy1H4lSBrUazrbyj5Aa
pGmW3fNmi6ldk9uNcDrKzZfu7AE/hcGZjo22okAGRs0v67N/XGTMmokNbg+yRyBbxbf2ZfBNzF/5
IE/h+fX/I/foQ+lX5vmdoV0KC1GyTc4bXjXXa0QSs6h2grJ9cUVByk5QT6W0USP957iWdAJeTJ/t
fVobJyMkgsr4bej80s5ZJ9CA37VCNpKVTYljaA3kt9GyXml3ZY1Fuw24qBFoUHgjKFvP1on1Ff1+
v7yJTFktosTz6qaxtqx2G84JG0jzSyISCGulUQujRKQTwKuHlVDBrrU8l1+3tBYFmNP7oIaHIukx
b0/DklgmsJCyl6n1uNPZRD76l19fKIKY1VSwkwx525CzxSGfKzi009ncJvdDyrFQCMRzq8zp5KyY
OLYyLngDgRxHzQIIkkulERRauliTG+hLyyMkOWNhMbnY58kspSPsXQT6Li7t1qRCTVwo2HcFWOV/
ZR7/kY4e1MPkC7HTKLxgPncdZP2wbbgLmg8epgCHQKITyi4Ao4e/6Suhs4fAvZu1/Ub9qlGwDYK5
qfuyQa/y0o+JjMRFqgnwBmB6uh8C4FYHqDnTRipY2fvHtIheS0j4T2fFRq3B0GZtnGdX0g6AOJjx
fQy2cRuOKc4vqdqTwbEtog5yQvQAQm3WT59NtrjIRaYGFPMmZVOQBQ1usTJpbvL4wgqt8B5OwfHn
wQUYRCysxcukZo4Ru/1KlynqAqs0v0Coi5VWbH0WT2v2BbiKqV6jtNf5D7qg1yfxaNx3qrKTNGxg
RHtup7gWkHrCW5t9by3bTyzi67MZp8E0+sCA+m4Ay9FUNnfFnLbEGqHUIMfiwg1XNE76TcB4Demv
9LlhVsnlU05KabxqnfLih8eyduQKeXgeFRfjYodf9NPAWtjTBI345n+EKWbO9kWhrb8DjvjRy/IH
dQ9oHTqMm1oM3KnQy9JHPY6FPcHh8e2ai+BDZ7xFmwX/97pmndWPJaYQrzGzw1RyIm9449mAVCXN
5wU5Wpdcelg2Fa/lOPeL2ivxGtly8XwqtMLXDogaDZHb6tyRg+rOiLtuheppzeyqLxD95HZhxc3u
VUHomnu32KIyRW9d8ICTPmRHVXnUMGR4pcCec+n7n+r7gpw4Y1m7DDk9Zcw4nygxtr57lE3HStpt
LhwtIbLVh9Db/U1xuhDgPEl4TRER4zwRyi4+5jzcB1DSezq6EURbReZSWqgf/kRkvUajXc+nyTdp
qAxQn0sJCRjDBldNv2NzRETjfiEVyU11si9+jc3lAkMBoMnqd0b3KACxiIk2B790+umb3YDWi2Np
GxFX+oT3hHKnOM+rmyM68S62DbsPRzNB+UzUvH2+79LatjnWtmfrkgnTLF4ZqUoWlOEFkvr3quN8
BsbFfLBI9RxNW6ptQ8eZmkMAF/z//JeLD2AxW61CR4P7KOk/Bs3WfXIMeUAw/zpfYCjwzNxHzOED
yNOfSj+uon3+wY+xUPtRUqt8wliWLYg5QmRkJZRc9dgzJmUCP6lUyS+oiB44XUgtALelTbOkt0KT
027d0XSm1D9HnyYGilELPoP6YFu8q5jP1pG/8Qt/gDc3noKANiXeQCeRUOUSg3U6i0lrbIsP7/5p
KaSyEbbgTmlPLB3EkUHFERn50Vus/wwxaSS5Q51W91ZRO2WHUv0atdE+jMT9f4uR5O7xKCghgaqZ
vL+/wGxnWSv9EscKmJ5Xd8M74DUtb16mZ26gnSgjggDDXINPEQ+NpHP1Y7+fnnxwKBjKUcN/VEbf
DuRPIT+0yhx+Ho5TG1TTfee0WE+LaqHEAPPVwwwYC3lylslFtD2G4+b6PA33oRAI8X1HwGluvg9h
fm5NcMHmatJNHGupqJ5e8OxkEScQrCbA2MViUH7vBGElUIBLSWaADGb9JIdloejYPVlEBkXV2kNM
cmtgyqxuUzi8thm3kdMV5B4H5+LgsERpwrcVI+2jyDMQfrTF1fgoIAJhOT9pKOoEHxQ0adosOMrr
EyC1rl9X0DFCb+z1iR5+5JBLFM80lFxodl7GG77Eu9TQwcNlkdQaQu3mDjkWCvkzz4mznf6jRTpL
7ugYjhvEbcUSs/3a+QgMUEjtc1rgy4Qpth/IBDuWqW3ig2HyaQPqGAjLIAXb+wodoK69f2z5FRRE
dwyJqg/mgp3HlQBm2JNMo4v0pM3SPF7WmVnlLeBTDlFTkMJAqS5LUB3DgcTQvPOxT/QLu9Hb3Ar7
DpZNHEn5bcp1EfvW9IPt4wIJVvPdnVZ22PngrQcrNjaf2E54UCM8cMhrsg5CQLGsAGEJdp6wOShJ
za5Lw9xZS/0wxMo2FO1ZtE+yC3mjt7B3c23EYAiWls8efHRDmSoVOCkGEyL+4a4/StVwyNFVS9v1
43gzeg+h0hAyv21HaRmC6v4wlj6FQ0ZM1Gvai0fr4IgR30HiYZjhY+2s3DFaMZ5d0piBal4km7so
YjIvwwSbQ4bsc4q3j7xTMs5SUmlpPQCzL+YDKc5ehuul4NGU2fYPQ+tcy9i9Sxs7QLgiJIA2RIh+
7Ce0xnhPM4m6BIyj2yBUazhBTwbJavirp1mbY6Kp9rd0gzR5Dy1cRJoyiajE2jM2qqGJoFyJtv5i
GMus6GAzx7dAnEu5vXnygsL3N0sVJ06E+KOZQLlmJSO9JGn/rcE4SIhZCNyDgh2p3eZ8ZokssJEQ
eqtki9+SX4hAINl1y676CZHU1JT0b7osUXkrDxHJSM9HPYuj6EglNl4lNrQyItTafPEkwQF1IeDj
WvmchGaScFeltVaQU/zaTv08rg/4NV1ZfOuQcuixR+3l3RKIzcxc1yr7JocqmVDwnmA+vuBPXMgR
gQSq/aKAVLxBO3DO7ijS74Q2JWat1VC+CSaa8x4nv34yu7qT3oSbxUpm+2M8+3PNi/5IxaEhcVBm
idRajo810lVaSD0RztfVo+WZJVlCrGm30qwPlLvPDrdDN7Vi4tghsdt+V3S0X+ss9mzAMKMuyD7p
VrCkzXO1HFbGVEFQy2zyY8+Qtkgxrmfjd7u22YbmAHX+o3XRpLinctza2vE2RYmIuWz8IjeNpZj9
vNEdb9+SujVPpjO9wErTlpZpNVqMOtomfbqF0MVgRtMYlSjGadyERfz88K5nJXZP2HrTobJc8LF2
N75dJ+yMQBF0zFJskDJQs3pi5vOVijieZaNQ+ZCqV59oYcFhk9XfOu7PZRmQjoWA++F/HrMCsHIC
PzVMYV5Fq5Ky0XtKn00diwukbygZL40oZXGjv6iSwEKnj0yzq2IlIud5c6T6Frrgrh6k27GY57Zv
Bnei2o8psoj50+oy9gnULqyq72MQyVb+sIkIrQ7y6Siqeue+36WVHVyHHy21GkUumc/TTNBTQ/Aw
+1YgxK8sVFfdx9avNG6XpEcHKky20lQJ3uHcdc+2SCTIq5zuK69i8+Iu4MQFOFdRgVtluz+NjbKG
VAPa7AczCLEHXe7VtUVt1CF+ciRaBR4UiVmbZRPfRBINAlxbSvTDbSpFgV6ZiqosyjTJ5ScClH29
lRWEPy6ZaAV09p/7sOTHjOVU3/9DsS2/5jLcLbvadLT7XEnHBOmGnFVnqPJ5m9VzKIr6jjIjm373
XvBbBX1m4WqPemLs/UHbkzS5HPqTB5xA7vHSxWYDc9pP2zlb0FHD292kTcqCgX57E4dzRk3TYsne
kAkFUAspi4fP6gRjKiH1iMH3nSyt74Ccn9bY4bsp7UDBKeHT4GjgqQosfHId0/ZNe9MNqh51dhlU
s8FL593JfRtEqykR+FIOwb78p6jqyea2eLTQmfsxPetu87MqspzogjG/3Nvf+HQN4Atm/Bl7zIJh
KvQSlVp3+rdJPDLS/wlfCbVljMWLsSpHKTS04cS4uL+glmpEeO5vrUMow8JyXNCULNEYNTnZHP+o
gTc3uzJXEu7G66ardpxp2gBKxMg5bz8zQS7zJ1+Z7+eZCpFkPslEm9z547ztz9vIfaU7uPzYH1Rr
CTY/vYj39MnsfVV9qdSoCC34UKyNxpzEbmcIOZjHmWptIUoPpcSXgTyIL6tQxOmkty9F6ZYmRRci
Fo6Y+e/5ZsvAMlalNxm2nwoQmwe6a8rzZzm2DgGqV4eaO/aYqmyH3c+Dz0WsneZ53s3Zk8OIgOQy
oWYJ6wridclhjDPdSSdtt5aOjzbMOHF3TQ3a6nuyk7Rj4O3EDcI0mo5xqjCtYTAM7KdWLomwxuHZ
7p2hjiB4f6O/yfo96ky2X5GosRmEVhgGoi8hiE/paTwplAMAe/wQyUZUJaLUBDj9Iv+1wJQQ3RLS
Zwy1My9ZhKf65BCfNCKzuweSfJu6ntB1XDyZmbleNbnCCvNYN9BdsCbXfPyA2di24dcFWAhzoQWK
KuowDEC0YffsYOe75sCy+NKo5l7c+8dS3DSZkkAnwwW3J9alfVRSdBhzNYMjrm9HmDNURwuayGWX
foeuuJ5Tk4kDDOy1KmNcE90Inx6UBIIE/Gvf/UbZGXcGhvpa7i/Tr/hSlNNfZHeLwpxVsdXLAA6S
NB4vj4SQltm577ouVjAZcaBGxP0w6ul2HTnhS13ro8qHpTU7lKMg+bYDyIaqh3n6UjGFsXMug7fh
oZm9acj2GDIhqU7ig/ZoVdIxfPhcTXBAYNoQRnYe9fmRUD1AqKKEXL+W5uO4AM090ee/G6AQHDz+
/d30bhg3tgxq2v9Cvdl7VM5aUeqzsXddUEsoPPVtso9Ba5EYpS0Bi+xe+3nC5St9pRHn+0xJoe+U
9lzMqOQG0LgN4twlDAkUBKZNiKkCD32v5RTEyb5DKjnUj/hMlwgjCJyaBbVFMaELJq9RYOqkdHH8
Ian8SapS9t2pSk8cnFJkzaC4IOzSuPbxzdN3woRZonhwFCPseDDmZiqishrV4QLwYWfYppbbtWeN
GgzAGbaRPGa3DWI77hBghje7ddEx3RNgYQsZXemp7JyzrTQO07kKZwwrOHnVJ0P1tYu9F9eX8FbJ
E9e+2vYdSjgRGbUv3ixI6pJYhZl4UJkF4W5yCL2Dn9+KwQLRmA1P1z59CvbiSDHEfOgQ8x850DOs
DnO4OT6ZcMg5IiyUx7csZw50JcCoPze2s73x4LC0jwv6YuRClo40M+ov9QyoMvrPepeMdVWdiQ+W
n7H+d1RD0CM0P7gCCI7HSnP5oK9Uf70rDLQTVLB6QaRQMf20TX5BGIBwMrI6P283NBNtMNZ9Yo3p
1GFrv6rvrh4jcqfYy/haFgqFIEj6Gif0azQ0Po/FX9116S57M4VkAj8kljAehHUvkLUG/z7beg1T
vLurBdpp9SH3SRu4HpucLCagF+qRe0LU8vK7Qg++GhU5j4QFrI5A7OqGKhVmBC/ABvvHClJP9SWi
klkw3jIQCO4QMwnOn5vUzLMB8LMtGcug/AZjP80uEP9vf373+34aXAD3vGNPeDEMBVMU/RQvu1Xj
cdbMn2eyTrEQPNVd79BBtsa+lO4k0yT0sKxb1pxmm39qM+ph3mYZynfPA/roRVbpqe3bW2jq2yQS
Ug2C54B6Sl81lWbhIbTTM5sVEhDSIqZZt53vczQZE3xH8gfBR5woLJm34nt8Q/QRmHMvFCP+TRSX
kjpUnnfgQBWYBCKsUbWa3fPWLJOZYJgXJJ1SWZnizwCSh+FKGntP2zn0yD3i7X9lDwFHrh/8rP2U
VvD5hJYRUwQr6G6hqhCOxg++6ndXy7+jIhTTwX8isrlz0YjgI93vgnEiPVSVH4p1zSn0GgJjM2x6
q00w2JiQ+zMfffKjegQMP8pIyMKIQE1+y7jhAXI0v+AdwsfSDI2PHjEDJvvqTRbBfdRAQSMEKJen
o5LzCOSTRlOtWE/LS1Bz1zva6awTzQWMqrO6d+it45wVPJptamS2WPERDGnq1mW7GpryzVbE2l/i
xN5Vs9AzF93AWSo3L1jF7vTAngdDqrp8BAk7XsQbMPaUz9AplGWUIBNHer29wYWJVy5oTjjI7nL2
ocxsxoz/n85/CXaWvspuIp1ZetMMHT7HGrp4cK0l+451e01/Gvv/usZbw+EO+h3XbA60dwxk9fVB
TQ8Ty7sNQhTqoFW73UfBM7iCV04s8SakSDhan8hbT9ZffpQ+pwA577+pqDkPp+TVIvynOd/tvPHU
qOYMOXgxPh30JazPecreN8qx7dTuefQAxMLGcFn+g+vh7yPSlkcTSoCPYssJ09LsaVDDcle33Wyj
lo58GmrSvT5Qbz+xQgZ/ciPyY/nnczMH26rJk99mMvjH1C25kibW42uE7DKHHcIVwP/gqu0MQxCh
1BCnGqpGNS6L1VMNDG69BHG4sF5P4gCtbQRdI5oozDqQQQSzZ5bu8pSrO5Aql+Q7JUiMwK/tHja2
i0PhqfIt2b4JwUs6gCsavhsxn9mTG/t7X8/emyf6BtmpupUOU3YbTRbfJ0sWi+YaVzViswAsjIRb
/UgNkdUpVQAz09f7UIbmppl8VwXD9GkCDpahYyq6YZ19XVwCFBJs+NpYMTtJ5C0NdWLqNfx2n9ke
oTqNvtk5zoJWwy+iRU41VenKjv5QkLac17sOdw0YnyIgY67QHIfqJePGPJCWG5yCsJ/DKHxaAP7p
wO4Ah7vzV3tYwksdbtbt3jgg0qGheLaKhMEB7m209ejicEVBv6hWYNh7Gu0GwN8NhIziYlIrAQSM
5MzRAF74wIGJiR4VaN1G5lhrcf8qJYDWP7LQyml7Y914ImQZSRr8fI9KN10JXUSp+GqA9TTLcmhe
8KieNY34U0Lz4aAKiGKY/liqF3KtG0S9+2TKD9dBSZaQAeyEp60gYqRKibM351Xo4nkuT563Tfb8
LMeldZ7xzaxnUkfXhdl77ajl63RarStsiMSsE6ga5uPJXbrffu3o6FJ5bM79SUeYNfXgmpdqbXQK
H18Rsxx29EKi90WhTdiFb/5UhpJb4rTXiS6Cq1xseWoTO1hy/zoKdvNghvydGjs+R018FEqfPuYC
3RQa4NadT7dSemHM4BKLQ2995HILo5Zd5eBeoUbxvlY8IaV2OqLoA6LXQNwwrMd3pVqDPH6bbdIn
D659um9Fw7pm4e5YqMddt8dQlO4XjTTkMS5lj2gKl4fRQnSM0fWj7c7gFHlfjMKGD6XpTjP89Sgw
NJz6OmjJvBjdJF3XasGJMgCyrW9vkNRgtdqlglBQcK9vlNfwpIpQbn8htvZxHrYQ89I/i61EV62V
4pm+NWV3ng6FP2cBS5wBFzj4xGiELonCQM3ww5kQvoiWbrPuVJvd4GHTtpxUWKSaHXfxFSKY++c4
FHGAEM4FRNPqEwY4KFzlakcQXWW4p7K1irmWYRz0RZaxJjT1VRj9jnuupFd5qQhvF6Le85+hl/nw
MQblqEl1pfQqCWE0hxYhl32dBIZbSBQ8a2caLILqc1CAkfRaWpCd7Fs0bZWUZhS7pSWaBIoIx6JF
Xf0w0qu4xdTuR1Q4XyrVIqYWYFFmnSLXI8eoaTV7Hzcg3CiFLIfsSPMMse449h3HQRfWB8LgupsQ
C7FRc8uCeyOlfB0R6OolvCO4dJAbdyOHwalqmKG2myfbTQ2CCb5VP5u0NlWcobsz1N28QD85gj7n
mFi5U1ihIrV65Ws/Y3kiIpiEfG4+Hr1HoBMyTBGTRkq1oXT3j7viwzlj2QDU+x4R5yz475b/3MGO
Hk/IlVg5TSJ0PkILf5+mCDCwOL9vsg1wfUGNZNhYcmq6A4K6acjGYv/usVFDY/INvrF5I+F4Vl9t
+vfRFPTdP50puFmlNm4DwVBm+GtzFaRGmZHV/1mZAnrTehlaWoulIV9jtvkqp6/cpc/usGeRsCD+
69MLYwIPTrUq/gg0CLcz7nifc+sUj+NeRp7nNN0C8q9M+9FVw1RRVzTXJKqnEPoPneFjsuWStH40
mWOlpIN24mU5tZC8IxPsbjiofsx+YXO1GVklGY52g2In3XaBlWpYLgDp0/mhwXD6vrybWNxTHcfx
3GE+fSyx/AgS0WzZg8+Q9nZssUrB1rXTfpQ2PnFzdwGACgdtLrdwErG+EpbxVJyY7VFmUkYYtF6o
gRH67hibxlb3LvxgXV5PmbzO5eToeS8psbGmiMUBdHJ5SEtSpdJ2khFd6WnhBREOy8ZKk/BrOq7A
4nT2tNrLIIl8dYZovxws+hKf9bT9IUBLJRXMDtySMnfPnQkHTrg2bYFTPRiiY+nh1gxNuoXP3Ij3
h7AMde3TBb9kL4zTRD+4KmHDE5/jmpTjQ/ArJ7kyjTvcn4knaibhHFeAoqgDNCX2bfitRPnpyQPg
F3sX9Xg6BLQKOjiQ29RpjSin+EALGYH2yi+FII2Xz+eGojBCF8Te4Jk/G7A3IM/+am2tzHTkcru2
MXzZEF303pZcMGx8umkyNF8IeiPbM5RM1xF3n5pj2jfZUbEv4TUg8xhRVYm3ppGrYCcZbL7wRwov
Zya6Y0vNPRsZPmBm0/4MZotph9DuqtDt225kLGr8GCAYTLfytcarLyY3D/H7DhdHHYZrxhlynerx
xWqirEPyDoubkPLzHB9l05MSW7s6+NczHP0tP/ayeRb9K4YXTXmPEaPjyhQrQTlBivmfPYJg9AXX
IvbBpXc8JAc0uFqMzMfooQOpLhZCDizYZCqssiAVRpcPY4nI7f+g+rDklglz/efFh5qmnkX+wVIL
giNGWcwBxoLcG/BbogWch6C9M+1YNsR6BiH3w2bJQX4JicqoukmjeMKfMx/08YSeOs4lNSPIC/sz
+MQH3b9FEFnza/i6m6oyfUWx/+d9q6ZTTL4dJ7RJuIeGuymR/RSqIFu0pi0LyFpBA5Q+2v1+MseX
RGj3Wf2O6R2DRL6ZO0OEITwmyTKPBzya56Kx4o1g5YkBLzr/oTqbk+0771Oo52oBMd7F2vH88yFY
19bkRC1ccL6a/VwP7WcIOgTv7jdehxabfAid4E33gbfZ5/I93lAQe6a/fPt12pSYHrA+KSze3PIR
TbkGpaw7Cu7lLUdGKZYbCa7gML33VgMN1HvsFJRC+q5UfX1p7Cg+dGiuDCpggce1wMtb7vK4vjxH
ztWfWP1+9Vc9v1cmIhdWqCKRihuUluHy4QIYzNUlf0kmSKNLuHlp8ZFFNvoHpeqjcmPflL9cRmH2
911W3GuBTsfdyhx5AfykjRTENemhvfJqZghtndJ7xY9p23EDnNO5TK+HwaePdkiT/1mKj9pf6Gst
pvxwfvLpIfcEixZYdYxxnHOr+g4RTHIUNUlWzLV13qy7PWKugx1ua+0N2Pf3/0o5IcdweOajk0KW
tzaKR56ttCYJEx7eI3p4zAgLAZXofAfBcmyIlmZuRA2ePa2CVQB7Po3ggn6cprraN/RBZ7Kj3hOW
BR2TEh8/nvqsyloCAPHCO+fECWRxoKsmHEuHm8ybFcjobw03Klut/T1PYhd3h9k8A3QpXIickNK/
t9G8aOpSAhtJrOXcYsSBxACFTlvtHKrQcqDjbsfR2Ud0cr0qSlgmjtAbF68jqoyvSGikoHfBhqEK
/TWPObJ9itBA4IT2E1HEkvOsIPz0557GJ9fYayqOWCE7B+GRLMrsPUWW4r6GXjpOeySqRaxB9HZv
eslCu0ZdeKbt4/Vap36+p43iAws/6mBPqcZeHTuFS+ICwrZfx7CLndj/zqkCsZ2ei/xaCVz0Ymqq
iXo4SnyoFDe5aiPZwEBbXbS8CAsqabCGm9ZAvTgHkwiz4Ks3FtG4wWii5H163uxtM3413e679KL0
lwXiDbKGgoNr0R/j0syz0D242L9T3OJkDUSmbBlHomCNIg41TDB+RlkGWah1NsxsIEW6OWVLLKAH
UmrM4wjD5zwTgn7adT79qE1TaHMqIKBIPLknxh6FKSvXkFHYcuEz7+mLmYctpv2lEgsZRfBNpjvG
kPcZr0GM0Y2w3ohzDfdRE/7YVTBiruMHa+IPY91PAdyE+Dn0vnnBqInTkg6g0jdiVHU+SpGF7li8
szu1NYIEcapVTCrUT+jQQyieqHRYUM+v+RRHPHB/QobquVD/jj7gD51kfHi+l5cvjuvsWqjAJfc6
uNZT1Ar5vt6ewKpvvI+16n1EjqkdcUMnE/xbl/ZEwgGcB1++gLnk0Z+YUgPqcGy4us5IHx7AAxzq
HsTAoCSDEa4Q5JhL0znKlWmz50LpEeiEHa0ihM/ftyCceNcBbMMI1JI2ro10nKvfYAE/7Cc75/of
goeUO3U707HV38DU6R+B3gu+/2AfhXZNvW5axA1s28mUQgc4/FBlxGNwfSupng/r05YCTOZpesw6
Li8ANIjSF2OBvqfZhATcwdQhfOsI3eW7OJD6Gyd+pAxj1o37gwr2XnopYzHCDO2WEPttbJCd2D9r
68TsbjyAu6keznY4q8ar2zdhjW1hRZP6ipF/6K2NJ3Uj3IC77zAt77MArcvawrB6nH8nPk0vwfi0
jOVNRmLLkiyR2WA4kFb932jJy6ACi17i08FfHvE4skNzJBtdWsnAas4N3G5vO9VgJ6dfqSjm5qaP
2K0b5go7Y1rX6px6aF0faaj2KPDpeWuQ6BIGSjggPHj10skCJfSGA2lIcbwBoWwwJfI0CNhF03T1
gkQGCX54WE3Swe9xBqo0j3l6+14zpZOYwHb25Y5990lpjGd72QRx6FrkkEQucx1EvS9JgTrDqg2a
ZNbBNfT1mkx1Mxk5CBSRyFeHvLUNdZSVIeJC1aQell48AxQGoyBW2RsF/HAfCGPgRE4yzMR/85M1
lTrxW2DixrC/JYFNzp1PBcsAQpUaT2iS92Af+n5myQUUW2ycSzqtQn0N/AKVQmJhzQcNHlR7ZjvJ
xBTM2lokHvYtPHN9KNsbVf+rIS/8Qx62ts5O8RbiTYbos4A0STX2X0Fq9//gRMLeFoP8WAzJUfW5
FaQtEU/gNUvBPYoPkrwgCVOgvb+kqR8bnhU86LxGCuxn7SAQgLal5bmLpu0hpgDHma2TZzcQ6gIV
j1An4djNZLseVEfpVFlLzxin0ePqv3+6RC/j3OMo/ZnV6z+HbmLEQ7WiJAncVQ4jBKrt+TgXBWqb
FMm3t1O2ZxIn4UPdrJlxj/KIT47NjjdocSkPIH7iQ5h+JC6nBd16j8LzhRaIz0vbYqA3QFIQEaL+
LV1qgW15/c6hFuydmgpB3PC9LS8Ea0r5L1seJ6uZ23JKebWjFFMc6k3kWwqjdSzkp5FrILlOI+CP
W7pH9JASebq+RCpiRJlqX2LtTa2hnZ3AGdmql42nVKTPf4MejuvSpDVSe6fc5jpw3reHX/K7B4UE
47QFSmHehZ6PXVnu6MgJ1BOj1bv7rRMiXXOKy6w/WnHArmmKqsWCWSvnGpmYrYw1VIkp7usCe3cW
hJXEOMn0xJOeF2H+4sHVIj8Iu7XXv7mA8XcpjZO3470QPS2Lm1uBS9OkhyGqKuxhoIW0yj2NaaDb
bS9qtK2VRxJYMONuRdwoPxFEOQ3IQWkJEm000dNW2jI7OG5VOBbqAqFwIuAOQSKAWsB4kutwx8JH
tPE6x57ymslY2QxO81l7o6qJhJDNVkxtkiA+Ea5OeMveNMJiVztnQ1DCxROIvQjQu5HTsjBNQwH4
7bwOCEaQQWd7zwi497nrXGEYCN0DTJH6sW+PiLD1fxRJMx1kjbDg/xxzd7UcmoNTOMUxpYZ+FvHk
1CpPKp+GHt3dGcmADw+rMM4AMqcGvoeSz9MCFsdrsIX5EnQEy7sXE3J0TDJxOgtyrKL8zXy+wPXh
kUNwp/5A4AVdBij+bE68gct1pIUFZaXuPj5McknXIQjmNSQIQZHTPmkpPwL2OOcgQ/Oa1pnRWxiR
Dkd/CawpHn9wfBH/r/5XVpMIXBUcleay47O2SGf9m6lJcEnCdWFjR06Hv2hpwmXHJrEqo+QMYDWM
fQPeNFd6czwkQXDCCH/qFp7f3TOQgQ+QmFYB9b+fGvRRvTVtgh0LQbiROig/saHpKUdUi8JG80Pg
Ff0IkgDPXpZL0JW67MdLY4IB+qVqxiyaeXe9PpjhD9zKLGkvzvlSy/rDFDrz1tDfW1V06VHqDr4/
2kZx+Yt3EgLReC8YJQ7l5CmbrnASy9E0laStLrIFF1T9STApQIZt4gPRCSILfWTBFJ9NKbmCeU0E
3LBOFxwzqma9cuufL31QM8mQ5/KAXyq9XhQGfDF/yGc8+ISfO09AabqmpSk2T6YmZBQHXhgUyx94
KoxSAPvT0nujkvhpP6L99eqjToYEoDXR+l30//jyaOOgxGAh+TU/QNjHyxOd/0eRup1t2DS4BRIR
bVhMiulGh80p5Jb+WqPqtdC36QS4LGWUOBZFHdqEL4KStMbblG0CyP+rfGEn31Zh1hywxz1N9A1r
9nmIocx3kJBZRNnmMSxw/hS50RqQEGv8zwCGa1yRuf6w72/OZBUHevUy/agteK2ivyCGxubYD9U0
lJZNaP5UAFwoWU1hz8tVDwW+t5n2GIbEPv6HA+zdq61gQWzGf6t2oSumbxhL0vFqFLhprISfw1vS
OLisGR+M/1YXl1npFGpekZ5GZEt2VwDAF0/tPiV44hqBxmzUngjlMRIsdO7LQpxJ/egY7CakSLEx
HS0mHmn+mshp3DAbubsTEGoZndL0PUxLqBIrMDmB8WNOFFamV7QkLX+Rlr0m4b83oj8HpHrZcBDV
5u98dBDZZcF0StPbP1liZRy+3fmREbMvUjeFAkSLA3iwsyLrRvQszKWQJQz3kPPH6bhSUVIyUdqF
FPY0yL6ZU3dLckUfMlMWVciAJU9pnEkrEX5AR5XztCb8TbBxjwBYFskfz6c41s0QLzHcc+pKinXJ
Df7Te/uQoMwjOt6HtiS9WM4NWwu+CWJovOBijaARpZAmIqgg84/nzUP+BMbbHYHMwoCem3k4WEFO
wAeQ1cEVuc2kaxHnSgRlBft30KDOEmr9d7s5hV8paEL/IBewplGJjN1bK3N/nsJt2JO0v0ZcIykz
vp6ls5qbaYZBelxNaOqmV3ORlI7dQWOXoBR8eoqa3Tcj8camVsqa7IhC/p0oyhDMXIv3sUCqX7be
2cjxlFe8jTWsmxV5eCDbssDDj6lCD3aQH0/URCnTOixswkQUQZZ5rH5YzBVS8r+szdNUfQZr3bwN
AmRPxTNk5Msi/mxymJela1wOeK7jzTaU29otwVkMl37TSYEoKbjpgn+USH7MYctEA0N48CBpTQjw
O/dLsb3hAd/pwSwlAp8X+PfdTlbFgfbbuRahGA+sygUSCWoX7FbhFQ7Pf5QzvKWEXv8ectHIzqHZ
E9yYts7V2xetCSlrgDb0XD2+WlJjSkGC5Qy76HM1O274X8w+nvawPpfXxGUT1hsBfqN+OUsg8CL4
ixEJzCO2lEJJ/1hz8A8GtyDv8lsrbFuUJqcJ0RQk8tZ7f0b07dsUtI6Wz7dCw+HTlvMlcxTBK5Cd
tXEVjPI9S+1Z1osxFl2OXVB18ThwXxI6y0d+ibGZYzcCoaSqgr9uZqvP9cMe1GE8vHpd8s/a2riP
7gHa5vt5eibT1EVyfAkIhiUd2uoHflSczasdSSsQMyTv71lsGflPLPHnN3TxyK7F0sAIjLaEw8o8
TFosxxLAC3FtyxxmwWzqcnitnU1MpjyJuv5kjOHZtDGaT2w2ONklUthjZVdQ8baB0PQ6+hcKmZG/
SGEqdeBjrvth+ZerOuIXkb6UDAQO26OL11Xi73b84LkJss4CTYj7GdyxxtYaJRxMAG9BmcfZVI9S
woauBba7mfkxXG6mZWqRYtxk+kl2Dn6UgSny5qnB4CeDksbiLyPnnXmEhta0m5WENoheZOKUiOAY
Y+YFG5XSFG1fxsIUf/TFW1g4BV4gHYcU4iiv5qanm3vsaVPq92FuCURP81PLcOBTONuao0WXzQSd
D4DO82Kzl2fbbC2HCNyubaYCugMXEL0mXSssPjXJjqGIljggLXMtINV7EkkFj6cJWJucbg9+rdPI
EF+j5Hw1fCfc9MM3DKSTXFni5F9Trmm+4oRVv+kn5G/f9ZFUfCQ7a8TsJFOYFj3lmg/53d+PFD1c
lMmP3Rwx81RVvfIH5QkrP85RmMm6O4Oe0Z9fhvtaJimUxfFdQPxNZohahWkFkZwhwoA0pzxeH4ck
gEO2nuQ+frb2vEj/M8Nl+5O8NyA9AOf8yG33BX2N3j98M90NzzSh1HSGLkDw3XPRSllbgEDIPTuX
JL8WPhC3oShL5ndPmbqWs2LSl3AXU/FUHNw1vcOOAtQbMY3C4DVyyHcLQa8BmKNh2PEV+sindJ+6
MwkOKnrZ1KWYv++T3Jp9NSziX2Ys5IECf57nSnFZqcDchJ297dnq8y/rnvSzgff/KusD4NQnZ5s3
hRWQ6ICZ0YRaLPSxS/rARInrLDfipBItpYeN2yWs8f8TC37BuzSQgR0Hqlf4EJp2M31GBXDHM14u
44wJEMU6Tr+sPPksm7/8bEyhTFNmMtt4PKGVrFNJ31Xm1dfrhXhrahYtTf861D6xtYuwtaNFHFEP
6oCIiv+vtA9CFsXsVen/VMMlIC5mENqJP+ds6V4HRlUpyXLKR0yVvzqpcrBBoHpDnJfc2xyzGe90
KjpfTUH1wHYmSygJM/bTO4of/rYr5Egi5b8Nl/lATXEf9tOZ3fX2JcfY/e2EqqwY0iIjn0bk5BW1
TRXE9wH9EmStd6RQ8wQeMmLYLQ8TWKtCkpiEdZXGA/dIMIu2msFK7MQrNhMWjhaR0mhUsTgB6b39
YY8Yn/SxksuKn1kvo/IhuNsebY3Xvhp58J00cljbn6ROiFzpd6RV8UTsvYhMzbOrxQ1CgtzzG8TD
fRPPQT3lgNJ1GCIn6n+NNcx0fo69he4OmrGG/qDXIZ6LkBx2mYgHAmGExhfbgsJkwrTH13A1Xhre
bCGsoqdQwYHywP1/S98ExVT4urgvTw/b8SYuvwkOXAWSjZjg2jDTBTOoG2s1umVu3BGsuy/u0pCI
AGN21ov7y/W09tYdiLy7JECJ9nQxL20Qe9b0wIhm3B8bkfJ6RP2kFQ0R2ftnM/QCw//RBylgsSNj
ApclxCvfxm59uHPrGHwb7w4rC4TXeja0Lik381B5i3Um7bpJ21itdo2IyhXtoyNexUYJpCiihecn
3XIAfG2qc0zNbZw8ekKmizdEXzG9PsOdCjWPkBdOq6Q62P0DM0ADLyR3dRnS5cZLMmmYlX/G4fP+
wGFqbQadfLNzfNlhHgW/edQQW9hpSNdLgXvCK1Y/TKkQvYcwqOIr70UE7gxUEGq4dSqftyXo7Ydv
Jd5QxDP269v/BqRwUbpT52qtubavcZ1Hfs5ioF7ikUN57WL1l466i3kmKVJFHpooiNyPtLOu0SOS
7sWklyOZZPMb0N66viXByEp/0wE4sXX3vBLmifUaBhTziIEn9broCK0pslXNE+UfQKy06tFQjKdl
g5IrnrTXoAZlllHaWqR/KAlzoPyy1gwUMZyJELFtaa5zv/cBlhzpSIKxHzB+ADsnE/yQ30YdztCT
Ed8wkMOdHMGnCL35729Bk8H/1aQtCkJopRXxe+fOO/EjzjjwhQorXtpyp8uohDWq8POJ0cO390PC
tVIn5BLIfNnmrtE72WT7skziFtUaNnqjEk7dJXp5eV8QgnvVEZDRQyad6lIAh3HYQF0cNl7yy2uc
Hp8K467X6RFoUV9K18Sjsp8Fa7ds01zti/69g/gUq6h7TVpeI8gL2B5OJaUTa0/a9WRPRwNcHS4T
b+OmxXPjO/riwsHCXpsnjg13XwpG9KdOEtZTmbrw9EtKK75demmvjmeT4dwE73B3n4pHfH09h9PV
i5RV/WNKxXJQuF8/X3ALfnuHLAkQ2OCy80kBW4FWgp9PM1ZxZlRY65PAMJOD4fxQ7IEgTqZkENgt
s++MxvjxxDBqkNKn7/l269aXClg4reNmf9p90XM5PtrkGE+Gj6aSriwEWqcwi2EsjtO8CQox6V9O
rc0ugaXJKMschoCPuwreLn+kWRGj6R7y0o/u0uFBquIVSEkahjeE3Z3ualLsRu6Z1p+uRDoXvOXI
F+8MznCoAcibyGHOiIEwCd4oOKsB6PMNaYvvZgTcr1GwzhDmCeEu8sFM87gL9m84Q+e20RwEbpLg
y4n/yAkB2XC0URnhfOYKkBO/SbA55Z9vyDxB8WwxL+t2//LTjMrejDt5vgErbqWHO2ek4ls939DV
OBcOM1yhVan1kViL4wZvFPJJJQlPeE+Rxla9U53gHE/e+EKrIHao1oicRO7WSxhrBvw+7qf6PZ3j
Oq1TetnKj2+a0HqEH3stbsnzUDRYjm6eObqjjasDIQr7c9V9mEWF22XrUHi5P2/luvCTaPNHyytD
UXMak7cLgJQynSBn8IfBfuWtyyNwIdm6N7us2B7eAWXiJfiHLsh55sZijIb4xF7m1tFWLyWKEtvf
9dKcq94h2XB+aq1hxd00V8G7TEU2HniAjE0Dh7uJI1rxh1GURFY/AIKcgtfLn3/aZTVXjQ8CfAUk
5tjUZEwUqsLNfG2MtAGN/Vn1OP/SIZd5floRlfMf3uBF4tjzwb/61R+bwNzHz29Ivll2E4A5hjZW
h+H9NtB9Ley/5q4iF3t5buA09inShfufad6SBe9aeHFXVuHVpS1xxANaEcxx0Ey7fvzdEQmZvAT6
CuOZHdouLmYwmJlQpbQzu3+sJC/hhWtse3/U/ZKVAtM5BIMJZPlCmzql9GzOXO9EU7rKYR1/MvlO
d32lYy1m59cL39VnBMwz2A3Rnkvlcz4kR0lOGJsMENdyGSrouwTqOaY+ME6O2gacWxLx857RI2ZL
/PzIVVwoJnC3EUe8A5dsBTKn9is05BD9VqEtQJWCsGBGYhRc7EAQycmQaG71ctvIG0id+khcEQE7
Yk8vpHZhoTx4Hr/szR4tp38ViCxAcxSy/Y7NCOzeUwGeXrW9m0wAN/ogjDJBOsWm8UJWgl5jkdlj
YDli5MC9l7mEtkLeKKkPfqKbOOHQ9uogmqv6kz4v+nQOiQXtYQD1YLqDgee1DJeqjVqtmDSdXBhq
MjCD5TtX9UVhPOaNWrp8JkAFwRkgiqsY1y4e1V5jen3FTeQP8CSSzpCALvLLgO05FFmgPwKxrUSh
onm/0l2J2CS2bVocq7o5ftWrGWvm50aqW8FmQQ8ivfwWtN9f+3gDqz7nMoGwicl93j2jZt7zNyNp
iRc9gv5t7L05fFftNPmdmZrQM61IXXj58rlGEuowzbhLYMT9ydysc1XYI61OIhdN/cbypsTXxGfr
NxDj3jgbP1LvCr4TXCwu21n1Pb/7Dg40pK5WdLs402LFrSfqHwHJhsx2ciMBZqOXLvDwsPaNMNIC
AnI7nczZ6OM6rsMDvnI3QV2w4cOptDYTuFP8yRHUFJRHeGqBOlG1ulQp8ThLFM4cs7OofGLTtbQh
FQVQtIjloOM3fQrz1CzqN6n+0FUTYAhTUEihKD47jqOzJYikzRpnva2xxhc2moYMfloQ2qbR9TEB
eHF9sVCdMaIZxKpp0IVFJLQpX5Go5aYYT/wnM4Bfo8SVp5PtqFPTeHpD4f2/Bhc+dDBfUfYJmKzC
nDOvyIi27UIMwDJPx/g88LxAkATqAt+amNeVfHa6TX/K0WsHdtB+XP7BF5syhNoD8cx/KukH+qb9
+8mlU9nrelCqURg75lqw5yf8CIkm5N32rjzw2Rk/U0oLTJsOrJf9uWOcoZnS/GaVL+RB2cN9unRT
DCHm8OZt3UOvfODdk+/jg2wSOtTTUdVxjspvQV2kKlfGQyCnxCzyr9s73g1VTWncWBPIsXihFXOa
mGiMDpUyRFIbmv/FgsNXTSn5/IphVJtK9J6CiuXUEUf+0Ut55VJJY3zjSoJPzUHv+i0aGItWWjiF
52aR0z2MX6AGsD+E6zh2brYE4MeX0qD2nL8CjKVvtQn1dxngKqpvHRrurv9p4D97iXeHfEL7pAiQ
ZhElyqAVtFafbrLxL1nV8rcz1HiDHm47B/KhM0Fo9DLQy5WfP4x5LKgJGlcBj26OPHLKmm8Wnabv
GlUPfu7ZSRJUo2o0EWqZAk+bvByo/JSjtN1JAnJ/7bl2h5nwnbXDd60TYAD7RblJiwxdk450vsAy
WThkh9LnzJ2EolK7Cf9Z3ryqNgcgv7z60teFyDILo+WhaRhNgN0QY6Ho+sTWjkmHzmAood1x4Iix
vD+CPtU73w7ez4Xrl0lyNwJ9c05TzQ3zGoixk7qchbRhyYo8Sz8bTOXq2be97CoArpbyAFWFeS3M
aL3Um4GLMYqKAK4Wo1/W/GO2SjdQCHFLNQMRw345KgCy0d4awXrOkRRm3XgcTPXGf/OGfXCviPLx
zIyqAOBeZ7NO2XYC5uKicNz7k2FdemwDBGhUu/TUF6nbNhNed8DdNNgLm3TIbqqWSxGD1aLijTun
fepIOXi9AZdTiTKLZRCW2/WUSkem3BuUFR54tpj0S9YgCtVlhbVljfC7YtUANUOfsGgmiXQq1cqL
b7r1o0qG4+ppoEOnokndwXIKopkmUACDIeGt1ptA9y/CtoLMkb2+X3gJyKxMy7BgJFi7InlvA/xI
iiDbwWcQ+E/XMKFyrADYTqiQx7NbhCZjYT5xX1dY1/V4s28pV1PHcUkZzbDPNXdC/+zat1BFdQSI
zf+sqM+A7eM8MqASR0fRuuIH6D7Odow1ptDU5hQKA5daIsZes432rrsnnrMes88kZWS9TMK4G6l4
s46YxJ2xRW6vEMWQS+ArzIrBbSW+y9xMMZeqo7Hsii+/X4Q4saSAweUTwcm3F8nR6X/ass4Ze6Ij
oUBllx4z1w9gyD/G3ynXyaDmQMK/d++CZENqvtUZuVvbhi71xif0MZV4B9jAixRle56fqte8Z6y2
EBTdLZ+BQQjIniZQG0Gg3U6QheB5LLPH+0gDpwP3G3jL8Dr+zfLP704fnpmbzy786mJDkxx4bnBP
nE7o5+MGyONve3vXrk+ejSn8krAk+gjneIT17On2mLvJQyTtjjN6NRbLcw6rL4MAY0ghs1LA+ggR
fyY+b+rfO8cAKdQxVxbJbEC4ZCWDFhTVVXKGCLkqAJddHBWKv4b6GoKnBmWtny6NLEMuCcGkK81E
hASzoaOXbsI9G9v0FR8Tqf1Ota3zZKx2BlL49miUROBfC/Ljs7jlR4OiaJgykVYhiPYtvZnQKgHK
99Wlo4WHWFiI+xbd/SyTEo5FJcUCr71G2wbezs3he/FRp+dAtPRroc2glX5csmffxT8BaCKp9R+y
7ebeO+/zLLNBxRs5Z4jppoRR0PzyMejAWLEYNjiVV9jDQA+HSDGcNoUNEXp0NG9evZXKE6zbHLRo
cfPkZkTBvWpFIAlKbdM1WzAJmgRBgFyc5JaXUetOdTonE7U2yvflV3RdOWC6aq+T8HK5RQgYdJDu
zFaEfRUZEy8rKfhPCG1IHgGKDy4aGOa+Ho3DC/MTknkNLvF/jIOLq17Sy/IU2m/Efh6SP9aUAIoU
fodERi8uA9BUpeB1StEk/909dakg01IS0r6sxyIdCHMOTNzcH4RnxUpkCa1LTTQdq313gqS23rXg
tjkOD0D8cCWEOJ29oHUNazHsJ0XcZSVa+8RLOznVKpjwJJbHxVf98wEiwi0LcCVxTRleV5Rjt2y9
G8hojNEtpPYHkN+RAWxftLNfcm39EofuED0c4x00otLE19WE5I0tCCGl7ockU93nlaKz+bAFaszT
cGy5yRwHhzOACJoJNW0VqBRKUBIPeKf11LVCvBIkQsoPOsdoJ62b2OdqsSgAtHx/6qRgVMIeGByX
Z0pK2kteyJZ2SalxHfKm2KjplXbfGAl5Wfz2uIWmS90ENarHF9k6YsS4gpkR6LWpuomsMIuHYzBN
Vzh/QNf59iVRdXgj4YOaPHUdbnCjpfXSNrDtmMDJAAP10UDsL++EsrN2ELRG64mloOyFJZ2d4hsS
IIdHnALKKpmiqR6i8ijy+inv7Dp/3lZ7/As+7eq09fA9SLwDLpjc1gjgy67JC6DJD3JD2A5VJACS
8kgkmAJunASMYIK2bIQG1bGS46bAzD8mmOFoMGrrZGLBrJizcILxzNHvN5BHvbwsQrgDIfPvxTB1
+FrtRqx1EFs2xNKfdrPH2oeKQ8Fz7eMe7mVDkU78SDUnR3oMoyExmNVJnuPlCBLJQnwevDCz+8/S
YCqIP2qoapAzMy6vEmAmd2Ox9MChOFjzjlcZqxhqacRQIcStoPYBR5Z04rjn9I5GFYy+6UcMKRNy
GxxwecI0f9I4V+IAh50uLK/YXxwoqKhSBSV3kDAE1jXnhTXjrpszuraNEKY7hWkkl6yktpnClAD1
8N8kx94jmFPQ2lmWUV05Im10LHIQERJiFehbDDK7/itfOVdPjNAf3lO+nQiUHIMbDEUKHt7Wn9qz
HWIlUVt8y45Ivw7rTfNoUfnWhFmLCFofq19n5HETP47Mw/LmjyQk8gSWlRhGAB+ef559tbqMew8P
oxSBgHzqJyUWEv9Uo6SUQ/lcj5GMV+xeW4x6p68MqXlS6vk6Fby9RA7pNS7X83AwWL7qwaqaiqPJ
x7/ci9i82LsbcZvdCBtwn0R5yMRnA4VaynvjkyK/9sN3rEQMx+nbujt7Hu04eI6KUhcBZmvTuLLL
Mn/Be4mHqxYx4IR+pNR6TjECqf0VDusLqYPWQmYioLNZHRVFDUAf78tUUBMzxy2ZhvEibxxWR5GW
5gFJCC0j8q6E56vJxyRs20heDlCcqxjBjgJTJyV4f7bkOXkGCM7rLXb6Pv8VohB0uE0s+dSBIiao
GW06IZ3aUquAuTX9AQWrv5WV1+VMqJxjMzTMsk8E4kSPZbBRSHsY9E8uZ4sXIBfcjRF//qshno/a
XKvq3tPEOPYOn+HoYdkjpF0RPiieQLIm/HJRegTUewwYmvLosHWr5i7PW+WvsLr22sJ8yuHCAW1N
5eYhsYnHQBKEtmBgAisfArjkCph5tV9OAd5qRujp7ZB72XYk6dcYo79nm8CqlD97LlrlBVvtSOjD
dY7TtvR5qQclw4eAtqoYvJ5yQM+4Bc5vc4nf31P2N218mRoLya6j3gTgN3nTH/42fstGe9G9lLSS
4jDtGP5YOvXWf7WlMjKpFp3IKrgVLQrwLdubCTGvYmLqvk/2N26RL8Cecq1bjLWw3HODw5DWIQvV
N1RaadVJ8qjeK5Ba0I69KxtB1uOJqcIPUrPUGSOnepzbxshi3LU4KZisXGpwn49TvlK2j60WwGmn
mIbuP2D9l16/4zXUa79zpOxxEHcNqT7mokPCkSDi2UYFh+ICEbwrTgU105hv8jj4pBWJ0efzMno6
q6+OYP+3LsDZBN5vbUGQxNcNkRRyxHd6ccHP0OP6txu3hfIBrsMutk5hz6uV5BbmdkMugOAlMOWJ
SFpBymn6f8+k4qHuj5El/YIiEy1wY8B7Xq+Yx9jnuySrQ+wUvCSh4DZum3CMgV0bq9T44nL+duEj
nCw53rU2oBxiCKaFAb3jKZcLJV3GcCnS1/sq/bX3831vGd01H5O5U6D/GdeFZ9HLccP6G0xPOMvZ
vg/SXtPBS7o0uURBWRm9QtLpJYuTROZTgkWVtKRkmDtzzNZbdp0yauFB6DPdBF72XIo20WaPibyg
6Nk/HaqoCz6zzCHenY7EBC1uoPQ3NtfDU7xApwAGl8JFJn2144N0+hq5gToHSjStNLc48bxvu6aZ
Y1bubONryILwudlhmgqKOpjANW9U9BJtgkWZxr509/j8egM/BgztHM9LU/71ouv2oaGDH77iAzz6
Bl4UzWfWo73eTMPkbBhry05RN513Mpg+XpqWqWYYd8tswnW/IIwImDBj1qMsnUulnNJoi12REzlq
z8DTfUhKQMUpKmxruQDiIdRdVkTYc/Cr5Kfra+SsfIYFBBNWjtqqD1hNTVm5L7wNsd1Gly9X1MJA
xtH5OBmEensFkCXiCP+Yw6+OJ8W9zjdX+5YPo/q3hm8IwyHEKXau8NiBFRnbkMnzjUhv+WWQ2M0i
yA3NQH/3xhz6trNb3pYxRsrApCjCKf1Mr4JuraEdeIB3TykvlSO6SDZTQSzovE8XM1+kvaz+g9PK
bgzD8Y/HCLpR8s3dNNZ4FUN6z966MYXysQnvCl97CeN/polMAYHg48RbwmyCtvMFPnl1RkpiRWyq
EYrkk1aR0tcOuO4N7gl6KkboxkUGwmgIETsK25nInLVj6wIrLb3UMtusTRzS6S9fwoWflPxE2Fy7
nBd/kzi9p2nGQJCwFVh5yShu8OqU3g9coOEo6ll55zbhfXdWhVEYuLGkT+ADQgISQ3mWEk2BtIOn
DEOLSektn4NajOZ1fpyPxI1EAhIRcJzkhf/RmUXMHOwP40UKoOZVbwByflU2LfxGZ5aSYnEFQbI9
5F65TdHJrLvGBW+Izq4zrgYxyDeNeuxcKmz4cLP7Q4mYGJaFFa9Jam642AEeAkXWvOIdxYiUvtW6
PNlPO4g8c2s+wjGFIxQmgPdrYC7q5CcQRY76QQpnn2OFKHKHaZs2y5mT9QWBvd0I4ccZYlZ423Bb
uiEUqEfLkwgv4z/j4yxKG5aqyl96OyhsF9CTvQbT2BVJCBnJ/Xl34RHBC5ms/q/jmZqGE/OiW62Z
6WEhU/YqOjtf/SRB7PnscvbknB8OcMITzFpTLWQsVDPzy0OySwbLKF+l//esKDB0qLcNVAlkaxb3
cYndkREHz/5yuHOmb4AbcNsMnmDFvTmq+X2cX7xl5f20xOrFasSb231Zjz5J/8GWG67/D3OrabpO
SMj4jpm75TZldmfEjglkNN2mdabgWa4o5EhWqj9UfmIoUwNNkmoMa7WnJnQYrzo1R+zxaqSTa6FT
gu9/Cx3ogpsh+j1FyT838wS/PrRTzL+/TDd+P7s9YdB+z6Hmsfk0UD6mjei1k8bQpdKCbw4beEFi
H8bgVEC93MG5blO0wIPZzt/jpIueb80K0HhV/84/x8HqhCMgX788lLHs0hBAW0dvtkvm8prugbTA
Aw8+lKhnTfbilPd+O+xbXBZieKRijkQ70qQnhQuSyCRoDqrTtsAQHfuSPSAVqFH0NSZsNInLRSqH
vCIADXM9G+Q3oly3ojfwttCnRx/o6BTW1cDTgmR0NoiHnHd7RAXd7PQrdChrxWSmJxeV+c1RZ6kF
X5/kebkxyXV2RyhS2yuUtR3ubWTo07qR4PsZfY9/I9mdG+lpNsJJXm32blBq5I6Hr8Ka2BDPvkPX
jTAz8y8cc4t8fMds51+u7npR0g61BaY7pc1MUxKkBfFoVtkr7SG4xRXp3/xi4+eg0Mb+C98pJyt9
GHSeJ6ajl5bx22RY2KOkkFSKmICvV+6MJwQ8fGfXvfwEKaywzeXhYa/+uL+T1tevluMfl4+WeQ+K
lN47dZ+TDP+p+vooyw+GsuRprsetxNQHbeI4hVjLeWcGQKEtuTjx76SoRn0AS6EabS0dKl5d/DPk
qRW1166AMIr51H+4of+4eKMaTl1gwDQHtopcndtxLe7rVTuQhf8H8FsVzDP6bSVTCVCF0qJr+6Ju
NG3Pne27tDlKNvAub/QdMfJmnCFyqU22RpRiE44XiX8aUSZRLhoIiMjNE0vHbTE5TcY3pWt8w/tu
Bv9yTga35CoBS4Nzc4yMfOFtFOFd+QcWqSUa8I/nmCpUKXybZkfGHswaqL+IRbiY+Wdld/+gaNDb
bL799gpba38hWpV16B7LlX2yi6yKSnJAAHlvy5Oe8FiUieLxgb/LtXcUY3KEslslWB9FU7fvE6lx
7ILBV2XcLbTHZprmwnfnxeoxrx/szaWWDhc2AyFb+2FEx6CYrUMyq3lrhiLbgGj4T+DS6Oor8PDM
wRvW/DTdLFnnnk3VjZUi0esRRiQXyHNRRpOjCm50AuC/Syf8+w2exZvhJh6TTV9mBknGeG0ZFRtq
KhoOp/8cCvjrhsKInV68tDDaaFrO+jX4ki/+rbhtqXwwREb8qXiCPqr6ZVGzIa1vol5h7Kg4K6GA
iYXLz1F+Gde7Rh2gICvs8izZ36xkgnDoCJE3YouLYKCzd+HdsIcaBEqVLFtwMXjZjkNx3Rbn7nMa
IJoY+YSr4GR1joft7gNjVmy2a0ZbCo186vlgn8xVEVSqE5eEQMJV0ovqtAoXgdtbaJmr7caPf/ZC
QL0d59iCQdnJLZEfjE3Rl82/WEFWDmm170NQrqGPP3+fVjkJrZMvl8UuRCaPwsRQTWuxp18k0S3d
gIsNA1PQXSPP4kbbpNZxEC9VDp5WAet4L5epCmIX9ghdC0FA4+NBtQq/qYzPJ7udciNqs9jGDD3q
8LNFygVP3w2oooa8/u1EnpEBlpqRYZGtlKTEmeqelQNgVDImi2gPILcV0S/7N4CHmpl74iI7WE91
/K/K7VfZvpgo3y1SoEjY/Lis7WIFkl/QEjj6WPMPL7ZPXNdicpH2Ki99d4C36RN3XCcWLok8fHsH
HtwulsQ4Rr7kpkj8E3Wbo6AzkiGDCrBb5G4SrOXQRdMThsyOrERKTVRjs7f/zq9CAvTj7Kk+MWnJ
WvTekyJklRj7wcSbdtV4ltR+7hWM5hzXxJBWpM6scwEOJU5ZxGaI+IT5RA2IgJJ9jkhq7NCJMUSB
C5AW/CXm6B1I+yRERdy0puVBLbyveYQbCUcNRO7iHob9SvfM5Li3MJa57tJ/0Ew6u6gbCIbodqLv
ve2m6AzvI1bPVGUAk6u4wbBLZPjFHpoh7lqdDdMzDpr6hgqkcA38/QHEOfntPRn/KOqAVM8+lFvB
KzpjQbyvw1xVIJVoQAA/dAX1CKSQGKiPWFgpnB6sMF5iPh78ZKDJeCNeB4HM32YI/9IQSMYfF5A0
WqhzIox1hzX6qTkGz2v8x10l9h9MxGIavWhR4m+oaKrHlvMlAz3cYVjADca4uYS5aMor1MHQ+jGq
n8lNmnlZIXWprQjev0m3sJ8yW9FleQtxPksa4mnj6XvDx6f30UkZFaLZMikE/clZ2aY8mwijPmBu
2oDfA9l6+RtdD0+Vz8TbYfndkZmxXJtVKyoWg8giUM7EuaSGlqOGVtggzaS54JdQxM1y7ilW4vvI
Mp0W3EaGTGBzAmP0K1aWXhZdNWQ8WxpSjIksyHhBewjD3peJiZxemde3yAsTxkaATlAx6l2Aeu7O
eJyfG/ht5TH6BMDkn0bnEPAr/xjnafHHA8nVXXjWLXRvWyaXnA/3HfiXA8GtKiHcadIB+yC6O4ux
lME5MI+dHpR7tUOR9Cq9+XytjP4s0Ent1cuPG3CJNU357JTi8tEEu8DFWmSFK9hZRY6b5iRWui35
fycgvASsaJrFjdv7lNHdVSSbRaZypzjsz7oPgWUa6FlRDgUpGQ37LyiTGWkZ2X4P/VEMBmqgYO+e
9Re9Kuo5YGeq6GjqrTJCiQ1j4dnYInVEJxBCBtgvykvNsvdo8ZCIosD5hcprt9M96FiPVF5G1Ubv
LrDQaq2O4OjCoBW82jJYVtxJ5ZjSgJ7sjGyGffZhnMYzX4SC5zf3eS6u6eHVQsCtiS+L0ZU6OoJZ
lp5BFk1Xxt35hUTFgJQW21XWDf2tcWHpAMZYcf7yR67rDLylnFTxivMnRUCJ+3TkmPtpSD2O2xAr
G5rHphGfmYrijLcfRknvC2b0Abi1JZFNq+I3ThH/fsTV/9GIvzY1JJJSIYBjKg9SCpZxGUohxZ4C
FJ8iZZ/tAZe3M6vaRCLsgN8rX8t7LtjLN8hG9X9KBN+8rE4sk+oVvCWGg8hAkO8VfjVRdhCoBeyv
WBBKN/GAdHI9zKAHN3aAaHp/A1TyKJ16fXUo0rWTaXiPmfRW8R6fs8h8zYPrzFNzEPTYlI5jTudI
EEnF6S0SQCfvzIncHG9t6uiM2o9xbK+K4yNg+LqpLqSvmLE6vXN99OX+YmXm12Yg58xrDlXxJo38
s6Lz381FcFCuSSwtUw2pZwEQH6j08BNODJPDfqGRjfq/SuYn8RmyjIo3PJU1eLKDHc7XlniW7lt3
GE18oKySdOl0QnxtNCj2tnfFseYaa97wnbkjQb++a8gNEwA0OfPm40hKGqFQi9RPhtGMpw/0Q3CW
Gb7HF6mzL267WcjQ5/Rm1K4b9/rB7SL9zgKrAa9i+Gk3Weq8xHj73tvyP1eTl/GcjnxU9/hKUBz+
0FMmvkg4zO7a+Jtqt8Q4ydtsNzkrUPl6XmQOWCKpiM+n9DRBQ4BeApzxtcabwKgK8kVBPbbpdmJE
4q64FrbNhgQx8CZME5t9jvha8dXoxYuczC0KkrXZK8sYi4T1YfvuvG3FjdyP7zPQrgLsCFeXt4y0
KvihPyrCQ1oWkAWj1p+lbAudQv9TDv1uFM6h2+F7CV3HyUN+yatXAeouUEH+MWt0rgDP7Ex1av+p
8HrLhKDfyd0FTTODGD0BbH5lEKckoL34XWDPwwVuZvTkkWehaEPQ0JKuIHs5NCPJ5cIYju+boeI1
L3mvBVyGDkyp9UWqRcRy/m/wpFNMcZd2aTEcyHd+uRfnDsht9l7xOfOrnL5cAHUeSUOlaXD57KAz
cdFRV75nsccY+g1t8TRKaJJKPsUTXRWobuTbI2urfrnQSPC8IIr3hJ2rNUkcmaT5p7Fn4bdtjGca
Yofvck3rzjpKFfoi8Bv8S7c1AUUndyWCw9/03IFoUoSVpTi91zVRfIyUOSEpZ/t3vgQkucLOn4QJ
SDbrUyn4ejTL+929fHK1XUSGQnmvxuFaug/A4c/T5QJtJoNIXne9563IpCFvUA7U8v8Lp1dAje8h
D/skOIlKp2D/e+xExTxEQ3pLEFnC6vkPHHaSntg01IZqOO5KW7QEBc6on7f3RdrqHQEBhODLAsBB
S40Maa15oa/166KTtWHLvEhwOEp9ktMUxPFaHqsbgowsPGvAXKGlJ6x5JDEggz3FgcOrExXl5AK4
ZXnbTuHTqPK63DiuZSiyHI+jS443aG23QEXKM8wYJ4YMxtvZBFbJCP9bavjfz8gVaNUCg/vMczgM
j0OYnzPMoSKeWLvJsbgoaMqWLsUzeDHRAsQsQakDtlsg4VbgifiMby4eB/rbkpvKLoQVBuW2qDdl
5CmGcWYKVSjZvGYE7rEUZLJghg2CSystUunHrHfWuKwQ32HbC6k7u+G2kQPFl8lfOtH83RHSnueM
IJ3RY+wHV8q7fhRZMo1kuLm2W+XRJNId+OlPPcVFGKRHT4U5vdEg8VdzT16rA1LsDf98tob/UXNO
ijWSok6861G3QB41GgND4VLDrfJNXAvwAJDi+qLOphTEIFl//nZSDPapyaDINO0UqiLSKbO5Ujyd
VlX3+bhBrNHteQ/VkOTvr2TJbe2KMsbEWvDkIQBCFJRyiZbkRBX7gClFBP69ecj0sCrfh37L0XJY
TaDh6jLrxaq8/15rAKeux0t9cE5DC+zalAw6xXbN+jert4uxrAsCef0dTz+NRwoltCfP1KXwFkfy
ewhxSS4neH04YQCuGD+FlTEHfHFV3LvsscFfJnjBo1L20CIBmxyG9WyHb7pIZNGrg8Dj9JgfNdEo
vO5yd+m2cOLmb7hlIW0uz3noinkTarb6ZkNG7dM3SnLPh7nCDF27ltSBv/aJTBKk4w1uEnf0GaC1
IHWSiwTU3qzbF8svZpc8q8Ro8cekC0RnzGM6kO6jOiIEeKMe7RLebEqU/NRlsrxeX9O2IDuXxCiR
rsg7jd7huBcgByfmlIx8yIRJow3FzektCajK++zkzO5CHWqjmTnsr5Km/jkuCNTtQhpumjatQbDx
Xc3ILSlHN7kejt8EgoSCDIf1ODw3OVYCfYaxf9dPG04HZNzlf3zLppHt5FOme17WfV7JrRfiCS5C
o5pze2GOvEJ/FgxtVdx0/cftLuEYIUXH1BFSZfslNRqoaMiJEz9G/phSSiHQWEK29op8WRJ0MBMn
WG3OllIuvhlnEIJoYr7gilOGKLN+fkDbRLsUfAFFZrv0KrwdEvrY8KxkTwX9lfsl0FVsc3Ln2CYh
kLtFxj2jT0VX5a/YpMGsnnxtpDkjoA/fi8HM2vM/ZXYwVPJDwl94IV+EyrHwyqYLprDQMSLoTVUe
iYZ1FpVmz4NR795rL6U1ooOm3XHFgU8RmwUne10G56UzSVHSirE6j5pkpoMhKTLWC7kUMXMkBqXI
3n140HH2qE+l0zWINHpBYWjOS+kZlmaJOWuqJDYxJdqmQchDbV2sQTWppNchLr4R9akdf0k/wCyU
C6YN2p1BnqwgVy//79m7ABIoWsm5ZMvjd+lpjcU07l99T93zvGRcyLbUDFI3WOk333f0Jtu1UYzB
lqFSewSJMJrPX6xqzopeWkU3B9gW71lFdvaMOLRobRmiwjgkd1iY1Le7b5mBgDTE81UKnMf8shkj
c212guBPbBfNsGGNaH2htbQupKU0WnB6Dt7TrjcVhrA6KZ0wN2jPTtFRc2nDxDQl0I9QMfNwT4Ge
H4zzXac0Y36BPQFkTptqATt74uEKmVZnAlFYJ2W2d/W2UdMWArVRl0SKSbPP8FMImordWBSpD0ol
QezFmCriqTH9hZ6/3/5Zbu5+ojuqvaVuc9g+aHNHmtZbE6h++OD410mvSNooSvCbRX49dJWGeSob
V1/xivurfqQAhSSne7W/BlREnjZwA8szwK7LvKSILjpaGuQQLG7KNRlGR5ywj1p71+/0thb20Lfm
ypWv3ER5n7F1WMgFZNs8Ts9LX7/RbRuX5fj1WlE1Z3jJIgF1JOREp+cfpPb4ioxlRq4bTo6Z7NB0
9QMACEO63giya4FE/SWxEQO/cOVyx4nmZgPDAWHjKomEn+PTJHzqrfHiFTt1bKGmrWbtkTaExFa1
qnKJCfrwhMLDEAsbeoPlaPaLrYKKSoqdFslfDQxSvfZ6tRoboe0LjAYjE8E167cC4msWW4gh7gS5
0syH0EbZ+6p1VgmCGYB87JxsFogdmE2kqL1U5a79sSmQ1CFqcg57Pj1A9jQZKyH+gKyCXsHVpgFY
nImaDw6FRrJ9t44280WFWNDb/jY41U7vujyWg6/FD+jWLogC2SCrczfb4zn1QDKuTRfw+YIi57m7
aHkSQQOVUIE8DmWMr4gDV8kHxyu9Kar3sxY9kC2YiHHtFMgvu/yTuXmv0g5MiIXUuu4Xcf28caJo
PQ+iDg9xtxgCLVsLsWFpM3M+oYZWhsEzKCrz/kV3EcsKuDcX/7boFf6nTpQYuFEdsGtFrV515ALp
p7RlfM1HOSavx6CfBMifgzMCvdvssi+GmolLyXtY6AJVbloKzQu6ucw9AHjTIPwspuoNuBM5IvSc
+4+Cuvv2r5zxAOW9zObC5Hfl/gLDd9TcPDC4baQ/hs7tZvOfKrm4V7WZJhgy7lA0bE0aBCSSmuJe
AV5RAr+6jnH9BUHTvHwKfjbNICfT3j48bzokel3ObOeLY2CudHJ+0DHTnyv0iyOkTnOCNpXRHlCf
nOQrY8XPBxPEPy8S4mcdf5I8AH8whvrL80sHuPgLS0M0HLNSnlu2q9pTn1R+E6F8vINkCDVbJPTW
6YcTfbNGA88AZil0aZ1V9O6v2M8DT8a277uRWNO9s9RSsBbJy6q/36lP5NU3jHcjw38rOUTXjHVi
4MBglT81czBkhOu+hjNxAkvQqck7XQGL2M+N0ePlr7ypCTqEAq+zEdYnE8d8hiOYzllrbavnSZxT
9JF3oGNcS7XBz4qxwm43j7pK193J6QS41glnJ1DmHECjm4KNihKPlgx7pKAQXcmppum0sN7cr0ql
+0zkV/hR1PmpIVZljxJwWBipb8cGdvPvU+Gt2/E4HJKhk/o6+ILqC1yyJA0kTXsoZQOJuVh+dnO7
bmxEtS4npG7Dxqt6aNIHOB2BDdffBwvQwF0ayc3pDMLUjthLzSYzWyI9pQh/OL+V/a9reJ4fpLN4
GPFwA8S+DtjATRVNx/fly8KMzDp/3Xajz++vgGOU9MVAj4eHBlXi6W7dZwrk1L4GqcoPIx5KqeQs
85VpSFiw/V+dvn5r7oYIR8PIC+xNe6dxhB0tMy5Yyho+NJhBCxlrEouJb39JYd0ONcvBNsL8oS6r
aZ4VpApNMUGtXITNy454SpNyCQwuXfUXFlUPVZJiMF+NJx+j9FwIopJu0RY7O0hvDqaFK7W5k6bI
J15MsvMBl8gdgyO7wwNb3l2a0zARY1SznqtAXc4aiemVKgW0ASKqYFpg3OPsi9RH8CYdxZT2ZiFS
r9OZYWJuFOtDK6osnSq1Bh1Rlb6xf6x2Cu3V7CVX1BSotD2nXoNGnbBFTg8b3jmId0TF0l6EnVb7
zsjvUmBYcM+YgKAomrOylQ3j7phYhRrCs8Mg1gzJbZ7t2gbj6Dk/Q0Alrz4lOswvnWi6iEzxHQ98
UvyiL9LM9i2gK6CgErNPt9cqGhxI0qM1qyVgR/rLICwNBNekdF12YYmFLLq/o0ELjFOjdcd3T+A9
WMXotzntoeG8wfy8KBouAAbGwEU7m4z2GedoK6LRCjoQB0IjfQgsQhS+b0Muq5F2Y/cX+rzkBt6U
H8fGw6a0/NbkLIiG83XWRrN33+KD00IuvStXSHAwX9Ho0me4QNuCmRzOLurUzXxECUqPgXFhqsXx
Zy8WOeo2gT7LszCJFPdRMXo11RC+jl2xrCv0/jBT4MRDW8uWXOmqRBb/KH6uvxC9Az1JqkP8wHDF
sTBkeKEubvjbBZzHbN7tBBUNaHfeqC93fNyPAFiXxQdyLFHe4kcOe9P1hdhLhFpjLSkOb4WrlFsg
0uAXgxAiNuvHNOvTTNmBu+Xr1j613bW0nVdz8DEEETBYAsNMBwr3aam3fWQdk32iSjqZ2gMkpU1q
19Er8rl7f/2ndOo7bJNrnBz+8fscR9LWzHPZGO+N+IFTgn1V1jN/rGg4mCxfuu/A3TLmTemxfs3s
AqIZN0IFe8pwPxopjCLH12cNHCzzzajgdNlGq4nKLb9p6TthuQLii3NV+2SO8Oyk+anNPJx9CUhW
rKEud55nW/TnfZ9yKpk9XFQ54MefAXd2TyRfmzV7OqwSMbqtW/EL0H1laPueDOqRb0Paz6HMwEkd
awlhAaSRUExVIEVN46suf8cpp/KBJ2FWPQPaHBhT7wCS7H/m/c30s79OWJtq5x59E6B8GLTSel5o
flSx+bxhGz3iMhSb073CMb4b9LBD2KS27hL3/uXy6bKxEjVINF4wn+ndn2hT0s5h1qrblfGm6fAn
pE0dTcU+TyNKacMN8rNZZBswO62P3/jzIC+MuW3089maqII34dXX9N0WHbCPFdvdhBNZw/cI+mrf
k9BfuDQcL4733MDmgwquNxqmxchHvTm83XQ4JiBs3tl5/MY6A4re5a7/vclu4GrdVGCCX0kiZJ/z
/0pADruOaoL/NQZL4ZoiAAtBW6OLdFwheF22q1gtE551hOG3wJR2bVtRjZFlWEslhxW2S68rI6JX
gE6guoNRLHFAwpek86gj3Xx981QckKtK/6KArBR2BJpt+jDQ28kOcc1bbDdo5kIij66yMeXC02Cw
UUSUM3novINEAmNgSBuo25r45mRJR0Gw5l3wjNeQcrmWayd9bmijAIBbbYSSE1OEXuguAAmxjaQk
vgGI9Pm9hz4SWhY+Zwt861F/jQcrYFqqAJdk7ixW4iymQAdKAPhkCZkPrLkO2pfhWQd0sk1EJsSV
QVno5ifvK1jorpPSYrQrd65G26fbVgq2DZgrH2i9gDNmI2AqZEKYEBJFPKLNw3XSrzT9T5fBtQpr
Thd6tPuswRQRqXXQPDFY0HawdAXWF26spXN3xHwVT6Ai2rVA+e31StzSEWdmuxlKV9RsytOMJVNg
3AaR3/7+G54ig3Fv9SFioidqu5Ntjog/LK0ms/bNRWp7hlpKLmeXbbtkwxLK2oEhBsdMCGpNlpGG
KGfJUi3HXA7JJ114zMSy+r7VsDyZtyBDA9j5LBBFxpaVgUmN+Ac4yR/0C8mPraKtbdnku1uTKHuF
EBAV7s0l1/otWL1FSYDpqSEND11Aj0PyzzuThhpZgGyW8aYENCAs0B75edowaalU7HNhKSdMOeyn
Qt74txubrOKbYAZL8UTka7u4zV4PIE41+3tUXeMORPwstxOzcbx6L1sBR7xNrkaW8jq48uen64PU
NXhSICfpKwmu6xHoyp8TiAC8fMt9wSVDSld0x3I60zL9Do7WUKmh9mmD53FHw+kbh3dd1PU61nc9
Fgp2yEM9vuMMzrBViZdYwV+bxbPYBCkvwKz1STkdt+6/ug5h+XOwDT/Ef5SzFuam6M2oIEyzP/HS
aCUkBIJsjWvoRHbBPb8i5Nij/aXbYYHo+rIU0qGX5U9Ol2kHtYD+1pcFyuHjbp+OqhFZ2+w1TX/E
Dt0qtZAnAVesqZ/r34wkizwk985PWvJTGvCOD04hbyJn55Yu1NbIMWk6cGqlNmnuKjFZdcAlDsBl
BtNL1aLc/Rcix2amBw9q0Wb2Jnx28sT8Z1XpkAEb2Z6cO9I8rgHsfj6EV8j20SZHCaqoSYXY6s1K
j+0Uqa+cSYYjSSVrZEiqJM4eI3pKAgvSs2/JIbSshzvxAdlY+WMaKWMEYq2p5Cb0Me0YvjiVnciV
b7knzx7Aljw4tibFIEAaqBuYwmF7XfVpmeSdY2uXc1vgxPu/nyU4wPkeUv8AuWuCMZBAua96n3lm
mrCpCSBPqbV2W2PKyrWBmQlTIvUf9eMue7TM2ttuP3TofBvx9vcsF+3hvQfSDsuh8Y+rIpVNxH5p
RHrU/XkuYrBKbH0UnZ9aiyXtN5g20Snt5UBmQtItZKlHpX1j/T4/Caym8eSuKncSvwB60w38WL+k
4UAvq6tKTTCyMNgGpC9uyug+h1D6zsYm8dLcls2DucmR9ckV/WCtSSO2QqaZfET/TR+mbshSwXSo
ncFbwvBLMcLkDk6qxN/KfBP0LIQR4xhNaBLKXHPidQnVh+Ch5wiVFl1OOsbA4D+bbG2G4wVSYNEt
tgFFPhC6suBWtq6qyCauSKj/0r5yVVh6JhM4sJ93X/yJR9P+bVv9UDq9W+0aU0g3zUD1bIEnwqXK
TCRNdhcCbRuRyYwnwRQzkV2+PmNf+cSr7/w+jvaV1Lo5n4tD0jD6WrI4DP2f3G+x4BPXTQtg69WM
9zpPpOHdx2tw6NkGuoYFy9nrZlI10jaTEy0Ts9vlGsZ8PUOdx65Y+Vfg3RllgpILRBcc1KTNoJYk
NUV16f+UqUjnSx3/OtZS9qiM9qZETpVxq+G8TEiFq5bPxeYP24x1SoWezWebGFPjXhcwIR4uGao4
IpwGEDKzsztrMKlq4Ll6eBva41mbWSD1eImpPFOu1OV4eKXFIDyKOXbUTwN9Q5751Dxq3oqDTNs4
srU3vSoqMC+rjjOsaWz3ikE9EgUxCyHYpw1sSAhzKPzx339qXHH7tgD7anv4mFIKRQTu1JuIa/sh
4dayAQzjBnPF29IsA7KUDWeZXs1ZDOAP6vUj983ezo8Jqxdg7EHvd7F3nOT/5QKcjqODjvM0Q416
Exq+J2zJySWKhY5xoDY3EcTmo6FCCG7N76C4gN9Fo+ZO9UG3Aij4ua3c1NgwGh0DPX7UlMBfxV92
Gz6jntX43JeFDrBisczz8WL97d+DoipdV0pMgpWzUk9T5kA5nbcVslbWk0oT0h8YXYTqTBPhTdVS
+LHdkuFXJDbbxMAhQpgy4dOm9NVoZGLuunyDf7iVmRMIjJ7dkCXVXG1tiPlNmp7IhnmorLR/j6U8
yX/YnxWrv156rQjPJhtQJcv0tqKSQ+6X3Yn02snnjJTzLb2GbPLCXtfY6wSen0myG7kXO42dZ/t6
0TP0bLCpQD9Oiy/fLK9IrTc6hH3sY0B2ffF+CumXcDcwzwuXRtwo7Ep6TABvYp41Se53GN3bIasC
NpeBlkNmS02YsrHe31Fkid/htlhpYBTqMU2l6wXSxtwLspnGIplwOuc2xgZO96M2rkcBh7UsfrEF
oraYz3WwHX3VBOkn3N+x5WVU95pAsbrzUEOoZ4EUsZJ0ig08jIaKkQib18V+fvdY6/KOBthqEE+F
us2bffTGNOr9hTmJlPkFlf3c1SXLS68fFgcrlStMDWvEpYtLdcfJvghiA2IlcDZug3Cg1C7bc/dm
NwuSnBqygt27MYFwbqN81GL54W9KahUGeFVjbO3PWnADbZMcQWAAqCqbj5eiXsE2EnLR9H+3kKKx
6l86QlDBdlzfrcZv/fJVuEtmbnKZ6fWUpbZvDOTnglk2mKKao1PtsA24Fa/JIZi3NPr6dtukN5Ea
CeHUaCoFQHJj7Qdnsbo6bhUVWVHZQ69b4er3Ub50/0fS/9jleILY59MmILz2XwvXTbNLibx6JmS8
/kdktGSxqik5HsVhcLCadBo3eVgiIxmrwPjCqkgP9v8JRHuE048iGD3OfrlJAffjCWwCdGrx+Xo6
aW78LK+y+J5fsGtn/JuDByKcuzjfUlq8R5mgpdMnS8T52/kr8p5x1L5jvvGu9JwSGnR7FfWMYHnn
2Hi8EGsJ77F9A4INhtQd5Hw5bhUxi4DRZechhixPDwVGqsr+z57EaG96qby4A+r4XZ5i/MoXVKwD
M+IJk4AktQcpGYGuQcDOAubqcvP7bQ1ySeVhJnVwIfc94ylT54bna9KhrmcQRmecgQlfdQ3NGaO5
twRUewSGrUComtgcfAumJ+EWUQw8xHM7giSTzjz8VKSxDn22g03Y6dS90Vhdcn0FLqItk/3s10rf
7ReZvce0jlUdwK8WItFck5GX0Wsp8BrcPFuo3QFIIZ1o5GE4lIMH/y7gC1oTQmjTfMC6UNOPReXA
2E7dKFaomlbUv9x0hfIdG1qxN3k/x1s3jZLlz4EVWnm+ogi7Gw2no2D4AvQxkT8V6n0aFZlj0l7F
6ir4E0Nbb22z98GOZoI4gsrYhum5BR2y/tPq5yxe7nRXktRCl8BG6Yrb+dLcOhSf0ptRY0Yd0AD9
dWfRQSgy7hPo7iwTsmtTSIfn68DyBZAZSJ290SJIX2sy/u4taehf/OGRc1MJV/cj/IFCmoaWiS+h
MdIRfnromcB9aEERwM6XwJWxxo/NWK+IbiusuUfGHEeJ85BM3eK+kvhWdWvAA1eJE2w0QVXgeHRM
ZoQvemXn7jsz55TOk0Yoi6PnJWciTdkv6IaMfao7rvC9Cr9eDloqvuDXazGCwduSSej2PDh0+Uls
y+pEDGlKcO+8am1sJD2l6ps8uy1IEjl1nUstzx6Bou75bOnDhdPBxf+XmrVHx4t69iF1/aCwwTwO
z7AJhxyj4F0KYCMZREgi9iqFqc0MC6uiHDf4ZWpfMKtKlamcAybpzqyl6hq/FpWy+44J9XiTJGrr
TrjoOjBgLLocMzU6vVgHKM8jOoGTCu1imFJxgNzOb4QtGq6Jcw1LSYaugwMLb/AOxjnPbWGO2Dmy
fL2soVCpNhmVJ9SrGoE7yGlckTGXKhLVRSbQonRfGeNNlyXGLermbSyDkaFz4qQA7zde0qqrE2pf
wLmJPp7rBSF1JrjX+frPdUOENOMBo2LK26vMKmQuWEsyspKB6idaQsmINfZOamBh++s/m/+AfnU4
8dmJOkCKRSonQZ3DUN5Pfba2gxH7uLzqW6qzKfyNxGzvdSGtrhsOBPAHox5EkKsrMqAzU1laUtEN
l7Zz4xH9+AlffKHDU5ciVwB+z36zt10m/ogA/RxGmJ1jZPe9/Vs0cw6g/AMdVNXHVjmaD5FZsATs
+8w/0zi2Y5B18hFOJ3BfpNsCRJTfQ14/1rSvBc2ldQ+W8sDOGL9HVjbIikiaupgqXCD/SbdAZEsz
nJbTg9izvpHuabVml1c2cjWGy7JZ7pTDHO73wWkEjo3R76yiY7+ozyY4xC2z0622y+TYz8RvXZPB
iUPXYmgRHp4Paah4X03NChRXNKlPUTZHaiwLGfGdvlK3kX+E+9D3digT/0BZy5s8wl6t7xAiLc6j
7WJGyOXOtZRiumNBuLNkndxbLXyI7gmgEofhdhIJ2n0ACELtaCQVIvVLj9FcUn6xTSdt5fq7VnQf
S8immgs4S9xUKGLfzYsnDSIOWGCv8SgyfEYs9TVpD7/Vxu8FZaBZttjwON2t/b6U1K2oZrstZn0A
/eeuZt79DjzcdmxaGTVDvdFjBIpM1hFxb0IrrFhkp+5H2LhmxR3oNK5LQ7TrURic5979Fuvmalh7
wOM9flHmDvchAxGkwSXgb/060JoYMEs/1CxWYJ7MOPWfGhND2FQfaV3fzKQBnSad7MFvOMPonoz5
Gf5D0sbe8QSiuXXo2DaJ23n9zXsBsTQHqyX5dzzFpBI0WYdUOPFlXytzDSJrFlGRwT4L8wRlbJVC
pxNvMHT940WSvV91qT0VJQ9O4fvJDwBuuyU9hM8YgvuuO4IeYilMwkZbkBkNwuvLYHIq0+/OTKwL
asQyt88hRdjT5olXTrw9bMqaa119b9N2ADOg+rj9lwEx1JzxOovC4vq1ltDIPMjI+3ji7Das20n6
ha3KTRV+7p/DDJEkJpFM0on4LwE2qVCPC7SrkSVH6oJGFT1uIZEMUd3CWrKBJIzyemfF3BHemYHm
nw/U3lFE1mJFopFdIWdjjrBSEa/8ab5gUCmoVBbK9nHzbxkc32+TejpYLyH7lkfjzyEegcdwg+MD
xBnva/MtavB8zZoYWybxeHhfyDxRUCI0nQNsqyruhcweNXDRXMRUNedXgSRRTnbNdxz1WkNrj5Q2
Rc09qL+n6Zs0kGYxDe5gUoOpPY/GjL5EU+fXszHWWtmP3kUeF3IG4yuq3kzOuZEXrKYexhQBAdbt
fpzpiTXBnSkZHpvj3ovhzMx2b+dsiuYS1bHyiTjM/6L11JoPKT5u1scgIag01IwnF9rU/B4TFi6E
LEUCbQ8lkPVswPywLqmRYPxP3zf2Rt2d0PsQrMrzL5sTfXaIdn3/dXbw43Vw9w2LZjAVxafVqHas
kRhChaD1+ek2f8OuDNk9pSqFrPCeDDcvkOr/FueSeZmNKbnY47pyi1kq1cS6+V2J/N09KPPA4B1L
S3m5yiAxtTkQS0/vkxsrLCzChzWBH2WN9BTDIpNpNFtq1qqtv06ANM2nWm4ZIRN+XOMrl3hyVTRv
reYPkXRGm1SeKxfKuQxyzcXQkZHTDD10VpFbh6yYqNhRsLyAWuz2/NfDegFdCLugjAKQaiHeJeT2
f0ZQa0UX2p85oL/Xw0eoSwYnUlZiYOSeRfOWwuXa3wq1jtRpboly6A1XjfQkwzMAxJknMi2cdtDM
takXYp0OuYFCUrFmGWHXY4fyw12ruRbI3Pz19GO2iQp8wapnM//Vc5fVraF1PNLLym7ZUENHLMSQ
W2q6N3OYpA8gAGIrazg6fzqDfDhVWqm6RM3jECF4/C8rwqIkp9oMwGS786vk+ppfemNs3XWfFGMo
GmVoI2y+KWK0qgmURAa1GRMt1Ugr+vRYxeOfrMJmksBxMYBOusOlnKhiKxQ8YnAd9wOb3dg7zBfu
ivXv2rt9kQha+6b4FHVG7jlSPHp2dw11CxIlOUUoLh84fubQA2PUENn+X224IU92+SBwnjz1J2Xw
jeav8/pQdTo1BJpBWu52LVXIGq9GLGEguw8rjW281hDy8UEA4ehUa0Iz6J8LQZLRY5wpsEFjGWil
vwuXJiPVYH3OugLmm+nJQIKnBI3+OPXfg1osgsGeCCBIS3Dr/QUyi5knOKpdJddEDLFlA87/MuGe
RvItJFGrLMeqCg/D2ymU5tEKY/fnM7oOkoESdRdHnLi67/o7wghGDB2aA2l63rvOmfwdGuAyeCsZ
420eTiOdYm7pJzpsz3gAJIUDF43GX8UlJECG1+iULF0iNwzEb3WaBOrFzUIy5cHtb4x2F7h9SAUN
+EiiKfNxhsSRHY3HQib5Wy21cYlx5yHNIIUI0vgPjsNx8WKSX8z3ife3kLrXzMEjsaXcby0xi29p
ljTmoOzcKS7D+h8ttD3fjnWq+ICDK91kGkVIj6hWvzu6Um4DGi/HdzjpYOj+KB0LhKqBCn3FzR3W
4oCe1Bs0g63SyWbnFWI9GCeBTCUGwkTo/B1d9FfDZMNxTsU6aYzQhTN+UqV4J0kYf485AYzilriy
ZMkZKsPTf+obXxt0KSjULQtjOyLUXgUkW7FSSzw99aw/re3CtjysH+mZ6Y2IAAHT90CB2O4y9iqL
JgpS0shxXJvcOVyVwPK1YXorpc+JyTVyRWvXun3yN02OOL6xi1oRGpePLfvb47znIokOioK18n92
SJK7jbhwHEsPr3pmqaY/ysNnYY4E2ANbtLetQVZGjvUB7kIYHV06k9bUhEiXtxV1g2ex07snnKGc
g7tRaQHKnUfJBWxbLA7ipCgU6J0uyKc7Mor0XfqEzqIL8qLQ9Tu0IVJpS4/+FHTngy4fjQBedIWl
rnBB++vvMhMlpUy+ONj1209uKU8jAGhoJ5xegVDWMj4ppCeGq6alXw4SJq081F202qUNcDec9Ruj
5d7ecj2NIJYGm0/258URSIVvfQChGziKNK9MJTMUkBl8fqGIcKZkDDMlE+AgCsKJ3dbqOVbdoJ8S
NmyVE7d00+j7GFh0lhRdR1slmxUFeVxf2WfhZyaFcoeSYksAPG/3Tin0AWPfCkHf7j8nAiwschGd
N9HFhqTvTJha0MnNJWi9MJT+MxCLTirUati2KNFj3gGv12E2rzwlc6j/40OiwbQfZiNlDR/NTHh+
M+U1cIwLUwu/qmz5WjT39vWKsbYIknUnv2VFrDAk6+qeMNNmygNtBmck9T70xxL+gZ07izw9tDCV
gOoDgX6+LYK3ffK0IBvBPkJs15nZkUjfnxX5lkYVSXdY5+IAhgVtA7cOsiGMbSGas/wgNUEYkafS
XtPTi0VAq+jGByOcisxKj75TtaZiK6/m3won76vvHEam4HL4abiKmmBRHk/7dBDvzy82rerVYq5L
PEqBY3eWMwBs1TIPKsyiUyDRGCBMviLpm7o6o/BhphrPFJl5OmfDLvrYBMs1Y/wmPyMLgQuo1gF8
iz3QZ8Jt5dR/ofkkbBIXbL7w5sO/hx8Tas+dTyPjJwjWehfhaJE2j1qwHGJVEbdvhV/Bz+HQ675m
XB6gvzykCfTGzrrPUQViM46mkSGPvq8JLQZwGkufDPpsDA0ninILHd9mGOiB5YsyTQBKfiwOsDns
Xrf9x1JsOOUzBo2MBBnL8oMyCwg5eV4AAo+txumxq0HT+/gRXPqzUTjNqCCWqEeSw60Q6A4+JNjl
STLaReCdp2b65xmZ/YcOtTyZ9lJX2zXVy6k1raM2VCIxmIe9eKs+KiGfmaWdwd3zd5mKttEc01L9
l/TSd/b1rlvGfEtpiQrt4Z8mCaAFasl2joubd0a8mBCz/g6Y/Tt0+b4mnpKP/dZDjhgChwQnVR6c
CR2E3luPA6x3C8VmeX5BVGAeKipJ7N7x0G2mxK76wYuMU+OpFrXugGWB19qUPH4t5EX1I6icogRP
f1i+yMYmjqpgLPNP1tsd/JCEO0ue+ivhRT5zkvzxkzJTDfFo4S9RY/IKPzfDB/LJF5EM2/6pytuS
uDVRYpLhu+gOCIY5cJ4L/cfJpO8Z8rIW9uF960eC1llMeKAHlApG44yETNYnfKObLTU82cFEEdQC
rqyZjDPYKCkjs63ef9sWG+N6Joigl22pgmNcaGFy0x/iTt+48cqrZ0NtHkp/G9OgFJ8coZn772xA
0SMvdRfee679zDjqanq6xxqGZ8yoZOWROiCA4b/leUDJHpnYjREuu6SupDMLjkHJHkU1rcKLHliH
zd4dWjMPyCFHMzVIu5zAn/LcEZM0So18e7lcUtrZhCucO3x6oMPDWdY74H7DZ80dhBTiELUnNOvs
DS0Ufk3nJFYk1cMsIhv+hwp7beBdTO2nLqinUJXaFrLqqvmePMeBcx86GvLqLePoradAbxHrlYpr
Jh7oC6Dy0UZFDxzisdLnHCtSVYOxgwqDkyyVys2zsbqUEy1uTB/iU9xpJtzrN+1e5xOGcssZxgjW
uRaUSTJbFn/ZYtlbOfoSYU3rA/2yMsF2LMXMsRu38r8+2hx0VimjOHct8K4eLaI7lYzXQOqB8beZ
PnHnQcJG0Sj4PdAIgYQ/MuzZqdwgswUfld3cp5WZvqcgsDC8/Qkf49h6Mzj69h7nOAH+SwPqLvEG
Fe/XYEffMdI+eQraAXesGSDYRlJ3qv8K+1Skx6Mq/0F3oom6Dd1TsHUUsPhZZbtoKgBCvVhTcmht
kdYBXExpAROI7r5gLyRWq3UE7DFNQcHdmQw9GSuX01zOaANEup/Eut8KFrixcoJPyxgpnHcLfJul
nyZ3mJUlxdkdTzWyxo+Pl3SQYACthtFJWSIhEuFHW7HOonIpmxycAqsKt6Jzqah6trhsz6LUFII5
Sniz0oiQZUTDI/S3+1YBZ/DuktSCPnwx0142ob5FlxpdUlt3qAJajHwFxYj6UWKTlLLpfa8Yh8N/
Hk7RibHcJxcPW+SgsT6CdKaMRROFc0WcylLyQaVd3PzH+8dE2OL2MQBqLspeQfud6v+iDIHz+/tZ
MFZBXNhHh7yOrFEx6L4yzaToZ021ZTgsJuLvXbUad8O5BVBivRg6FHiB8l50R2ac+KgN+JC2AEIP
c5saiCFNSkhy6D4aJd0NraCv9hRUGcNPBSdL6GU48BQEQgjuOLR3tUhvHvhMKfowNFS+XqE+hbh3
d2JfotScIWOjdo5CEMrIBBJPqVRUGZ2CXkYL/Fc8YRi0S5uEAffLrjpbvBIMQ1m/SenMM1h0BCh+
DPgL+/aRNqEGoG6Hpmi0cH3DfxC+X+fjPgNNxFcxEb3Fn7cCshtmOPihFIO85SUdhmYiLvHOb3mE
l8+nPh44Ic3qADTrWnqGjOqPGgtbUULaWAewltJGp4GSAMSEPTid3XvDBXxns/nukS88pqMcd2wl
otIO0p3UFmWQM+gLjl4NXQvvMEWeyz1DXshoxAA7yV+JD0/LCO6kmnUZtj1N1jpnrQOV+XB+r8De
pheXMsUVReAf0VnDJi0kUjOpdQDB6liV6vq0M5XvbLnppmowNrtpwTsGhR/MguB4yhBAyvvNrN0P
g3vw4Kt83+xGyY12Wmp3NtnVVlCN8Mx07q2ZOTEST1NP5noYPOE64PSHfprsudoXgynlppm4bvWu
XrvhHGtmP7NNpgR9ARSp0JlhAdhBrLLWR6OPEV2i1whS7wjjxoYAAVvpf9HXURUEs/IofCQRl8mh
kUPwdUDp7veQNAD74Zp6FTMgmqVNSr/gqE6tura02xCbtFYJUbMUZDF90AMCFzKQdJ6kpVWlB2Q/
GJiww87DISojonUyCj/+3xiRHN4mfkYIjOGo1OQPtjvMeqLgmQYB0TZKGxBlXz9+u9rM1R5pKe99
VGG+ipoki/ogsxqnUyBgLH14h4hfE/DuYyI7ourBAnnOK3vmlBmwWYELiHbuTHL9zihfskdwttJ/
a/GPbyHBVOg3RvomdOY4lAsbTCzexezaoi+uhgNkdmoWG3RDhw/0Zy4Ntteaba0ZU0Qa53QvbgsD
t0oOGfzShNF9PayLXiJpmHKCADOGs1gZ5fZcHSh26QhEvYzDAMpWYSUGsGcb3S1c9bHLAgR1CteS
rrwDMmCKOcehrZCgRohH7O2rsTNHwNWxHXdfmj1J4sYjf3dwDfm4xwdBRtvT1ouZ9JkussJ9Jopc
r0818/FjA2h/8sL0JqSaWr+TELFF5aGRaYVu9VNkmz3ZE7lDeA3t+xGFBkgbqfVkl2/Efd0hqgx6
jKgO+xObcupcDqrE8OT1uj3FajmyxHUNY1fbl6CsYN29T2UdaxSq8qM6cflh3d9xJaGV/VlwxYkn
fSLX9LFrVN/5/NHUxwmIwRqDkXb/ZhUStAzv0M9i2/GdRnQvomcE6fpnsxrAPspcNL/YCNAdMpH/
r0k6svSbXP3PSzgB+1i1W6W+CcjJmSfcRJbBDWhCEiK1xr+DPwWqwn8pPdggkPX5NVixUbbqy4gA
gAlURh9NTf3trMYn7NtcpiaI/cqmeJtNpjf3ei9BZ4cv1gncI1QZcK0QNXn7WTq+Xm73yOmJty8x
q62WcOZuA8w7MeVVTt5ROfkkPjDBO/P47jTbNfIsjBiX7Nb+xgyJGfjW4PwhMjVzcW5V/LGdO1zQ
ixMMh6hXIouQXQat5urWY1mKGNYWxpgb3t7tbKzGI7mP4KPyUS4/aaLU3w5mnDrMSSdyFWQDoeyM
mDXyJ5mLPMgJ+0ngDXyyxbhAFPB8wzH77Nz4GiFm4XEnhmld/4lulHzDVd7PyEYtEoBrkgutOAAP
weltVL1h7dGcViqP7l7ui+NE10hC8SZibYY3xIi1/f+4AFFmTbJx79sfAFORT4FXV/S+MZ6HgBNX
bClH1cLjrBW7WAJaXPvJLwcKWf20chQlH85bKOTZKglPmaIUWptjtasASKpezyI2kLVIxlxDN9Lq
Hyuz9an64Jg42mvpNSEYmIyFelroF59OUDDtdC2JdBuh0P1N0EfittbenTF10bGkxQzcZOzw0PmX
E7DfK2EDRypxsY6aaBjzK5rXT4C1lieSWcQOnO4WCcyTzoqW8cZlrQKZQNYUOYdVhfOeTT978+i1
PrtF07yM7AehTaits7DJxQHVAQRw6p3aZnPQbvfJVYDRTOpNQOgal2RdC8zx4bK3HnNytEws6bk7
YThCaDm9nt0vC4T7TZXZGGT4YNVvx9uJVxStWk84mcaz6ckqDnFUzER/qWRLMX54f89HEvxH/oWh
+OFI+QPX5dunhQ3xStgZwyelu8G/HZHuiPQ18PBqatkuHc0rmfp+qsBDk98qjjezKbyCGdF3htJQ
adtMbsF9oLzPIk+PrGSUdpoLEkCinFqC2gJHlo4AiCXMj9dN3+RSEOYa1nnREWOjA+kKO5BTe1i2
UX85tIwdQ9pSf+c/7UEQIo/XbfKecUJjMEBlyYOc1w56RQQ35t/Gby+BfoXpD1tse6T5koxy/21X
RjxXP2CWnCm4AZUTNL/YSVo2r2wuuyPrTG5gxqj/zkKm8ykFFQG4fATglBaWrx2JF4XRHywSMcZk
DjcQVZOs5ebR1Kw9j1Q8/giYwUa7Vdbsd7YuNmo7tZzqYk2FOJEIwKnA1CUucD/d4Q1R454KiE8s
DL8D92rmuJHqyEUcayGXPFjt1hrV2PovjS73cd3yQsIYtxmoD3jvTuUAQ+LNiuye5SsfBu2WtDm6
Md8/D1sd+57oCwgvU7tt5mKqr/8Y9DANEjo273BGa9O19pBxP5dhiPAsg6URu9LzHTPjfcjputBl
KYYDo+VcNYs5aYuPcI3S5j/Wp4Qc/lNgSnPCZw6vHnmBiRY0S8A34n5XYYd2f3+sjLewFq6R/c54
8n5HJLQj3wbGvQShrdRNV4Cjuh6GLobzfmqrCFpI2rtU7BZlT2kUMeirZBkr2r+h3xNGypb2OjzK
8YBI+IToJyTLGFxwKAXufuCuTC1hhlyNrUat/UhwbZ+krr+61lesNNwmeTUha57TROJewazDGFSm
wv1KtltW4B9oxNIaV0y2tHB8cp73etflB50afsp69GpY2/Ep59cTMcyReCLlgdSAvPeLsKvMUofT
OGihQYYQfu0PxCWdGTAVLCiIXY1FCXo3amNga5zmFc1rcnLLVWmYyVtJeHQG42pQWlg5T3X6BRPy
/6XXv9mgc7q8LwljuWhoxFk9PCK1YHEdwlw9bX2xc/tvYzqY0Fo+zD21MUjMOzzaatkCINccAtPl
LZDK1hCKfcksWFcJAnSCzL5pWeRCvKkRu1Mi7s0/I7Z9Le+xGRs+QsM4UKWINb5cXKVAI2J8f/Fq
RXibAB9PvUEAq3g6tO3QmjVig4SiE4Vp5j5HbGYwDJU1LNcPMwpbQ2CHGgaI7CUn1ADHptlFiD3D
7vC4vJCMf8Aw7NaidqCyqRaTtFnslb2ntczlr11bvtXyGuIBfz9RwHzQc6sIBATvbBEIu9mheS7H
k5tOgOomXgkyspC1yV8Fm78cmllSjZI82l+Fr+nguHqGDMW4Eaf311p62L/C3me4OfDAlxKfnDob
2g7p59R2vSqRGbv6b/IlU7ztqyPTga4Uvq6ksOUUQh/d6AfOnKmNRA35QWPv6cTxtSwNUsLUK/qp
fDrnReiSlq6wnLBi6jKG2vmSmHgRgOHF5VgBhKmaIqbC/9MjXDce4JNt+9eID0KgzOv3BkzDlsbe
NHmAhNnqbUDdsmbBOcE7wTSlzVgQfenA+JxheOq9SNmw8KJSiXU/dWIBSFi6RA0Xb4Z/DLkzKa5Z
di73EK7NDQvwlbPMjW75pUDcIuNZB6kiKYEubyouvB0ujfNbOrjNpLeXzgbhHp5c7iYJe99K1hSY
uEJtjVsCKh+K24Y8dmTvzezG/egOvqNFwiLtFY6XZftClO4B3SkRiXMPbdvSbyo3j727xAzEkJuL
t8lc4b1G0ADJVhUyNf4Fz5jlgGaEbJKePTR5s7I0fXhV/Rq5rqIcApCHR8uvwCrNZt6A+fiqRoEj
RCuZEHU3VSZOL7OrmGEOxFp9jFv+dnX3QZZlrxr3NIwkDz5pPYpzv8opsto+/b4EzTCY6sYwg0k6
DZzMjmhb2A4Gc+83USkYyvi2KfK/6/OKYNroVxlNN56SK9plOHsGRfsBCQEh8CeWYAJ8i7gSJbey
s3RkjhKS0cCnB07sgXqDqOZG5WCYglpXTOQmI0YCt/XezlSUj5kcwoZ5o/GiDBOHk5v84pzvkrgV
VjMNKPlXwBwW6aLJAnrZC1RrD8e/is55BLC65kmoC+9652rXnmliSy4QEC7kX3YUjLfKuS6WoTs3
sLRp6vzpRZUOgSZtbHeRWcXS6TjlQsRPLiXfaSpux98/D560i3urqjIwA5ZmdGs5LrFlQcd/s+Bx
il9QFOkntb9eqkIIXnKC4tN6ODZxNxVqOwkAIFpv6Vt74nGbuImCf3RI7yEviL/2672HQ8VhlidE
lBd9haXMpS+iBSqPY3ZWc2O9cKoLXyC886o3fkqG3RwZq/M5rCbAg10LObebbhqlWk4ewiLWRr1s
z3KG9kHvLn4R1RgBCiUOoPphVocZyKskjBQ4L8nrgzt9rX+GXzE6fQ3pbsbvlK6NgFIDwkVs8/Fs
rCY3X5UytLWRMeDuGH9tzpe+d5gZ2CZvX3HC9ao/BM5HhkoqptRg6DKREmW9umsbKE78E+8gFSoV
HzMmt3NCH2LmnXIyFr6CLoPwtEcHN0Kc5ZmE82vT+v/vGMRC4AL5nYxtOuQ6DN1etpcrNc9o3iK8
XP2GkbTC/38InRj3v48j5Ifm0zgZkLGYGPsAxv5lrimYbtbxZ4dXzTUUT8vsjezNFvQMqZ9LxVzd
SgKopzdJ/FormiaNlivLHDfpbCs39SumJ81dcomBFO41tj8FieLWKRsqHxB7GQDqt/KvVvRaUw0m
4dHS9ePN1gJSgf9xCNeFicqlHX/rDeAdCVkx9JhWQc2TElQKTIgGTkvqBsqs5YnKfTzsyKsve2Et
ej5wC2A4h26xkKHwJpq0mQjm05gXhwdr6Wx4WmuBjYbMYroxNDa7RS9OkcqStL1wNw7Y3mnEMYJy
bVaSgazOqTP4BlP0jdnOrsdmKlboQ/zuYrrIxrXBQlksl7svvkdmFReW4hOsPbnNkr4krvAWWSPv
kQkaAaz/va1VI8c7d7fqSSmTujUBjEoRhsMLTrlmzqQWnUTS+bEL8dZ5oQN+Yu8lpbQeZe4Rb6Yo
aBuGVnOVxQ4Zh3xTw/WAP5BCI9pK7nZXxTOEk2KO9UNrs/TUINGmnsGfRBD8OnXw5RbWDBvBEpiU
F2pdqVcobXxLFP7qJVvJl7/+AW1PGZOSxdd8oJfEkQ1GgTONGz43VTE+bQ7I14t3RBROApFlWhLn
+0hQ85uZGyddMakmr3XQ3ebnFExfOV4xQPQayau+7aBRN4cwM7IT7Av+NR6jclvbuw7asGr4nF7W
HNCn0RT7OT5L19ONrN2s3gcwQjESKyJ2+nGNRNh1+PwngCy3/RPZUewIraOhVnDmmS2H28TdxX/n
xjIe09+DVPQpUQKNSKE5uiTWLTH7Mh+njLckVSTiHM+RJ5TVV3R7jtEA3PhV/j9nUJL4RPr/IIkb
94PrOUL1Rc4uEzffl0HoMRmimnJdNXHPoURYoZqc1+nWjwLdbvzKWqkzaNfVmpevHbrh4kX7Nxaz
JwH5zzZmKH6BsYAHuqjHGuSOhghJuPbAhoarpWTs1aDxabF2FU9TVHcI5NkNb2zLvVfVcTEg4r1H
Z4rbaIEEzxnjGrQ5SlMwS3revben+NeCAcSZN7SmiyApREKdOVGmsFrLkxbK/yibSZNLrI7B3mwX
2nw7TATxXSj9l044LyzuKohTz1nYW3rDG9cr5za+f0+pzsApr87aZQJuftyhJ7s2hvKNVYnMaMqI
JwjU/2uyNd++3sAkmhrCJZDmhpSTbOXNi3+4+ArTPicv5XDnJt8ldArNxWkYYkHzqfj4CjKcbI9y
gNgCJ4Q1bGz3pqPIqXslRiExrB8X9SUIiDHddTemAiOusY3zndKGWcUAN9Lw905opPCuBTphHnn/
CZa0wAO/fC18P2/9FdK9K7ctDOrhkbYLEpOv9SQPpHrUnmQ2k76/ewts7EFoJuwSmvEKo3ifx6iC
uBQag/pmGtwD5JxIQcP02VbNPBERvtxc2qntzGXv7+EFFmjTKz2IrE2nkWqaOA5PlPKXrwH7zlSV
/QMk4MzAu1R6N0jppKaPhRR+mlaw6gvYAKpKxb4NZ0OTsBw/73yl3LXDbhtAQU1kuG78JNM8u6GP
Z/+QaC7nr5a4DaFZdd41IXDBC3BSueCDu1b8LHqTGNrPR+xZEVroM5bdkqppEbshn3WzGrL7WesR
nYI34ZESJf4sLngjpOKuNKdb2kfDP1ibkyvjc9sw1eKaafFgbSICfDp1h+m0Frk2KySzCGL237Kj
JQ6dbNi/FCxakoKgC4VsMyXxGbYGhTwowGz9XGvMxEV92uIdyghaO3cKaWe9E3g2Jl9SUKCBtLd1
OMimFNLa42dxy+Na++HKEIxkzw4TCDCaof6645CfNEtxsdblAWWP5dhP08ib6hQyTQGmdIfOAEv8
YgG1HFElW12aqfugfzZWruVcZG5LV18r9hUlkf6NE20g7HRcNKaSaOwviEuUDApaqU4LeQSQNexx
r+AGR2ZHz3aNbbgx8KGuuq/9oAmJsd5Bq5PwMr/ko0F6CGargp6Bl5CbC/T53V98Enyk/iDFVzvB
lLkOeGRZKZExdKXCkUS1Y2eB1G+sX8ePi2D3zVd9gOt4FEQgQIV/zelc6bs97/OTflpXmKNpiO3z
pDTcnGDu1uo8wA6lnDxNIZHC/YtRbH1nQrYKgNao7Ko62zCwuQ/0oc48GvRVlyfjq8oJtdbl7R0W
DCgSnYNsVPBILDH63gQWOHriC0KQXylUGk3X//+Ixd2n9q5q3uxvUelrTQHbLuFe60DIC9G97jnU
hWf5cu81eXAXzjkbaW9EBAB1BmzEXLXOaUkS3C5azi8+tCnKNMguAD0Dvwr55jpymHHG+h9jPxft
to7PwFTKiN4ma8tkAPMyCBBQmO9QS1x2AqTqDSf/mUrwrdUqWZJ3PeaiqJkZVuKRDEgcK4Pfv2mk
bGC1tENHwTPbKmbazjdOdaLFXx/G679cvMtHjscFS1Xr0QY5auu3TB8cdLUZw+FmHnZcsUAa7l8p
6+EKLJaDjjW/g4PkDw9jywOOvE6Bv1GkexAwLffwxJT5L143AJUnWDetI7zqCLF4fZ29I43PRaZJ
nNQ7Sq2YYcJjL2ZzyPs3iaZxC1VeJ2KhZqF3aNdLmOjUriRw67CwwFSpIb/fng4SKu18TLUwrSLD
4NYcDv51xYiOtu0m+tdGZ19g6V7rb8++R7heSGaVzFOErG4nXNm9T3An2gkwu8ANoqOEh85KWtdB
Xzqm45SYGi7TJIqkWUctFGYJlQYCdIYqzEbaVCZQPgh2PSbHmGzmhObWrBFtUHszp6X5IhVGFObJ
JjcS9MVn49SlghVNkNpSaoDVP0BdPA94L1kYOqesOCZSDC/NaTwiMILKii7sjwV+/9tukNiB920g
EFE47fsx9EERylfCgA4DFoUJgbIL3uh0CWczbuBXb8FyH3zwdXW6i2mSuI2PgSBT2XF46ZRABKSB
qz+I7/NIjLs4EOMebHevyIHlfP0RBsEbcdTAhmZ7JUEHKKuURRsc8f4p0XdEPsyKv4ole3bLsgI1
2j4qEvqiIDtCEubm/brCV0PWQyL+IGjdqkCzPAkAKDoq7+F4ikW1FSZcxxQtBDD6LMAPEdu+W/rV
m1xVMfgN1AwWFqDUESQQPky2Uwq5akBMe0HWyUP4rLqspr5JwmXHVxjOanJ7bP6uAIrdHQWu4RZz
W4m8xrxodldO4pQxURgH63SoQR/dWdLydaZtc4YYaJpfim0D3QhyJ6RhPigiDby+57S5aXgYarOQ
WcmS45nw/pAOM83pTm88jCF/45CODsoD5spYCrhw6mSXxDsY13k4v/sPVM0wCQK9a3nTo0bneppO
dS1Ji2Os3Vyu8v9715dMj+sUoHit5PB699JNKFauAiyEutPpdO9uZC7PoxPoophRo+CLVGDD4Z1n
eHzq+A5UUvIfVfBF9xVMqHG89P5rzvyb67Y4gYSLQjIkkt6CzVOzd4QFTFO8T5EtJluPxQ5XP2XI
XEx80RhZE+O00PagPeW2BdxSYSw53/izkUAY+gzMlPA2oWfRE+9rzHY0bRok+rMz4v2m+8pxwsfd
oE7XA/Jz1BsOPWrCPB9abpoujl9TjSD4CRElM6QHzwusmp98TnRw8i43c/nUzEhRLN6yHNAHc2Qw
2+0hOHZ/qkkPlqw+dhiHibx91KgZaA1rFMBdzOEnJjmC+MDBQzNJCjxens1AOTT2YfgoJPvUnU3H
+roau85JycD/6CmRqcv84nxSszyigfI9PC3q8Mw98+A8cdazvDw7bJFYGGC+D/FODTiBrhagKUx6
2nx6mJ3hnYauuAq1GlmAX/bQ2k/kaA/tC3SscXcVWDgoAGrhRnsuYnocxh1kGD/ZWx0CSTe2i+l/
MGGM97CatNdWGjDQEouhac52FaopOOx4lqziXdVakWyzow0wcvDnZYMB8IULfBAyajxOUEjb8nXX
EGkgdUtB/LK6xNvDgT54v7XAIbcSD4lSRJGk+zHTKAlxzkhPyr0CefQHErUhkmP24itlh+wHoMuZ
BqB+/XbWDmcW3TqguD93D91Ehu9r5a2VV2Mn/1tbLDiNA/iCZ00jqEd54dLu1XmaYmiFWxCuhB8P
Jh2q1LPfwcJcM7Hwyt+TpEme1d4hnOyPACWpbBcGeOgbwvWTSA18TofOB+CJe0HffAuS0/BCuemY
AWyRYY3fdLPMIUMb3bYMJwfnaBNsUJtR8WRb/LcWB1CEh2sqxSSBBwdDmhHaoY0qlymp+B+wY3FG
Swn+spNotN24N4UjGsNGoyzV4iyzdEmG2zOtl1A9HqkAASaiCTx9OaDiW6A9TQEVM62zMizU3bmZ
Yi2XjyIx7quIEGMq2/YIPyTS3OLY7oVyiV+TcYX9WaoKEmLpBPU18DnC7UA+8Cg2R0ujEULmgX7B
7fet7buBRQsyIIxJv2iQGjznWQZkwU/T4v9k5aC/sMtwwRUjbI2LHOGdnWxf7GIJt5dHcYLRzppW
d7qFBX7G+W+JWC2H6BxMEYRxlTt/wEYFocTsVqn5l4OrIkNC6bKN3ifm9hGpW0lyYIi1IjJJLMAI
MMrCFzladqzy6dOszpQXGRsIie7/d54yX/gq9WMCw6IL4cdgvS1vP21NlxuKTAmnzO1pDG2Chvwy
Cs1a4QcJQm0D+zVJYe3UM0ep+AjYyh4VLOO84zBg2Fv39PFcwkBi1OeQ6IK+IvlgDt+yoxnfv+4e
iXkJiokajR2uNfFY3cX93dKRKFA8ZNK0T0yCkbdOHylhKmoKPppJsP0jVNSW+0DDqWZ8Zhxc/Kvx
zuJDxxSuvzGp8kdRUC6AT8W89NiSUYPqt80FcCvv4rlCi9PHJ1utFo3Qz39EW7iiH+kAtnJGINNC
AotiW0AS+EbxWUFWickeLI3OSk1UUCXSMHiiQ+o/qTjUUh0SPvlRcqtByWwjFV96HtWb64rxm350
5AJhNQ+/vyQKGiBNQGv41WuD1AoXD63Ium+jfK9xeek/pNWdlxyQnpZHKCCLsgCOgqoqs97zobCf
fLwy34di7vaC7TuPFKJg6JFRwNfocxddpuXpkqJyQrY24KDd0WOrc0S4upUAvG7zsjoWXlHo2MQa
kJZ2d+iJfUH8LabG4OW1cuezkVn/kfN24ZYU10gz0ec/h9p03MYu5dBUoip8bjyHGdAiq7ypPS+L
v2xrbKlukBcwEPpgyI/oZsLtJL+ajTBS7lagnpvzBxVhTjUH0QLtuGwUpHTdZrOZsLkSOamgOsEp
tW1Fi2idSVPCwtqH2l985XCAS2tFKMYXs/kksCXzoPflPzzhGnKYyGkulKdJP/gVtZkAoSWSUt1p
2HYM/HfmLYxC1lJ+7Kxvde6xL1i9w/cSe5aOy+5uzMGIhPSUOruNJLQtIcpy1D9xj5mYrvPsqQ9M
rSKY180sL6Dgwf4SHztJmEZwtvdmPMKuSOa5urE/zKVe3SYxrQPxWGVFj99v/cpn9DC4YcEDJ7Il
I6kvpddjZNgsCIUjDQcLmYIKk96dCSqHkLDZyqZPTJEl8LwMij+ROxxVeFhNXCwTes9EnNtWr4/P
hLQ06Jlev90MBTVrfxGvYV7JKDTdExQUpbKsYXgx2wI4iAsAp9N0JygyIOxyiqNb9vsqXp1Ypz/7
M9nZXekM/rGgDlrqKrvdkaXdo4K28XRhLZpsZkdfC1UNMQHh0GYhPrfzdrqUArYKEiNL8xs/lVig
YO9UN8zbrdS3DRr4tN4A7Me9gr+T6DUYQLU3M7e2tCHIyMWX5tvU7eofGjxdfnm9w8tj7bPRu0d3
kB8NxHGaz/tUjEJkNNhasbpLorjF5cmfttvp+kSPE5Vv1kShaeDzHr6MBvod57Tmu9irLsJJlilk
4g0oAd2jXpVGSIgXeCqe6loZPVAbEerbf+7Ne06ApVU3QiaRZfnlX6hoEBHmW2+GArYbsp8l6a4R
aucow+nkvS11CaCxvz34TY7E/nB58SCyQ/86vuNfCkUK7F+kW78/YOFDFwIvGf84w+iTfxpkb7vf
wJQmyiAAlL0/KQoKblJDgYaZEc4rOjJSm5GihPOYn9x61V4FEzdbcjrXE8PzdRBvUmcxtAasSMfA
wbCpE4wkB5sN55thh7ib/0NhpOe3nY+Q/t6nV4DnHqsKvPAzU9OzD8tofMNMP9LJRmro1Ewc8qnI
vtaNCjKNh0qwj80pmUdOkrvb5c4EkfMgrtTIKIFilzL5F/H1RzX+3v8KcYopukVjrFNB+ZBBPsS0
PcVdHpREWoWF572EtvpKeWdTyT6oCpgwQstXVMtcehCRkjKSHyfdn925sruk78yEJWKRjWxBjpWg
eXOurB2HWuVV1zTX8aFEe5A1qtezALS5cXzX0a8bkUImPrBnaeYvInICYz+tdJqo/089B8QcpQaC
cwg0vVS0koQUx1txVT3oLpSp+s6GrgLKhM5TFcGKglR2Ea9Q07UdgL3IX63SneNXofpo/WjqbKqR
/PcgSLmMxzwQvvyc0X6U09Z6bh7GlNw0vGR9fFgy32u97pLWUSFXD3Tl4273/n1LZMPBHlQ5Q8Z4
ufBXeo8n4g/zeolP61UBxTBq4/LS40JbNuLVNypS/llMEeLlIJ109T2jcWi1wS/MjWqqWovZdlDu
/sqys3tl6R3O6ear8mfxBmx+8rSieACVbCGq4yNZkFMO7GhJi9M6Pwenh2y/nLuk3xxApLbRRVnp
RmhGwOr6y8KX6GETHqND54bKTzub244AgFejGxLHBr+bSWudJPmLIN5bd5F0itc5unXNLAmPiFBS
JYGG+jb96lpKDCXdYVeBp6J8dFoSrPaWgaaxwSz2OV0AeArBbyPmDOrttThtZqrwjaXSnPSWTSCz
ADP/8qdplglOyRGai0AhXz6ibLYzAnSVMnWgeQXgrQ04lhtnGOx62aJB5IN+XCxK1FD+ef/F2eqf
EDKAkk5PdpqVcVP8BlJAXAjMHxfmhCYeBlpJscGXl8hMRuMsw4BW0auVAa2nFEjKIUPlpCWhkewi
cPRlf/cvob9QOd+3aUpywVIkbEvmNa1Ki7QTWa9U/QolhUIA0ZeWpxj9q3SGuYjQOkXlIi6k+zV+
kiPnY1DRaAU0cdqWEfJwI/xiGijVLSsHqN9J/bxfdPsJORjKw0eQXsOl6Uzs+uYOXp6f1eZdAheI
u1k9ATFMtcLDW3Fu/ebO9jlmJ66BvABZ6Rm0m2ujvjSNWINehy9ZDXFcvQoODt023coguFwzXPXu
bVGhlvmr6/HxdfYAtKVGGItbWM37mGBcSdlFE+oAF2bnytmHCfikEO4+lYsQo34YLyUPk9JJOtK0
zA/T6dvvYKeqx6xxO+I0SI5vz2uz9k3SLGQwarNQ+g+J0lVUMG6trjMuYD/chNvJdnWtDAfZQJvM
pj2xtet0205DDFaceslGs/jh/DgVfES9S2phU+07ciG3aT3ZV4en4pdD2Nlo/G1nVIdxUTQSWVO7
cqqKNSA5kasumasgXJLnQJR0BYABOZxD7Woo/8I04SiN1zRqk4/LqgydKS9gWZMMuMirCdhGhA32
pgMkKLgnfgNR8+5CzrDjM8bHkZBhRsNBFhawpcMRQ2zYgxJi/JkSMEpwG8wRq0sfKt6+ZJlYUvkr
XYmxaXxmEi2GSzSP0f+JClDHAN/3glhcOBjwQO4tBzrtf+RIR9ZbnMZEluB5hIBcI5+/fuvv4L6Y
/jor9BgUa9BbAbr953G6i30e7t4tNzlLMHMufjDBxWa04+TUuqI/dlMAYmQ9Yr5jsfd1iAhMcvOp
d1W/oI9TQIQ/Mc+5Ni3CCEUc9rLrY1MutwXCjYXTvR5T+RwTYsjRpaZE2tCl+Vrx+2/0YMOGsqZ6
NxOLt5nMhzmpdPxYla1xbS5AsKHzXdKGgvBaPHaxxM/JBePDzpSBu1CrXkk4FDmYFvoFdb/kudwU
9krNsh8u87gUYhOjtZi+/8Br+eXkUGvX7TiXzS8Q748MkeMDZA8mxHn/gKsKGzqGwWsU2pwWYbXS
JI4EUhYYV3sGvHiKWKvdsH0OsMOpM+1cvEeyZvujGQsNyEfYxc4ke8ssVjzzg3kOZkUMfgiQ69iC
yofdP3NGEPvmtfe89ZI1gdGiU/CFQBDcIL8HYmHAuFDns+DjkoCDsxhgTqwLt/ZUc16VYStYcWs1
VeHWZqrCXki0DgJ5LipnE03jwqNZADK4a7DGC4pqyxgJAdUBrznAmDmn8aiYL1eMrt6QsqBZ8OlD
gPgGhCtTT425WAt7QrnluR7iCWqaBBnCV6OmCV2HTkgotFAe/O1HSJlYHZ/EuMp+LN2mn/HbstrT
GWVNdKC9VfE0kGrLCN3rt0SQy6/iA+UT0nq0KemNhwQa4Wj8N7i/s7topQbbMsOnE+PGbQcisX2I
GL5wMzSQT8FoZ6dcTqO08GRSrw2dwkL0wYAK9JqtDI7wwxEw2PSXrOh2JnQE7xADCnyg1QLCdxah
/u+CdULeJc69TSrAKDUdnFbKo9rU/5HVDhOQ9kHfmeTHKUcmST5W7LzhK8mzcBvBkBCUDKBXgO17
96/kP9VkJMwg50u/vu71pNGCXWFbw00b2u2cub72biqGw7jVHK6ZkGTfT0XJvk/juWjk3SPxmGUY
XPFzivauIweiaxtAMJSfP72BVIBGmSKRyGx9R2UnNaQrH80uJZDEcHmqPO7RuKgvkndA1/YOUWRc
z3j0vJQ75ob9BUcVGesALQaN+D8HSu6cca5ACTqB36dpQSw6DHn8QrWRqpOQqR48wRWDfnIutqJ3
hiJxhBwMeAPV4T1Hxt/Jjkx9AYJaO0FSM670RC7wy1VtuQlFNhpkSnrY8mp4sPa4ozdHrr3KjbT2
Avj6vGEZf4lNmin1E9CAxjFGWjVWsKOb9+xRsssQZWpIR2baNP35Ns6LWk+MMdUhpW8e1h/g5BIm
USrTAqp0bLCQ35PXJaka41kvG5+RoKhakwCPctwQJ9Zkf5GZ7iA1BbqZes0DJyqrQCKxvYw/fJ2C
XkHika9xvfBqKm7Z7zHuPeR6gqYA0NgSR/TykWblEU1YiU0ESyAUMhYO/G+vW5IopSSdd8CJ0IQu
p2t5if+Jx4eNSuyq+MVWk+9Uy8HnqSqg5FLwyxmXXyi81Q9Epl1DPfHPksiweMfUHfaCwDfHdyAr
/cznaA1cFn4votzJ9YZhMsto9CfM/W8fu7uFAGzB1aLUEDP/1NEgaQiVaGFT9m/82V8Z1QcpCwsS
MS6XumI4io7NRnnNCpMeMfVZRHCtUs/1+0wOy1hSzm9PFpbGMX73RCdzgf/aKazk8YIYaEU1IZOm
dWRBwkTiq0suo4o83O1JPuMIe1LPl9d3KusUnKWHhrbO0Va7FCsxKjtWLE3pjelHDgzdngSEIAeo
10yJotOX/jSgnC2VWPtNcFBP7Q7heExkOM0gi1qmdUcP5pmaWNb/u9qMEzIB30Hqp4nS3xib9rRR
IM/N6wjM8sNpd1MyFjXcoP2dDz4anCMkVIUj8f+jjuqDQD2QfyzPibn/MmHEoeaNtFwkDe80hkU7
huTeGpyIGwS0yzDewRcBSIHXj2rhTsHIhP0kRgsOfNc9XjUpHP2VzagbYlLfZsyiuGJlAL69PgtX
ZxtJduKxYtIuWw5tbG712ALfD7c13WHq3eBt7tOE/4Dvv+cZBccAKdgfwUYgN3M7aOd69Th0Ny+i
V3mD9Dsixlo6LS7KaVWbmebjLwrP9rraNp9UAlbrZDgPFhGz/d8zgokQQ1e5C4bYCoMUyZTfK6Vr
7zppqeQtUusDUmWDlSpTOcA3KuZQ1wNkIDBjCIjEh8+FrqUJrguQ0yxDFiQkPcW2ydU+bC8QuHeW
1wh+KY91tmr27zoolZsR1iPg9fADNScGNXxeJeYJni6EGizPhTh0GD4ryi4VDW00ncKj5uvqwL99
12kil55uV/EKhaIjD2rDZKOKDIcc1FGTfjiwh/SiX7L3hg27Cnvd1NSjf3G9isOOuedDhULkxUSA
dlkfz3gRt0CudctguUlLQx0EHdCvordAl2SI16sVdxGDFHMWM3oNrFuWjaiYQf9JZ30kU/q3EbCm
IfJz4AM75fSjPbYMB2AdYnIB4uapLi/5sHQ/EofRm+Zp2Kyc+f9Y9Iqw6hjtVKbzQPcIB6B70+S3
76Yyz0Cn4NYp+OX0ex42H4FHdBxew4NOts16x3eRqXEMY4UpTfBUO0fiHDN65rPe4vk0PqxOK7DO
cLCgoJp8r488mhsR/C9wDpw0oXhz5N/43pQbXF8aAP436p8pnpCAQh7h1Te92Zh3ZVmqrKMQgwac
ue6O76nF/R+AyhgZ8iLZAU4Nyjo50QHCePveN0gvq3uWGlfGY6x9sCQAhGaG/SiZETb+mi0yZQmO
SFfrnLpTwSGV4/mIhUvOzkCgzBrq+Aw6W4Q3ca/VSyQoBCIwq4Yy0lHurkY/5+8pDv0iu7ZdCykV
WomxuoaHkH0ZmlrORZKChdxxt3id3vc00lkTg0PsUB/7ODxov/u89twWDxDCvTF2D7Mo/NWGcj8l
VGDXq+G0FGYUhoHi5O70syjHTUvvW3v/9tc7M7c6We8bILsRxGmWH9bX2xxpiGByyZG8ciEpUK9b
PD3s3HApQoxXs78tpxzFJHq47TeArsjtZFd+E9jfOykap/K79aiHHCl5PBS4MPXNTX0ZrDWH1NK3
x+h7IiiZfF8HcDW8VtdBj2ioMkCvT/xo7Yk3UnmH37Op7CB5T0gaK1WVhNffAZjM3Owxg7mPPlyU
Pbor19ibQOzBs/V8oEsjS1euSxRPc2I/xHutNS6ppBbDibIXsqHsP54mv7+CB62OEocguB+BM9Hz
NBx19r0GFPtZpZiz27EthsLVHCc3E9PeG2mqu2PERB4L48V06pEBCagcYoKrj+sqUXzIZ7c5HjTb
VaWI63kYwEAFzCpctROo5LY74Rkqx494g9JBDzTpW7dC7wF7zzM8zFme5ZDvqWLrvp9r/VmnGQ6s
E4qfZhLODWUJKvLd474cnFY8Nq9HPVAmp+6b61ZvMQTANrjyNYoX4NnV9hBt1qC/mLngizQ6fBET
Aaq15UBVx+7Uotdn88bEaXgWsbF7zyyjcpPGxgpsHwjU5zF2pib+r24jA0rEF1Uq4h2CT6BK6y8P
ASpMiiTaQ0TsF/1dS4o/rKQHFTBp+5yPfB7x38geVl9d3/e06tKP8PZ8d4XMrIw5ui4RNpVHaVLR
bDKrDC1huOlG12W2o2IyxVXnqHxM9hhMtHb3DJRYGp174XUgqwyRrrhVXMpp+tC3i9wbwu03ZejF
ZVFD8DcwTpXfVqcp2b6+FQWLeVneagJeUoyBOg6tYcJomxBwhMzzU0MF7aK2NxX1WlUoEYKXyDsd
f5T9qMTFNeey7MvRnt2MlvVCs7pjHePUMfh7+GgQoAVOP5NfCnBlqYVZmtumy9LwataKsWlJGTAU
Fu0cg4YNEJuH5ccT8PjEjy/cBYl/2S97Q7/AVbBHh4IKBhE44LFg7hLLHplt+iSNq0fehYnoB2Yd
o3ywkxje4o/5KFdD8dig5s1zqdrg7wDjmEh6JIOGYb4x0qm/A7ZD+Yu4oRO0hdQCRXVTNWksWpbE
cAiQYKvMwyVgH2xYH2GSTDoAtdq2bRf2XhZzzVHAHgjq9zNTga/GmKH5DT1sulWWZythTNRncl5U
FGADTkseXL+4uN8LB8vFVIDkW9y8MqI6Q+y74HEvwGhsnX04o7HyM2RzPjWOrqR5xWFbuu2l3GLK
xiSuEQBo2iKq3mvKmVsRBpkeK0zy4ZURBPhO2BKL07R4TiGcRw/sNZY2eDPA/ik97kSV7iAG/f8F
DD43BckwNyYeXAx4MNP01naaLzCKxM7BlToL04JGNyGNczgrC+kjIAp3Ky2XieRYxOFRPQDtGk+R
t5PImzympM8AxVdHbQaRkW6I9m/nbDehqQbYWj1iO21P2equ7dDhN8FroNW3R7LRYukTRlDDhl3u
OaZHB308y7OLEbG3pKhCtn+FZLVTRqAtuelORI3SLjEZgKwIdyc9vSEtXiQOBQWfE4mJPWMqDDwr
T3ckuZplP6JL7Eq1AAdPu0KcfyzJn9kaP77Urp9ou1bXDORoEEhzcGqjgnZv+oQbp9POZyGCKa76
Z0E9VY5UEx7L3sVy/gL1itkZTVkyeA9eeoS4Jd+IBlTOvpYaQsFqPon0v8q7ha0fC9RWA7GRwYTc
ORK6GpE5l+Fj8SrP9cdG7+Izu1eDgCCodAnB57rqLMiAzS+TJzVjD3mSkpJuJ39N1agR1IrjlSNq
cV1wWkX5rM0PaCqiuk1pD1ln8nUIRZluXbruyKss3t1mp9nPe2gjJUR1+cHHTKcbGE3Y0AciLOC1
ES5FXfu6PF26jZhIe9/+r+pVi5D7HCLGnkyyZ76GUVqjrhdN7PBuMkZ4sovrIEiI266dLJEoMw0U
an/YF8G4qL5D3kCOmezWQTtOXDuXS1W86oalxTZCtnadQH3DwousKH1ZGfdXi058158ivh0Wa5Rh
1xE9YFvzgn3yRvwCz+EFsS91hrp9/yyfXxkGj5re/WamFZrp1t/i3GSQcVBBEOZKsQOFb9iCV+xq
IKpTZIKS+AHYgsnUiRmhNm4yL4k38GlzXOKBmdtAOwO85+IQcHgGFOP0P4TbBI0WSJBbQPEQdHY0
WwdRF+BtvhWqXLnfDsA+5VfkRXiQRdtdtPwqDTD3AByzfj9M3I2kahsYFyxlTGJNh5nA6MI8JEw1
yyvE9MUciThX6fkkQzgU6vGV5lwYtjn0QE8sqQG3qix5Cs+D1EHaW8ZQEgwa5pIRq/THx0Yz/jMY
KnmGot72OzcRPirzoR6caG8fPvcnZoaSHaRGilu3KSUZik6lYDwqQtVr3ON1QmOFwanI8VCFqQvR
Hi1aCu6m4d1Mi3BxkVedZZZMeZpyiwhWYSVI141ONCtmiMa4dYvxipnmvjT4RUbgW1jFooTthefw
YvRdnWlTEEuMw2xAxPQzUaHV5m3qD1T3e992TWzrdZHvm3IL9pAJ3vexVFbPF0/5T3bxcR6SmRLr
QBSI2HryaPldopNJESIyzuOBDxxWtdQZSBw/c0SDcp0rvtg1aBFdiGEcRuL5Y+9PMy8EiAGAM4eK
7ksNMSze4aYzQitlApEg+CXLHTcm94LBMOiU/TjH2yK2ldgYn48l+zLqNmYuM/vtxL1Gor8vkUYm
lfRrbR+QofMOFCtUz2n7ia2KIcDnjUA1Gfi5OWBMg61HWfETbGgiOQMPKvoWNL8Anb8gVzEzac/g
UkzA52nBexjcLJ5N/mDXP6qUQogPZO5nIakcL6F8n15I0QCkXVKSPASkM3ijKAZzvbo2ByJTxSSu
fQ7HsVPMw+9hcW7EFONsWW4eDEm4XLqKxoMT4oYsD/PJNQ5+yfrnYHiOZAPOZ+4Jzpwht7q2N/HQ
lXI53JSXRd8IivLEoFkIBuqQ0DvplFjhTWuSyb3L40UiMFHdAqI28GpTZa6N/FGU4KqeassmvMAx
LWfm+yNr6soU+g7oQGasAaZNFE/x3OXTS2/QJ2V2cLJCr5mL67qgED7eb9GRDJsUba8hyeV27gFf
BP0k2vXXrLF0mU8J26SH/lOvjg279T6/YZPlOcHag7Zbe3dZ5GGdIhbKn51lDdRjnKYvfi4dFkU9
gdMeubFjeZkCSI4126EnfaWVWILMwxlwVjAYPV5ZM7xmX5slKxUbJ/8vzqjKTF7rF6s5urIyvxSC
HQFiFLtiJgkxxLRXFhwtrptpWVOeXTG0A7VHB5e9ZPDQBB8Ze9gMvKBiyIzELeuEXEzNQWB/RzaY
0PoprNaa8Ln4JVPBRXUyA1termszn7eC+Jz/EWsEb1wdbLuE17Ogw97VqrbNYz0jmrkcX/ZFIgM2
nZBug3F9AWejtwz/rtOGo0w0BVHGAQwBtEbFke96+UV1bqEChLYD7iJRPMLDV6U1rXRK4KtiHrhD
8whp6y20zuwTc60TOn35bgEehubeKTO9bjWuHrNSfXVhvo42j2E15lvfuspxK739acN+yKNJKkH8
JodDPFvQJJvcw1jwNBpqbToSIqgE5GmIyKfu2YyfSvVCs0YqkRN4VBLDPL7ss9T1hHXYjlQQrofW
S4d06Bglqho97fEmyClqgzx3eZdG5ciZ3UYdCD7cC8kK5r5ld6tZMQaek3UkA+1NMoRSSH+N7gBs
cof3UsW2jjHf89+mZhqLxTDApD4BeAiTnMWVNuXq55njGvGzAj0P/HyM2N77j5qp57dIzaIfD0Xv
HOvj6yS/Szq/Cqj/QOJEXYusfLgACjncHXv5ZDRBuxguV/4FzSPuw8LUaetH9bL4VfNhKh8yDI+H
sYWszW5ZS25kgF9lZZ38Wg7QhbXtMaTHRlm4DdAvRYbqfpYpTqY3TKP4ziaDN8sgyngt5bLNeIBH
gJgKnseHMHeGOjbcDyeWZKKY/MJYn7+8IxYjhUJ09Ng0zRFGiUxD+MtHzxDmkgjYXHAr48cQWAYn
DR5q3ucYHFu6PP2+1EB6C+gBMGjtJavTW2kxwXUHfKAAOvo94SJQzx4zoLUd8lUlksd9rK8kn8mo
7LHAk9poDijuygtji4n/hqyYE3lMZxmZT461vmntHsKf4V4jcIsUi6V+8qsrY3WcKK2ElsSz8mFW
dhUvVcMA+KBdQ3IyI/tx3wmL0TLa8sw9ygmAG/SQ+MrtOpzl0cLspar/UQ/X89vRYHTtGLks9vQa
xmp+xBvUYpUuzFgn5r1uNxj7NliSWwPPOYJXxCIQkn7dFpudPOPnZk60d9idt8VWgkWLdAU6M9nC
4rFRMToLnQ8V6r/3eU2GfqMIUrKAdMz3sSL/wM7wcnxx2pwohb+5P3mxaOlkep7TTThPjtaVCOkr
QzLK4d9Pb73fnfiOH4wFT/0V9n+XzCcLuTe/P8lGIXWDoT238Rd20sr1oL4dXn4QDqjRv/PM6joF
N2ZIhITnrrsDSXtlgh3zga6dy19s8VrioXsK/hJgv3OmfuRU7dptuqrjumrC/iPWEck0HIfxstWp
jbtT30lST/SgDRTHR4nj9Fr8VtKc6q2507rsJaIxSftO50aTbNuYhwpmlzZID51tPkt9P5BgivQQ
keRQrPZrPuB7wstGrXzNB/rfNcTLqSPQ4O+UM4u7sxX7FwvQ31GuljI77dkuGBFgJIMrP5xchIy5
I/HWczHRzfCk58SByvJcQnl3IdtkK6EnwKehpcY5Y+geStpvxQz6dQdPxld/q2JfIOT0XBrZgGq2
X3cJAcqbWoFpEf4ZhHLHwhGX3hhQLyS8UYKJC1SbVGzeF381tltHoVSNORdLhr1wIewCbvKDZOoP
DVefQxMFw4c4RK/55PJC5PGeCuUmW9JLktv/ncJZbGn1Q0/Q8cN96RRquLBqNeYOm1jgh1NJ+jK+
Ug1I+bW5K+QZM5Jj4icQGYests5H8+TE13gYtV+J66UG4dCEMwreamvqhND/rdKVgqczH6xNKE3y
ne9eSj02euM4nj78oEygt5Er2YpDgQoKy4Err2jsAUgkxX0jvL6qpfJUf1O4fzdX+7yiOzaAwX3b
1Mt++/2FY9jd033lejBu7MlBu8qVEsTDqPE1sw4DYg7j3l9xVyjfWnQnQEy3TEMRGPHjCf0wjd9d
1Nf0MFiaRYRT1Xrc0KMikY+wLqZoTxmmshF8wyLV0rG9ARUcLSc4odR3IUWwvqVKHxLt400GPgPH
CDCFREtyHaqcSLrAX/qQN97LUKD5QOZyLbJXaL1WGFkQK6NCdzbND/iWt6htGb7c+krX+8HwpaPr
oavE81pODJ1BCGzLzJshy3fhEbJAmVAW1doJsx3+0tiUcIcj23x+jA4noOwWCv21tKiK/u6VfeKm
BYNV6OVSegKsoa9cW8wJOGxvyTSoEwL08ZuMWzV9dqU5MUu1Orc5Ko0D1r6EJROaE5vMVAGNqIVd
2nX0ribIgY6lDvy18xbiSCqyyphYgaIYEOxE784um/QuTT5o6wReO33Wnm+QoH/RMS6XLD1uSKhz
a4YjEVPF4WbMfSLvfPKosTlPmQM9cM6BLEqlbQmGQOTHbmcKHAyeIzE90RK3DKEmIVFafat87DGt
UTX0bZYrLWIjAxoavFDDDzKzJIHHuTnO3Yt1pr+RGfF38aHK1TicIlkOTjIKAyhCDbePpYqpOQG5
Cm66loIcgXNU3ZOyT+rL5vT4BVpvJTy8Ln2nvaTN9oHlWhGOl7ZaCSwvXLLznM1QX5xyD1xkfJhy
f4Sy4mwrG55Vb6iTlbSU5SR6U8paO6zWA895BIKgZWl6v5CnxiHPRMKGLJARpxCN2POv9zFLhZZi
K+h9t8u/OzHM0jc4VSu0m1RPM9AHmFMoE6nhgcawZEs1rg5toUr/jFFLFlITR5bHlodsZP6WIk7z
6MKY4yWBr54PlKnZQWoDYyIVXjhlAP2XL3WjDBb9xjvFfi4RRjF0RYFC6M7o0hKvTVE2eT4J0VxQ
pP++FSRA8LVI+p6KzXuV70/06BUrktxa+piKV0ZB1QtCeMCyvk6xA2VfhC3qxD/NvCwYLJkOOi2y
W9pn8NHW+Ljv+5sybihF08eoQSGV4Md/QMKEbL7GqlocxAbzGzxjOmCyu7XG6qukeJCfzVbizgMH
TTVRvmUa8/9d9lHmUn72086jI3xVblr/ou18ok9anmx2zAvYIVZZNB0nqBm/2dvdlWaCYd0Y6g6k
R3b7hwqdmdbqfJPB0EW2uj4Rr0TQAQH0/PcNRigxu+pCrysMryynGm0WqNEaGnoPpc71TaclKdh5
nMjPFv1zuHhecWxUiiZZJfJBgJii3KC/BG42R8/HwxH+hjFeRhfJOQcK+vSenZFJbvW1873jua7I
1WgoWdOfZNEejarKvN+FUZhX0t5/r8yLqdCQ+SBboEUxXkaqlKcNbzN7zIeuzgv7/w+qIMHb+bNx
5s9bgt11DQr6t4gxovXS2h9aMy9Cvx4tXxioanK118+yKwoFy0f/xJ5W68ecaZTw2/Bzl4IEhBkL
n36erBT9wjiXr0vV3NYJuLoM3HvU+m0rbYqfDTMgGkonEL7V1VAzNWs6DAWd/9ESsHH45o5f4O7K
V/acl43hE+OgfxliWJwiZxQe5GrXRBlVWCfnoL3ZjYHLOnQ9VK8ChOFony7mnYIaOAhqpEbUCDvw
8hWuBvBhQqFRTKm4Y6uAbaTcjDAoBRXpxNyGTzb6lX6HgAZM0ySX0zVfOUT6hbyM8KLfRKnJWB/a
MTiN2av1TbRXLuM/2lnHDO7QZpTn7/JcxOQZD5JK5skWtf6pzjhgBsoNk9EwA94aQ108ARHhRb+m
cpom95cAcEVJe5ZumSHI+j1S7tuHVeH/cFprUeRng+qROfpduN0Hc28lAIivAq1VBE2/qehIHP+P
INa0rJrHZLUMp7RznszZrF67dqbhczyTBlUFmNV3gq8eAPrlgPm2TsYHTkCAJyrtBWvH+0HKK96e
GEf5tM7RWcxnz2Mh88XDCdR6GgoWiHuLo+0qOo/s91NrF5G3lus+nCu71gWeiOPgo2dZsN0mFjyr
9hElmzWe4wmUmSpx7ypo33y8RODX0Uxe3o1hJ/CXrSuPz4Oit1lSIMiPcr4hghegHH/kGncV0cWB
oyZncbeBEeHv57aQvo/pCzbRogLEf63XNiIqIr6H9sEZuOZVeyW+z6YQTAkdHqhlN5lydf8EBQiq
MDXaVHoh59fzJ13DjVXl0+ULbQSNELiQBGEo4QmVlsV8jgdJxxUkIn0upesIoBDcxax96t+/Hwh5
zi87iLXZvf5qSxHmhb8q6FiY5LE5zillVJfIOGLsTPruCjlSDl5RuXwPjRChT0pAft9n7/ZEuLJX
MCeGTpdUwtq3bds1+1fpJtHCeE96tSPJ6t/Safj8hmsHYJokbWD3Zs28RuldbC3VrJumRxnUiZ8U
/H6sfMia7v6OCK7fLFlnU7QvIvWJa0kqVET8GURbn0/2Hr9wFu1JHd36m/WygtDQ3yZs5ghldoup
L/bOqB31cENoWPnfT5mJHiXhIr8aZBcDvRq65XVhuKZNa4uLOKZQ0l1PUG8G71NYcE3vNmuQymp4
CdSq+K9jxnACi7ADojXAU13793yTSa/xaX6VEO92pjyWcXar0AQNbS0/wB5/j/ZAW6KJgoFCn9KG
0N/J71TSecfW7kzRxSQ4RBHh3h54iGyc8aHRy/Y0EUwPfAH75fwXxPdrWMhC5ryYoNHdQDfjniGz
0G/T08NMOMz1HZ+h3k7pqs/M5sIeugE6uv1El8iOVHXHnanwmmjVb+XSFjFHyqFUrNrsyV/DhvWR
RleH9+b1bWkglqERTQRvBbW/klcGe04LXGNsoo7t3IL83Dyh/2+3L1aMEHHqBsTJCUpbM3y/u8RD
tk307TdZfavapui0P72NKx05VDy4J+FNu+ssmBf33VHVNBn+gHgvr168KWb/8ib1BGOwDcvIRNnd
nXow/swv6RpYTQvsrtrYebw8KZDCs+IZsBJHEcrC1YidLAMvHUN6cBcUG3FLdwKgaU4P4We0rlyx
dggwmu10FfRY5Gx4TxmaW9lUmQ1OMCzzB8IwXrHP58ZOHOFcEWB7VEPnKe7bYIkG3vaBNd7Lz/I9
n123K1NUeDdmlVCyPUcqUCYKF06zfv8whHW2gwDcJrnXCUFK1oUgweetNWwmUG+RWgL9DbefwJtf
R0CBINcn2g+BnYkjYZpluMdcPscroex6soijT/r/OMVrvOIUeK/F3GJXLFnEduOv3Id2vHEZpT2E
VWlQNtHTxe9LIc1w6t5Mn3EOg0gix1SgANGQu1jTf8fGXO8vumRfHrfbe+RcsYXZuq54Grpqcnvd
a5frqbF23dZm5jhefEajtahdYOk1x/exxtuzL41GWxFTo6mDrFgsBpAfkwLselbzKrfeOUEPQodD
K76ZLLAYUDs/zgf4Lz7b10D1j90mO7/2gz70Gpraxv5znyVfqYKRTfVsKPAnsdtG+jjBwH21tl7C
AF1hlSI03jCOcaiWcZAUBVYoTyz2GrQ+Z968ig6ee3/i12e/waHah4sdoHOPseNZA1ngunOgPVmD
Hhgg2m6d+UB3qchV7bF7w6nyxHfendL9/TFK4i7bFp3/jvylsXPyAU8kYvGA9oTccUY19W/hJ32A
7o8gN7P79f+iIzOHm33mkDMKzZz43sCCfyETzcnGv1msohUXkxWyaxVgJbOkY9NjaMBAiV4av5BA
4TP48ozVhxfeTaE8fHEsB4Pjg9FTHcN1+Jx840yRLBfuutD0KWAW+NU1g0u92xCgvefIct4yQ6F6
wErhZY1L268xOotHzIgLy4V0M4GhQATlO+CDlCHdHjtF64z5TGfbNMKkocweUXvGMRIXXMTuTvLw
EhNO1TSLpSgns0xZaeRmVyeIO5l37e0z2gt+uMqI7kxEKzzZ5aJur3PnyXGCMB5JSXltw8WIHd4n
pbWZBqMjcHg5Acbq35hS9yAVOe6tfzSzpsfj+EsqN8zW3dP8ZSSsJNNhsV+dw+Z96UpqQihcugzF
M7JQHYLPL2p1Diq+RCElAqKaqUl5BkeNYWCxN63lBUkhfmTzqugB5YqRaMBlumBK/8pywxX9Dnn1
YJa6FN6KAg5LD13SbQPifqeKgMcRJ2xGi84JkEohzRdqP41RxMFz90Q4F1KCooioJIK6KvpyDTI2
oFKp1BOH/ncDqonePG+vJxbkJeqRcK3znQzmQMhAzimFzUCgqguk9h7uNBaAXJKaFT77aWuQT4mw
rdts5gYMayBH0/OKDjySTpP7S+QnrF0IJ3u8OR+xoiDYQzcJPZrI6r/GzLyV1Zu7EAgB27H8ldgI
RutJt+RSE2gjVM7JouPa9tSeCdITJuKV9PyW207tbTMEk2qQnAmuDyAyQlxxigCxNGNhjJwRkk6e
caG4kU+mCfmWT+PCPJV8cGA/Cnlp47hQC1jF1MyRFgDHV/neDQwKfay/tFahbvST5l9jjHJmlkBA
3DE5KHWtCpx22uLR5jHClcGIcrTd7crHXCFc4cU4+dqzU6ramlyJJVL8MhFTqsOb+yFzc6By5E0f
P+Bn9/BhNis7g58kbhcwWSWhFs1/m/0tfcqWr+XGg+2JgkztpPL6wErl2Gu9QteYpRKtMnPIhgC5
PSRu8dQlCAHLLS1n3OWChWZXkqhaIQ/8Hjhg0cb+mgfuFg3cnVQQZcf/O/0psXhJR8pQ2zqxsYA8
ftdUHPkJ/CBDaMLi+bQU9dI1p2Gqmyid9m8K/X2hHxRJ3We9RMEbmsGumQqx1iYgDt0u1etgNg2p
prx4ZGYs9Qpk3PO4wWpB5F7gEouzHYKKbvcDih6LYaazrcjl5XRySFhhdfDn4TV4In+C+gHlW5Vz
58LRAqCGjWjA3Ac2rGxij1Bl3RiGfZhnxxcfvrVQSntobUC06jA3Tba5YUryTF03ZT8gF0TM1kcP
3bmUHGElDWIdPzzXGBQ90FABQTzahcY2UM2WvP4fsNat6nBmX4qEommb9yF4MO8ecUaLReWzrw2g
OFu+RHAJxKG5PJGoVlPDgprNul3R1tzQyoPUUocVhRTex07T5iAQebSL0DjYQ9rKYkLO4Zi9KN45
mc8T1+wao8cz3wnONbJgOdS8XSmwkGnt+swGTYflTwoXf7bhC1lbhO3SQVNI6y6cau8FWk8b/lCd
ZGsKMyip9Rt+WBdl1Y79qiu0wQUUwEoro3Uc7Gxf+3d3U2mIH8ahbspeQrnqXgY+PUH8ehiP1OAe
ILHENdLQlcBRAE1+pAWb8BP9mHcI/1hWnuuYf7WpM/QFunWWg1Ve43OBpo1n6d52oexy+VGp+zHq
4nVtLMut8+KhkDaKbpJmf85CUTbnDuJyURFzFqtgYYzaVik3Hes+qAoJ2fc3Z0Mu5BkPOeQaOlYI
pAKnqz6P4myqh5m/BfRuOj7qkj2ZZP/vCzNng6//gmmC5Gh2FCtX3AmR1k/ZzqaQCfg9DY9d9GJp
nHkn3Ep56rMYlZFPx5yHF7oHyezYlklEg7U+9sTclyZHXZVL2nGubUJgnzfVjQAv2/UqXlhu4fzG
rmwA0CUuG2p56oSbzhy0G2To5YcgZj7EWRUcepW18OiugwhRtZLkVEM8Zve6Hi3YgvfvDgbRYBdw
debckoVyHR9zmeHzWuO26DH42K2UnKOmW5OlGwBkGElKbcR2NozCb/fZAVJqqacV5AJf+KfNCf2u
BDugCuN2DmXlQv1L2WbPugPmTu5soIk8532VXOH9hvv8cD/qAixW1ES5j4OSRdKV29KvWmhorkjY
OS+Ln9CKt3aFZU/O+318s29/AVWhu+tq+PMYJF2pdvF80jQX7pi2BXoPBVoyJglPuxFe6JzklJBg
cgbA/TsL6Lofr/jBbC3xiMX/tiKkLvd9PyStlyByLt+l2rgvs9LHP4bcgnhS6kLnQ4XgfLsWMt+y
bSg55WDaDczbOGMsiBeTL02NIf0NgbWKnm04AxH71l1Boq2QRXkq+wvwximQ0rwogeQIYMgbnQo0
+ieGaIEgHAwUGK74+uHmFYdlDXCzZFYKsCXn0jOTyubrno3V/mdSGd8Wu5USpKnQ6pVc+HEc5B97
n72g/BhumiQ5voyTKTjoiIAlqrO0lHfcj/VbRMkIImb2JsxirZ+FtwdodWogusnE7vl6tz4YkAjX
VPQNiWEZs11yP1v87QHfgEwZcAKnGGIS7vUxZxcytZo8fyuAsVIwzzhHBjAw5ZhTNq2i1ZO4JKd0
A+cCLk2Bu5XbhJbxqwYdV/1XKisQbtynWdN458f1cKPykz/sYn0n53b5JOW0+qTL/OlKmZXB1q1w
Y3DQHPKpdK0LhAsbbqqZBQr5FZ5nPx1C3nj39TGiAp4btMdZ6gS1gvF9SnVanl/sUJx5m9/vFQA2
6MbdqMRM8So02BZx6u4T6QILmd0RjY0YyP9tEXKBWk7kSyRkfgiqkebqvwQdPAZ9Hq9ZKXwyKLCd
/V/zZQzBoMSmV/6vQcRQhGiG+C1C+VQsn81KBq4TRpTtBGM1Mo++3HMTT+7tQX+VBPbY4MBc5Flr
jfCzipR0PTOWejAhijLaUOonetxkuiF9rxVoj/scjDRuRkw5t/qlLw6p0n4X28YdO7eoQeVi77j2
rzwBHnFWzPQ+7HBTJTfI9TqxBY0lY6DgvcYnu6IKb2IGUNi6VopfFD3Ud8jDETA918deZ5djyNsD
aBB9n1v9wLmDtc482sUCAMy2Upw1uK705nOXifYC4LL1waC2b5pHvxrtD0WUyZI3xJVOjHWrIFLZ
e3Ew/IxnUKiHb6+mW3Xg26i8kYpHVvKtPr9H42bccgxL/TUfZMsCIEJWBvdG6XXQJtVNPeMYL9X0
bdaOcUFSUR7mcDtRBgOIS1a1LJzGMZQXsdHmaqkN3ZfAsIn1q0Jkbi1eJ2FHEMC/cfruCOyRfQ48
O8zX8PEt/pEnrDrgFkLGGJpsEf6mV0UDHfQrDLlPn9E5MG9kEAbLUat6nXq5eWrLBLSjXPJ7g4cl
ZYvXE1BhCGkHYdFRF0nYpJWp1VvF55JYykGcY4+fB4jpgUlzpAQRffJEe6hnbDKUwfdtpMUXoh1Z
+H9eQuLGkZSuEPxV2NoK2tRiLjQZOOM/sJFfIRlQ5sqvJt7zUjFij5EBKbFQrGInyODXEMEGdkq5
S9kAsE9344q+wtHKwutYTE7hDgnVVU6qe4476kYzsTXJho10mN0KSvvJNOWWHIFvANNJBLFhYxXq
r2pK5NwR1gcYecHIj4m2Z1snW2OHK7G+qYu/MNoAYAgVCEvsyX1dzi+HmzXwte7oDqKDfvIZOrUF
4C3cQh4FTKuLnQMMkbGAgzX0LoPDBJqjLX1JCeyzoLpC+PKxyMVGpyjydD3LJp1Qr9yur4wzJiv1
/fLGZ187m7/pzGVlJRSt0rdyN6PhdMsXKzNBEoa3fxd+d8O4h4dIuqS7tHZ+7AJqStevHiNmeJJz
LmpNzFAd4eFgi4xXkHCLNStfMbWgipt4r+JMIMKChlQLYoQfXaqQcsdkOzxJxuvJ+ja4lYDQoD+i
k+YFQDoSv7NLBqnUVAInjf5wqK1SBI9McM9yIjVMvjv81iVTYp4CfWF7HNkTh7onYlfrJNhXMUM2
7rUJPHLHSukj0CXKmX+P4AjuXjB8fKU4BXlfEzkK51J+j97MXna+IvJn73Z1fdB//mqbYu4KhTD4
PalNNmYxVpqvljD/mp0hAmgkfJ/j1ehptFifSxctC20sjn3PtjAsCWuFt30S16+9baXrrq9OtyiV
g9d/zVWwk1wWwAN/W7GfsvKX4vRt8okZm0EF3jJd3kQaJbfLbEuW7OeThQ4vnWHfi9se1FLaRTxo
d7loclgiCMpCFmiMm1+TfJxZKkULMQyTUAFZkQbT0mzYwaMLmGdsNZTBKEQvYahZHBAz75TLvyLU
ldAzp/m8w7rye0VcHR08ns/LGfCerqvrFmGZyEGeaj85Zy7XTvIwV70fVSaJDGx9x2p7+HdcnFbf
SNBxT7t/W8bUi6VGvsfQutHhweshFE9Vs2fkaj8E+m+c2l+o7G79Q2iz/P80P3QH4DSJoHABLE7X
ol70nnrl7L0QPQ2GtxC1Eti0G7abYXwSCKfVHX67UgvvCFgTW9w6aKmdleI7tggezLpOBQlRJ5LU
8LOfaLyujiB4pjQEJRU8ctU49WATSwyzBw9QpGuJ51VZY6QL/mcG4XmJWlszed1+NKGItBrTnvUL
rkOJBV5KKruCL4rIT6sZYy8XXqiWPKk6cRZTPGkyxQiLHeBwLmP/KIlXKsJsP5O368GtAlbpDQT2
FFVQH8WM7qSvrp0L+fKxN4SApAJ3GXGCnB4u7JnnqEUR3WQy+zOeCz0f/9FgpOplRG2QajsifXxQ
UNIQi9tCJmGnE24ns2rRqytwqSCnhU3iUSZAxjAWhxw+X2m9dUjj/2SW7CxSo5j1RwrTlNBiPHi5
Y8uD5q9Br7AMkACx0rKQ0QPtYytHwp9uOhHzaI7y6Lqx9SlDkIPJGHedtus3/eX5oUIE0VG+JZ0F
o2ZNaCE0TAx9T2OtdfFlP5IihabqtIjGaeEXvHsH9GTvx633Jx5J8hKPatb88nLfPbCEDtQ++1l2
jHajuNMjLtM8D6/6XvhkMaXTXgUWEbacxTwUh9wRcnASummmJS003bmw3NIZh01S4yh2XgwZajqM
laZzOh8HbITY4/QV1oHgpzOHNYtmgPwH7lT0xRnvCNcYUtGyNTGn7J1vg6JmhO4uzC1U8FhmP7dY
mnyS61/yIUk4uPgwu6QeF80x7OzeV65uhUwWNJse2x7VHKYs07VniOdcZaDPErKoa7fxYa4IzKKf
bFBs1Dkha82khgqxtADRcI0oIhL0QLJeM1WLezlSuQeONyQV2j1w4EkWa5ldJH7PHa9ijoy6tsU6
p7DxfnfKHKTHqaMvFm0Stopp6Sm+joO+Gf86cqkNOkHwpBIE6L21zOO/qHF/cbiS++Z3as7WTTmw
R+GuV2QrgqtVJbAiXRbGNwsmGwjc95A1DRH0stw9APb4CTSXwg4Jx8okOc5Sy7ApziJtcT5luUvG
4jti89KMYVzXNXSKYookH5RgTetNcILTckekrzvzuLzwjdEkUhJxL2SxSR8r3qIYfnd2DIWr41L8
8TBODxN0T1g0t9YbUybSUUwiBf7A7hPjy8QE8uWK60dbi4kRb/OKYC+NpZTuhBb0Wj2lCRPNaUjs
eoEwAOe1HgyUU7InH0R3Z6+nhUnmb8ofckHQ/kKcOHzQW5D1eqLPBO2BpBxvtGTZ2esQPr1oyhCO
xq2dOy4vv6vTektpF2doK+QU5B2edncO5XZfA0H6g/cxiUiIaQynTbZ2UbZ/N5yEzOl4toPuQ070
h6Zkkps1oscNAVE1o0sHiBSS/mz/x/6kM2/KTyIgEnXKLKBCpDlQ6E0fwfz4t94mE/ke/hJ1zhjv
CabomTlDabJq1Y+Y9PTITZx2vAQR7sMwjXJ3z3795FPAdgXUjBuHRHPzMd44mYzbMRXYU2gPMEZh
ydbsqmc+x0C3cCVPIwonw/TFIQlsrl6/5QnLgcC7FxPeC6joeg8HR77jpbzlbZ/YSox3k2yznjFd
JHTi7+/m+Y98ExSw5egIo9NyhdvibYQTqtDF+l48ennI2Jn2ZKxwt7imqy0EJqLcA0D3/2lv3/Q6
6yNEHPCqovdplG9BN+xBmkJeeZfOMGd6w81MFcf8zpuHMcoenZet12vuWRE5zdFEsMzkfuf/Moxz
Bo8iwSST35mqGrx9XXH9GNZYXhWhsWpAa6uUr6Ndaf/P7tJEUC7apRHzWXeZj+kKC4Dgrg3w0cd2
dT6Nye9ou86vGFCVvefI6elg6W4pRdEZP1vOJ8PlZVbpeGT3emBRu0877fihWGmHRh8yo+zpTaYn
fUqyxyFt4IETgBqS+FBPWbX/3/OqXYXiPLybVDtqxnBFB0YbBWIrlHqWaVf0FtzC+w/71u0u2Gvo
5JJaBpWL/TsoerXN/ltdeKrC3rSyb/S8MZPNfekI7kAEHPfl0nS07Zxr02AN9jATgvT/BpECvL4C
j6W+0kzF3DHnfs5hLz9lmP28qX/GaApDVm6ijJlmbfo1/8DZYyZNCt3SRtAyH6CmmoWlAe0G5M3k
Kf+w7bQ+e0EYVlAjWxB+wrZZfxrG7K6btUf6/M0gdOfp8MCkkPduhoCoNtr3KTlAz3+3rvEJGFLy
RdNPcTnoncjR4IOwZjYbgG9VpDL2fUcW9bEF0arLm5NWDZ0f6VIKADynR8CKJk82Lt4Q44MwC5sT
udqjT4aLjdix6fHjBOJlVh6I7dNwnNZB5XC0rOID0rZfzue0zk+L4+WgjtLEr5bbHm34jgYAG3+V
oaBt40YHYPrN6j5xnqHWhUXOqJkhydYfV2fp42Pv3VmsDoZ2TIV9kr+ZVDN9UQMniAdbIuK0wsw1
xw9BWG2ipnmG5A3d1Sd2wZimgwTVvop0Tmi3RkiWGJASpiZk4l9maH8hhGLR/D0mih+T0gMrzQYd
QmMubdiPFRSzf4ov8IMdyIx2Btw0U9/H4OZHPEM8mxB3HBjIEPhd1zE81+wvCC00+e9+YvxpJ+2z
iUVk54emf/eFcZERLjTFU+cY44NklrFKXZAAmDRKeKcAvGqOcUwp7BifIrDZdHfKg0n5hwQ4VE9K
KHl/55E7bBLkY3ut+XZhqK+vGKPIF+3iS0cG8OQRg6COJRXC5FcGDkQ7NmbCl0Uwb0EwtZC67Fzz
3N7YvqmYPjsPnivgIR2SNRaS0ptRWEz1zHhExKPtW+mMg9mvf0l/aq/gQtGW+tdPyF999zDXABXH
WxbSY5HtBMmUtjKYa1kta5ARdvrAOskt5UmlpPm1xuOBwOxDtjMZ5+C1ceo6+6ZISHy+Ou0sr+85
lzlScd1VXQsz8cq3NMVqh+SrBeXIM4cSaaWcGqpNsVCPQXFEIzdK20SkB461d68da2xwovJLaZ9d
jtRAmBKQnB5UUi/fpKiF2iv1UKY4xOxl4T+fgBTNdDVgcbUaK/sz4JMCVihMSMGYsBCYWElE/57q
WaGULlEaxaq1jt2pB3HF31tXFOkHXFQVNabVd+5vsgauuqGlahulrbittfWWbPDqkL7+u2EovSTT
xvI2Ury3f22UyMPRXL+0pjEoKtIdFiObJrM3yHuRp5Hkw3sFlOmqQ/R8BcU5dqptyvBbBeRKDiUC
r59LFMU2a24zQxcfTqedx0kDI3hx4Q5LE0kUKJ7Y45KXHPFNH2iRf7yJRSV7NYhJA6nM7y3StfnT
3oUaieKs/dwGlbQDApwLR4RQTpwBRlv3KLDT4QLSjbVRVSRiz94NL6+AugaplCPHTizk33RHM/k5
0Fy3c9hyS8lXGSmp69H+qnoymOkHFjzlAhm9J80TN+XGHjTnhVLzF9tvfhj2qe0SO8E2r64dXlit
+Am/fRKzWCBvXCxHFCer9sixShBrT4LpXR5bCDpsSmH1wdRpvzQAWI20mJVzPkhgjDPJUiXcvyfZ
QecFllk9PmjDikXuiv/czL1Ki3++St9+Ykkkacj8c2WFgaRGXYvxpgZ2zgk+ns1jz3Bn011FAUMu
73eex0Zs7Dz9XrSaSDEbWixBGF2CysbjuNjiskTympZI8aDITKZ4M0x7e+sqlXfR1qW3aph+Zpqh
gqmU0sIxZmKpU7CpCaROF4bZzQIdhJUTof4F14OTxgtUWe32I91TluTg3wkLd8pO5Y8FHf/UpOns
U9oTRq99+A/UIn2oZ7EDJRwIzJOcKk01XnaRfMaRIkKaGfn0XTQs9kT77e3Tzh6btmaxBiTXfuUr
mEW0ibSRtvJVQ2K3bBvRc0augB2KcSqqPx9oaDug6B0YYUC+kjt+/CEe0PgHKHy64T++DGVAx1Rv
60YemKZDUwYIehUNYiltQISi0vcYJWD8vfqfXf+Ewm9zO8sP+/HfhUY7UAmtp0Ai1gcyPCvOK26m
ODvnuI5VUDydWzHFlqg4j0fpAVdsvL6/xHj9B5DgpWS2+b0bqll2g7pFyQm4+E0omDusy3vHOTeS
+Dzj5j/a2bHb5ocXyk98JziBCvB+/BiXUx4EKMzngCfwqfT4g6qB7p2wXM0xc5pYRDn3uqwMTq2G
df5FEqtohqrC3LHh5KoypFfMJF++mjq4tjyMsRK1e61rYlGYxUoxy3WoOQxK2VsumNBWFTQqqRFa
biz+WYdLWpsCqv5cYp/HVKHBXUgyfEduvNB3CynoBONnQSWfbpmKSB4Fy5/wIECa7TNgtoB8Hxm6
HNOM0GfNipLae2cn141hLxV9rUFM2UjHSymMByi9C2JjUiY5NH0EFuNAbsiDQbkjGFg/vC8cJcCw
6F1NvqrEpmcqz2U8k2GSea/RCnIrzlxDur4HNYimvB6MECbFoVZkxP9zF/TL+RSzKSCPW6CLx30n
MxpxA1eqPvkdjsvDUXs63raclhvKNTW8TDfgn3BafW59WupbXDsvt7pGuT4GicZIRyF1HAfVMBMV
NKSR9sCsnUaMQgWYHoBmFfTQ921WB3lRq51frWek3y7Oy304ZzMii8HpRgk3pWmtL52r0vVN5Bej
SEgKbpU5kCmQZt6sj0sHJB1XtWfXAQ18+u62LkLabvOya4Cz0bqzFj5RncXgw14/9pnMruvQdNSo
iQIIZc+nQI1iaHC7OCQdOrnV7vLrkswslmTPWKKjLxMvB6NQD5jidwEpdkDAhKMJuH/0p12nTfWN
25AP/OjaSvOcvSf5dPKribgGHIHucbsuI/UTpczx8bPadrQI42UVh/8W1rb9Alyv5EGmkM5VJddw
OjYbTQeBFj33VrdU2kaZ8oRrlrtpcbPifIF0g0UKaSzOhd3AOjfnYDKEW3o3oaDORQP1O3dtlRzM
4K1z5A0M/WpmtLmf4w4kGGJbR+kIOwpZCuX+n1zUzjWxOh7/cFtOOIXmySFc0dcULkhdzonPn+Mf
p/+dIjFZsxSTDXIPpT4+5d4MmpKprhXKh5TmXxDzhBXBCL9uruNH3/saiiYgyoZvyfn1r7H1thDu
QsgkWMQbzwSaRAscyKRdLwCC106k50ZcbSNGC+JzECgB/Hsi7MtJoKjCTjTW0W3Dbh1TsKLWzOCt
tBWbgJL9iFnE7kP27NjIgCwuTgDrbmf69WJNRf+1sMpmJ0Lb71QyEzHVCMODj9etvdCdCEjLNMcJ
XNT52XHMwxBm9lbMqe3QFcy/NUYxBzJcsmJF3US39kjUW8NR4AF8QoJLyCrK5bYOPaQcZbFEHbeQ
87ZL16YffFb8aWmUdDE/47qM3jM8pFD4X0NUFU9Aj+IREV6/6oANFE/CtQ2xaRQbaR/Ag79s0fol
YhR7crCr+NYdraeF1X8wzw4Nnr5lX/6dujgWkxogzb6wLBLljCyVQRks98bTyT5k4WQTvvKREKzz
aFiN4SZwdkR1WY0VkZDpzgHch+qo2fPTq+j8Je4jKC2hFpDhsLZsNQKMWT3q4QLnyxccEeSrNW+r
2liLcGFAUn6KB/QSI0lVwIMR84c95njlTXnKqpZchJt5ntUA4juX9h4qWgBEkDGU6jiRF09vTRJi
pxMHdNYJR1IXLyOmxgLRFXln59xa7tez4Qx1yvV0hRwFpUTCXmXRzegWDIWBm2fmzy9+O51BqToD
u2J8iY15yo/Iakxm0yvNCMKK8G3qbPPRC0uT4Hw6pNpNDqoaoGmrQWD+ArwU9jQPdsmfj0qRiVY1
ai+UwUGZZ/6j1faVSDnJOxN9TwlwDLXMMHVdvthZ8SAV6/Qcw57SX3d83fsU5xC6ihg2ZRRWoTjb
rAehOvCwBKwoPDqLsCFBfZGi+hbnLdDEMDJ8gMFtFss+D8UyxcIs9JPFeoOgwTUSs/U2npMchSWx
c6x9kQuRcnykO9jyxtpzYjIjcnW4kYvKaDuaakblO3CAMZ6/75oR6/Zd5HdObNCMSW0iI+nWrCu2
r/XyEmer+BddZf6kgsMvMTXmYfPb0KVbV5BE2Rdqfhp6oygEswAEM5CjzoZ9SzLLSb524HCSnl0K
4mtULs8YAYEDFvMRZtVlALXLuLnCKBXnuv7HWn+n/3k5KX5kKNob7UcJQ3o/NggR7cnWPdbFCjb2
fr1yXLAtYczBK5A38HYuUDHWH8jl6a1TiDWSAoaWy8echlrcn4y8lc2G5v7L2RL7ipALiOyWyj2o
9fvI5ZFlOaj1/FhE9tpHuIZskM1TZ1UtBLEpXEPOilFDFTZH0yR9LJaBJoAY+4699oT0vjF+5Yy3
Cs+cMb3TV4oYu10X94agwbuBX1I4NvBC37HmHbXLrvGPOZb+h2RtPN6jjbw9OjP3aZjBsybp3SX4
xtq8PNFuDPijLrHnJqPbiVkYchbno3Q9uW4eV5OYBiKAhX3Tg5SRCd3bSmidsvtDo6uZBaS2Z0HJ
3aDUjbF5/XZXZyvoBgfWhXKSd9IPECyj6srOGX6cZfv1KRqZ1PqfxkkmJsUlivOuDyGqTsLxSpgc
1NdkLuVRQfjIfE8j07lk19rEocw+koiLdpTq2uZaOL67WFqYvRzxkR7L+1ci8W8OiasZc6/M9kf7
QA0b2Brrbctdcq8RbtK6qtL3nmBHgMfyqLfmL6BDxZADD0II5/jzkxY4o7/9CFhEVRNb7d67I5qc
YYKuYWoaDR3Xmq02K+Iugev0HTEvQjescnmdQr7Qk+PaKE0h/e+FnLfl0/ZdKA1QA35NgtWA+bMw
y87cioiOD4Q2I2sxec/AqoccX1fwQIIOJng/9obduGEo/3GAGqTGlCiTuho51k9qPMvradzoGKrJ
igK07VztdwPepE00a+BaryMLzt2nGIz2qzRt07hYHbipV87lB6EuKXHHimau5g7i38EExom6V9FH
T+4/Diye9+J/sEwnCFTYpy6HYaZsKX49GuikNlRm6yscCktxBr9pxKwf+B9ZLwfYDoa1VZJ85k2h
dL2pQCUlU8BNmOSI+FJSnUgp6b4RRtLLGXp+g6tCCS9w/22r1xTDcTgHfevXsYGDgAl297kfaJxv
yTQDslasN+e7wL6jq6bJR5yhCa6tKpnCf3QgQ8B0ibZVaRXd2z91vk5F9opf4k62WwFqjqhX3hkG
QspZUmD/Wie9tTtbHaRO7u7HEWQaIPmdnWGVEtENTw+ceNs1ta/jGH8lCYq2nJmJA5vP8lvmabab
YbG84T3ThPb2svlXcrXaAnke2qwERFP45TC7QAEzmjaHhLsjLFkB5PpnKQNs0M/VWoOxt48tfHMd
W3QChqktPiczAffOOXGSSTWZ1G+dTldoCaGBYBbaONFbe13Zab5tZTY4sdL1qfGAL8NP2RjZ9rhG
pC/SxKE4pvHYNKuDAl2eVb5ergi3KZs3jTbuh58tRYP/X5heogS5Xr97mOgvJmTQz+Avri/Cq1Ib
+3dLLwXAif40fRKEI+gwaMHhpKFLhYf3y0fx3t0PPlhA14qYpkOlibzllJMaGhXPqG7C4bmWZMaj
0azUfGSOlXsJtwrAiJvUnd/51YDIcIYXvzblFtVnnG/DR1YvHnNv3wQJX4JvqoC8JvvUtRBo//uF
GSaoEVbM+2AzTAUYFBjIqLaJaJDhwRz2c+d0oHHRouOsZOrSvB/g++A41hGV3wfYsrM9cr3ZoSXJ
8okFsJz+1IQEIhr7ktKvTvjNep8/7pnW7jPpVXgn6NX6ewOJUW+akm530bIQnOTHaxO8TnCHzagj
GFsuW4tQdnulNH8jY39EdYWYOROgAKIrnFXXQ1o4OtdxYUlO14Uu0PNCmn55h3STn/M6Lf+r93oi
NOH7uAfLHHD5PbqeJOGKPTHzskQLF+GzLHcwPZNgSgFyGxEo1vual3GJhw7EH9VqIRO/JPaBTMi4
afpowVGPKiau5Dff/Z0CIgjKcpuQ/zxFSm6taRu4WCbQ0x+MrwTOnENNVXLbENpXJOW0/VEWUj60
PIpVkx6ceyvMR+TdnOTurlVmmcU1Ruu3WPE84/GYfnYa5aW0F9InZDuScNMqoP+D+Z2PGVljb+x7
ZEN6MniMvlKzMfJLx/pnwAxrmxn+JMWPaW8jPN8UbZFY5UCF25N73O1qBQoCXFOaQVSiAtIA4b/r
vVpymRuQGs1Mcnon/m0Km3tf/cNp6ml2Hnxw7hE+itSlHjqwWfXLo0Nc2T1sZ7I0NMUcVxBdqYSg
nvzOeACTTeYaJivCUJlfFQthtJ6LXU85wUx+o2YxzOTxvQBNV7IraUzuDWr6/sV1YjF0NiikzJsK
r3UWNg5wKzDDPIbAmo3LLpJBEbPxGTkmkRFUl96J+LPHwQGHlr/E2lJy2NDT4ux5VUNFvaZ81jax
OTRVxzKAqUr5VIjFTJdv7ggMtDHOrhpKGD8WIo8q9sgCSg5D0RK483JIOojfanTebmgzUBQcpZp8
95aHGbM8D5XEWOL8/sjxTUW/jOxCzD2KLdiCfSrXu87StTighVxFGhWPgNnWqzaZnn8P7CN6Boe8
j5+ttpFDct5irnAqWXPEObGKo4f96R6Dhb3qafNZJwAQED7Dgu9g0DNpOAByHjDgJl8RcKDk0Nku
LUfl0kthuASy8CobkVv+j+kCNhc0aMxhbIsWVugBRBuYv3CV+3O9jx7DOmeX0EiWBkIdCC2ayRk0
5ABGWR0XEZZOUVaBm4PRvwX2Zp46t/rfXcTV3n6a8+hOA26A37/Zns/gfAZizu0kufcsY3aR1G+q
un0pxN8hgBw4fxItXxn3pCoXDzgSwaLRyOum+tY9B8YVhIyD7huMWQa809VcQoNRzJuIikK3c/q+
gOn8nuq0bkLKcDe5tZjZsMXLvXhudQiIuV4XMgLbCK1v/jEia18HoibR2I3GwtEbELppiyNu5vNM
3rrkg745EfJ8McfBB1+dmstBTXECmP5uFQKVZZQSVi/aO0/qgPVY2+irxOsU2T/7ql0jBZndcx7I
JoFcojjYQ6LF/4bQFAjUfWKpMoInuTijx/j6dO+pYcxfcbfjzJlRnsMtp0iQcOUwhNO6PgSO0uZ4
jUJZ2jpMJtybSupt2MM3v0CkIiHt4wKjRA28nn3PYgpvsqcsTDeMEC+1VudlIRRh46PJjXpRHjUR
wNJHa/LCQAGVppmw1P5M7o0JN0i3YgoCFXWwQWNyj6Rn6MQsQ1lIxsGNIeN/bjaf51opKbsYve64
B+zSaRHf57H8UxMmV9upSC0ATAqu4wduINwrtp6la2hr3nTrxHhffhrdxbudbXGfR+p2Hfmloz5A
QKGrrLB0LymA/2Tce/TVB4Fjkrg3KygLAodHY512dYKoqRCSPxEdEe8YNj3VCp1hbV+Fy0K3zYIQ
7kpBZHGbhO6qC4mLhHIyemMTvNYHnShc0/eNV8Ria8mZccceLna6ZaU4HqigehLMbPihA3pCJUWz
taNfG0ORrBGBXjKsv4Scmcs5lbftZYVtUd5kEOEHMsR/wc/ls4oN7byt3Oc8+OEaXcwS8dBVkiYK
JyEBZUf96FZzp2nkf+PyIZbdrENgaFQkvEhQlOZNt/xJz+glKYsCadQMqD5HH7+a+lXsWQ2s0ydu
c6/0pOHDsdo7ajOmwjnVRAU0Mf2QvOcTUzz+li5WLmS1KgLyP1uEoPjh5r+ILSTHhcEoKJ1up0iI
SlVXZatYfmlipBWNjcWXpM4Fb6JAG9HLP4e5ndjPnM7c+LyH7ESRZBkfv8TWW4adWFqQiBxVXE2R
jnwAG2QezoVsT9DvWAp2h25hs2V/Gc/hnoKuFOfl7vXZ6CUS2pD/pXn+MNEXFPTlagDVX1fLfgO3
W+aWmkxk2cZKa3aNY28F4Rf+KhaG/m7oSMAaTyn1t8b2q6F5T6Y4cY6UjHNT9pcTCZ8Qf/DqPmJR
mG7ahx2rEFECT+zFBVHX719PeCOJElb+FEhwc3zjnYHe2BCe4ZU11qtA8T4z0dlBBFkeO4eHFi7q
pXURdGY11uzKuFBlE7jhzYfB6r18fRIwesZtNm1nFmlE6O+eTRx4/JDiReJKjJO3GcF7oFCRI/2k
kkZibSt1cl7wThhGyJgKhdzPsvF3wDTHMd0BD97C0wMN/LiMZPDE4DMdVO4vvIOcN9cY3KggO8xy
Pc1mp0oaTam1hN0sY8SDkpxfXFi3TOmsjE8GWoNKfzN3GrSWP662H0tO4AIvyWJdI4PXRahoilil
HxMzduk9VjozTNORXlkHkiY6Qo2Hgq8BLB2FODlLs9gta6KjTCOrxDa2OcahVjLh0G1TI2bJGQg7
GVGGK9ylDfkX5v4OQmxR37nPhKPGG9QU4WakxcKuCt4Ug+lplvSHYCGNLh2AxxBYsLNGFI27VXYH
iHCCpm6s3VW2pj7IFlBhvPQn7vplcaskYsPN/pUA2ZitUraU2Hm8BJPdACXExRHIR0AsHC4s64/n
D+FGa65v//iFJumDRi21UcI2IJfgNFzu0LRMAyhAnJ0g0VWC5Ka5XLAvWPZrsDUekWR4rmMiLcUO
bhFhTfKD/52WQ03GSu4vPlSYe6alZ6EMHbHWMUd7ZPX/k5tBoHuNHTWUzB+HC7r/m4l/q1r5ud8v
mnzCNjqAhOX6e+7dymBKwMRS5N0ifcSYQ/Wxp+ysskuPcmkiOQwwwXKXuBbkx9efGvmdlbWXB+Mi
7pZLEZ7kxugTcSWWsh3lFMvYpqH1SNRS2LtOWMT0oFWxOZd+yeI0pJCS9D9R13GDluBo1AtB5R0/
w84QXGnbUTnKgMKzyA7C6VlXI+WsfN5jON7OCTJVzsdPUSo5hpXM4aCQumwn89snWoUlHHeKkho9
3pdf5i+iwoYwS8t4V8c0OUS6OYhC8KFzPEhHxteD/W5s7h3dqeOUxMh9kb1qTVTl2I1Oeg+tqWSQ
nzV59brnoUWVTYqlbbLnA2ahWmy96zJ5gGfBio4tXGYbzdXeo5g9de1DxljluoNcypPC/mR0BMPE
EPeVsR9PqzN7YWuV/fIZbwWLqyOcIruxpE5NoCruQNrSuuB5s7Gj1J4qv6wB76F35CAEyd3KrGRf
Xa6bvpDNl0ht8lWe2YKUT4f7vn/uqtgu9DXqutdHEAicWrRgWdp3PU+nws6AX7vqHjy4pw01GtpJ
Z6QakTNu3vMXGWLEf/WtFXLlS9aunItnaoYQ0AK5VZVuDA/vposSg3rbK18R/vE7AkK5ISmeRQVT
1bovHwdKczdiPQ+2D86xKzV+ae5lSK3InYbhwOEGTyOKodB9LSLyHKuV2e1R2tUmknJdiyp5S3O+
NcEPs53UXm/haM5PgQeaZvEhHUn9AVd9G08Vu1EPv/O5R15uKAoztg/o35nHbokJI9tZHuObtWy2
gH2ZHevOXm/J/HWLewkJy3U0nl7+0IyxSyNK/dgoiZ4jrc5/GlsyUT4XoUBmDyWG72h7bvIBz4ci
4Jf1p0Q/3mCKznzGhRp2HAipx5aUjb5diDYAFa5/vVWydU6tyikaENkWzijyQNk/F997DdLnHnlk
l0lqnkwoFt7AZ0LBqRFmOn3tMTgn+axz3skJREss0Wbz03+XRC2Y4ay/jRgElwZjYz5LvzyaGdZs
/qp7L8d3A021UovT2wmiYT+kuJd+vgmsrdXtrx5uR3bkroy+sYSTTl+bGq9AoSspM5rxfILI5Vjc
+4EGEYWZ2moZbXWSpuVrFToppSJy5+9/ZCBruRIfoUP7tiVn2u/ZTDmbPwLiFoICxAE6898hItIS
L5FK5skl3btVUb5xRM7GjLPWhDvTh0NwhiXgbnAciE5Nt3P6HLjbrqDE1b7d4pn8DZPXRILg8EE/
djVEb8Gv1i1BYzzd2w/Xo8LTHYbeiwPmBhIJsysj5ij3BCOfqeWOvjWGVQAmFhHmgIlavChmHpqa
6+bWGMpQ1g+WUxLL6GW53/WVpY1q2wmr7tgPRUb4JWbBGe+TJtsm/UGMwrrqUIxdb+MhuCeRStpx
y3BAeRvRfH/1rfemGd7uLbMUS/kld8s+zxzJXpFEIIbMpryEEHRzDqYAiSbh2VWHvjF3FrDvW/IA
GaCXEnQXUIX29Zz1qc7TDpkB7/qKlkbT+zpWPrUknstzPXrSzG8Q3f4iBYngsUvq272h5aynq82p
7ND583lRZB88oHZcu2Z/dP3kKETyKvroK5n9l7qqEhxz3rrwPocj1CcDDW6sNkmRDz3L8+aAJ3U8
T7lNl07N/1wm4pa05FoUVzr1aVdicGXukGxgSrcwisl5L8pYDshIUN5P8pMHgUEtWSF5N49YmDO6
yVBDxY79AhixOQLT5Rz/IHkyKCD/wXdHUuMOE+6NMZWmB6DZUI3wcK2qSi/uCcjwJ3k5JtXeGDxK
JoNb0WfZ1PYrSK2BQecxh7EkQbQvsFD4pw5BSRiQMVaxcf95MuLHf7o0Ofgvqtdtxm44DUMtelMY
oK58XzCQ689OQ6CyGE/RsBy4mikib6LTa6oPumjL45yZ+8khSvD+n/3BUz2282xn58LeI4SaQQTW
+rhI+n/qxhbSoEs66zymFR1aX91cR3SI+MzdoT+GwhFxQm6C1OzBFucZfLGPaTIdgEe4MXm7PnDy
mjfL5/fGNT4JraSFV9+gfguJw7XfvuZgtel9IQ+4QuGthlaRT5LWp9ITKpKDjd7xPbmKOJj0qEKR
CoDsHzgMn4hgAZoH9sRG5bDgr+oRz4d/FjBowYjF7J7c9iN/MT77ZyzKNphqneWxfcEAIc1sNLTi
RkRDs3QexOANruz/7Q+GSrvjMgxrMyr9LOkuwBXS44sWOZJXEB0nYUKl0PpPyNjL92zJfVbrhYFa
OySozoStL13+QAORdxrkM4uDrGNii+VVuPYV5AbStEWQWTfo2zhr+1510iC8LJocqXex7UjdKU7A
5zNKoFz2RJ3PxfQLXDLeJ5tuZ5L2Jp2aSo2/Vf2fRqhnU0cUases6fnGjVt0cjBNlU+TZ+laKuF7
DSOs6xm1DuJW2TQG+KIsL+GmetTRVrSDwjLjEFUJ4LyWr3qzAtSgu4XAN7/EzQOdJ5a5XvFxcAbm
J97AmxNZKOJeTajLOO7kRJ6wFILH8zgPPuVZP54BUhY4vcuYQQhJ5b2rpdqa/VSDKCptzpBSS5ke
ksM/etunVuNcoyQ+GhsFYPlFaSIRlRg5f66yvH0eTlRxHSJbFeueuuX3gCJRucEamJZeuMi/Kmyu
QoQ33AOGG7BFouuIR/5vO6UGUOADejsct19MLiEnkW/cH8tF0ocSPcxetPrhMQ4W+77U0BBwId3u
mKjj806StXHgy1xu0tD0tFOMfAVlfZtEAaS5/dzEdigg09sQAtquWHtHN6XR/79w7a5o5sSiii02
DLCm1Q3BbXfywslW541atSoqmoW/l23yidBXz9HRNgjFOHTmVnHeHZlUK1iVriaO1uxhsrE0zdOr
HeRwUuRkGpPwzW5Ibnw132gLNByaV4k/MvxNOHC4zl3mxvxsxNUbGw+uWGYlCmYplBb/EwJXbDun
3BAeaftYU7TkApwzjHiUYZF+1jBvf0F6kJk4unUXMKifXSR2fRo1lmnd7jO83CJ/zIIleMSsBNl3
BeFd9tNEtyHKxYa7YEnr6OxCY+LzoB7AelayxrTW+RMPDT7+nKWscuUoZ/PDf+y7zsJtxQtKgCOx
gC+l2DDlN6do+zma/SaZu4U4Ss6joZAOqMnDHt4sJOkE/ML1M+4ZJsyEqh88nNztchMQ88pCpNu9
NSCTd0OUI3w5m4jbbhroMkynygMWItVZ1BPdRZk5Vv9hjT7JARATQAXx2HM/1dl6+RwweuquS7bZ
RPyuY7glRzyt2A3nbZ3FAyrE1v0ab4fRuTxEwB2tSspICgikUldM+tgaJpa1AsKaWQhiT5kS1Nsc
AHWg+8hA2bXfzyAwsL4l994ZaQb0wi2PRq1kevXjaeygRafKNWXrVlqcB/BYjIZ9Hng8Rt0LDa1Q
AVSVH8biKDEc6ipK7GhNLN12qLV6RPr1B4xInEtTJ7qZtAqQYLeuRXRtfYCjMXpiQs/PWXL/uWIk
Uj+YN21Pk0qU9qKMD/oo1Ux5p2Yg5KCQuO44UlyAXno5JOPu1EZDl43MhIBr41pnSc7k5//E+Co3
sRdlmHCtsgrGrQlloES/sxYBL0zEQANAXeQRys08U3pre5ZSmJ4Ms6CWEDvgGTUdiCMClVw4xWYa
TkxqaO4J0yAbwbyMySZjn8c+/D9l68PbRH59/x8VH7WAUmMWx6qjrxSDqlgguJkiNpYc/rYCyfqV
4d9dyLbd/5fgI56IIGSjq8Ib/MJEK7tl9R6sVcXvFUwzQA97SjYe8skoitn0o1Qjt6yKgvX6LwLA
2AW/vctn9qKMteHnC844dtKkJenoSyuDwZps5fmDvwc17u+s6gDHcrVHpd29wMKbZPq7FoWBOnmE
lzM3TEwaagyjHzmKJSqheI0BW2ovAzNhtI3Bqsk4IVb1cKBr7TAf5SU347BJrFRPf+kXbbsCpDaE
XS3hPCG8vUM+hJ84yeHolte5AaN+GUj4NiGidI6nVpb7IlOeEdxPY4h32jZryAYN2CVQfzZLOJwW
AC6WpifThVPkQLnL8kQ9OPTtziG6UVtrxPCteHy1/IjKY6Qu7J1CpqT3JjM2NIy+Ah1sFSCM3MqF
M/1xJkPN9X5uLiQhXP10ZrhhnQiF2T71rd3CvD5AiKS2U4h7h/ZsXwN39+TcoJnmjYNvMsAMBEzg
w9A+CkAyHfg6EgmQXLkmgWCcBKOnmxtNMwR+C9wZe3Un2D5K4aaNKLKlzyqkNz8rvjfxQkIbVzXX
ZWVhQcuViAR2A3paAh7YORYCG0XJpqY+usmOl004s6B7zu3qG9wTl2FAGLVkrP/h6rleBiZAh0jF
sOOFahR+3h3dRJqbKATKhCOf3DeaCKAnbnRZu8Y6B+8UdGeBPpOjb9C2PYaGj9CIWIqq1Ds+r3sv
C3QceKTrT1nr2tI/O6IofHngfbEShkaO1QOA710tvHW+WBiDYi1zhApHlb89rhufiHcUsOhMOFtH
EICLIn3mP7WIEQKKuG42v55imLgMxMwU0vdMoGs7bzLmKr1phbim4ShCPxzeypyxgqIDrG8dHaRm
poYkoZE0/SYdXqt/RFdt5+TwleUiDa6Wg2ocfes+PjBrECgNcMU69kXr5rVC8z6oXu5kRk5xXamK
vA6irNi3y7XTid2+Qr8FwHHjOn+v+SXcpI4Fj3bqCfDKiAJp5H2Nsy4ouPJCO59RBSznlbVXFYjh
rwi9EvRJA2SMnQs7v2HLcV8pKBoUY2msX8+9O+9Vd0E2bVj5Z3Mz6GrctZC7G2rWHIPEICtho14W
HaJ/7OV1C1Z4c7feiMdmkhvk2d6Cbr8V88uFmgE3SW3py3s8CJORtzWULKqHSgBtcXIAQ0bT5GX1
NrFED/6fdR6mCzq4AY+cjfowPrWunFeRWdWvEEgQbg3WVGrPBIBGxmya7L2tM3r2N3wmjtv7HBAi
mFQSe+yEWX91RzNQ/kzE73Nkspi/nVKFIZD4sR6bJrUjpZEq6hqzsjPALYnkAMD5Ic3XwOs1utG0
pFgZsI5PJrji5NqOx5TSmd1gWJRt59ws9BQt+s6MjJ0+zX77/iea57UeKWFwHqJ6K9gOyvZIdWg7
Tp0MmJMIx+JW53wJF9NA6W7Q5wiqgPN+jaPdvzaNqDeErfncu9TGUMqpsmsq4DTdwnHDQYEitIx9
1MdtGLN76VHvXyp00Nk/iKqNIDrTOigPVYoYZc7b/IXhmGD8FtMxKj6de5IsabLrF2znRatO//KF
VTpZl3Qpc23R8rVpJeA5P2lUgk5Snvn4eN5F66oJcICllVj+cuP7ZSLlJSIwJL8JalsZgalDLzjX
7LBABIJbupAo8r/Jdx1U2WvBWlG2Z/jE3ZqnVucCBoidxMyxK6ad2BsoCcND+1qNTzgBiKoGa6hX
XmvBOMXLkk6FPzEJqogExsBpUhisO22/OwihIYy7Ur2NmfBG18yepIQhzQvpK4T9z9fVKvUoGd90
No1AdGELI7xeDhTQCa4TNVbEE+Tw70dCNkAi/LtiHohKdh0845uICAb6Stase1KUw6y7lLjD2ZMh
bLzIGhfZVgVnFV+V1ROo0OMpGmc1f4Ni2SxIy+eVjY+5Sl9sCxD/DtcgvscSbEWId8FxN1l1D6sa
XRfB77aoK53Z1sNWzsAIfTVtnFK6PIBMWKsvn3rsKPv8UmfqDgPW8+KjzMNkOgYLQQpYlEWXXqi6
6iX+D4ScZuV5xCEiIYhfdWWeKa2az17bpgHx1McKrNN4YNMxRWRlwGvjqodp8QAgP5oItBE4ZzXd
wGf0OJJjhGeMlYSfUJ/A60m5vh37xUEVkBK9d8KzsIi3xXDiGD8e36a3pWRczhxwhwgU2GcGuE9T
Uv7FGPJictqWbO5ifVW+T4rQGTF0hmRd4zWlGpgDRLrHucfATQ1bCDEt/2DLbWQb7KmBYXSMMDRQ
m6cCq2H9NgShqz5ly7SNd2c9tf2q4ZIuyPXbWlqr0OgoapxuhzpBeE8rQ1iFIALT0hRMI06oWq9V
j9koTQtEsc9pGyrCHJSmtfW4yeqj618B1RIwWZWHSniSeol92v0LDqXsxQKlcYoPT+cyfrbtz5zv
o0E5iEZ3g31iiKvGbdI+Um3/FeiGF6d0AHnKnzJY8dT6yj6NMeSUp4UB08reIP7tKq27yZCiqrd4
/iRPjg3GSdQEJpjcVtBy6U8AtxKFX7WZyNoO1GnpkzUEG1PfE4coCwtL4JBNZ0gihcZ2Qdd2Vntc
Q9uGk/bbp0dkOAoB3YQtdWTbv20pBJT82gMPw4TwY2GrcFTUkKYKIIfU4KdyGqqpxhK/wbtCVH7D
xke1ViEK7JTpVWDwcCYNkXFyew3uoqx+EFXOKQlBW4RvdZTGEUAhU56UGNVGVpGAvjUKX0N03ibc
UCbSzL4z5AGiNTsnvU95LZLBJHMQWOoYkyj7RLxG4IkHYMtfSfsYBCivy4FQrNHqbJmgX9tcNh/x
ox0OHlB1ajGOmEAG+1Pylwg5BxOyiHav7FxqXlsuCvMfx0A3peOeF+7N2P0O7UHfNmnzj5KpUSfB
7ym5EmVJDWtkEFcEbimxQEMt9ZPOjSBkj0aOanx5epG1wb2ykntfc3sqkShcPSqf6VdBrk9ENKCr
m9CHysgOSufMlLMBc5u3saz55sHXzdt5qjflX+7rCgTlo1WZM74lCdOx7t7PfzsQ7jRKnyztCL/J
Q1IiNoxtCtWQB7xfrx6/MBKnYEfnje/kdrAxL6KQhWjfF+epv2cBGK+M2BfqaADTUAcmPQzz9O8t
zca3MmOFg9ioE0J1prHDfMlc+QkFDKhs/7qEdVOwgUY98Bnq/MwYROXoNubcek4Ag59eumG+z+6K
NBUFASZ+h+RogtNBTZvh29TJq3WoWiEB5GVvsW2WAPOvlqLcb2Rjd3ajRxt2FbegiXNQNcTAYJLa
D1eobM6HRcLcZJXOEXb8h0e+d/ZxS33EjXOSIqVXTLBTM0xO0GgJ867fsrdgNGd6RZa+tuLOnAqd
llOrtQvYDHoMKfshT4Vx6+0aeJAXrunu7Ax3nYH9tzLSsFpu/zoYbURXVfK2uBAQ74xjQyOdbJIO
3n2uKUU023rpbotjcgRI3sob1dP3F8oDeG6eFH6JLPhC695tcoTPND/uoKY4052GBonYWrH9GKq2
gTR4rSU/maNqiFHME7eKBO3M9teXqN6laMa70Y9vTbPVL1sUKyWkxh/clEfhZCkMGwu1VqiT1wVX
NvnLGu32w9VWFdkI4lrGIlGBjWZ58AeuX8prbFioE1sjDUZ8jSHS928uYzpErQjCBI9KecVajZaZ
83JBdH75jJzIf7cv369Pj3EHxVIR4fXJuLg1g7Re1TU689NfQw7ZJqCQNnSmx2E5wjDpFREBb/QK
c0jMX6sdKHC0YTyRoVZcSb32fqWSUTT0QmTN70vZwF/3cF9DCqw/ZsHF9BVfMwjFmWVHtDjFAFZB
SS3wfOy84i/UTGxmXt8nheMbS+LDX/qcHMlS4QiqAxrelBwnzbXNrxjeLXJkpkPexczrmMVCi3/r
mtU11H0mo7Dazu8kr+CQp9vdW/D7bkZ9S7caOSWwd/EAb+r38zOMOOFRgupixSi/bgR7Gw75/+py
7k9n2G8gD9g30LK/KPjj4QahFIamJdFR2PeUwCsQXpr1sXF2UeO4Xy9kv8OTwN465ECX9zp04KLI
dsKFNZlV7TRWKYiXuL0xhWS51xT9t05uzgsNNBOdrv1QH5XGJ9fBdH9bsK2JWMICTF1Foqb3fEab
pB0Odh8+G0fSUJbcVTJuaZBjhJE7ck2vQ4vXbGHVIN9Qde9b92XO3T2XI+b2eIJJC/BDvbsSkA9H
pO1rjlQTNsM1zELdJF5clHr3iDGcA23WlJS40BRjGayxWPoSbQLHXHPnOcnYxFZi8c1UNgjMWjTC
pJaz/qnwCv5RZN+F731QkgaZk0xJRAp3vrEmIGO5cV6Fiw9I4BZkfkLe6L1+IQl2JD46R4CeVgH4
dAM5z3VgIhUhvgmP36jtUudg6yM1S7nmJ3kk/JcdwtrV2nsCJDKDfmZOrWnvx9knQY/TWMixvRCS
HJ7GcfuEYwFt6WD1rR8Lyixm+TwPIeS9oGwKXQxgp8U7cw7xbkmhQI8UfqbfV+HxXvj28IgxZFZS
KOQEix8ehgHXU+Ro/yZTC0b3LK1ComfEHG7bSuj2jR5O1Y4OeLJHQNiq+bBgFFj0oKXOdu0r/4c3
rvoZRF26i0mBqV+RWl2QMjWcDqulXcRj6to/ASYt0PEsm4L9WUFWAwzmWQJLrBq1VyTbrTwTNkkA
DBJSQXiVFyxE+02i9npqZflgLKlrTH/cJuVFoFRDSLwBkaZePaW5fB/FI8Lulqrh5M0+pUY+r74G
Czcwpd80BMOsmCeoJ0jc+M72ZL3Rzv1O+VIezctmRND4D4IahIZZBG1zGFNGO3wemMrV+CZOGVUY
cL88gg4B+gF5SZdrnn8LCi6FxgcUH+XgCDJQAYSr73xhkg/nGY0B3GiuyIphxQmtnTQclLWI2Oyo
zoaC/O/C3paRhmhckltXNJBXI18tqU168YiuPupldSTXhIJISaS5RhYAf00M3q+l7sA04PMfNXbs
DQiPKJbCbh9L6ZUosxGOgLZaghEQ/09Eb/GshB3nBHHkGkED8v3+ZPII5kyATjTfu8YHNYw2v1D1
U9okY65Mi+Eoo5BLe81KiSz+8hmigVAy+PZBcFmwKdqGy8VXpjIBu4Er7HE3EoHrUZaYvenhIfwb
MwRBidGBxFd/clvGcHdzR3rxfdttHmi2sb5WFfQDjeQ33cXLFA8hqglLbh3TJUOiB4DdkwqAHI4r
06X+zKmv4FGBIn0W7EDr7w/GETVmev9GjspryM/4O1d8KUPRvQU/U8MsDdQpZ8bhZ+aVpoQezo3V
7SN3lxX9p3PilgTf4Mko4Du5IbcdbUgDxX93/pDUWCo2alndaq+JGe2oG2vKcRVs2ROnhtVCtmv0
vs9otGfqfI1JoWkulNbAE1uANEaXW5dRA/WrxD+Ec7i8qOua5onTvnXNiVJPH0lwvMV5be8M9H/4
z2VgJ4A4N+QLdb1lcK/tu5wZ+KkgCaaB/fyvO8Udl1BRJ24rxVkue1UFW2vEfx53rPZ5z1K9VW4c
lUQY2KbJ1uI6JOi3ocSS0HgC+xo8FrVl9wwxXFe7lCH5QqhQ97p/YHONBxa4lEg6oZEzxSJU54iZ
Ub1SIacQYPWBdXR3QzPcUSG2eUDaOA3MVSURaKvpdgT6wYx6rwbpirWwYXQBqzyXQ2hl0EAdShIC
jke7Yy/m0qlpcpg4tRb3ayuXVZQM5iNk8dsZv1Pui3WvIu1xr5VdoSB2yurBjqVOSN8cI7n2V05v
AFo4PWP4p0F2rE/8rbZRJyc5hS0DBZuwCoeRsG8uhytwPoa33IIrkWp4qGX8N07y0eZm/AU5xNMd
L3+5oMJ9p9+eNYnTzu2GxdndQQvzWYexLGMuYIWY20GSxwoklDZPZ+UuDzQe8swQdvzzzgmdBzY4
Dk3Q87trTgjFxTKUhLUKbUGWk5Usn2FW0HyEfIC+9aZGlr3wcNqXZntr8FYaihoO3hpHldXLZuBI
IMT++sdPP3aaxEWug36HcqLO/rPuMMzd3ZigbT70tUnyEeOWIDcHfoKEHm1YIX+un+eY+xtVokBx
Qnv5hNvwDI0c74v5DiTiOimMzuSZqkyLjOxteQHKO+NQQsWcdKqGC97XelYqneaR4rVY8zrIy0wR
KoJcqBpG4JV+6dzVscoYwraIGa5TDwDEXUWUhXrzufkzKbZrFHy22yaxn4zYn3kD8+/NO27f0i7D
LCKZo5S1gT0xUg4Jrc+mlRkAfO1gDh7iQCfEmdz5TimmJIOcSsYg7PPw2grEyIn8aHGsiZr+cm27
kYQxKuL8V9wyt9YO0EDUlEAR/dTNosaUF4McUfDWLxy1+92BpWcA8XusHBfoOV5Jit803WbOFtYh
Tw51zai1im9cwT1F2uALYMHYBGVxIJ5hOMw9qluvZoMSGpHERj0OanymnZvW71TU2AcRJ3cPI/eI
REjchsuNH3DzID+bfr1ryLj81QyfouOfL/Nan9JZcASobhlhd32oFaH4pGJiFWVmSYglm2P1B5yF
R7gtyU0shJhkHhfQCtx+mHrDrN9FGLXwMXnsnGzsKTk266aIJOFhMlE39qWPw4hLfEf/IFKTudUs
2U+W4nVgk5n1LPsbccYZy6eV9MJr6GBakN50U9hmyy3+ZEYCnj52CsYL1g/c+uzVUh4OtzXOpOpo
EY4OA2P+uT2u7LXne/6sYVNpMAQ62pMfqA7KqA+/phpiVaUjXFg/x6so6YmZRcU3S4Q3/GsdGGyS
HmLu3imcpk9SzDAtYG7fEwtZo0NR0d453FUmU/qFlYpZR342B18FIPMb/XpDyGCOsP/IdbmP0h2Z
8uHGEozHKrMLLv+2gfwvSg0371GPh8fTL8nwWCgGcagIaIauRBxV787OEdGBziAUGjMbEK24g14x
VnKIomwv4ieiZH5FdgCHaldWyBPLUJd7ZX8ocpL/x/VFLJegRkjrGGKvnq92tI9szr3TM92EEwvC
dAoyTYF1LF60XTbgBaqxbO2QXIBOk7sdgahen+zCSDGusCmABTv65Q4j7SIhj9wsF0zBP0v07s3m
aZo3D1q/UAhoDtPQO6vvdt6G6LviIG7kq3p8PXCMobn5MEMDd6lRh3jTLx8g4usfLSsOG/DVpiij
OUshtofHXPIL2Ncdlcj+UA1PVyq87C4muHl12mH8YkAY5HQTtu6/A3jmSCAODbcLfkiz3pc2ppSp
0+Hv3SrlRzSJ2XXPpqyg4GyGlKffxaf6tT62AFbg8JoNqjWgSKZ1OJRqOcBYLZZO+gU9TCQakmId
FL/lKi2/xNGWAQUv8sEr2JBPxXJQdEb+iSWr5IQhJB6tYZgg58d7vDEnw2OwmnJSEeXhVRNwbisg
OmfMdBX1DbycUEL6I5ap2I/7G89Mcyb8b78qwJKtnR2R8miAMNYQt67uHufR0qmfKjd4/Dygftn7
TsA22yF/9ilXXpEwhuBz1H24vn/U7j0ucRP+o9syTMiJXnqokRS78ODbxwkpLRZh/yCpllRcm0oW
/Yf5Ey41TIVZ/R31bK6K9KMdLpCATHvTks2LVdHU1aIp/hEShpbPnBvg5rv0Jcvc69dvo9ZfGwGL
23ob9oomZZFtibPR0Um2sIP6SHMnbeOpfwi88M7s6alhy/JmK1t5rc9GAX0S7UfPmj378xCOan+P
JeU8WwhG1slf8hh5d3GQorbsTJUpiWx155US1rTVheOlzKoXb0zoydRqKrcDSdt2tXh9HLKK//8L
aaSHJZkWQKO2DDW7Dtk2v3HXmvoG8oqJYZVo219fF7UXH5+MoMKASlW4nB50jLXV/0blH0wJKxmG
y4TuwIEPOYpxn/5anzqWQyF46l9x/P0virjUz5G0rHEsvnU0nIVwF5oWkEQu1876S6fAy2hM5d0Y
vnkYcoCbKlY9efwG9ljNetwuXSS0Z/THctV3DiQPBrvYQPBrUlZcOyrORjbhtjJFPPUSZVTz4DV6
KujHW8mp2OfO7BZbsvFKdichM25m9hV4Q5D6WTtcktdgo4Wg+ZFZj7u2LjCWNZCoV6BX5Jzz5aZF
wkEXqf3FaYgdzNAQ6dgJOnY/xb3+K/XBgCCJLYsp+USB0yKQfjCGhJEsJSssS9N9+e1xEUOPFavS
yoayEnF0kfAAnrq7VegN2yi6jBxyePa+BpJ4RPYWMhGJr0MdPc8qsGJTyw9IF6enrSNOpjQxc+iG
OMdT6MaCIMunjGdfyKS8fakQjI7Se+JoBaUS0ST5L4dFJynxEoqzfAVxofYlCdfAKrrdJ71IAGR+
SIPbszbEfvr4cxpwKBWueuEpQbdc4cAcuC8DhEfNlMYLOlFKVf2JvXSdkeAA5/KxhWs3SkefdPqt
FYY3BTLoOXkKUascZZ+3z+r/6vrFbVuCXw/fL/GvTuOSQfKIFbX0c9ekJVne0VjFq9fLcsbKqRzE
HF7d7tSsqTDZ+N4aulng279XnwHRdiiD29vtc4SuvWHGMmcc3XsW4P/RJG3YQnvF8a5PPg4qUfqT
+ZXUAONB0k02RUJEokWQZ9mCi4K2iMDJfFmA6rHgyqPHHxwQcDTMudiJ+FBb3WQPf27p7jfJjcw0
ljRfqXLDIj/Ca/w9tEIkZVJFtBaXes1+icud0ehmmc5+wC4o3NA9ZudS3DmMpm2Vp+f4/bH+h8bW
ElZGIQSYU3uLGcELzEdXMjmtb38rLcyf3RvgxAf/MzgdyVEWjaCnPJmmmMBbOsI+eK5g4vcMX6DP
rUSht+06uViJWMs9F3RErEv1+5BffCOilL0bQstmOhDgAmHPWnRQj6H875iUaATJ6lsunkkJE18L
j4SXDJ1LoCQgPHG6kmiHNOzJHe6KXPz5eflqBeYEMVAiR24LJsH3saD550Z84KTk+7UD8vZ6MNYO
noXg4HZIJVFkBvE0mvGAOILSxuZtZJhLXRmrNPmTs+nkHoQqzm4Uggwk0h3MNeM+7v5EftIhwN3P
uv0YHU5rTvzNPWb+BUU4vVeK1AG2uRB/h/N4X9o5dB3wLmCvrxbU/3SbZbZnZF7ZWnHcU1DzlgZe
WC1t9S/8i9sNZoiieGvAkEShNvNfk/T44UgxV/aPOVNLVxu0xE7NIAv/YfqlaC3N1MsbNXz6iHt4
3rLcZoQuCbCvKdkxwFUxGsYIZWkVGxsAwK76CZ1aD4dXFO9y4XZXOca33HDnc7kw2c5BqE/YQBkF
D5sw2F00dN6qf3lb7hbEoTSSVyGcBXq1IINU3P1w2iiJla4LZgRdZw3uJyfnXp91Jg78X0dxdZ6L
W9p85a80cJEQT2EXf1Rv5dWWSA2KIRhmsp6cDRGUed+rThTsmIQMBBi30H70pzF52pJUOQLv4s4p
EEVmAm7T/PvZ7pXkoF+jPpAT0rHQvH2rixpvKhOXoldknPDAt2w/hcxb3YIH1cZn3MsnoHQBf/HJ
VR5m3FL98PRKMsz//uH5RmoY9F+DIa6+bGTdDYold8eYFaK0y8tAwRFd6rM0l/76NpLEOUS2+iil
Vg4Uicy0WzCVfbtORpdpiEarfXLEszzVd3BJ0vR1wjNRIAji1Ditd71OB8U1b1SIjG+COXcqSqay
h+UgXn7ec06NxAH/ZVeahrRo0c1IxyRVDr4ApD1V6FEyau5v3rcyd8ZADiVcrrDFiul27Y95ABfD
0ywy4qjlW5EA4/BX4ed+r12xrjNAvoLrjrAtMIMpTojJANT9nZXQmbvwYL0cJePuWGCdFzCP3gxf
6rFCPU+WZdB5hIyGjnkTHYvd4R+Niy9dPt6qHTu/WtDPjOe0txNkDMJBA6632snv5RYkcpb+UvrE
+yESOPLe176TC0hF0otBMRXHGrAs0saJo9q9XamIbLSbwL5p/JwVS42aqBqXyX7yvBjIo57UQdnG
YyLad09kcMvF9vIX8cmbeyM4trvk9Znad2MHt3q2cqRbCzOADeExmvEFwm7UVq1kGhDuiE3QyOn6
Ze1qGdkuXsXBy2UrZwqMiq8Ous71NUdJl6NRERcsu4IyygicaTQrBJnlgHXJ1noa4mdxMiDCFJES
CYeBFYICRDU7RNX5oDYl7AaBNWtSnPaeWzmWaUB3RXREL4ZlghniREfgku3r2WZFq18ziut2Eyt/
Cw/+9wt2SiwSEMLncsPmELYTVPLPrv2E2pWKHuZusX/LRPtZK7pEPEARRWwNN6bksjOyPpdmrMFg
lkV9vZ1IIFPRZ627+rIt0OovS4WCAeoiHcXhMJ12q2k9Rrc7B/mWIbAyeEBlFYLIzAiF/IsxtZEW
Q4HAbWd0U5lGsTS5fYsrgz51jL4B38WNQq3mfpsUyQ/48WIJYu7XbCZtgxnOLjzKa99bIjNpupdi
KSFGuCjJvFuyUrTvAX5WoyScFHnJs+32psNrg48MKdEIqVnrUUNhVf4PIo8zVjUKl6brMqqCier9
LCjLXz1QfBrcU4DN+YP2Kj4IizZ1A9VQKWBRv5Yef9tUirrDhN3iq5Fxhf3vSB4E+VRj9r7y6Hrh
eCsoifhrLG2ex0Zb/Rl7ZLemJQiGeDCLUdx5yG89pITVpQ7jW/cGcO4OIkFXqPVFLZkeMccA6jeL
IoRQWBI5HvS59d1La628IFLpQk6hYtGh9yELp3HnLjf/Zbv6R/AJPd7NY8pdqRBgdoHuhSY0MPUQ
SayNnSWc4rZNDeqzAQjiGET+nUx7FJh5T33IqaTteYBq2VlL84mdqKYTOf+hDyIdcVXEK/y/2BsM
9HKvUvbKkHFUYFmAxRNHjWWKPpICj4UPOxUtBew14MiWddsnWh1qlDgQ6I77nNC8xkrrU+ODoiAc
pMPmsZG7ghOU7CArK4vecG67vFjcTqJ8jvi9xgS3zZ8OHXVhpXG2JqVUckKb8ng2hisCP+XHAlwB
zcly/2OpivpnLbJVtBgCbBaHm8LLo8uMeGS9lz5J9/9ezbNgfN2B++T96LvxqgKSMQJBYjWPRYGQ
tJqL0mc2qBQc/ruSgBQPnytiXGFPG0tBalXSicfti/puyEbJvOgng9bZTrVh3sj089omE7KXyCPx
VWzto624YrtQkNE0X3aP2uECUviHR/fUr+LWf/UvqqjSvrirFV4GNtga9FepUVGXR/RqCzFVX2Ji
SUl9SPMjV7sQ5Wtg0edIrDBHAaMoofSLGhF8sCIQuwB6RY75f+VEkOfOmrVgzqH70238dmQudRK4
Gywa0WX8eKF5eAMk1/icj6eorgFZfnvPkxHtJNkgK13ZwqhwSDO7vuCMVAYpkpNo87BkmSFGOGwU
+wbq8fPfKJVzUjRg2a7qytCbQxS5Ilh0Kgv7bfNjDnLM3raNbRRC0TDvvyKUC0zEI1yF/Es3bW2I
P7Koiva3CECsNekG600E90vBiRpjeUAvPqX6NKoiPUd4dx1/UxaeRslPq51iZo2+OPWRKQXsEXZN
urlcR9XJkL4lgDit/fsbspF5Y/0dKwvAZufv4LnLdri4iV2T5UcIucAjsgc9F6oOtchrWBjXksDO
5ITTOvTYhurEzPbV5WEjbxnfBKL2zPpt1Kw7UhgSuyvNQle/BoncpYEYWCRr/enOXDEh71J+CDkD
sQH5ES6Qbud5I7YdmqmI6DwHpgFEPLPbSP7o9an9m2hDCLHoQv+q8imDk05MglurXKO6MYYx3BDH
jWeABGOS62RWvQJXYyRY/9K+ci/qYzAMQItJTKN+20Ba82dEyx1EYfhPtw8YARqHPZikVSqEC+Km
td3O872/aTftVgMuHUCCNIzrW0U0SL5w0d9AY0miTLpBZ8JgrK1bk6tpvZZAi3JjvLc0Jqs1OrXA
Ey9jv83YDwxGNjw5HAgRPR0oNiZCDIayRGRmVj2XZvwVHIhHTPgz6PdwJGw/Q3F3TyBc42BpWEZ2
48hg3b9p+i0qQb5yvDAs6CxW8us7+cw0S/iqrbX6Gmyc0XZIqLqUM8px26ZWP42YEwwMwa/YPBb7
rAlvEcjHWlraFiDXZgvlcYikN72sFaiJs7zpDfsjOQ4YbJus52PB+IBC8cRveWDWaL0iQ0Bq1vGg
VfwRVqtizNp/Rqh/SKyo4/6Vx84VJRL45b9RREcaD68ek2pLcN8iUKMU6tZk7TzcgJ42WI0c5b5Z
WlWH5A9kcE5h5Qg0EEI3uaSgsVeFUfCO/eMC81nKJ5ElQxjxRcZmKJRKVbvzGljmXH7st4L0h5WT
5VpCEbDqd3zm0WkTbzlI8VvtOdmTDy5OckU0m1QYphJMjTIQp3SrijmIYoIWkqjEA00+0LMvKuCA
3XhitMmgHH0A/28YiTQ00PZnGSjKsdenz/5oZ/QZwC3LZbSlE3vK1Olz/rg+2kdYVZ+/q5XTU9SZ
dnltIh4Y1TuWK6uITv1b/L/kPyMl18BA1jaLmj8FUeMB0wV2pCUqFTpDXFGsf5f27yuVzzDWU++O
tJTpKPHBNIxceQgDAr2tnzDVfSHYAknTYKHW+bwM6orYKdqIgv16W4+Ui7MFIYBBS8/2WrLgwcjX
mTIrJtRxfPbgpasNE10qmbSCv0wdr0kHDkqldWT2ftyiPmiM4UZKt52tviSNwnQW15VqiEULKH9C
zZaggPqGcnIc9F5JiKEhXyif6LS3cnfaEud11c+z51b3d77UTSLuDgrfDvP/JDAqXWZ/sF41tSo8
hYmDHVD6ZP68zgcZh++AlMi4TqALB/fp2r+b0vUPxoidAuBfDQAUBaq/f6EjZjSfX5oyAfnTzsB+
+NLq4L/avkGWz5tDuwC3+dsmxQDwqFEbnfNsdo9z+Rdhd6Rk2JXJT5rJxlGhOSi9PFwC3wu1Xstw
S28y3GfNn9UnX4+J9r8Sc+PwFyDFIeeGWysMkrb553hhjqqiaMJesLJCAOglc8gTvYiN8d+Tx+hj
zO+nnTXYw4lsKaaci7ogcto33d9wFRhbYpDZeNa4JoQXqW0KZVAeDytDaJhOaI7VQpWHFK32zQLy
4oCHDKB3QBgSEPo2yNPhT/SgR6udyPzJXgQphM6W/Q/6KpbsnmvYDjnXOZFhygaSut+LoM1izw+V
jyrLVONa9DfwLAcVxV+JuBRjWrXA0q5UJtZH4DbKWPR3jmN23PDtMRJNthmcaFUSv8wLNOhI9nX9
nOB7VNT9KklG05m4wtDkQs9pi+s/FsXp8jts8zc97BpMP1oB7BFwPggGuMCjlyDJ04fVQUlPFIGX
7UEPytSnAYtLvvgVqO9H8DMP3P0sAuKhWdgaANi1aQKjaNpNpku8rkEjH6sXbgljDgnbFzPxJvns
CPkrhTJuI9pCy4GnlPTqjO8AIvwG6e8kU3xvBLFHXe9/9FV/2eO2uXAJLdmHhI+5NjMIs+j+w0tc
AB/YtC1qYY1cT+jPza0DGgH85LNj43Q57DDoMldZ06NioDEvPKtGBlcACXGZqjTr2woOS7sJ1CD5
6YtIejmj2N+3OYn9TMykKA+l/hdnRZ6V5Lt5eMiKSq9VdixbSWfN2Zm4L3gbxvyjSKxs5A8BNpXD
SCynnnL+AFZsBal3J0V8v4fjXV8F0HI82UDBPC0Wr+q3QLLGbMBu5rXAXcwr6fa3Vd2DR73xOHq/
l7XU+9P+jiqa3AcwmXeIUTZO9nik9P+4CqdMxywIfoC2B6Y9JdgwdncZvKtnDVi3TmAbFgxn+TcV
V35yIiquCk/Snd4cyg/Z5ZaxppqCxqBUBqzICPP1NMf0HqaPpUKdeOfsY6FsJoJhGx2nV4VpU91W
MYrIR4dOR7OvVax2X5fhrudtdPEOT16ZGJR8A4/clfXG1p5Eeno+jH5egePo1hQbeU5EasXHyWA/
qH08t8G0GSQ+sFpnOrhIIpRM5If0XdirRiPP5p9MlNb7o2X+mZ/ElH5WdSjuQI3HvWensRwODjuD
xDmGB9FlJ9Q+5vRqmClSicSeZUfN8RFlzlVdxf+v5nh14lMbJWJ91qPhPzd/B/UgNQtMXAG48eng
x3MoQnebuK0pd+KmL6jtLBRlGBv425evu016UqduLAda5KgCC6q+LAE8sRrd6uyNYxbpHPjEGOI3
+/Tt1j07VXfRfx63TB6dNF7TaYo01OpokLsLyapH60pM510Dh2v+13WJIXl54GEh6R5zB4IW65ZO
Gy+iprtbpPEFUmSO+R3OXriZfLqqUZXmoGY57+sgSGa97BlafB6uMxrPfwJQuH8DN1cgmuBCKHaI
rshVeKrG7FEl4xBqraL9w5AR0nU27+uueLsswt6SAYgLbk0+WisP3s65tmukx58VzwlYsOSZJquS
5xQJHHRx3ldaECBw3bwMvKWq185pYZ2HlDLwWHmCryeSlSofUr6NNhbDJrEwVtDnpCpGg/XMHzew
rUVd8363+G9W+gag3HQjKJJoYrbsZPJsh38VgeJE2AVA1NTljPokfESp+SkS8OW6xXPBNv0QhGcG
JyBsGIiRfOwPr7Z880kV4J/qZwqkRBbjrqr4J9A6NzMq4sX7vv9SzrnuILaeUuJ+wEOC/A+ja2SL
PE+b3w1hl5DDQ1brIlAJ4P2Ps2TXOB057VzXFtzYPVIGK9FEAXo7q/zlb0EGr777r5yv1DsGuCm/
utj7v7QRz8st7H99RCmcyNRpg6UZ5xECFkh07ugv86yqWnOvUdAo8VmTVJG3TjtF5Uifau3giSZU
kbfFGhNCa2Lr9xGupFtlGjl991oRUghcyivmemfm9K8ghhCY+HYUItG6SMan9o6NDmOmKgH+hRIM
VpRRc/d2hVOhdxz1ACA0MfeZznonyMr2FuE6GQtETi7e2RCWNitZNE93pDrgD93BejQvggkqbq+C
fAKxRsxPUNhetZVZvDVKCypf8l7rwJXruGbbJU+D1xTgYhx3b/fnD+s6W98L2tmYB3t/sOFdh1gW
aFpgaFqbQ9ZlhPzEeBy/R9YdcC8hNEsoHUh0EOGSsZvnNE1UFE9CPiVqfpnS4p6EjnHKXZbL8awR
/3cNOt/w8fcrg1GrB2nlY/yAJn/G1rrILAsZev32LU0KLwsy6eUgwtFmrYWjcs3cnFqDTH6O5F2S
PqMZJroxJMcTTQwEjLbaVSZA0s87kMkNK9uUv3VWbBMdsGQH+6qFJOr6BgQl+f1r4/Ye97cAyEZz
zQiEpmQCFJ06u8N/yuCGq6LOsSRdjIapTM1EYD/Vkh4VZsLXxbRAxtHniP0QcYLt/1vL+MoeQ1xP
H9v7MKOoOoF5Z89QmjepXugeEKlTbKQW4lhD/cQcGjZ0/3dm203O9hNVZ8THtdFRvrtreq8B4srV
E1ql/9CAbA24t5v2eKI3Gsk9IrQgKXwEKIxKdz632aE9GknbGZ1wjCioIpK0onMlzEuxZODjnmSk
35QFOc9ytsa2G9Mb/1p+hYB8NXe+nxdm022r7CN234lS4kowGDpIgeZQ6K7QuCFdIdV6rRoaDG95
mqJ5GTnjwWA+IjmhnOcv3vi2eJAWwOWjB/ySacXKfNnebtzmwxWPOzQAau25DCG1doehLz//O7sW
k6Zihyl9hnNddEUnIFKopTjBlTOoBetdm9J9u1J/LMemTv+B/TuCoJ92vmlAwXZ22l7sTSNwBNPx
KleZ+sLHjEa71n/yB3M87yS85pUhE7jAn9kbO+jIlIco8GnIwcbH9owUXFAtP+TiqOhmfdmjLUoz
nCHb75xot8nKFn2v1P78vPW6ntKYQ0Veu1Q1MuI4kxIJZX38aS0//VzB0PfPsiRX/lRgoiXU17n6
+8U8fnhTtG8Q2/+iA6YchHzZQhmM45ozEZhitGnycsd0JfP50ALXYjhPc/BnIg1S7Y6SDgXc59Ph
yy6anJkrVqplMEySZ6+OL9kbLdUpvZHIQePYtRg2F65rhOnhTzcTW2QZTltD6hJXzhFuRliQJb4F
CgUfNhLVDLFe897Z30Gw5QR2chmV2RWJ6rW5XAdTGhkX1nYBhc8QSUI2ceg1uFEFGOgl1MDck7Ke
DPZPmmMRg7I2P7pp+j4fsyLXsDeTYAF7sg9BUNxyMrSmolJ2LlxEiJPL4fQsKty+BElf8zk9QDxz
MHb3l6taKaY84ugmnXn5jGL37FmSZ2l3FrHLQeyQP/vzYYuQBgKCi2zO5dbXiOY6OwLXgHIjKD3v
4MIoarkCI+0qr5d5TiYKE01rnYXowg91/wicvuTSVo4jdFitklAJIvcIFcDiEHlSHW2N2o0wJWge
6SVXigN2waCJe1L4Eir6zanLRk+mRknFFbYN1/Pda3lFWUY/x3tFr4TGUAlzFV9bN2S9N8jJUkMx
Bz+ClvwyzkjLZqxwH24O41Sbc6YUQaGFeyxJY9NuOFqrys8wEXJa/+tx1eqjMcZY/9mSz9jv/Hmz
gbBDCjM9hEYIL0dsFBArrYLCAu+2Oi61vxM1rYPxB97/j3Xz0YK4xGl4M9Dg96p1oXwGqDQYjte2
rK9CypvcmECH9eo2jLOO4DU6Ih4kfPMRPJuvcfW3spXXnVyE3pduW5s16kHkaaGv+cmFGvledsxa
Q2tZHVa3nMvu3P0O4BSLmUXDmYu7jF9zwNbWVSa+OuMQlh5YmIUVjEYdplKiOOfuuVP7E4ctOGco
qyEKZW87Hjr96NTBJkvojFh9eM3oC1y8pdnkfAeD1UbVAkXua7dRyOBCgHq/fhg8L90W4Ofk1Rbj
XpcofGxTGB+grBWY2lUzH9gxzYVEbQWI/3RqYCuExVokc0dIKVvpAujf9m87IO9yZ80GR85bsa3q
b/lr17oUvkBjPMA6nURn6UPGFqzczYKYPJoU3PFf6PrjaIpHWcvTZcG+tGxG4ZDBtwx9UARU1cvo
yUZV8Ovi2eOqDoTnq3XEq1ybc0bjI94+QksRRiDlVzVmMl2mjDPwvmrvK/gqn3/HNi1BXSNWrNTD
JhoVQUOD3M9j0t/eDlbkHP1X5eHUYrTw3hKQ5Cswz7OgSKN5x3wpvNAF3ftmsD3Zkv1yn3ClrOix
ceEclSfaGwUa+bfdRAS6a65iipUEL+Aso6Bpi+JgibS3cmAY0bKzKKKMS/k5WcfT45TJbb2Cl9Bi
4aRHykG1Syad3tOJwyPNvTpz3cr3wpFxgs6GGAjJ6wi46lvAR2dLhcP5zatHifBI2QOZahvK5EIz
QXs3dVc2Y7I5AysgdiwAUIMVVvZmEoJW/mDvEI7ssI6zHTS0l2nqDidnaIDy8/aY7nk8jWj9GsY3
9t976Ps0mHEBRJ1zZE3/rv1Bb2NbMIbAK4b7a+U4xKntgghN4MDrSv6XXZxn17NBMD48bpJ8IC71
8MXWp2A49QvlBoPvoa7ICOZC7qDp2y3tsMhraOdfl959khxn5jc1mjV/2CCjuoi+5Oa3RGUEWzJU
gg2wThtlYi6cc7pTk7Fy1snh9U9lIqfqdfywPyKhV+KSWQai23opuqFAygzSaLMc/DTfUOpLbDRt
MgvXXFRNyqNR9sKVHgnM3zBdII97gAgIn6JUt1YD0ePx+9lSuOsloernt5G1hzkU/iU/rdgKPq81
58XF1VtNTvEL5HrnBya0FRFDQQuhzyU3gzb0sU+8McKpgxMQV/ci7NN/+meTJ4WO7/pP5LpdK6OT
IfPiTlQJggb9V0KPeo1SvqHL5+KVhsYCINr7mpqqjfwPIc/VUOpbJ+Waswdvf74GZKtNWoWZLWsq
XwyKtObcvbGjvnQeoiVR+QeBRh5q1/5EDebPIpY8MtI69AR2+FHI27gAADs2PAIN2SSQorCByLnz
QXvldDvJ4RJWhyStPlOszHZp518zH2SaQn+XioYqGgesRvZgTca/B7VdMYvKtut9OHRnZ+1EynhD
4PlqWCId1QrjRala1fYoNt8jYyWiZsjQe7rYCqwgKzOX29Eglw5V691p1dlgm8iFuxDUSHTbpmLk
36KTGgEm6pKodTbLqdygvJjoAGc9wfGnXM+nuchESkgkignxqnro2rc+NyKaRDoEQHsah1FkDvKa
bfiXK3O+PMF1cA/oaTX1ea6wm3RRomZrhAlmeGMRI9qD4GovpSIAPuBdFqjYauGR3G2XtTmmWwx0
opk3d+xEY4jcdt2xKJujVZj3tM7honBPSy/vWS7Q+4SNYJmTDVLfcRyrjfxmXnhOC7gwY8YnVuad
9COMYiycGVjTl+rDyhaevLYRXQlcGgwb4Po98Kgcb5WyATDEndSTxiodypm0FXFAr6VGzkLSQv8d
OhZkVdocPksEqKqwPXwIOvM+FH18Q2PxdPN9zCM6TLWAHTKftsF7MwD8etIMVmQPY4mWRKFgaiHF
kkB9/H+KvGE4SA2mwA3SRJNifRYb4h7DRZy9gN7dQLoODGMGx59G0OwSrM1zZdnpEEfTC4TutpP0
dlXQ3xPqaIbwlZhRmpbTgeoLKN1ey496xySYR+oaUJ3ZG3x+TUlaBRtZYqb/RXOBWumHd4LJRqx2
8Y6gxRdVNJq1z0BwCYb0R9AODRYxf6HFZMxfNoThJkzozB579qDE6oQ9xMbdSmP7bnesMMEp9SC6
Gect8G9yrDdtWgeAgdOjpz0D5JRSnome2UhxLlQkwXqfbDqhWVSD9oure2072n6EMm7sfxzAVSS5
LdyuWNQC51azVi2H4oXPkuy4sjCwilup+kHChJ8ZLaC4XguOBrPr+rr6HJauL4Pgkkg2KJipy8rk
tnnMHlixJ1QwVrMjjZXAL7cqV6dhOQKrZQ2vYYeTjTqRZB+N8qSKtVG0lB1uefTvPGfCcpQyGJTy
A6oDUjN2veyMhctrH8A0rheathMUKajuKULz6kVii26hRI/eO1PvcNPtVPJnqu3TPwzLqNTN5k/3
Dzz2CXVzY0DJ/CrzNc1hPPGZUhaF7i7V+aGezIFDND4g6gToSQI9ADRKY8zqvRW0QGmIjpqRxlEr
dOVYLghoGzLXdzbMnyIcn+SVylB394zL85+gid0SyvEzXUXBWy3p8zKfXEJwfjL3kb9YirYa5In8
FojyZqdc01Ah6L7dVHh7OpaCzSRvkmkadfJ2XK9EV8to9l8shJFrypO1M9bt3vNXh9yxpFIMj7to
nGd4QWJZ9bnDBFstqhj0a1rWUpgNjNGBM85kZjGjIL+obQpSFvDggraANIrsIWkkzucgvkbkLSim
XwWKV+C+9PE8i0VjMrP8bVe0LwkTRlduUKhPdYvaeZIIW01IUtZE8ZM0D0v9MH9ZprFa2iaOKyvp
OU1LGYSL9WRTL3b+bAKtyxsWF1eS82wEJz5ysmZMkV2np2sJQeuOqPWBRjQU1SNFDnAIFHkUoR3v
NKNF2R8VmKrY6TG86NELvq7xQh1yxSnVBLxGXyVZlgnyuhm6LFVFE2NMlSpf6Z/8yesEonKqNyyM
IABwEqJalGmO8y7nLNaFJYQj9r/DPDqyb9Q9E8U24RdiJKSjxm09KkATiPnzB6MKti3aR4EZe7tv
ScH7KwF7bLf6eSYEICwkYOrn+rPMfJsgR0PLV+3U5TCEEP7KlfrPefycc0Jy8fEkagTu8Y1Ortsl
AqHoDaEXmLwd/wKC7af4Qd9VYAQnax1hpjQDxXHyWmtWbpNo9l+mTjjhMJDQBcYFXeX/7bkEP7VJ
VoPIOrRgJQ70ag6tL+B+sYGTOLOawxOZ2ImVmnNWAlJOOYKdTvd4WJLR2dnV2jKo8BNlB4D76XYm
f57XQPbOvJnp4mYWOcpzWinsMaRyS7PbmAQjiKNnh0jbjklYgY1qIjD3sDcP6oXbx2qqpB1FJwBa
ElcUqz3b2YrfJ/QbrY5z1M5nEqCb6BouS8eTE9aEsdfzZ3urJ46crYu/ni/vyuahFVQqq2x3W7ub
WMXSjR0hdsLBoG9lgYTxmbaPNHKr2JvOghI9SmRcAfHXV1dX3CVx2MX4DXV52CXF6eOh0GqI64RT
f8oGoZ7S9nZYvCVYhcgi7/nTD8RC/SUoDoxGviDzl0W3blDsQ3SK8MjMHl3U8lwE9LLVoIQ3cryR
5OMIqK9W+6kpLlzK7a6RTRNUZsyujn3dYhjS4lwfl7MRIK8VjaFZg2XtZsXMy7adVB1X1xAlvyfD
Y4KV2dCXniAE/f2wla+tMs24lmvP2GvH0IrHD/Uvng8xnkAHo6HwqsG10SrOkADfLDJ7R8GXPJ7Y
TK+MLGX9u1xx9GoD4Pf5VmmHjZSMY3lsmSdUX9DOa8Bh3ZEqFyEWM9YBkUC+rbRvoWsS6107zKqu
bBYQdD3IYj8JiYj66tzn6eW2LX0wNBOirT5KWu4DxDm2Eki8VsvIS6J8p1N5lDtYnx3o3sPbg9PD
ZpONKcLqSPe3b4nrzZKCLqgnBE2b4RNboK/ctxEm8V2HsYaYpZ4KZ/NP7a7DnjMm/m4/b0LKc2H7
fmE0low6dpgwlKdtgR/sQ6VGoCcggf1V919ioLfPjr0hfnz0pEAX4EtzPlM+Ru5DBFvvlT3zq2Cv
8dR2XtFeLLFAB/L6kTsbt0fWUzprZxyfiubfoGC3wWXIMPru3zUfwGq98+tJEVkIYlHPpaUMImeU
rbLnvVYddImZ4gpemiNTDS/U/1VI/EilhqK5Qe1mdpTgfzrhzTADBkVO5zVkAMZEVdXdYpvFVTOC
ND0Js29KmOjFpdY0ZWrvYrSvS7GGWHGKmxGu2LZPL5tFxXuE//pLF2nwiZsUJYAu4CgO0jWnjx9M
uckRYY6AsYIu4ptfmy5PBVvlHsDtWp42ZrglLPHPR47Aty7FW8Msloxy+F2e8DT26pnj9mFlt899
Bjz0NlOTWMZx8TgnAZjki/EDuDwu+v+rw917RVpAQNQtvP3tSgtTIPjWsFuRB0yOKZmgBLfNGO/g
5tGdEHbbHCAlHMQ91DAwT3yGp/Y+CHzVW1ELSFprF8RiTpcQQPRsFUouTM8J3Z3cDNFV2mbltEuo
CZ2FjYQqBohHcGrCgFV+ddk20wzTz3lE+rmGq+C9jVGSo245u9xeFWMdoS/XYnxcPcw0JxVAUxB+
ruVa0qK9TXHBgM36KhTZfOeY/ENeHF5v/5suUtm+qV9LA+sbLoUXAjIyJdQSZnY0fjRahP7HVq3G
hbDKfGF1KTjd8QxweajtFA0DP43E+jPAe4EbuQvuaxhLg30yA9ZXFPSx+a0e2y1Ciz7wcSA9raB8
blldfNTOaYrIrZwqgaO6/aqpIU7wQvSd81v6BBV6eRJP+N+aallU4oNO327+NvvvU6tSuPZ2LAxv
LZhNWv83+F/BPc3KqPqghYB0QAvv/egK+o5ZyA6Y3ZPk9g3SP6T0Sg0mYkoJrnhU9/jUEQ7NHRNC
YCYglKSSVocvolJ+6iSoftTDzmUO2cTzr+PKkav+xTWvX5aqYzs2mddKTXQlIGvScYFeRcT2/56h
PzOuzqqJCGdooGnDfT3FinzHgptIsYOQzGITYqovzRtm7EGnq2yD5nSyvOCu3EOvQzwy2gsKTA3M
22tFHRJTwxoChkRMAf13nYnDInCEvSG/+EGNatJbg5q3Vu9+8A04MKX3HG0/RHw7Q43jrIf2ry7E
jZhqAgkcMHQ/aW9jzVISQaCMP07qKW61BWmyU1z3a2hAZ6cb4JvWqjL/ge6/Pav8Aqm6F2IYgwhq
TlXU0hJj5igAIiTShFDyTUXI/tJk2lXSmfL1XhAOX1gIdiIzRQfkMBQh4Lsw856N6tOAFgPvRRlC
Q5Mo8uMOsJDptdNj/wZkqXc8DDyny8nTiCxvZA49KKJBCM9KWF4j1ByRz/zxUbP5yv3uGXzzyjBs
3hZT6uiPwJKzAmLhCuSyIPXJwkiy2W9WcMkuTBelQYgSYc+0G558LNpNcpCxxDQ5HiopIfOQex0Z
Kkh0x7LVe+IBxfHvvmF3ozuqpOYQA6Pqu3H+2bnlHVbejChJV5BXHwIXg2StGjFZ9jOonlXmcGy7
gqk+81IhEulk6D4XAd/i/3ijuXHZ/MmVeCJCtU0OIYIP7P9hC2O01ajD0elRDkNw2AGWqLFKc4PH
s0P0ylEosn4itFkFb+7EAtfZE1eZeWID6ulSdMOTyflpcUnauqf4mevz2idjbKRzFaoXlvK8LAJu
ay0imle1uLbNqpKPa8OWzxt9mKF+oV+bXL4ft55iwVfwHQfDat+HicrIUQabe8FqTH4DMOJovbDf
gVYF5iTf1g71lU8GiWMxCl4zbr9aRsQau3fYqKdy2Gjy1gpeYae5QznuwOGE0yA6QLbJq27ihBoR
g3FO439A16wAqSBhNCNgwiZY10FheHCSt3BdosxaljDKdYeF/O08xv96pBQaX/qtBSTkQUKBHuIm
2diVqYWNFdjsgYcdCgmsT+reIOMFBx19EbznkWldrvL2Pt1VUxayYhMH+c5z0+yYgHjssjzJ60CZ
INw4aDelwFAF0hT5Tp3d2MMtDWM4NQnw88fpRyUFjoBpLCRGv+g4yImpKTYPEwvgGP89Wz6oXO/u
KFs56YDlvbK61iGGzg8f/R31o5CIC3D22fEkXy1AO0GW5tNoHdoEtVNjb8w0vgowZJKnA5jRlrg3
C5A36TTV0y53gnQnZwKtIdZoxcK+evirY2hhnPXgdXRs4FKz2lRyk4hjopNkgeO5O8/aoc0zy+Pk
SIIh0HFN3w6Kr0hH363idN58yqtYGLPz18Lr4L0+CAR9ynUV5Sc8h0SfXiPb1eOSIvnS3mtjGgFp
wPv+FztoyDbBUAA5jJ/mtbzEc0QmBLnw4Im4KdDab9fEDflNlOTZXrBWNy88mvs6eGuFS23W5ek3
jomYOSFp3Z18fG16QXhfqESg6v3JUIDguhVT1jlLO0LgvVdz42vIt5g3bQh20A1FYdfrh7XfdErX
lvJIwESTKE/aTptfWShGSpAHPazbakMfhUwOpEfOucS7yuxsfHiPU++CeawxyVtJzTAtZwNetrPw
DvibrZ+H4vXfY1aQMT8hsgMTkGAn4oaMSCM2/f5rDIpg+iIJ2bCZQeQLjyezsJVK3m/ezE8Pn8V2
3a7xUr29T7wGCSSFpXGGFFQnYCBF5DVvM2MDRsX985o0FWFWpNElGd5ngZjUfEcb39AAYO0lCZIK
c6+OGSOExKybaAfMs9d671Dx4UOpkJYQ5MQdsICcvMY+LVD/AGcFIqJn86mT3HFqXVgtmxE5yXT+
UV9Mg8Yb33Nwnzf42tJDWrQugD6ua+LWrpwF1fQbUmKkxR88Q8LuQ0Xlnk4AbDYi0Jv41jH63J2S
APmEL3+82p6xY/6YILS4g8ev9Q9ynKMj4pjvgRrbqDL4aZkDRO9pZl21O1lbPII3i2OQ3lOMqOjb
Ks7wAY4aoWW/uaWCutT0aW+qaoKz6ifeGqrWcX+C4sv+pYecAuICrRQTNbDhOVHIAm1ShmAmRQrz
eUXVjFOtAjqjIZ/Kily9fXNVkODTJSUYUtsZNaEV8hjadUuTBvylBHlY+QfHGsckkrqxLq9+Yvb/
RBQBknc54c4bjcQ/zFaj6Gu2y8n9D4XAN/00faWWhjyfkvXKZ9Uzy2iGG9PNCZwV/jDqRc3eMRUy
CTIw4KjwyaKiaq6hUcgyKjLSF1Xmlm8MfW1akgv6FL1Fy7XDm/Xn4U6VQp96q8/StFt96pzkcRBV
jHPH6mDZ5gGlnn5pWAY/5Bf818zAnBgNmh6rqEypH7xOWyqr0s9GMb4ouspzedJMSK2SqIDLGDae
FyY9xMlC1vPX4L8zSlUTIObL5ym0kQrrVLmzcrL2OY+MW/dV/L3GEG9b3ZuciDzG+uvOV8JRqil+
zdsiCaqoXbOosP+eujQegjlaWUEFPxMYPxORvKcL4fAbD6VsRgB64sVK/sLmZlrFIxD4kv3oFQGt
u6a3UGOfLyRBCWvulET1OHnW7CrtHeGyA4sFjix6CuWg38q/AglBlZjx86tpp+CeH8aPZCCtEcpx
sEFk9kRqu8Jrcg+tXXMk3Bz0o095sGr5RmoXpugvBQ7f73bDpniSY4kN3uBlpf88A+NRrsaZGvs/
k9BaWqLKvFhFcNcMeJndVMmoFXq9QEgi2F7RmQv5XDk5hu3D5gP5mlwafcCI4u5eI5ZhcA0oZIjk
F5yNqm1qIA1E8i5irYvS5U5AaqZNOmA1fjJX14YZgx92MpeDqVLGypT83crMX3h1rcqnepSZ68mN
gh9UJckNRWs+LoY90u5d0U2J98P/Z4rQiVwehA6AcZpARbHYm0zKBIqnQihlL0UwdLIZQ1Htzp+e
aH0xDOGMtLSwl/MSt2jN4TjW7QbhB3oqsXwXmTOLPTKJeNezOaL081DwfE15T+w/tn3A4R/8FDKc
3xfl3bAngC1k+ZYzJ4FkU6yJ+C/ErDId1aLM936yhCsopLeeg7KMb0IPI7LBaws0BnbBEWdHVxqV
i3KDr4UazT3RiFaksVhCSgeOCAB8qm3Ee1oCed7bvroBg1W90BY1jM3RwaKnqa80wpmzdSKZnL48
aC8QQCWBr6RiDFkkb0SXoo/aeWn2h+QyRnjUzrfEF08GPZaHDM6uyctQ3CBIIz42TdnAeiXelOg3
uwixdfEtKjnNMuu9T60KOC7Zjj2d2qawzET/V2UFIODcD0heLghTRRgcVLBblQchAfsGRF44FlOf
IwY0d68viJOhYzoRpusP1wobbw4Dj/KZYaTagMCUFoMbjCd0RWrtirpJNKLwKhruS31Yq0VCfuTM
/MNnTJwS7vTQrXIoUL1sTK1Jrdu0zNQdsfoyZw2ox5g7AvdltVL2aU4/rHFFldrMgm8c7ZDYrCov
Nx7ocCn+dDrO09nrZZvKH2jXZSJDqUsT6p3a/8OT9Ni8jGYlohynAHVlmSRpd7ruZLn01KM7nnjS
HOfQ9P7iUviL3hxXxB+tL4u1LQJCvOWJwxTgPVWS5tD+Hek6gyJSCfCKJsLt3r0PrYyowgJkd48D
EgoHrYRnU74CE4OxqvyChluNgA0u7BR0IkvkdoQ6DHDin83TxGYInatXd/JPLEuEUxEUvlEjCmDt
RyQma0SKP0+iOW7Mpoa1MbQ8yyJmRzbnb9bzivebehrV2oWpxHVe9SBQ5QoJ2OnzBcS2H3l3bVUm
5zJP3uhykW3VD3vUA3M1gnFYqi9ooqQaoZCV2ud39LpIS0kWTdhqa9yoYhIOZ9PKAw4cenpt8UX1
XUlcrO4d1uf8HGTCSpRrqVqJ8+cwPlWxHdk9lRH0VZTbIA97+d0lO9bqfY27G+e2lmUCoCX/jhLx
QGKy2y+Te2914FnqtlYBkSZOCv7f3NIw50q8UR6wj6i8EH03r+eUxxYMt6KicRl7OfTnGQf0SVOl
7vJ55O9Vu0KIi71APnlLh0N7Irlsm9CtcdRnRlx21pWkPQ61IY4A9k+CSg/pA1CjpthviAf1jidR
z5eqcQC7thSe5i6Q8iA0kkOA00A7e+BEKJr+sNmsrTn2lJ/S69fGGqD/0mrl+lsyBvRNKA55Uv5M
QlWXDz27rjd8GtFOrFCpLEv/RWRh7weAp02n/UbLGX6vQB+WI8DA3Sbfn4srKoIRogcFrLWMt3xX
069CdeS3Wq4ga+sw1IYu8HiR0uwS9tqFC9L8q+xm1WsU/YifOjPt/kb7wDz7ZEIs/hdijsotc1cF
RNpWBdFanQI4tcnH8SnQfsXgBkDHUaHsZtSAEyvAMDlrfGL3FiFojofP4RyHSjlj4/d5G588646I
/uVdCHvqgF29HD7ZRjqzpF0mmBqVIuVnwVzb4zCvvcHLhWeJlJxj1dMIuVSvNK7LGieBS0c4ocXI
oZPPn1BQmJTDqnQlHW/dOvfkxtml6DJK0zpC4ZIafuaXLM+XnU41T63M/6075oe5RPbUdidbbpgJ
avw9auyH6agXfSkSGCyKNMnkn9xnaiWCPnf6qfoLX6YgG6/xmDXVI2XkAQ/4q0Gb2k7vmG91Vb3D
vOQdrRNAd+UnMKJJqX62o4laIPjATpN0XXhr8kSiEYaMJQpgggYqXFHur7aSuoIEPbNhkQJELFZU
LMcVnucfEteq6AkO5WvMm2E7MfsRGOQryfHuqyX+cQ9syGxiOO0JuIzW4GNsEjE/avcdSd0uQmJj
JXfenGCg9hfcXw7WzDLT+LfHzB5yKp8gorlOWKAUVmRbiKF4h6JM4cMXPu12+IOe5Tjoxu2Z5cVB
zuiTk9UFlnrON44M1QrZ7MTZMeyBf0t7v/oRFFd6hAr0My7hKSby/FOj30fDhahda9vPQR/x43bv
KdfqlAtxoMREk3Vp5n7xA05E1lc0Afo/WFWiZnt2myHUsGRa7wUxKwd38JgzvGvPn7BcQUUFibXc
ePqIxM+zkNPGLZgb1aWAeQa21+jmFhP0M9MvmHH9QglwojYcHbtUWYbMgqC/cCRHqCtkkSPQB/mv
Iv6cANbPUIPpYpQHY6P+UNGddkQiD3RXoA15r7ZzFAGGOv1WH6ARh+/xk2PjpkFq+JrXlZu8ePMq
uOklTvtSSBZeuotz/afF/V0o0KGBn5Jv66/PDDn+FRfQENCgX+cR/zMBi8vWIdrmOMCw83txdBin
dPoa2EfgPv+2RptPas/YlPZLLAlR4pnYbxCqYYBbbSYY0nFCAn18c1CPe7ElmJwlrvepLoqqhiw0
dLqXrU2maIRRdcsV98IaXd4FBdGPa7w7N7vvePCvaPPNV1l82CAHlyrmk3qpZm6f1YSZR7yQUnxf
A0earPmjW3NE7J0BGH0nv4R50bWO5yyGc0qoCQgTJrmJfD6MnUFIhDeps6e/myi0FkyZpAjlku3k
p9TZ29e6ZLOK0Y/QFIybNphUoVaQ+SdgrWBCwO3xTZKAXbZSv2H7tTRg8god3RW4yhQvO35RsF8W
wkoj40mDlBxbAnev+40nty0xXmN2LbPW2UDzRn4PyQOEN6uUQWeyhKA59WDW3KJbt6SF38zLkYmr
PlapkpERhulSoqFwd/8KDQ5iiLXksiIMhlKG8U5Qk90UTipx435jNBdV95mG4MFuvhc1W6yOEpwb
lv2jUwfBS9d+KupyekZ2KyWdD5EFtfDD0n9IgafI7+ifPDYLnZynxSmbRJ84b6sre+uWlsF4sGA0
rVAVrhl7qC2Ao973icnHFo932IYSKlHfmKGZesBr9mjAToIxQdjzKWgRFRkSCSiQDEvzyxpKxbBP
xtn6iP3C8LfUx26oAw8ruGQTCQeNKwz+kaq8j0nu44gJICyMb5doD/SzgP1OBLpshAK6aUVEByWd
f1QUKStZzy7FGHxa7anoFXNCTRh6KhITnH5uxYthRYTQO9xCM5KtlKqqaHwpu74YMyb3+cyMGHvR
qipicoadwqyREM4zz/6aaeUjz039c716EU5Bg86cwvkzQ6fj+kHVAy5M/CWucowb7epjkaA5jU1n
F/VzWB0d+pQO1Dx4UnAWO0tDlyUWpmHbw+HFVK14KnnfOQVruuLcBMwVAnGkzRqb4uQxnoOfvj/j
NHhSwDpD6AXP0vf2V8DG6DfUyaDEADBskr53su9Jn83RCfJRUIlgDsLolaz/h+wR2bm2IiXvolAb
CDD2PUasZk079/kxLP3kPIUv7CqYxZzyA3Q0uVPaagMgjb8ExpjBA6/tjs2QxH2R8gr2pkpIcMct
CVwAmpCKoTSb1J9JGdFOipEsCUY47ifAN+RL3yhI/YmR3/aOvaVNi2s0iCYSA89FK7vNIxqwJOJK
eG2ZxEvbLoSNtCfcTBidwUND5uQ/ExPBh1mEnXqoJn3X8fXReNV9i//mAhx7K5dD+I2avzi8BEdy
wa6OXCEWTj4R/Tot3AElLfsm/ymGcVqjFqJOu1TZDsFIVJXFia+b+Nhx9svAFwtRBGiupJwP2AAu
HDRMlNsYLdkAtkIr+Pwefe7JBIr4xFEy81Gw/vwgZBx0lgFg5ksFvsvoNwX0VsQ9CorqQT48Xq/t
gFIUclR2By2uKV1lrto0SQcq4/48xtmTlUNTd/zH4q9UVzOqc9e7CCpaqT9A4a6I66QLmsdLk1/c
WZmInz3nkmo/kZq1oexabh3JaXxNmL/9ZfZ/Bpwf/L/YaV4KpsbdbjVFEzhM0xHejeqFfpFSubNY
SdI+lGP0Ruf6QNQbLVH4cN6Tb7vuK5tVahpuCLAjGAd3QAUc7SR4sAScVTsDnWY6ogSiS8TagCA4
7oJEO5oknA8I0xPvA7V40dHGjrfJ51CTj3sBumpCn1OR1j8mbFK+O/QjhqocDBbhRtGOZz3J5t5/
n4Jm+AGbAmaDq1MJXtmd4IvG2cXsqCiElaQ/qmJpMa+PSpPrRERSijnp1dCQAmMjzYrU77KVa+A+
upCjyVnuGEI9WZJNfUvX6lgc5UL2ktgJmAIiSFL8jxtuzVdTx93cJnXUgaIZAFaKxBWux8qIvt27
js6ME69r59pxtiTm+D22PD6OfZhGQiE0dgP3QiU6Z3CNc76sQVFLWYlBcR51mrxsx4Vq6vRxquGr
3IJCkdcf//JeByfT+4n4NcFiazN6xIaub7nUZy8JkKANqNqw4hC+q8DFCU8HgvNC30QzC3WfOa8L
WUTCklAOghXX879D8BGF0hMKwmzeLH/NK2uRt611x3o5L2Y+JRLKL5RxS3KmcEE8VBBoNpWTVI9y
5U2zwHJYTbFpuVCtoD8JrePngqhc/0sW6UiK/6PMlk1moT3UN2gO4NQoQKrfsZ5aRRX83xcsDbC4
5OPRK3XjFhb/Gca7KhMS/50cZawk7bTSB6CFEqDgBn5MantEN/VlHQShWJMaIVTNVVWPOYqRcCKT
okdRqdhRgM7GDR6or5RpMH6+JhBOj2WQrPd4lcSdGQbA3BzwHc9YfJ9/QCefTNdiH4/AKPqbQpbp
gpAkSIWXc9O9/3YCD0bxf10dMm1INAzj+in1zg7T37IYquGu6i49arOHHpmVOlOC7a7ijX+Fz0Lf
N8WrBNQuJY/HIViq8RM9Ajr0QzKVClxK5dHEqBA9+7xe46bzHV7+j0MEAfu96k7TEDi+EqAFiAph
/TfLobniykCK1DNQzriwhvcPn0R+KEyxxw9HnmjKuT3gKTeaSANdqUQzW/E1ObpbE88gvW7kVvIw
JXU2hKZhK1aQfVo/yZ+AU8JOeZUtmwq+ByFUvgJU/DmGWRgACMn5fvcgfnpisyqzt9XsM+LYFwpO
XeU3UXpfGMiJC3VpbKOaIF7iQr+ejnJcv5LwOJPhiT6Kk02zCZBDL67wqQpt+jhjtyD+y8XrQbak
T6Va0wozyZvLvBFFa6zwS+A2nijn3YY0nUPVhMEq3oGvZ/WYuablM0Ek5Fj9mKu1sC6dVSE/xMxw
AmmnkB0hJI8J3Tgn5F6MikD/gfHamFHoVKhkyzSVkylHg2Wuy8PzOpxAOvo10B4ReG4+4eMnaIwe
xh2kzuSiKOvN075WZGzGBEBVfDf4L7fA2aMlFss0bYtzrWcVc6/zmDk868ZFVI9mYJmmot4XKDuc
yKj56WGeCOLohEt3oOB7OKWhtW10a/u2fyZiZe4cs+zVdrrNr7ORDJVLIWrebW0kj5GYHt+rKD2A
MB4tweOaBWHmPI0G1cv4uBkNSdXhLl6RFxKNBb7gfBFuNdRu6oqnzC8q8Oo0o2NddMkmahhNwwrv
nHH/ojG2KHD+6qaOaZpZN7OxP1rSkFeuzy8ieuDgkQ9ojwWXDDJcOxUXUoHZ7QD+VSpLjXDjIsj6
NZRXPr2bim9Pws8tl8Eg+5IJWiFQFmzYt62bsgg0NKZ+T7bJyKZuFhM57j+NsD7Muaw5kEvoxn0A
V6GQA65QyMt6P4uUPpbW8kvuGj0ym25TA1aWbWeqBDsxSJh5+CkMr0EC7YCAkm/hbd5oLilt0wji
NLxyz9U8/gUJ9EZvorG50Iv1v/a2WxWCaKq0CTEB1MjBPDhh0SaJyX04GXzDbzurjkihNGXK0QCw
9C2Lw7LDweu2UN+pRafb4GG9E+TZaTrcqZL+eqvoI2Bc2XFLq20oIqficCTEXmrQD1OKjLOV3mW/
wnWrQqkL6sRvEXjuxdywt6fV8LSau5YZpkazIOjMNaxRKRG0JP7rIw1pQmvBKRxx4ZaRDKRV1DDr
uQr/5RyZ/RMFC03fpGSbdTShLIZsioOxtow91WMP/l4gDiXCNqAYAMBo1hNrZU50rais7hX4vFEW
MbQO5UavxOJ4IK8CtFEK+BNzrTEA8SPm/IkjWexJ8y7hoybOdUX38mAhlG2EB20M9X/4QI2lD8wb
B8/dsw3rXOYYMUVmOnLU6Qb+6tbB3RmAs43V8pern0StQZMo0hzusodUBdqowgbIrXbcsG8zmAz6
PR6i99y0DXqJL9QP041HqaE3psLJd0Gd2dRV6TfLA4CrNIpJMAqRqcV3pbQiWPDtaNm9V8NK1DK2
nP+ZlbXWXc9Q6su8IlnwOQk0KMk0c36tm8ba4UvE4nGu5NixXQzhYwZapiH6PLiqF9rSA31meOyb
PbeQIyd7mv4fHWfC7kMXHqD4MiF11Ch7Y5q4wva09p+9Unaxwm5heGN2Omz2eVt7mYbRHYmFith6
dSNcsmgyDXy9CKq8B26I2fSYsTYXzNWz91+28LFLWY3GRr3GwvxphMaL/BKgf5r9P3lrfH4dg1HK
zTlE+exmFTz+WEBMQ2nopj7avj4IuNo3btPkAoyb+iadxh3+UwLDz0vgNGR0t60bHPtC7DJFYrg9
51bgU6CPBXoIkG+C9O/+YP0aBVMh/mFoqOfh9E+8coQsK5NQS005Lh37NnOr/KbK4iH3IsTMY3t/
532Zg3pkDuYCya0VzZPg/jKYj5BOhrTVmZkcp61im2aOeUePkBe5dM9kWP1yAjq9VFbmMcMtbLX+
Aqm16lZBUC4HmlRta7DmA4yF2vUFsSW2EjC89xU8TBRl+hGC77wd/X+w3QERRprbflSAOvecyRRN
FdtoVzoYAcK5FgwAcGMXXCJ1+plSN3D2tV5MNIYaFcahBkoKcSPsmHVbB+A4bfV9W+muDa/z4svY
+qIKfIjIlLcuum9lN1lMwAzO2ytxmvJvgHSY+17EROdIg8YLC+hvp7SI6Cc7CJFgee/EbgraUfzX
YQS7JjQmQS4hwxnZ8XnARwpmchtp6zoNItvT4O2W/7mIc33ntZLKC+LBMKKcPHoEDx8TLwxhBWAh
d3+Dk38HiqWs1kj/1SXzk2ZtMtaZrXWjYwwDcg9p6ozDbd+OJ84kZPbc3XRxYrO59KGeXDfwQw/e
pa4nEcFcOBWqZwXmKeuDZG7s/ZzD2teZExsD+RBX74Dr7Pvgi2ci8+mtq5P4PXVLX4Xo8vg7bO/b
kLcwiqsR62lNxirI29I0rx26ZFolyfQK0Nsa8oM7bDKPFGIn9Hvmsp1GN/GlV8qRxysexWWo4li7
elC2odmLx1JGnYBpFgVP0w8LMEuDG04ijrD/Km1qgVhtAoguzE3US7SL38/FYgZvBkqJN2cgXgIN
ijhozkgSLlZyqFKxefltN8sw1jIwF17wkCyfW3jrMSFQLM7JIc36Q59qgNQuwQM3djtCTZnFgwxt
J3UsB0NIuB8LJabhCOkw0WUu1LySnhtv0giLddF+zEtOdBVKk449ycyUN3Zsz+gsDqwIyrSvDJ7P
GtHAffm79OizcGUMtHDdI28tLePvC/VrleP8QIsSYKSZM1yEQWVYyM34biSb4SL83avE1pquXpOR
Fk7hdx/p2Cg8wfhwG2Rvd1LHvYBJkiMEQb5R7+inZ5KU5STf0AZxVbloIEe7HWU15z9bll9HW3fg
Y1D+4T8KiaGc/kkJbzFqGZScNFFdkwjz5W7NiKiZTE1HCS4XlPi5vAZEHCMSPhctZntTCeOQT6rK
j/vfVCYqE87Kq6Qnu3BvADP1hZv57rcmMi9Ka7VWBGj0oY1nF+zUBgm4ePiskg8CY4LsxW/DY5pU
CExnLapNrgbkNvLNbPNICI3nzHnXubGxZ/kj6G43QwRWcYL1ExOd6tDH31QbtyOZSFDyojfmM/0I
5D90u/hY8D4alGdtyNiPQTpUc9CwYUYYWBnSrMakWyRxesWDj9W23AUeyKWQDFnfrB3JjySCfJA9
ob4TUpe4T+9EuqBVELlm5+wMkgRCb2TVAtISTa1WeQJyfZydqUNenko5wtKbCoBCzf4l9e2bSGPE
2yVB7I+7yiYaqn7682yeBTM4iTwcMFbVvRPa2M8GIhQLS4efYXuv77Job+d5SdceQils5bQje8FK
cpXj6Iv9is/JySZFmObf3wC4Zp8C6GYzmPWiqvxvviO/JrQ5wuPFIpkjkp0o0T1ZPjYf/IKKb8GT
PgMrEWsBE86qgRK71Upupp5cjeh8ehiBIb7kMZO454lKMq+TjPujbYa73Yd7RoVaRJtUbCUHLZ8T
Fab6Rtnj7WoFM/2XKdCQ6vifu29smtLnYX09VQishUi/8LowRQowqUpufPD53sel9Uu6yyQMb4p1
rP7XDU1tlgcGlCctZioFENq9DN4QG4xSRzbTULbBySz4kWmvIUrEs4zN0IiV9cWb7Ef5A/VYZjcR
sJzyHWUjYvwRzXUOwSgR38pZtSJpN4itivg/Uu1mlXSN5q4wFiyNsbNYBsNtYogsLV6gNA4atnu3
JPukvBbKpqZuOzenOSLmQYVlSFK/xPGKC0ogST7LMjbr/FCR0xN8atarLjEoOp2qB1LEeDTDffqi
jOKrM7Xqo43qKYvihyrv2E16K43BDO9LS4eHgtseI2V0kpfs9v5Hgd7aB3YTq/ABEiR8tRzB29Jm
7pZGFTYBouu3k1+QlzU0opG/tT34OfSu5p9OVa6jV/5Jntrv/RnLCwBGoYRxbbC14KGn09+kEjWo
zGp+GZZIE/fKVVIe5+ejMNctmd1Z9doEtNOgFlGw9MnbdLWPGN5J5MM5C4lwGCvRQi2Bdb8OIMoc
I1mrxLC5L+IptMgAjOV6d9AeR/J4OfpBFz+r1kojtyy9pYkEsbRKKgJLIrhd1G4rAQRsf693csHB
DOz4zRtv0Y6p6NUf237qzhbbtdtYoHpCHeytqYxNIo5z99sWNbH0WeEOCHSCejiimC3siiByniuN
ePh4pE7ZhY33MWTAw5a2gCr8pFEj1UUJpz9pxGVCWUCtsg05/81AcyaRKe55F+pyJMj1Z2GBScrP
/kiCt9pL3TOEbgurSEcr1vjCZ2DDRNnsa1eqV1ZNZ7RVxgAu0Zcp94ygjIKWPsuNUDJIQBd86Tp4
VZ2Rmhncs6szix5K40CkHbIYi7GRROMEN9okm+of+u8Trse/eGe/Ov9UTGsTR/0/Y8V6uVGUgLZe
JZkDwaybhKFC9/wNrnoc29U+8xNat4fXF/7q1pUBJA1LF1kHbqnr7qekzWoY1M/sBSFwTQYZSe+T
EpBnY5RPWAMGOefw+9byPkPEB7GlxoJrMujhMA4EkmPl/3sIHM3RXWTDjIEx1PCeVPd+wKfRH3mH
yoh/Iv2a6LOv1mVdoY3882zm6rHpFrZiaoy2gPfqzUKW/OZDAa6UWQWp3IzVZwRcHOM0UGlHxEMF
cR2HScTOagmHfe/zWK9nKo53l6UwTmBjJrh6g/knDEYZoq1HG9Mi9b7wl7inAeWJGb2Yt3wbOiEL
0XhGicZgVxItxeHKFIgcyjKC1RqUBK2nNiRyamzwbAE5pYfsFaz+952QiYasPVuVrwlkHtZi5GFu
ptvORFKY4pQIxTgNIg/wc59J6fbiljfyCeu+2Qk+jco5l1Yr8IJ7diQlyEs4QpTsvaXPxotobb36
J/e3yf7X9jITYXjhjVT/gQargDLlclKlfDXC6MDicaEzP1+IwDSK7NNbWTZidAkUtAgzTDM5pvVO
4Yy+IX8YQvwD+CFvLggy55PGl4AUTddeeW7uBOWbsICD2doDvoT2Ok4ywEP1BdPf8HY7WZqmpoev
D2uWUeH4J7RyPnip9NLo662rlwMiNRWuCAVCHukPF6GcCsz+i+KbfO+5AuWqDCgDnJpUXvLi3AIT
07j3amJ4C3CNbM2ENA+5QsQI98P7EfAf8tOH7JhtKEcFDgL6FGgcn22QRXr8Sby6lvbrPigkgUdR
2Bfhul31h8rxBCoUmTfGHii0XoOeUq9hU1QcasVg3sEspJrjXiwvcd7OOBBPhsw2kBrgS5nwfGwm
Kky5ZYeAcTsW9cnC3mZ6cGz1Ofs9rZtZoWWSDenwzpB3fuK1wmTXAea/byp66zH/nQzV/2TaPEmo
u+gj6wKcgDyOwQF1e98TimBPJOSOxy3BFPoSfQ95ANzmXTn4GHxcBgiCbLBpaAzhGFpv3TCrgqTd
3AKp5i2GKwIzJDsxX1W+IMI7zogpGfE+vHOZITfDEdq18LDhUr6iE1ltiwmRjEBVVObG/5+jfOaF
LEfpfIe2wy9Q2U6PNlVpaGXdgSORcOGBMZfAU7QZGvMbM0lQw+/ERrFG9LsMCqcixdToCB2xRuAf
7J0vNnTSPXLGI9EHBcZxAhv7P7joi+ULdc72PnQ6wuyZXuNFZLoIxrik5zooLEZeS3Pdzoqf35lC
9cpH2oAUIbX82bi33KQS2RODO0OX09cTx3YKeyu4v0tWSpuhWHsRFDb38U5N/3grvbUtlZ3ouLHT
1nsEJER9yrZRNPa4XLD0uPbUsWJcY5ndiZ9zp0gfRU39W/QogTFJ6+TRbDrJfdCcqpj4HNxbuFCx
5kcbK3gCuPOJQp+NSVorcd8cvkodCPXg8GFh/e31t6IyY9fvINh/IU5jPVDH3E1RKdTdWxt8XHpB
8GrkS5gWi53Uh1EuT/iTCvq3vtMNg+MQwMg/y7P4McnnaNSHXJdHpPPUBDwOcjIgKQhyXjRUXGCx
GDxmROtcM4Kv6wolK47VUi86tU9buhoXZXEsM3APleFaeECCDcs7Xyov8qiJMqris0g1g1OnpSTM
83eVfXh2CrPIRGyMnne/zu78HVkDWFBVjcl9yGvjzLzjzEm5Dvgsyt6nl7TU9RgQQRdwLtcPACeS
GII1DH10yBZhq8jb9HzuAMzDC7VMGYE1ci58uOwuG1UKoKJ0CAmVIbykp9uXne6rjvWuX/G3u3Xk
hjNJ1FH0QwQfRdxB5wAk9o4j0cVJmE4FnFrLeQ54YzCPUfwJ1G0s/O+cfTwotcJ4f7I9KWe1JQkZ
JwqTmEEgR0fWpkO6mZPvQbTBQ0kpAh1b6jrfC03zJR1VSd3NrhYyv7sEd8mnoOVJA4uFsZ1+jjyc
RmCFiJ/A7HVXbGpKEDaFJx80b3iezqgMos8u/OQz+6X6XXCMKybYmg+vv84bLvOx4rtdk4v6YbRi
T0xfKByOdXC/IsTzL+/8yK6LEz2EGKLSneY303Au5FFqe0sf/sKLwkrhV4nIk8g8p9tFjWpo62YI
iWSzgbv1yURTP6ipJ2Xa6QrA2BtqlMcSzUIkzzi1CdymMToThRn3NjKwAZ/8CDpdf+xL7MYEo+Rd
bEoKlKwKR6+6qavAadA8TiF0zVhelj2MvrFJaZ8zBER+GzRA6zTwzi/nzTKKkjo3ZtM5kcJ0cHHY
1e3mIXIbCeZbcS4EJ2OxlqAXYTJ3Kh1JPzaERBA1o2JjdTKyWbgGuOwdKp/ifICvZgwsGcZk9OP9
iyVOR60WVVSNipU5ZHCkK7+mq5+1dkpLJxOhv/AwoGG0BHT1aOFe/Xb6y/Y4eR49R5RBzDeCch91
1AsH5V9BprUVpjRgyPOKQIQtfiW3fblEhe7KpEBAc8wXBSGAB8lkkwpQZtO2K/4DDPKgQHNQ3kmn
ZxNByyGZ7bnRWoq60+bdxZ0o/I/koZjauFtY5nGd1u+70DsoAUw1emN0WU4S3ntItJJZqwJcmwiO
DbZRNbfmh99sccGkIYOw+KRtPCDID+bhQyMpqCpISlPCyvWwa+dV+U8agx4glGgMNVFmQhKqB8Ni
apsmcSEVuV1WeAWo6ZjwaysRJSHDqBIe+3DP7r+375Cc/Z/Yy1hTGfk1DFCbC5JOG/K+7tC0qSe0
102o+n4Id3x1JIZz1Fs3RkMY/FJzNHdRIlGxpSChdI9NIHfCA34brFLdeY16h+fL8kovmA4sfUI1
vzM3rog5d2gUIq8G0BGhzbYwqLqc/rS2Dg/aFGgMDi4sXIjq2Kxh2BFNd7Pqn+RKttIISK67h76M
+TkkLYai058zwiKTp1zjXKI7w1TM8qQHUgJ6Ziot4g9TusVEi9bmvYkmMSKW7FXQCnYvyrtxcXKT
MHcWUuIMcIjdeMx+c4LWNpHEb1OduAxJ/kekEa4G+GL/FVFqq8+h8aRpXIB+zbv6a4z8ZDeFtJoe
oi1gtnX1W7Dlp3CpNtxndc+S+GSrs5vVVdpdDgZ13ZK88Aez2CMdcODvs1L3ZD9p5nVIr7ojKZd0
g7dg+rFgw6uiDUEo91oS2l+i1h3P2qOGhsQIOcqqsQLP0XKwJkS9MzYD+ofVsZtz27LO5SZcRn9K
P2i8TKjDwo0CsKZHccjX3HYfgPA5W2BY50+111YK8vbfujDQ4/AxEgeDVGyV7vq3XN3AAjCk55/9
6XWSYj6BfchunhtURmOXQ2coRX8G8Hl85aAgcZMHcEFTDuwFKNbBoB7nu1KP1fKniNPSUE8PCsaC
uZP4yuMH9f8dWnNQX+n7iBlV9o4FSOVsGjttrmm2jsId4VvAdgf7nbg4k3XLpsBA6S5lIwApqou8
XEUWO4hIdYVkKS6CFyZ74LVQ2pOGyGomEvJq8oE7w6jknCw3hGiaklmqmi4BtQQMBEpobUyZM1O8
pBevEDIKq4LbMDM317R1ttFmaSE8Bej81ANAoreyt6gu5/osMt4rgKf4hVkrC4w4IeBlD666iP0F
hUPi10uWD/hNivnCBtiWV5i09B33+p8OjSdUE6X4ClhpV6ub11g32y8MoWS9EIkflU6Mxx7WNFAN
1GRUCIHfJpO+u0cv9XEofhypX7tGztQPErZX8zKFpjUZZqRPvMYWtP5rhaliDU/j3phg+7OnaVxx
K+52Kt2awpQ9UnVha+UC1CiykDwAvlAhyMN4ONKsqU2sTKjdg+2h3c01i9vIRSvW+pejtv/S/A0C
GqK8M3VLnevTeq72Hm0xKVJ/vFD3Tc7/I26Lk6V4BspJuBMcgx49GBIHBudQDLAgdS85CJ07bNm8
mfdEqYlXUPPZQOj35xMrEKqAuLKtrcRW2jF61O6p3RLSCWWKlXSxLQrXDCENG5FzAl5X2nYO0oyV
x1+lZp954h1imJBeLS4X3ZpA7XzH3p9eAPWZj3Jfq9bF4+G/+X1ra0lrWtGFjCeY+gQqu0txuvkp
2P/jPpk6dIcIKdZeMaxLv6b2GZfoVMeVEDlxCWrCBzKh9D/anBioAQDuDDFRLDg/3ksyLYzTwHzn
neEJVEvlmaURuiIVnlCdlgKcvLv1XMg5GNYCeUjOsPbH+5J7BjtEqqB9FYEEXzOXoPGr2lbcjEjz
TAITS58I23inBS28Gswzh2euWMrVHTzyhak4CidZ1LVXldQhus0IdQQWN71D4Q/iTYpbVqSGeYEv
ZtNmQ7Vb2joqMWUMZxwWPzfR8Dwxy5CbISseRDMFL25af5oG4x3vmVMFyasKhjqrOyAj2sxzQdN/
gZlVRCAtqlBRJgAP57z7t5eoMbL0ut0mYQv34mjABzqJQ7y1EARGJqAdARI8K0Ikd/goQ+sk9GVo
SmkUuyrLrLUfDK8l6LMJisrURd9qYO0gbYDWhegBOWFxb5DQnMdtVJEuJHOwSVVAP8JCVm+ylnBC
u30QCr5l+sg6uE8Kij1paiTRRpirY+5brb+uw2h2Ql1BZH2ezEkigzlELq5g/F09waGgKP8Oy9N3
i5cmOssA1Bm+zbJ8ik4ZhsNp1Yyr8YHCIWsswsgA6N++xWJFF6Hli8KazyF2ZP0TTGxuxO64zLvX
yaffrDxP6Xm3LrGFQ1CO4TGQKGgtVSCLlu7c35S0z7Fwz9qNCrke4gk/YMVGkR+By7KpCCd4Iokq
zXqvfYbDQ8gnaX4PaI1F/tE2p2B4Gu6hyeQCw7uXjVBi2ynUHfr9tqbVj0fTj2NfJcSmnauZnooc
Pfv2t5ZO9Upijjz/Py8jX/99B75DDtdeycxpUqFEuPoBaePKXRRlD3KgZxghprBMVkAw0kxZJH5E
aUh/VBG0HsXOuEUCQ34TaA9rKao88AFe4yPXw7yRT5iIZwHETuUxi7WVIjAN9aXAmstGu0rhlE69
EmWnxog/cH8cTf1skj6Jirjrz+LZn13Ur0pBKy6eFVBoQD6yWa80gnvI6r8dJhUOdgyvctuoS+Fa
7wLoxsugM84YKCZdYePhvyFMa6KhMj964eMaG84sySPkzqPxa1qMVawguhWOMnVL/qa7HS1cKe0c
8pf+3cOri0UrhzYbQRHDH+Iabj84GL/fymQrJ3DNQ3uu1kL5kGij5yALae8LNzy1iYOnFK7T8Jgn
3dQJXtbqzO6aq794f2G4HSuNdmF938OIATXw0vaBlGs3ix587+ECvId92jHXlxclirlIYpkmg+RV
yPqyA7h5X5L1BZ5UBS7A6tBTl5hXIxAtPxFhWkMQ4/R/lHfuFHHy+USJFrEqmdQ+w0KMMDc/fqUI
z/UM/1WgoEzJbK39xQ0gjUg+hU/O2E4ou+TwiSpOYXOSnJziq8Dl0ViHZeqV5q8tAicyxUuOx655
GD8AhdCf11CZUVo7tg6v+RzvjU1RIeapUAl1r9u+703yvTxovxD/rNQcWG/GE+ngr3p2l8/+KphZ
b5o5rxieUkyjhXSS3RQyXZTzrO2ztB9cYj9zpr/+zt8Ezu927dxM6T+qwUkToOYDFouRVBbtI+ej
GkwRMvBgN0o/r9W791rk2wE1RCM55rN7GauwhcHFaGhDVQddhOPC56HJNkUv4qi9fES3Ig+3ttsi
yp+bYOQTJSSB7qdim+C2OGHVQ6dav3eU93MaLe55dQeZqhLVdqA1hyuguTCfVfe/5kNU0zHRmMeJ
OEEAbHda0LtdkyZCBPmyu3Q7cpZmfq9rAvJt20Z+kDluSG8wdN47CG65zqM9t236lQ1DtlQBbAeN
A2L1J0+aSH4zxo+3WgPbxONRtthoGUyfP/lDFBS3rJAAV6c4k7ubxkMn7sBClpMmqkzFTIa4C8s6
mHOINmHmgQQNUxzOKpIMY01fj0hVYslC0hHToHzIgkjdv3W5bbhDSHnifgkwQ9YFRFS6rUcOSwoP
5+oFa+vMrbXODY46/rDegmzG9dqr0Xpsup4LXyLzhazH39U9YGRUnXHzfMYl75UrglVkN1x612QW
m7BRgI2WbsW6ZA92rWQD4b41g7GAqw7b9cUti00/ca1EAGWXfczoHg5R2Q1uLvIR850fum7j2v03
MxoM1AvK/2q6urCF+MkDKs915c4Lb38EpHcRwUVKjluOc4ZakzN7ZdtVUcz+u0NpS+kXWVY7BNCa
l+i+5vGZLMqr6/wiMGoT1gbMkeVi2CxpQJypUkt6kMDvGLKZ6AlGp8izaTO+9bWiq4hwkWcRiNTN
F+m2Xc44/sOmcon7zhP1sAuhQL1VBeh69lHfrl/FVgSUJH+MKHf3GUbot3ZJeE0E/wti8GN4VoOx
eYjr2tHRNVoVA+hetNgrBXTVhGDDQL2Kdm7bwcAn6BCcdsSr9JMYjCrZmgfEWpgCKhfyylS05ay+
+L1KbzX8Wd9hZPhuS4Acl1ev/krCq5bwseLuZu2G89ffgvsJr05EiOGYlMZcZ3wMGWOi8hl2G3mR
hxf2nag8G/Kn1mEadxu7jtmCsEXXNjXZz4IpaQH3OY0GHNtHYm0Vm9p6SrDjBW+GI7HbsQcApWJX
jvSEh4ihL8ZlQBP9ykmZrWGEnEqezWrFfUKxlcyTjTXlw4zPwcZSspEYUDsYwqrCqs3H5xUhrb99
+SUITJyBQRMAogh6yql3o9LO2eVy4xtaF+yTtLQ6wC0n0LZT8OEo6cA5xbGwNu5xGgcyVJN6ZOVg
0vW1wbZVGhwbEsWcwVGZu7Tu6h7DqeEftHeeyV1j532loeYL02yr81r0eP/BqCAekyra2tBKATmf
xCX1YQ42iNsEQwoyYLp33t4xJPZPWitESitGQnMFBmgWM14DMSUEtVAQD6CphA/Iandyl3ks6iRP
v7PnEPPnJWJgbFXcuRDG9vFIgN3GpoGIiWWFkuYZLU/gE0d9gdS/WiyI3c2PtyfVnwd0fwr220W2
Sy9Go4HioKRVzY/b16B6wZwu+/jRoVzzPDXLOEeSLcMBiripOmJdjwUoUIZVyGPEfnJtVxB235hB
HvnjLKBtUqUPuHWdxvY5wCA3EfrKdzoSTS7vvPgEdhDn3s3Xz+WXpjy8tL9s2CY+ADgK89TWNyVE
H9cPcdHZfYcFrOJc81ubexlEJ7P5lxJfiaAPfBE2xHIbXlqjspS4jx1ACGorJisS4jsrbywb2KYv
qE6SZWN1PWcKwezgqanZUJAlB0In4P6lFJ8M6Iy0eF0Aso+UBW4sPWEIzsRZGzJ3z/yeBeCnQHER
mNJNuMWekWd8uwjcv1TGMgQxSKGvRWAuTbiYaAEmwTEUHW2uBuJBGtawsMeQ1oPQkENAW/exsuuE
VZan1xUOmUc2/eZKAMe77I1oiK5jg3o5p/9iAi/hdt5bxZ2NPlAOYvEY61PmN7Hn44V4bc1NV6qL
tessH5ev24Pgofhh5n03LHXQzsSwX90Xv9RWpDiSCHCqfjrWQ6x1AmRLw+8wOfiVsA0Z0Vi+jvOe
PyKki7lL8pUnuGGPgD1Cp9lyrPRdKqGoyvrfAoaABwx9e/+zKKrHzX/O3DQ/zYbhHp+w7wSSZk7B
997n/n3udnQ8HLfr21TkK4As4J2O43nRMQ5NJJg73vyOTq0cSNepKMOEau4yI4o7YvoTpaFUIWAA
PCgJFiuzmBV/JPg4YyYZ1NvcXZGb7QRbUlWrJ9u0OIVFS3yCoPXmC/lZD28vTd9qlLIOW9FgIkIW
29N+cmcZzKoFDZIDViWrRBxqjPxw21rrHAyO1/WNOD+XDKYvg4Cr8Zh+8kTbCr0kFhF6lM/jw8tJ
xXRONWxVw2mY53xNnPWy0eH6O5ARvF04g2GOsK+drpPiIxdouzUTm+g59L7obLOtFokdhP13tyfU
IqVpNh8jFSz1SHrXY+wDlZH2OtYz1aqOJKPOwUYV9OFeOROcV9vnXpHCw64Y9R+b+LxvQdDFReNB
RqFjL5n8dgNj/p14Pv4VyqN9ahR8vy6RgX/mOgl4bxNBvAVI67DRNl3J2JTu6MP/Yhiw3V9RpUVc
pINRrL6YKFrnjjTjxMESA6+OHfsOmEjjWs2tcGjBkuZazrRrYpYuHvW1MtzzO88Vk8yr+NzqIqi/
JmXB6FhVA1BzFdqDttOb8aMoMBr4aMTknnp4sJyqdr7YomsfhZ85ZeIREvr83EZCnPkvD0v4DviZ
F0Y5U0sVDAu4Qj2Dga/d4x8dMEy4myw9v9hKs0v+WsINTu7Pl3uLvk+WKOxSkcpeVii8w73ZM0S8
Sr1496AJ658a2Bn92dytKlTqvtyxcOpQv/KcIMxTMhT20Yf9RQL1zlLY9QnyTYenniRsX7DgYQDH
gDncWCPKgEjJ6ewDbjv2JWN2Hrp6hm65/sofvXyXxvPzuBDFAX1TZFjw6924QHkE7m9d2udb2cYI
jrT9GNdkGXh9gWVKqIF0slN1UsTgXbbMDW32svGZxhghSwQ2VLRDOW8y5ajeitC7NjLodnnTvBW1
g4Llv8/prquL47CgutY9HCLrhycpDqBQkxRxJosdGSOPLSVeKb7JPD1PwIwe6frR7qEvB/5XiK8G
WAg/HtXAP2G/bWSCxSrMEDexK8ZnUQU/m3nbT/97mgc/Q9Tz25f/vcpPad/Bx3kn2hqHUxDtfNwd
KiRwSC1+428oT5IleR3k3cpEPIiQKzEZauaUtFtIzT6u+wkOB8Im8Ijgknj82OHwVXmfGbBQZjQ2
xKjHKhqswQPTyhAfGorwa7/355plxy+Tp1spyQAJVauaLy0n3u7rTA5V+0ImHrwyx1ZgVihR68dP
dlDIZpNN/shkahEamxx4vg+LTSBxS8QmcsHwxfX9Yu2snhEQs/J0jvWWtvDFPlA49DFJCKEvUuG3
iF+hNbl6A/tmYmNuWlNdpZanE6frdWkiwIDeLSomt7GAA9hxA+Z67pobisE6HFa5qVPW/tcs7BA1
RT0Iol79ZCnHtVMtweS+NIMAq0zmtS/4AU8H2AxyBszFF0dGuz6K8b0NWcl+TkG1l1ldqjl1ySIS
DRibpYQt0VksN3eb4oXYr8OvwBf9DAEaZsHfjPZ5wXcnkm/hBrij49P2jhiw7yzZLndZSB6Nc6of
2yde1qsTAZOKz88Am8AArcTpQHYb1D1doImFMK3xVuG17NCgN6EatnDlM7EkK21tXkeNXPZ+HBZr
5O8uxfxFpzdmdj9bDbIV6XzDFasBsdQKZTJQOx8/HjCFEHrbDe87/liMKiStMyeQhRAqxAfUW94N
mgn2Tz4FCbNTrkdoS6geO7Tu7+rdM/uQpkSz4PH21xEjHayX/l68Tq+SJGYqSARB9cEy77SnPKsE
8IJRPXQLHBLjO6g/bHSD8QgTcEPrg1y2RvDTImWeDeHwRK7D+wWaQmwX/mnRJo0kG2HLTo6uIVUl
zHzuO7QXaN5JPGLWylK6x4x1IzXu0a3Mr8Io7QRHIHgOe/pg3iIM656OdpwKU3Y7GhV9DAaQkhHw
o9POydVGQtLU7riuEjiBambHsjupyH/dSPJ6lSbCy9tpbS7frMiS+lI7BxK4kimCvcbGi30YmOmD
3Ptwm3SDPuphLNX7ukVGcYCgEERlRMVkLwufOOZVgXK9HvfCjJsLG0gqOSfjWhZLeEhx6qPVefWb
OopKy1AsD3MeESepFpPcRYkc4+k3C+JCzecuIsbHFMl3E+Ej91JR7DEzHycnVgGNlOGpLhGcaWyF
7S48jdO69C0hJ6tf9PwolKBPaQ6Sxs/NM3zqK51J1xwXDVlS8XndRi5pLuOmPzDatAb+aJ+XAjt+
uEJ+3J0Mr+GxRTphb/aT9fhfm2SeVAtcEKTbrzY/j9JiWHFPrh86+Ycc/kXoD5RRdGRKpv4tw0j3
XcbPR1N8zBgnN10TslSovx1Y/z/fp/7Bdji+0A78mfIs57aMEqDbaG5MJhkBjaI6OWbXHPkJSp5s
eCBm7BUGwwhjfZMKPIX2psDNt7HvgaippeVUMTZDF12HzQEdhbyka15s3i0S+fN4APMHqz5Fnawg
+iL6u9RGwfHgUv/vffXIJsQb31KbGQdrS9qTHDvsx0nXgWqQIUTBsjDW0rrF8QHjOF1I0Ns2M4f5
1uXPiWzdkhVb1AwmFg/WOMGMGyHyHLjaPB4udzNpypJzZtVQORhIaTWY0FUDIws9pQXF6rBOhZJY
03KHmr8YlPADwq4+5gFw+0nPcvwc10dHJGymNFSxHkgy/NqiWS8eM7O4a8fcdfbzJIfjNZcRidRf
v7MsWaREt/0MfvnWJr7oWIXFrcJlhoNCkXPrSir1H2Skn65xZzpukepyuQvgT3BaS4u3qIh8iLGs
kRUwUXnRBd0lV4YfIfXXlVDaW894pQJB1A+9MdeoTOFYgvB5FQjNkSirH1ISTEhaietB92xG3Gp3
fJp5q/ZDE/TgE246PQ97D68NFhEWDQcZghlfE5COUMWxbEE+eSlR+JM81dEEy7SIS2aCLMLTyZj/
2Ig9nciDqglc4zRtHfNmxyx7v2ugCbn523WHZYS7+yDHzMOf6xsO4Go1rHfcX+7By1ospvi4Lsxx
Xi9dcCbiXFikWsyNmD9RO0csfXqNo2foRlDu+gA6l5QhDdDGYoAbMp8YX+kSA48EDB7/kKs15E6X
pfQ4zZFGE5waxjUBvWTjkj60qJ5aVvrPC3/VRwIIu4piiCbKtu1qOf34b3kew5QGDbdfFGQxmmMU
ykfK8ivUyfN/kYoXbVYZaQwSXH3ZflvrMtr1S9v2SppVhuPAi1A7jxv5UlhHjUI854CELBtG3Mu0
+yEfdwAewLy1Y4QYCslDkASpv2p4ClugoACW+APXRmulZmvxNv+sZz6zltPrZ7s6MvHORZDtCtwN
/H5dtKYcVgIr+30KYEk/68h93vh6DMrZ/0cE6gxFcx/JJ6yTrjHKp63EupFC40/Yr/ZJp9YbAnVW
i3gzYOcmc4t67bxkD2rIwC0sEokvIjLPWy29lCbZozXJ+G18cD2jpHlsJhVpzTfBd8wEDRTee+TW
w9PBAzpqmnoDIYfJ38rQi4OGkOpgzrLL/K80Fae9Zv1/3VMav7Sr65V/tffYhNeL8pz0rVUqJYOw
ocdo1oX8rJPFFOyJNEh5r6s+64dUDat6tLODTb+V3d2T70OdNDMNW2QE/f7xnZ+vm7xHXGI2GBkz
HLtzUnpNBXl1dLZOaWjsYE8cB27mTo5u9S2L/lW6E1qdK2e9vofvyRZh506ukR0UhIxhsz/ad6IA
ZW7vgFDS5MXZs5/vmEPvuXDhcpqVOn0juFoclMMkjVxfrWSoxK3gAaLiEpKeQDKOzwmcN9lUcULY
iu3ECUWWh4NwPnTBJ3fFykSpc2Ccv9u0tu87gAiFDAsYd3Th0gXzZwaqQ+EwnzAo5G4pJ8hO70x1
a/J+E6p6buXGJ8DiRI/PUgZqWtGPNQU2xKddN0RreH+mQuXv4gYayv9Or9TDOJKL15qjErGA7Jjv
l3Jck4t68gYk7jsTfhjIrSMeXrbFjgMB6DnIuptVObS0RA+ZTZ4pRnEhOp/UvqtXd8PhsW2oiL51
KzR8ye0o/T/vAfRQOtRO2D6KTGSVXc2NRA4KZBuyYToFt2au+8lKXT46zLKV7k+FYHXjN//YGmYR
+rKMfnGP23PRIW5S/d3kJh1xZ5XM4msE8EC0Lp5fsTtwvJktvnuO9+9G5kOILceSx1uVd3KnU67R
4Eha5aWm9UWjoSGR2UBbvO6tu/TENQGAcCMd0NUyrQXQ/L5D4sEu4nOQ0CroU9SzQBMzreebp+hb
KcmbRvTlR4ok+gqI05jVSpaQFgDZ3HAyX0wC9U6+3m9zqmZfoM45x8bDNTmzrVdPvrwBhQJ71h6s
7IR/zCBlNaxfKXs68QuNSmLIoYolY1KTqVdkJwWnzgjGIDjGvWOFHl0j1KeNnOIe9NztrRhKEJ16
jdfEMCy3j7dCj9w4YGUXiKGuu07o/z6bxut2FU0p7nvaHT4+Fhv9F2qqMX8dOcQ78IFMTYuj5RLg
0/4QMQlIENwJOp2NDYiivuzXg6dDBTgcKiI3OWiWIiAZFqJqQAvGT+2t2IUp9i0mCFhzTCArGQ3V
YBm4f9xaDN16F3UE58eWXp8I3rvAN+lH/iEHnoA3xgVGsQNYunjkKFob3mjqchLinuYDpKKZgtfb
7hx2JBaZFQzJ96p8ZBpChkMS/wX0FQVZcZqbTo7BT/2WRi9BqAQQUnnEk/FBmPJ958IqiYLeF8Hg
6TeT/514o9kyO5KGUdpB/VQYp3GliuDZ6jwNZoChwWrD0bxDX5B7BcMMqLZeckXgWV6/JyAeSeFS
N9lz7mbBcef2gFwsMZulxXSfsBiWWIaBYAX+ICM13VkKiQkn2Av3kXQ9Jou/n3Yv8kJvvaL62Nrh
lLCPDODKjDTR5sRRCaww8gcfwyQPtn4EJlzrXGoduVik17/Ohp7h6vd3xPzp7M1kBH+AlkOqMVNT
cvGukB5htsL8vWYWbxYwkphl70YaBQSlv7BlX/qzMJ1utRgkGPjPAKhSIncm2gBAf+0MEyGiWB8A
CilfRSarZtcwS/2qn8pUlpvItbkBelE8gSufnZ8HB8Rx64d7tjvbKvxaPnVM1GgTvU791D78hJHn
80TDlf9sUQLxgaiDtLCiywodTaWw9u6WaqMiD//pw1MOFX3+E76YBzy5eda9e+RUfGE4MLNzS8sa
VKxg8lqGAkMVnOVOIRHPoHi+z0xOF6B485WQaZQDYcYvJDuVafcZYPtYqxN8fcq3sBcypjpp0+Sf
fcugTHLhCBG5TmVN0WcnBkmkflY3IANyAVPZxaAkIdthyYkUBBCdVYpu1yKdasHmTCIZ5QB4sr2+
KY/0CDqdLG+4mTabTkmNjTkTgbEuF2dBmLd7O/wpIERjT+RtHEx3UyUggnxJeSVqGMKcWXKO/O/G
0oVHhNtC29pjwowNEKhYbApsJDd69pKujqVxYvNipJn6SAx18NQapsjIQX9vcn1WUCsI6BnKvm/p
/7O6bn8+mH3t1jfq8b4+XihAtoFUhL3glrMs2hNlVahXH80cUTIfon7TGa4XSrPoWVN7CqehG1TW
OycBS1rM7We6UVt92JI5Hwewh5VAqtRT3HWuroAy4g87qeY/uBkn673fAksC4n8vVsLeUy/v4rBU
s2LisGKOoJen/ZQT/XDvN9st2uedgDc6LvrT9BDZzo1nuNBHpXTqj09qz2yKaKulkjFf72/Axojj
y31aUmoFWiRj8Wdy3djLS/Cx2aPVnfC7TUjxtpsTEbGkTp0qjgKY3k+IpmmE43jPkWkzja5F8hma
Mn3tK6e5IIpdXjykD4jdMUUG6ql7eFzYBeAl6jbCdUwQMdlxA5Yocftj2vfepR6oYp2HdtU/K9Me
txOKlOOBf/g6OmWJmDJ6lIYzPBfLAx2GTGkuQbb2luIlcMreT6f3ID3qVL/x7MliWsLeDbHWV537
D+dRCFm04k3DNqWyKTLFI7v3M1393Ihxub9JMI0KZCdsz9GD/d9QVlzg+lWdz6+GKgpH5+/xld93
dLyIXv93lFfoju6wwp3ZZdnaDc5nlYN7zysoaolWNPbsVyZ89fTXxJ/GQXqPbjLwRBrpcCJfpfDf
Fv4AHGPuajxEoS/GXDc1K0Bmt9P77fvyJ7KsKvJSXHmxquo+XyKbKCa/Fw/t32YWzNHguSiuTE2l
plq6sZBTtqey2/dtEHeJumEaci5sZIK9kQp4rMeE8AEbx3yM8xvxWGFxMgO5p29t/TcmH2mfjJ7Z
etRxjAH2F31rOlK6fQxFgfJoqYt/P44VpIltwpBqWs+lFeFuTNqTZQsuTHu/G+/bkA49Aagf4VK2
49xyPz3THiS+ainUwIvUfUgLRYLrkqB5kdXVnLDaup0qAUBEVPe4PNU2e++XdLNOf5Rt3THkldIy
xV2o2tS+IzXzYpP8Y04+Scmk7KK+ncg8y/bvOXzqjpoPj3t4tRCTdrb9r5AHZJhU8uj9u9SaH5sG
6v5MfmU86TlpAksIrPngAn79JXfvol24+4H5/oajt2xHcrvHADPkaDdVgLrmcO2hsjfZdt+S55Ub
PPJEHOVS7kwVs12H0pGj/adlMM17qMPiJqLbqQSzZwhQzY2AFJVO3bTA9DdXDCB+yxPxB70qeJDo
XJsn6IBqWnxwvzVt5R7A666Sdhuw/Yy+O1p/MiAjpCPfRuNU1J8xVK3Ftjf+F+d4pVbprMkpLM6n
HJ4bbZa87zqnp4U3TIFsIGDW2qnzjiikriWgn8mgp8hZOg88GfEAgWkrWrX/OeY/dnrdoJYpd+AS
yGxc7fzBOyolr0s1MDhnVDLopR7yxwIwfErNVdqywjkSSe5agafLDkgXcWdQMyZMmf9V9XXrkD0+
/oLpfegTjsp0w+tdHtsl51jVcX9L0R6pNpceemAYQTinrTMMe7HZJ+vW0cHun6qevmOjbSSibCsh
jAMTuigtmz9tEx71evZUSqP2iZJ90njIqVdlZk2lFwNeT8b7W/rwxktprEdoxKwLPY0ndDZCUi3V
u12ZSxDxo5rUjGMGJqI54liLBQZqNi8A+2eS3y5haP8aPMI6+DPmkjfCIPT0OgpY69lH6U/l3XvM
ZhnhCnovd0kVCD7maSrsn1pFhwsAy5Hnt3GXeYaBniQgy4EWmN643L3An7YMVxWaDnSoJeL2icmK
yvWfVRTfj5RSD8LlP/4MiMuECUgIY4QGT29qGo1oP4Dn+ursXyitFvPPxl2CY1pAgHIby3+nKpnZ
1DAlVoUtkKFfpeTUwYSjrswrrEDJA/sFBqf7EpdyRdB+ol9jbyF1LhY4tRAvquBcEtPNdFpJnCaU
9gX+K128cEujD4sVoW1Wpu02Yi+RUyHCPdA6IlPSXE+ddb0hKtLngUL3lIkDWEzmP3n7i2Twrxgj
xVBBmq5pDAJRfVMNRcviCEoPaYpW4lC9pryS0APCyZtjkkH8Co02dVrVTcdrUd5rtwgU4wBpvJA0
Qa4bji4YTcp386I8MLMA6SXbdD49RBPJdoD4RK0fKacYpmrpYSjjCe6XPqXfgFJ/8Yz6Sgv38NTR
p14gXXN0umrT5XTINrnhCaRTEEIoeDxapWe37WEqQpUrNc6iST8Ua2gssVSSf0vDKiTqtInbZcjq
bIPFZu/RZu3OFaBGC5ukRtMw6s1UkRVXmr7dYrYQI7riF9TaBASJKyQ+j7zt48Y8Ln6IfQPTsJpr
5Pe0ITPuHzXzxSHcWKBbPpCXE7Vl7qjsod15+1K8Tg0wblEqK76OrfdMb8HTuXMkOJnUlslEjGwm
PNW2UfbvGlOt+sC4HvlP6AvFGXY45r88kBJmFglUeF00vCpwi4MxLQBhYH8Fv7h0tq3WCUZIaLX7
Yv7wGikCHVE1hmClO9JDvQ5KrUPMgidSfgp3uBqYmE9klKkA6SI8qtypOwr5WUAlmTVX9Q5Eo77Y
m6HPYPJ6ET6Wt4MjpD4hFHBfLq7H9rbgY2plX7XHIU8O57mb9ePIzBTG3EU8FFbWUgVokXWn/0cC
whGEgnsQlmplZqxeEnJtxCvQBgS8yt2abOAciTX7imGfM8/oWH9DiU9l97qat9VXXato9NERqFfX
2bbNQcBupLR0VhpRPm+9mFag1NC1twSrZJwn/nhQsQqth07WOnzFJjNS7O34yqLXOKBzLT3AAYal
mpl+gmOuDoK6LHjiAE6dt/uM4p4uy4DfucjDqKuocgLXpy0Cc5FrpHHQQe+wWdXvVOlRU0VKfm4E
PMoDYyBJZw6yZM7++NoAGlTcpJHw8YhhGItVfZTPCWAbOZw6azaxkxV3DCJSzgD2o0SvKcEa0Yen
6TXQGwT9K/3v8ngmI7P0PmqCOZU4BPcP20+Eu2sEkIzIRuGKXMOEl9AtLY09tGUZvlo5AIk+yZKr
EHneDDezJQEpr5oD1iK0M2Wn0xfUyDGJIKSBQh4oPnAwv/D3wtwXd9oxKF3Ab2Xw/9WUwb5wt16p
uO3ddbJRCQ5AikBERQIPBt0oegD7zXEoP/o7qkkEE6bHA/LfWvfuri8OeG9b9c8ABKBcDTOzhAYr
b/k3Z7VtNBCgL509eh/xvE6mGAzECx0xxB4XPaiJrFbpK3RiidHg2bab5l7ggq0GckF47MxVQvP0
jTEb2P2rbOmlHOASrdjIwvifet7DsV+opi5Bq9U46/1wInhLOGq78zY5DJva9Djy6eCcRabkshQ8
fLsHABxSV/9G5Pt46Gnl6i9NWaGu1CnEJGyWfSnaRzpSJfNcjkDlIb9Pq0cdn9fbbCpm3b3nxIRc
er8AXSSErHZ+msFSsqi6yYxBQcpRqZDx8n1shFshP15mI82qaONfZ5Bwp1IMtFIZJv/6uRScNyv0
3XBnwDtVw6AsMULQlK/KoX/OnYAu8qBfLL/tFIxafAQNEa38cbtKA1YGc9PcpA52XLpQwFDjgUcd
z+oSAwe+YzhpbcnlHteVEGxzG/yDl440RnAWcZnk2+2gSmTaD5N0JNyc6lnddmy2hCMDVUIn7Cfg
XxXRNk1SqVbgtJtY8ytXAa1Na7G3rTFwhnu52eAHGFOpp4CF1NZlewVtQZuUtgdKdk611tj4zqen
nVYQqnHw1L/Sidazic3aPoGizgdZmIGIdvD5aM1sIkmSVdXc3fn4jvoK4sN7rZ88aTleXYHebAPZ
hZhMp14c1Lx3Nxb0cepM2qXMIYeFOsdA8vZ/eqUPRdNcpW3PRQwa6tV0HXBJPZS8APFUpZM1u4D2
48+ubkBLQMPlxYV+Ckd6dp/HHeoen6zMaSCvG6WdCHmVlFd/bn+IWa8dcoQQ3Sk4vn0x/sKyuMyZ
j2pbkfSKT8duVATCFkIaeHOiwHCFNOraOyJFoEbm56/aZpK2uSmYKiO5G+jNFamwujHAoIL9ue73
VgPpabTtbCqW1/pcbOTYXqVwKspgz4YGQp/HbTI3q89v/UeMxuz9d873iyNzFGEvoHegaM11lP+t
Mm7EYRDK4h8Q4Uj8XbmueFNvfQTo5BabPe26PBbVt9tF/bJPNBRinQYXxL+NWcQd5/RcwwCOgOH8
0bY20knBVunUqDEhsvZn0GLVh9IgLueR0FqoJnDCbzHLbrvT1YlP2cZ24n1J22mCvXAK6gLH1Ujm
FCVXgfpAenXFpmN8xNaJeMrOKq/erSr2hyAHdYdG0a09wVV8KL7tktUUIodh8wTfvwHF6E9GiKrL
bVshisaxIRa3QJAyzFwXb0N/5LH+RWTrfpRI60qPlDpZMOf5Z+RYw6DtpFgqztC4e5Ia+7u78lk3
KXWGZ5jrxeIy8hQQqAYVtxKiihDnVFJB4QwQvTfqFRcbKrGTV89h161LoMZQ1KnHqMM1PppykAKW
l/4KH9xROlZv7mn07O3gAG6ySywdIwyJlVGwG1ra0iB4Nyi16ks/FoKdE8h5YcbaqQda67ASY1OM
eIXOWu8T4GvSFx2vXyN9FJdnEJRH7ksNSatzFXBoHwl4ESOosU0OXxu9W/hknvLf1WhVaOt7W4Kk
9lleUYJEA0DTIWbENnhyL1vI84yxJiNXCm6JY9mmmErXXwPG8ZBnMXYAigOghe25rBE+fZTTsOFy
A3VyTGjnEm/SXU+ZeiQgOiFnI4o11vKdEkIH2lZ+WUAMlL096h41aoo7y8L7XH9fZd5fsNMDQD70
yDEGP2XKw9wSfzs+Vl3lWHNgWZWcdotiEnPpasn6Z3H7lFLN9970nFO+pBnz2yeXMXVk8N1BbONA
tLNJ4QTFmajZwcXr+ERp0vXGrtkrXbprQClfLwrlyOOHNOpchoDv3IJbD6p5p9ifd7ejXBdWRPo/
YcrI0dgV7HVxrF5ApWj78ZckXK89xNlsR3Z4Ju5awklMNy5aHv4dVVGLQ9ciHHl+iIK7Gi1ZYlfb
fAMcGlhutgbxCeT080OtS/yGm79vcX6KSty8FVVzH+fInhzdDV0IW7JfnPbZeOsnCHHNeYmjLV9i
FCgq8QvrcZDSSAlWViXocWuNnkdV5/1DMe28RvQ54I54q3WcxSwWcoICUTdS82SKNE2JPrBzNj/U
0CjzA5C+XzlvCcmZm6c4nywcqEEQgaKXcwME26mwUTi1KOoaFos1OEGqCEtzo7KVfPLodCi0sOGE
wD4FqYHbHRx24HPeZfDrm/5kTf4quLISA3ArcHbcj7V+riKxzQVvEsWPBio1QM1w6uH1fnEdHPDs
KtL8g+MwmD7efMHz2QtNimiJTiCkDjSanNhZqBibj8ssrJ3n+F1s/IBl2jITGl13GKG7XeGuRrqv
EoxFDO6IN+E2TU6chRLWsk+k5CESnBH0IzDfMKHCnv1HF3ECnXj7UtOryi/WTqYHeSCID88z1QFT
+Hr508X/1rsscnQh1zvaAGJQ3ahUSP6owSj2+MKacUPrj460m/FkfZfmX5VYJNnG/dbt+d542GBA
y2Oye1i0jruP4HxUr1nm4Ee0mx+pO+jptmCFRUEhq59rD/vEYzY1iqPYPoeBpGDRWYQUy0Ta1qzg
bQGKje67Za1Cecgq+V8BjIUJd0Me2zPuFJF7Cn9DZR8pFjqdunhF3Ip+xVMaoqYBvdjekmxZ/BmB
nu+2nbiRKreS/1avO8FgXv7gJlOvCbp5zXNi9iA7XWb3IJz7BmlJK49p7KGLEuypprU6ZvcOMs0w
768Jf7l/DjKvo9hyYZ8hQ5R4Ezyw/SM8+Z1XnodIcYNdqrcptZcZAYko5tJlmX8at9H+i1rN7EVR
XkjKvQDbk4cf7sjNbXNCwkv+v4YQczE+yRoXn1ifgBaccOYOIAap8yjO7jHgWOS+KViNr19TCFpy
pugRMucxuIlyddcOs5j95frRHRe1jR9Mv0fgmhsGJGt00F48Icl1Na2NjZtmCTzKVCFUL5KJT7EM
8j9n0wx6xgcLJ7mD03oWCBKjxvPLVRRXKKhjUhX8ENCdV6GmO6+sj5drH6/YwI08V9SpgwWL4HRb
YIYGsoWp77QhM/oNOHCwC1HhZSzzGdXDi6vZbOqXNv+PLcxycPK314CoIA+Dtp+s1DEKeN6qxxag
FzLIY5QUKNV0wCk9bQOQJ5eRmqLn+fE8kPsrAM0olRjHUJvnP0dKZure1UFZyB3AczgyTrc9Tca0
hQIW0ufHRvwr7bJt4+L4TZEEavt7pXc+l01FesUucNZcGUHBdzNck05xp1XJewVdcMLRA+BLh/lQ
ug/TcBGFzR/fRse9xsdWadx1xzrg5t4V6VpNNlNkXUn7Bl/wA/+ALPIsK+325D8hiKjC59CVYewC
8lJDHaBVHT97hXiYV6uFJybzWv6wcwELM+qmu7OW7lsM8aWmJjW5VAK7lr8hsZsyj1dSsfW6ynqR
kPgpGiKgeETtASmRutVjAOkDDUeYNgzBpWo6Qnxwz7w5P8+d2iCgUbF3Ywd9C5afZw1emtid6adx
YiewnsCd1BNJqj6A16mQYrlF1IhzI+ar80Ps3DpyWaOgekXEZ9TUYVO4tkFI6feuv39ooa0azlPd
saxec33aZJ9LVLACl19j4tDhRG/HenlIZBLBNxWHDAg6RvI8zj9SrLvmP1sqIKU7vSZL0Xn7BsEA
Gxwja4bnx8GsMMq+6LL2hHykel1DUoNByD/NP+V6TGQ+j8BRpGPVgdtAG6c0NnP0Dm4SW61s35RC
u30ED0dzLOkt9rTHe6VfJRMUWznlwTKOXcntpAQREEttll+J1ETZuc6Xozxtj8vHefHj7i5drtcc
AhdsHnkWFhLl6JbKUNrQSBKDHym7ffiXyjpkPxqKqFClzsKFGOssOdWQJCmFX7IWAd5NXOAAU7VC
gPfe5IciJlCqTCOj0IIX/u1Ytl03aLqZK329bid0GpqTZWsN1kXdALGK9QjoM3d5gIApOK7hkrSS
AOZm6L5HJtqZnbAFB9d0oOk1CrxOwDvVPUil4FnPcmnBqR3yv5hi/YPycMSFQlM6knrveTl1hvyn
+7SJcYPT0pNVkp3MsMD3xT8LkvhAW7q2uaCL4yWndBAPQ+1TMiMfdJK9Id15ZTYEoateOnfkqo9S
h7vtDNfJEWtNs4mYIxHnn553URR5keC1pzihUuHwaDw3nSHdfY0SaAW8vXA464DBMmLJs798tK0X
fJe5WiNGs3UwAE2MT3ctlxlN6E7ImsW1+odAlvqtpgk88V/LHS9sz/qUtEzTBamRf5j2spAe2God
eo6ZdkzktNAPS/COXMc1p1vk+WL+xeNF0KA2X7yiM1hHfwOpvnXzqHOvHeqxy6kJg34eUTf95pv2
7N+aMOaUfSSVpTKjYi8VJa3hhpSFa1UrN7LjytRreEQO/k7O6ISeAPeoMtqSfS3AkTytkOg6/r00
qkYFdy0Nt9DTyzqL2oYeYIF9qqiK8PZH3nVBUCytymtqzMFaoGqDonHZikXdSIHOY3f/rVVyFfU9
TqUZ6Sab2F6sfI2KxKlZPvNIWz/OkoKGo1mWWyHdUFvt3vsHBIlWEhabUigaORb8lRB4Q/kkeiqN
PPxyZ3qhSGvq/Qpe+zH82VL7CKpxsH66IOIqC04ODFLEWdgoZ/1v62O3Oy0hLqD2dc9ZbiEqtHHk
jlCDAdVhlGTK1ZydAqQ34UBIkuyjAzILDvnKN/zYc7NKVvts9SLsHSdC1kJMD36P3gZ3tUpTg+ZM
XMU/VDLDlbqy1QL4HJFTSzqp+RVAlsRIcfCNT53PqPFd6DgrTmDsY4l4izhS42UwY+T1gR5pPWaq
JDza4XsgYS4fCZvKFKLIlJ2x1AekHjP2k3okapqDSpemeFl9NMruaNx7bCLD+pRv0qq90bxt66Fw
4PtfpTPuYoG5/bvb3EGaPQbG0Z2eK29bDoxtRuYBhrZXqZQgduLaCYZ1Q3K+mblgpyqjzQ7cmq/i
hQQHOVM04k30eJgJHfrfy2Jc0f6lpITrxUmkck7hd8n6Lz2J1YSGiGc/khbLGwrUgojf8HOa0NFr
4ocXD6os6UlouwiSsKvbkgKQLV1M2vXz5Y3mJO3457BvaepioN6g7XzZVfyNYDZgdzoIi9OrUf9Z
WLe4pPyzXDXsUYj2oQGn0/tFf/IiApaLkmNgjTr6ffaMK7xXD17An6YTkfZxL2vqhlnECiVnb0tI
cu7Yd/sT0q23Sg4EICGplgwPF0lPcevLTOdUfbxSgA2bmjqCcGiClp1lJXjsWtdpcZMJzJu1Zf5f
e9k6ab6q24PWhaK6nhWDH7CUsZXupGtRfdeCH348FfspOZxvEUYNzcO/d7lgZLngPAfYHiZ7Vko9
XSCUs/oSYbx6WpLZ8qWe3ZohI/nB1rPAnPmFT8d4sW1apfllg/+WJTMFoVFXnfXQyXNoBVI1b6nH
ifgjqONTFhk8JN7Mg2JJEOkRR6r8CpLwhfN4SoHo/El7H6ZbZUjl5+tuSWE3zN0M4C+tRdU+jE//
kIzARAD86m/o01idacp6AKQktRlXIJzgEucZDOQzbtYnqaOqqtc58IuE36jLAZwZt1GxnZbLbeYw
XWa+UfoCKw5T5AK5YTDsxVEJs71snl1w+wiyaM4EfKF9DW20c35s1vwGUOQkFmZWtvpURgjBplyx
66AgOSo02kKGFWTsqP0bu/aIgtMJ7EsU700Ih+2ZydQ3JP1/bj6nPWCO02k8l7/G1Cnp2QDCSOXI
nFKlUigTElLeD+Fnxk6yab8AVhVoF2A7WKwc5tBL3+1purfLMI/kQ4y9v3pAshHVtpmOjReQHcO5
3W3Pwte1ppD36ohHyE5S0bBzV7OCwwAzh7pk1Bjyb6V6YNhVZv22Oy5rkB8BKx1e6MxDzDUepJ8e
vph5Ay5K5/ZtxOUuXWfVa7k5QSmv7Lkfjymojgj9kcdMxCQUs4VJRtrnvcSRBKGOK8wV3Ir7KaP1
xu4gs8Jn5LRgmFy6N7vQfo+5jR3g8VXz47p9kiAoz6dLgu2Z7uG795OiAmLdnyroiuvOq5iYElG3
su4K7OhudcOSdmUH6hJKrv2KS7ewXsQCTbhyGYIPoEWa6V5Q7WdI3Lw6uMRvmGYtjN1euAdsjVyM
6f1okI4/IG5O6AtYVftkoBvGyD4REVwyzm6pJASD3a8UJzIWOgAL89Sc6ZHPCz4cMH/74d38YrGv
K4rIQuRv/Ra/habwqkd2nbojMqNDx6TQSKWZvaV0Wo5zVB5st/vAyzFtQBAI3LOB3yOa/6c/ucL5
sGhDcMG6OFaI8esf5gb6zz3l4L3JmHLj+ivboQwi68ZoHLnoTW1ouxCJNtDeOc7qkEwHLvsQcqy6
S4KH2XcnRwMCSOvoXETNzehfkbFN8XrfOV5zYN3wgzcZFvacbXvPE2TqAg1anjGJld+sn7dCqYQ9
sUxfgAsQSsojuNcCE2OUq6X71ncSEkZAxgCKk/OAAfbJDayjQRvjWTsOwlS1K/bw4DLfocYtW0uy
4DmpFsfp91ZdRgSIvxTdm7ThSHoLrmEiBc79q56iBTAXohOE0H7ZK5uGrzrC9IvUkL9KhNBKYIO0
uziybfNviZ7y/JkYT6XkiWV/7/do+VZGwRiRVlfIZMqFYr0AclQ+bxiLxfOg9F/S97sEw0GiStDF
jOXV3tDl4AcL9j58opUjrgZrtz8qGjgXIAmSNPwCssfb9dnSDWFKEUDpsNGcxlSHu/V4IsWkY/nH
F2PzylNUegvxJIJzdzIk/vpZ8Av8KJMQa9QidcKbiw0waSy7mzJGTruH3ABjIuHuvZQSeCVkV6dW
oGtPHl++TphtC4RsWTbnj9SR/4mK2RqAypMQp/uOnANoLFVKTNCJVMG1lzJGzOXnuC1H64smktIE
32+ezeGW1VTsN2DA+avsS0Wwp0kv9SeorHDYsMWYBz/1jdlkzHeMTo71El/cdNoh6WmPMDL6103B
yGg4Moz60AdNCKevQVya3c5L07wPxccycPCMbZfJri3XFdb19+p0TW/rwoLuzJkjyXZ192W5h5jv
XAQrcc33PTtswx6rgFwcnxrrTcKzzBMKgI4OmoScedlSd4Mn8tS+C/V/lGzoj3vnIiAs7c82wLYD
pj8rQ6OkT0W5mP44fqbNNg7qONPirED3baqTDl635kZ2durg0Vf34d1rBhM5kiqKE0n0k0DIqf8G
1OY2r5AvdxwOkli/9TXHuvY0W2hli0INHqQSCgaiG+gClLd4l8+ifsuwJfVVZbTU9+mHrlyesbSB
SC7Tnds8fBjEPfnt0W+0FZOG1vJNlyqN/k3dxnriJMhCMzXNoNgsK+NJA9iUlXRVzJK72W+D95+c
nO/Ymzx/o67gMUjZ9YEALuPHYnU0bAtLsRt7El/dOlmUG7aY/fZDDCtRoHWtWO8VtMZrdcRculje
LHfRkVHstcdm3cyE5hs/MaIaffIpf+xBvNXb/o//rNPK/ZWZs6rduMeuCyG7IMVdb0keC1+DVw2i
hrRss9L6Z8uEQ+yYXDvClN2RqSu989+RCD7PXR60ydF5zNAEK70EXq/PLwrBoUM2pB0FHVKeqWma
mxuI85aJ58f0pOu+jZ8ZmqfN8lWW5hEqUg0aT/9fwJSgcxKgrhLISlANsrj8u5oEVuT3MLE3OdTd
8cSojNB+F+HKajX9eZewQcy6LFzW5csHNB9XvuaSUZW3MDGuqdScP7wlMFToCkDMqy2jbH6f4cSy
vlXwZ/EKl41XAZ/t3m01zvpwBmHhNgDQuYsuaoOCKFsYEyv9G9tkUhT+39qbK4wAH7z79udhVSeM
a7nwqK7pjKHjUiuXYPI/ovhKTRmZDsHLfHfiTTkM0UAVvfBHw6ZtTFS/Oge/uTjl+Q/kqZ9XF24y
DodldhmKypB/N6ORy5mfSgNWBlMnp9sQI271uTV4mGAa0BbBJEDMpsW8FgJazqnCrlooYAf4oA6j
NCka/h7L3grzGJ4FfbMre/jEotp2OcdQ+Dm2wxqikP00UN2U5gfO7GFVfP43sr7pcMdj8y42Hpkl
E9zzA6JF0WY2KgYbMAIjS28YvlWIax+QbRNjKz1YDlBy/jbwV2hpcvd0dwgyjxwE406wJBeTtuX4
U58XBBs0o76DICzfu7sJpjrf0n4A0kiKNFhhWF/86BUI372cLg9nOsL+3OZTeQNvUeVq1R3bmGgs
PcgjYySTT5iIFXIVHE8kvgWpXJSGSk0ZEmx7VKs9KNwGfPXq3KUrutMOV3t6S0u6oTmMghuaHjFj
1e4Z3yirKVrQ6QiPasWTsIg31Xh3y04CC9tervZxWrdWDjwPrDe/E7goQ+wsDSmfctsff+mLJ1OM
rRUMXIzQRa3WOG0XNgF8tLOk18Xmkc9CsD37xMe5ez9C6RT5njOr8s8mY81rJeWB73CoUHL7wWr9
8zNSDw0wvNZyI5bICr7iRg4ueLEJxv+bpLXuSRO6bYrzkJrBG2Wx2C86+TMFXBpIbx4c2pKQEo/T
dZDM1EvU9Rm7fcgz9oEGNRijDQypP9jKn9IAI9UwLILE8O2iYROODT6FqaddMQRN9wJqF0YLWLoR
3xP49c4OJpgj4H1DLKNdZGWn9S7fSK0DdMZf+sVD1mK0wtdDo425PKcMjHOb5SDlc8eOJlaJSkNJ
UcOZ2Tx/dNdj0Uki1tBSSZYunDbEUcTZgQMCIVDIJKfegSBxmw+3Od4/od6U6DM0sspD1kyjIei0
bFbZJZQOJXQhkrLfaW1+JgFWNyxii7I49I+7noMooY6j9M5Ge9pj5I2rA+0rUvGiOmCjA20EpfaL
ShlYoisko86/sm82WDfeujGDyT9WM43rUy4N7iLI774EFbgxp2Wp+x5bqG5FKV0QcYnUSXJVS+9c
IrXxj6zJrr0OSJx+4MF2b8RkdSHQt6mS9tB/F7yVu612iFqwIQAIsckGlZYn5Ht4zo7eGAGK9Zn9
NTCS8hj/0g7zm5SuPXCh89MiD0u54AUOONz3pv34XkwkD4hzmUorOXBHJun6Bl1pEsvsr7MTgnwf
MtCAq7DkQDXckeg24cLR1s3hTyG8Uju6sirHvcVxrpVVsSLZDWazLHzZXBLXkiumWa3h0Gbv5jd9
VhV7SnQPuXnE7Zg2RMOSYYbPreev92sDxvqOtvw1awu0WmUCYWNqViawO7wNUEchMNheScFvf97J
PbtJsz+X35GwmrGkRalQIWXEXOYTKbHbMkzTv0ZwYxMUKrpgVNqlTkOOrvkAtN++AOvLE+gEpLEo
v8Kkg2WhqrZpt8xfODLCdQ30u6odZADcQ5uA9BGi/1oQkG8/sBs8cCvWw2UXsJ7QULNDtXbPsLLV
eKFUkbaS94snQdndTiVtP+FDnkjZ3C19dcc0PkR6swFS89YwKaazqZNxK3lfW9qlm/bv7DwUxv2B
ZDi0zk0QMn56fnxA5BN+orKDxsE9I3sqG2cv59I32mXkmzd3ooXurNBtIdeDEWl9Kqo76b59vNa8
3Wn3RMp3gwOhHoM2cfIeBevNZxw5ijko51J4D/FA/kIELNojSFPT9UCwkO0itMO1lQqglTAZcpsS
5GamYH4uFPuDHK+gZPwSTGMLoDGpqP0crrsv9PhKdIXlXTGjRchlMsm+142XBeG2KdEzGMIC3n4l
zBeQwrg9azs7/fg34646nBQxiJ3Oq2O7FYD16w9gP3GauMQlSS7uQ9mne7Q4MAPunDtF21kg6+84
dIUrfRTQFZsk0olnN0vCbVl/gjERdQga89sivfrupEr31aUcCNI9G2AYb/HNohzqTvjbKK438oH4
60HcoCk1VNU8H62e4dRkuEmfNI6TOPooyFP97H7KkeryRYM7s8WdbbH6OH2l4hZPSzfI+9SSLRvz
obiP5hJYcsNUlzeAKhA9fH+QpqEQvYulelk+UrAo74bCYg5ZYo0aux9HbKJXJ/uhHmdqHmTt6b66
wQtB5OdlMwpKDOaALX71BErQjmms4N9NwVpGqFGRi5pEu6oNUt/rUr7Irat11maVQm7J4W6ZSqN5
CpKUcgsdVDJ+WccbPjNh3TmW6x99EKDnFNUa13yzoqvgwsiLJtIlBVqi9ZXK72KWJ8OuGOyJrVdr
Z2hrJvW9FJM/BxjBxaSX7f9VqqhcMRMybrgCor7msLc3v11JGGegaN0T9kOM7g09xU5T0nPOds72
Gu9qJTiJjgicUk/Inl8nIdLdUKaKsopBEi4Tt6zao1aNdl5HLP0saAnEGwtoGdk0NKuSopLBvipn
gGivhTvZ6M6Ts4uZY9xUJHgme8eCyIzgJKIE4MSlgfwsCM+1DJEgUaYUJvBeNp3Vxdua8bwTaLRZ
OWXXK7esT2xSGhVoH9+TPlvSUN2llVp/96hvj5nqcSOZLNxHuV1eXqywFAP4KLB5lZ9JcKWMylF1
OjuLpWX9X0cA4RbiFONGK68EsbVu99E9hzv41Jug9AOimpQ7BU9rgCsj6C2lNBBRzsB9iBpzwOGx
D8RA+X9UoKFSanTZpBED6+E4C5whC8dySBth6GWDxAVF3OPDMTULu6Vdl3FJ/U/2Kiuqeyjhq96M
IjAQltM+RiNSXS7vnXX7I1wjqtBvztDhPC0ixAi/+TChtV6usXTCllpfDQ3TaqFZQqc/mmWp+Fvv
d+/jo4K1Nc93anXo+IbeiADkk0xoY392fikR5anhSn1s+HVovYYq//aFMDeYHhdcpKFc9aJGybV4
TjlA7e2mNzXS7JMchDGLmFU6olEMyJOdAFr/bqSrJOlRK1PEBnplBvClh/STDRuGQjTaxvZLLXYu
MVW57DPyDBMYOGKX5I1B35PsLbK3/qBZ2yE5Py4bdK12EahA02pxaW6z01nmmtF5UAhSVWcL8vek
WHWmXkdDah03P42RUTCye/5kDqXA7fYLBiGslfoqoTq3WFKy/VuBz+dpiNgxeRdBoHmqd4SIdCOA
RBnFajEoOHC9Hj31K8BU8n4XxPNeeRJ+0hwNSNqy3noyLqYrVC4apy1fW4a26yy7bN09JH+Vymyz
bq+2rhTA+qkVKTEwTz4+CotRPzCbgYbQZhVGl2IVeyYOFaZzzUkykh6bofKB34PAaWARCph1m03I
za942k8VEpVWTleEnusFAySu3KhC9mnAagpqysfnYCBm39o2STh/9fbM1vvvfWvS8IlskhA3cH/U
lj+pEmo22Q9yclDCPcU2C3n9Aa1khWxc0+5K9BguI5eT3bZP0I59r/LSSN0mgIIdqRxSFm1UBioY
GemawMFJ25ahJHuDmg1SGfVveNqe/ZW3e8x6w0KvZvI9OEt3v/b00GUX0/PL8cYsrlNP58y2Vgyq
IAOm85IPiqyN34BFcxyuWXn9A6ZRYnUG6i3vTdGMEK9DaiBoz5PTva5CVTnNNH0n5dMXZ5j6Zixp
pcw8n0Z2JnVG+fNp6uiYtJP/vGGxs+KlK5CSa8JqkAn8o5gDbkZbu+sQDrrTTMIrnILG1ySI76Ra
Qo+HSN5d6j9eTBx4JrMNCad9yLJJpxm65e0ErxQgm0I4VXFiB8wmGXNBg/sknFKMP425QpYiNKff
bKWGCF3VZjTtvttQUvX0Em3/M7XlORWsraUjR29trdPpYJbsb+TTHj2Uq6Vf09EbrUHFe9i4qyvI
dhExl5MLtlkKDk3lnvF3AdbL562Knb5EGerD01yxnXp0AXn+Q2FLhPSEFZClQG9NQLcsbHrSVAwa
o0+axtU1oXfuZfs8j2rSSPfy1gTTkuQ4+fKpt9c4+bb9D9Ku0cr+2FlWeuJQdCCwXNDcnMBFqi47
jitAZgLfFbt7ZWEIiYFEFKho/bx/jqkBXHIIlsb7K/gtihgZUo5ksSvTiBAzgQ6cM+/kYsv3RjwU
8BkNQ9ZJq3WbsWSyQGZpKZEkfdA6niJ8G1rMla3GPKV0/whlgmZy0XfFMYGjnAmscNafbnheXiwW
5l6iiYmgZ0LnuZIuwxu4/7NKmNiZOeaBWEwrZ++nDaYhkcF/jz9GEjDIeVL4eX8lp2pbJT4cprfa
1oBprEIEXcl/cuXg4drcLJ0c4ZHfWwf8VJ3q7GM08JVGE25qBuzhJ05vmy1gQQORhHCBwEtNtqkZ
mAbO0OSyHgAJjBMQYdnbbzvRJuvfQs5kwhPJTUj3fmZcTbPvDKEouh9NWdh/2e7MzgYGnbr4dWAX
o6E931K70B3VB9X5H7i48xSm5pwtS3hUM3W6vAmqNBOOt/ZNCzqA04m5FltJne1CDpN0SQT49O32
ySDD1MOr2O/zI103ueyWejsqTOQ6WCDYOdM9nnPj72JXVVB2NvakWNlg74dMVboYqgQ3eUOQ9LA2
HDa7DtMY064/GfvundEy4ZsnpgjXHOpkuGhHH3XpGul5M8okbC/mzBISfJxCrr/J8aGUBmS+ZtVX
p9YR6lOEiXESHPRJrwT+3qaQIaTP/AJaY8GLWfGk/mgPt4u48PXR+IKKaCC6t/gpUm15r+jPec1E
sq5esC8XK7aY9OgXdIitOnrx/isZVmU0kY7QclJx6JurmH4tkTE/WkP5yJCY2anrdpmZb3DGqASD
7mg8TG7D51p0AzycfGpzbbK8SR5gvDJH08A3jUqJEPd0clYLt5T7fuC1jJojKKcaOEFD1kiCbYI5
vmsgkBjB1RTUnXyHn0VIXSsf7/NGegJ5Kn4Mol5gVT1u0TbXZQKEz4/e9tncQPPD/Kkt/p0MNDEU
NrQQzKGZjyawtsHPnq3E2kZRK6bMlJig6hBBabnMrT6iu2w5NWC8nlrL9tbpt7EadW+42jGLFZiq
sl2fTkFN/hpOZrdRVUTxImqROcOS8hKARbuGlu+50ou50pYvJtspxlV7YgMCaEkTfaxuy0lCFwTn
UsGQ490PKYrlTb9F9J+RCxcBge3xKnTiMscXbf5jkFeSIttUVGzTMaS3pE4GHP4NKQJfIIsG0Es7
T6RBb+XkxCPRhOYkAcOy/YOsMoEaMu6tqiFCq10BzbwzsSkFv2po0Hjc2Qm1Ppqa67BWBbtBh6t6
LMJKQ/L5En5QDwWcowA6MkfzX97qzeEKiqWlruPFPsVCkR789Ti1Uw6MLLvMo7zcm3+OX+EDi8bY
hflRoXtrDrLCnhNHSlkqSVWn+afclDqkLbWnprbnPL6teRyATXM5Dbs3uByRCN30k5eRiL9Kct+Y
6Byx0vM4kZu7fVBc70s1T6dVv/qfSj0RYAWAmQHzSQoqasdo+SSloLYSDH5DHYnIwbxG4bU8zLYo
Y5XALgpamDECyyBYmGqNAaggL5OhAymCCEdvF0uG0mIoXovRNqj1HJGcS6Q3XiShZvO60qznoeXG
V+px3Mco75V8ZUds0WUwIVKsuxy1WKTkxHnzBnPAcO3A/9LIa4hAW2kWunhbM/sgJClz84Uvwh9H
mYXkXIJyvAHT/fkgf6SEvs26xTdIfarWlWm5E8j4jiBh3MCHnC1+B9vXDaz2DbO00j1YVu5p++Pp
Z4/85zxWa3BK5ZN7tfCMsppR8GQfR8PwKxoQiDAUY7g0kOf2/crgy51MGHcu/+JyAdo8kLlljgW6
aajHzk6FyHO+uP7snwQb3LWQc0DQUpByiX2EWSs2KJ6WV+X0ldoW0/3+BvNlhrHLqtpg2FF1QMbg
sTyhnQ7qzKYrIn2PxuHts8dp2oktslQMavGKacA5TntEsZPrZlJ1KqfP4CN+03GpmjLj/gMIyBab
bUl5B7bkdp0nLMHrtcqy4dogXzxYbJHrPjIFi75PFBcYiIp4Jxq0H2lROxOcneJ4CNrAZ1TacGWO
7ulg8myuaYapmjJzte7WVyioX198PzuqoRd3qeNSC+PlNeNH+4IeP4UDc7R1nFnlmc2ZJAT2lR1S
h8vCjXPtW7MMiZPCDVPmhVp6C23iUYBnk17NsQSPolwFhTDacy0hSDsHSgWy+E/ZgApztYNfG82S
APkewQq7mnSa3n/xj94DOAk6Y8Ef3j628pYwfc48HgUJKa27lpgjl/QJvYXtm7OZ55gIJCEY+NUb
To6QVTZ9bZNjpIGL36GMPvEdgYbf7SVnf2cmVW7CHgvCV+/K5KkdOxK9NxsxZPrEd4pwUAAMzA12
r6n4iql12xLJlYkvzD4ApLrBHqCkwmvhPpA1ydkZZ8YzfTijWV1nAUtHlhIQlHyaG81cUzhGEWtD
wQOM3IwvGMX4sNs4SXACYsj5iz8M1v2DnEIoJp2C9cRPIRN9JrXNgL8L28mj8qnKl8IIKly8QWW7
EzXvLfS2RLkDlDI9cZ2aMDgr+qtCFsgAlMxgU2lDnbktCp3H0NCAZp98ppfRvQRm+w4pBmukJuBc
Jt5mXge0Y1Oa8i/TF9zBhwtBVhgwGfqx5TGwYIFFoHP6wBvi2k74LSFU2/6LHplxrbaaZHS5FF/l
TppCrGZigcmbTxVbAO5Nhq9Ghur0wZzEcfuqOuao8YrhoFxMmmWRjqD3OozZnX14pI2X4rSvD4m3
KXy8L9zKluivNt03hJYaKxqOo3tDAX+HiLcRnWPdVikzzziLvZlkAnivzjOwNmr3KssYnBmrJYLO
6uViQDDunNPSxBXAE87S1zwoOqu5zeTCFVmaP2Mw3U3I0zXYqFXxKmFREZTlgr/bAqSSlja0iT+j
ytWA3xiRkhWsI17Mq9h90nUjKDHk+OWD7VZcmlUxi3NUUXFRLfWRpvoeTZi9VcTAxWnz4iIHrqz4
SKgXFB/XzU/HVUumuFRfTnSjJBf6ZNkVjEj04IpK/kwt6rUzozQUb41dO3coHF+cl240mvOicXzw
zhlfKxFs+gXLDSXZmw1M4UkjYXBelB6Z8cJKAkuBzkVdbNUfBGax3AlXIqljFfGDnXsZJ+slb+jZ
5GV8ibdyF7GKAcggCJmVI/9ifpMM31qfwKCwM2J8yQZ5qZ/Ihy1AZhlS2xBABSuSy8ElSCNRBXu2
op5Ie0YcmwrZkFBlq6pntigKjSgzCesgGXQ4cnsqCLTD2gRQc14WxO/7lRYPUvTl8jEu+s1H3wNy
Nc2Fj8ZRJXe5nZ1TKCGliJesPLLXou8quH58eEfoGSTb5KCKc+FTJRjAA70JbNbx9XqtypAKgqBN
A0x3KVLamBXqnLpljxSqgAOQuiYJgVhom2NdXXL5R4eDSNUIwuaV1B5RF7JMgv4ADWLmOpUGu2k/
DAs7w24++P2nWucowserDLSf/Tg036AOccwkdGVucs1CTiJmetg2Om3g1w5grgfaAk7W7Hb8JvJY
7ITf0/Igf/ihU4uIM9tqO5V9cnL88nHNRJCIiju19aWalbEY7OZ/jU2MC0L2Jilo7gSJmy1YdZDt
ACtMOlAy6nIX8qDR15vVdYkzlj0l3iM2REj1EeGUsRg53QOfV1chxCBDbhSrTs3KDC8OfqIbZGv9
Jz5J5RjJIy7i86T9TyuAdrU+zDUV19f7M9a4YK0TCEQB3kHSiesyd0If2vSUZ7krtZtu29bv/zzG
QxSDlzKy7epf3ou9jXVJCKHCyJSy+9naRPEsKIpiLqZh53wPF7g6qAtp8hi5M7VcN4tldK1io4Qx
wdp5Kl1VH8QFFATsKNKwsCtJLC921KMK79Odaf6MKTyf/O5rMKUBws7HOtovceA+sXKCtc8bLiSx
tfi8455sB4fh20oKOx2wQMBkIZTi4NG+LPBoAFx2bexDjMj5cHKOpwqahbjXYzOsF45KVf40+XVL
7BWDrk+TAZIDB5moUUi5nDSK7hhjQVlT7BV6QLaxSH7wCfLFrHXyk9IAaLQgpvJ7sU1749qqK5Pe
OROZ1SnNmb8gBBqEwUgFgRK5kGxz4oWs1MGLA/7U5eXTzYHSngbWhKAy9mM0RtX+8pIFEEqTnYGM
XEFh85D/ioCUcRBKenPUhXZ+ixYpAZHLO7iD2qx4n6M0KFnRIMAtmcSIln7AoIXUvaghKG4Tp+UM
IUQrI09/WekHkGn24uhlcgsryyed9ZXWPAo1GdLZCQ23cLddq9IsP03dKHw76/ZEZ1X2aPyYDBI+
RebviKuD78cNSDxVX3EaBuMn8JVupRPCdsak2JjQYT2t4wm0HtsROhX9I7KEyjH/e2K89c+aMoj2
ZgyaC4ITvGIsenhi9lqRnwt4edwJ+T4Mg/j8neMv8R0srdPYq0uMCVvnQI0hU0jSftDTQ+T01ksM
UlHAuP5OjpQm5zye5AA2P1bI1AJDcNcO1YgPKcwHUGKKQQJo6xXiJVNNkGoq2t5D1JyTNfpT4ZFD
GD8Amc9rmAZwgDCZ6dg/KSviCB3YUY5mwsZcOTB1+/nLig0MFYHLHJll8RuCGD5rRZZNLmEHhtV3
Utkb1465aNzqVplGad3P7PD8n8aTCDWe2OAakAJ3BBkHPioAQ5OMmvNOfbrrAyBhWgIx9LnWRBVE
VRWrG0qRzVZkDoFzAGeWYvuSil+rmg5B2QT105IEOp37PYqCXndklKTCGfO0Py4Q2SIw+QT+Edxj
kHfreq3dagEP9vyEDkWWN7zL7or6hBQfIVgJ3U+85WGx+6kO5cFsNcnEWcB6Kv3lkk4CeRaOMSHE
KnZcsPcIIqVirmics/tJoo/lCtU7YS7v+FSlgFBDdj7wCoYfPnEJl368jDdU5hoM/oXUxKpBkL1H
uVdPgUzNSpo8auGvztUCS3b6BFOkoJJquVJejK2q+t/SXj0you87/pi3vcvrQIWpAyGWFP+uiaet
Xa9ozWxSst4hYE7ZKypbHhlEVnIlr/fxTgT3uX1H9Q6pzSYpRN73NVxloe/uxBJav9MWqMfRa5uC
SM12xrM/xevthDXMieBiSkYwU7bE0dPZzocyVsOSDcCGe6CIWbMKgpXGRF1GfkjMQsY/x1stq5QB
KISfdFw5l3JrtcX9wRERApETmWHrRYEF16j4nmF/cxPU8sdl+nNAsHPtqKPjSlki7UgCwSdqe0/M
DGS7bKwY/OlHchdsNIIUmgYQ4MMjC46uIY/wvTvsfjUuz+W09hUydaLKwZksTu7d7kGomQL8p4jm
P4fQjeiK+KPhAOqpzVac1oXZQ6r4tPZJ7b4VYliQuqiBdwAgMQUeXZkwup/w3fjwlSgwJVu+7AEg
Gch8G68DuKJu4EWy8m0sXsKmaOxlo7GjWlgoR1IvfFnespjeSgLFN40oLyHzE8x0cuypr4r32X8I
ocL6k3g0lAtwmvQu/9FcYpX0ATMsL8M3tWAle4JYKZ+FlwL7pPJnmkqgmNCC1T8hhWnk0nDT1XCB
t7b38o75AZnsXN6RwjFGfngRvIR46UaIrXHcA+7a2uIxIjPt8kKRMHxgMbPaJ4cEeWv7J7kr2x/x
Wt20KvCBMnGeadvONjxLUvdVanfOxwwuOQLsVetwCWp7oFpU7+VB1t/gkvd/EJg53UU2klW2piWE
Lsgc2iSKE0Pr0e5zu+OX/CViVl1KIdVMb0NTCBsKPdPa+RJ33Yz3NyouhaWuUCY8muj+8IotvnvH
nl3RgdCKRc/SnARePAKwcm0eGmm75qJ8dr6DlhVAlXbYHvm4tbbzhWFQa0eFY3BzeDYXSU6R9L6W
lyo8OjKgN3Bg6SpqBalK1WGVblSBAQald1c1UN0VwUpb9WYj0EYggva4tyiW2RpES1dD5g7uIO9O
KqiAE/G21Qomh/meq44LMo6H4DiIZaISt5hGLof4/0xJYla1/6hE8oSSdRbW6U8dCuQo4hgfZfqo
LYxkEsKSpO+1cUSzG9DtZBpyjIYuXBytcleJ60wyJ/zBga2QrZ+a9MSRMgA7/XjiELfe/6YZtJP1
RO8bM8YJdBfACbEuo8sTcJNqhxJ49Loay0KE4Wei16mfxa4j/WxiALPvT2Ai3fKr5IgbFJSuAR1t
J63ULTxi9FD/ZHKZ/MK8PQijCPh4Ntvi6hZ15KbOka3MVuElRE8otfx+uV0D6iuCIATYR6OgE0VU
7z/K30oq5cgO33SygHkf0Z9Re9vllZ93HNrFgpImxHpbNNOriZLqEjgT8xLYUBsKD2k4XJXDxpqX
ppxqkVXz6GzIhYJo39kdUfZ4EgHpcl5GgscBzc0FTlrPPfmTu0J9STsVu5hjSFy96yATrhe+gIJu
GvhDuTP///F0phZciY1UZD4plR5/R8uyPec6tDGY71G6Xi4MhLWhiDjIV/iDsJISoBjCj1ndcreA
DPwcAftkbNvTYCjblQmBRKoM8A+7mXIXasguZH+K/1AbCD2IMH9RL7CAsIWU6zYIQRrngLItCtlP
L/MIRoq6kkwZK9FuXBVLO+abAQR0wi+/5zJX1O0AaFijM/kaeHbAzDQuu6DcuPGpeRD5v53KlefI
VeEUidUIFt6ZJEzI6YyoYv3idA+sa4Rw8ijl8b5PrdcoCu7PnTvWdeQy+fgxvjI8DxUWpRL/zNiZ
zTdwB6SDMqll1ReD7hohdruRjshSZ/Fpb+gy4peMTI347lsnYfdqxTcCKbio2qwDcxccBMGYwZcO
2WMm/XqRkywjCTOHWsNmiUC36rgknu39e8+H0WK/Wbgt4EOg8EUS9nLNPhHLhN6BbTGNy538sQcj
e5ZcaebKPCqfY5QcgajDU1aJUZ1pJja6bAcRgOj8MPqN2yFkBCkxS0P9vY/o1CT4d4Fo18vFEc2r
NFsxZD7uWao13GEbonqL6d3z1m9CYQWonCxpP0Wk1Ehb69JhlXQiQXUGIAn466g7WIT37j+bEBoI
vObSSKfe688NI5GHInDRppo0YYwWB7vVfnvzARx5UEx/22YrtnqZ2mQvF9M/nOBofrlEtlws1aNN
7FWb2+m3MGFI0XM0pMReWi+kiH9iEZ8mbA9VoyKULi9J7RGmMBl8x2kdPobBXg3w9poznyjx6RUb
4WWcauHxOZNKOcprbXSORRjRr9xBB4nKxRxxJ5vbVOBv6d21V527P/4HwzEgdkyoDkGbD6H0DtI7
D4j49rhsXeeOBpbBnRe4OyjKTsjZfu3/eqhMXqP/BbnSU/8h/GCwzFpppPCFN+NrrHLOGP0X63j2
2jNQHBtJ5atHqwhLNMP9oMVD5awLl9NhQFSAGrdH0qOEujvWQybXBWIjjJY3/EUZ84LT4FiNymVk
6e5KgVTwzZaCElFi0o3cGWh0PePfeLVwSPPDIDI6QyT88md1Z9Uyj72+NlvFSFiDwc0NNUSeYAcJ
mUDcwodLtqq4SxCi9LeOJIKuS8jjBUTwamHCH0WJ8kxtqQBN/2Wjz61RhWu4RDkeM25rvKHDiqsc
EXJpzmwvdmxB5hdXWFj8dvcaiPbrGZM0U0rkkUSGRqbWVlTcStUvgPlM7fkt4mLVwmiB1aZ/8fXp
hZ2La9997wctZ1b1Se5I+rri+UotJ2a5USPJMQZCr6MSJLsyNMR6uwfTVD1VBWW+hFfZP6f7UWUU
E+Jv70ngpz8prmRXkBW3sCN2biEehYqbP+UWxCagIWDt3qZILSflfVMaR2u/JwP/RcTxm6hEUE2B
jgWngl5O/+0d4N2zeUyc3gN7u7b9/2F3WeRkHQeksl56KWeDFUnVWsSl70rN2AznGSrdnehgD439
o1EDOkBqxXB/+HejqxGtspJqcQyKSWH2ep6b77V1Tx8NajVCpj5UzoQZ4e2Toa7Q0+Z5gNhpxKon
RjPAdwDYLTEk+XqI6MRxdWJ0IUci/vTk4OhVsc2+t/v+z0Z7sg2XB85EbXTPRRZuIRDl7HmBqTma
9O+5FWfJISWWTJ/NUgQ+tciys/Slk4IG0aOEgXa01ueljrXcfZOlixJE1f6zkvZJqvJFBfvjArKO
rS/VdO3F/J+c9BFh/iwSoLcCCvze4AutfoU6XpRLEIVRfoCZKSq2cS78a8c3vqZMf6cVHHcAnYTf
cPKyakZt0JAZ6rMs7eOn/9phNS/koET+Sjwa/vzoNmg9OXlHk1zCUegVwKUl9EuhJds7mYyZkv1B
Os38i9YeKOVcBn3+xvp/3yxztE+RFhaGfr3llbkCbwuLpHyszts7x5uyDyPU6SrjFA+0EYStlIki
tbso+2OQUpTYaGGyhr227lqc7u3wfTKEgGcHgS8r5EhqpEBFnvE/G4V+5ICYZfBAxKUGUrJANZpw
V8yD6KpuuWJLXP1ibD3Ans7FAkvir13le595KOMQZoylp9rngj71oVk/L6eikkNcUpw0lXt8Y/w8
iNxeF6A3BnRO9poyxc7xOFBmm4ozMFdQM20o8zATfPWAcCK6j+yyYpjakmSef6mqsn7VR8tjIyoL
SOB5Hpt2tJq8Qq6LZYPcMGU/7y6rfSxijXo4SMrSXhonyHScZGEhWu+ik9S7/lGIc6MlkB77Kant
6N5thmuN500YpuU949Te7RYMJnba/QFuyotoqkZQZ2p6Yym6SdBzAR24BXACQA4WUNC6I7M2CweF
wBt0fZBj/3B2FbdZh+LzW6+9g/Jhcyu8zwoS1h0HTITLsJ47ov9OBCd8LS7cPwKEUe2atlhA8Qqf
4/C6e5gja0eT+Pq8nRG6rRXFJO6vPlfztQo87WFMKgwYXMaZoatukjVyLlbtvJiZoRetWuS3X8BI
1p89HfXARIs/0xBu7lJ6gqBbrXwL2oj8rIpUu87oU4dCKYLkEuicfA77VKTQtmCqDn04CHCVzbyu
CsxDxde7CtapiL20sNRVKEaQ9OMxh3L9v4thlPlQ1k+lx6pKuGrCBuwWPAZLe6Pdx2mF7Z2yyYL8
K64ku6xFuwhe9X4v8celv3jAspUBSaaavBfbW9EFfh60ziSeno3DdLoamrfxyb3pD1fxk5I29ZwT
Z3T7c5j0HuSdwZytiMt9VsLcFzERGCifI4CSEFKGXxOBTm87ouwhpPlIrczc7Xpk0nfU8HEsHWbs
g8Ozs011SOyeHLc58217zYE2WJjxOW4VGKuGqBkQpsMarhplX1SymCjfrYGH1U2fI5+uXnKZQAgd
t24VI0Un0Wm/vN+AfRQQ/aTnrXDcPezUG8ymIJkDjjo9LWMnZM/n67Nc4N1Y+HRAJL7NF5Q8XPHi
EKAIJZc+2TCxc/pf0wvs/GrCppOEbt3nvoM5iYwbY269d4628wBtvsumkPZcDXwanwSac3jZeOKE
sjmat9BVSElRnJCxUH2qqFrwCtma31xL5CKrD/tLKJOwVaoZhbOm72wM2jOR8XFloMM56BesJpOa
fPE+DjY65Iph8YQoawTCtY4+xbPg396dUK8nwSBlIvhL2C+Ny2tbZfhYY9Y+PHZ+9gJNkSJOCs5X
bofnyl0ZQ0NZTaOrtdhujgxbVwpJ3cqf0xWtmiSVOL20dKP/hjc5PAfjqMCh0UP8UcWkhZc2USBO
9RovKXxv1PwQ9U1SpHS126VHxkg7jKJ4EiioxVs8vkYfAMZA1VUzcKuiy+cjmCMA7CWgMLqt6XVZ
5B3wsuSZo1lxRZPOw10OZ/98A3wy/UgyR+tDWMqIzyBziLudLN3tujf6n2CkBKC1rVY9JMhTlgkU
ZmW44iFqCP+//1bjLDWZuWGb1QAb+dLdPe+NWdR2PEFKVG9BxbPj46QjpwyO0Zn7/lKWFVV2/K9B
0uzcfygZ14IPY00Y56PMdKzMKs2+0wosuZE34kvgVh/woVJjHXaLBWMShQ9/1exFWqqia8RHHJ+W
fuIlrdvrYd/zH9U3qSjfucgr299Rex1IjLsh8Awiq52sSTmoD/mg6yn7ieYteMdxJYKZ9JINiYdu
VXKr/S188w0NwMt5hctRzgWHmpFFKnMQbe0k/2Tf8OLy0bQNWzX5PHYkEnie6D3Un97gHuYuhdYr
e33xzGkU1++4p12kREQquIhf0q+pbdZWAbjau3ZtICfdCUuYlytDE98MPMCM9MEv02Z85yPz5Chs
X/oM993w9qasxMiKY7uhlJVhodq2RqIQUpDMPkeFBvEy0nMiweixgSo+7GqpUOgsRGMmku4NxEE7
3I3XI3wAh5kKWu3YUhLnAxWyYJjcndw8MBbH1suQcn0L2PZBPrp/LFuuqKWYlROQJjbinTjA5V30
LNjN4gy7uvO0X8fNcpCXElOjXu4fEmvlnwNJLitnI6uNChE0YBLKfPEepgJ4WwDogO1vcmcIx1Au
ko4iCt9mn8cghJx/5vdYDMyal+vToRoEuWoVoK6zy/9yC4uag3pOmd8hIIbhAuDH/1ZscjcIyhlt
CzwPEQiC2gC6bTqQxxtoc5JRGvEJmtJPvCeCE2N4PHC20wqGI2Nm3MqdZ8zR48bX/T/l2ixC42B+
15M5anL1frqYigRgcf+E49XCESCUidMWyKa7yXmLJelBoMMXqyMrlPDS/BwJtLmB2xySUkkkpshB
rFTiaiR2ZXyHSMd7O0AmK4CXTUuFjmdGyqW1F8uu0sT3IqX9haU2HDFkiWs/0zGx2lxCKZs3LRKX
E0oF4lI+74p/G1hhfQTBDh7kwgERm+BixL9CLJ9CLeZFUXkahfjGl8mv77aOhk460mF9KYSmZ7ly
L6Oawe57valhC4zoNe7L+kP5DoTTG5y3nw52mdhqf0aNjjnBk2w+iyXEmuRXskMoIPEcDCDIlOfj
IBM09IM+gNIFohVtVX50xNUn65ZbpWRwQxBZN4ozpicp/kB78RpQa9E4TO1fSej7mevqHCNc07Ec
zlZOQpSg54LMVgP7I3bkp6WG/8rwOG1b/ypdTtfVjTyWEobdHB3l5Ep77GylWfUHLE8ugczGwoY0
mbDBc/yWiR/iOOnLVqjdze3tQrXoPAB+sZqQL4f1oM056ai5EIcBG3GEjodGz6f9CQUlZOQxh7DP
XJQU4zkxkM0jwHe/VyhzZS13rIEseN1EiNn6jf+scO0zlLz+IJY1r7NXj8jk42OxvAglJpB7gRzr
0jsJKmIBJ8IcifVTPrM3Q2ClOvS4/pmADOwqf2mcEFnA8v2kooXz5kZK1b8GSB43sYfg85RFI2Xs
LZmKu94Vec//ojqB+4ErxuMchDez2ldxFt+BDOabcE8nfvn3If25D58qMy3QGFI6Rmv5wQ8aT7fu
CRh9xQ/EGb+Ru+1rk75Iwuzy6lUxdQi4Ucip9YePhSCalyCKBzmBdGilgnJyBAGaab7TfFFooI9s
HYrSLYoxrl+7ZhsJ9rPftz3N/Y9arUeYuhqCFftcr9u8v0rRpsEvpFU9XPcne6QH4sSN0GkR3i+r
rOMp8end9gPch00Yk9sy3XcKyNIcce0MUbubpN+YlzI1A/DLdHgdKwqRm2A4Mq/QQu4slEHmy67k
TgAo2AB0sMD/XHPWm3KSRtCR1v5EDy/AVgBKcSv/hCY5eYycvERxcbBP7ds+kCuw5YQYX57Bc4bw
lswDwZScleEG/BnEmMoZcgAwEtlrIb7NdtvMWDhmUXrSrHU/JYK2sTTW5PYVruHJzSaq9rK/NyL/
Uuse6NQhk0xUbwxVIXXM8gLozsvkS7JO0VKdLM9p0z79FQR6urCB1REkmga3zc5hjNeGZdoJoHcO
vlRf1iHbIXY58ngkq+twoNMsiQ1omYaERD+68jH2HDZ4fKAOcvux3EU7OQiy0QQ2srp7QHJ8bzTn
Y+8p8o0Mvm7z6ab8h3kDk62IVfxzG2CAHjiJVZ7AlcCoWfCa9LLcFT/1CTd0MezTODMUgjQ0KrRw
5vQPJWAXyDxKJTSlE6sTMXa9DaBpdfMPKfVjkg0XG8iClciOets0siX1R6n2nmOkGx/7GWRTNmx3
gqOgHN7C0p8B0VohX7ktr5QLKSBP+4vWnz8uniKcFyVPi8bO2xMS4try615iPs5Vtq1RZcKoDEK2
TyvUX7+vmZDfbdm1xXNrLgmuhVENiyiAXQG5tRLSZLahXs8NKvhgeBea9vPBKcpJZU5msPlYymut
fnqLangex2j5FDpbjtlJqS1iI2CCqCIFx1Cx21tJqqSbJM7aKXHO8egRdrhyOI5SZLCCwF3cyl86
QTawglzoTEeD0A0xYBqgcFOjLqkWOpftOmOEou0AZI4ofMHScFV4eTYGKJi/MtKLqd46fPywVatx
JcVjFHlHhMBadH5OuyebeE68sUwqPuDNv/pwJdHmDWEB9rK/JGZNyDnY6wqM8cDItbl7C571DIOD
3jpGfalXetl8BwvxHZLItKE4H4XLdDOoAw3fwR6/MXROrywj/Bbfda5c5j8e3cRCYeAHhN7wtz44
KKWGC6YIwp1XlRxtP6PAwbVnK6n7Kh4koOa7T2nbHJgOwkguNv/3NFIBzfeAOSmyN/Csh6LxcmXI
WEKR40vApeRc7yCVIKc9nMuFWtcxe/Hzc8A1Ikx0wdbNEOfa44TGV2+KmGFaxraYC/8tPw/JJH9+
q6LQMGDfyfYPJLsu404i0pJJVvVSmbVx1beIXJ+2bPMx1wDUT3TcMrnNLBrE9g0KimDkKk9izEcR
AURFCiSHXIJKNQGicZsU3LuZt4hEKDnKn/vTRjX/juluTXSFFBGqD5SGDMc86VJ1OPdbKSzVe7Yc
IXQnQ6KjLRmDxBeVIrfqZxyR+hd8nIBKeUxXYHRcpKTVu5dR17f5HKWveA/8cxNokmjayOpZ5F5P
vSRG/yVbxmnfKMhUvUl4q4NnMId8Rd/SUEKTkOLmdZTGwJd+KTFLnmaay6fetxwHYqh2ZTYDMrVC
Ilv968WxnhvQ3INaFLI1SJBD3PH/j2JSmQMd0gikjKL2+MoMIcQ2E9gXsLD+KvYdK+EucEqKMKG8
CYI9KrKD46/qIS1Bmi+lYZVXoUbaG+FUF5ulRUVJC874dM5FJ5f2s4UO0G3FturT69z8E38TXSay
rtTv6AeSM226ImkCgdpjc0eA4adW0yT5E5GPGRGsGM4Yean5LZ3C0LkqqrxGqo9H0x85hBPCwu3U
v1AbcouXmdpBSu9NdFbvHA4I/wj4401W7uK2Jtxs9W71vOV8eXNCTUzkalEQsebpyc9tSN5QsbmU
tKQX90UT3Do+YAu3UuEsr49jC6jITZlIoxyuznJcQqkmkeF/umGp9Ugn/8zjOIsPMw71vFRK/hK5
erBM+sCHq18d/lB4jv8qwrEXnvIFOkAtZX0Ah34o8/AE8N49m4P3i7N4+f/mOiLrQn5SYrHzPd7c
/IaBBiTzrTbVz+/kxS+0EMY1lmy8V0EZdDmDEZwsH8/s+AE9N3aXYaAtiBROzAPJhFm4A/nEZxQT
4fu8QHS4keNItYOLhlxr44D0whcrOOH+CJboOC5kN708+kKxRRjqdFswVRy713QBZDyt2rhLPtgH
rr4E1PzJtyLTmkfb/yg5pn7Eu+PckZcEFfkwYKhGT54NZSeN/njTEHnafDizIfeAN+STsjpuPIoB
Sw98RtCRORtlo17y6QbSGVzr95BiEedjN0K3xXGPERj+WlmyESdh9HMwPEiJ0DfdrcxcdhtLbwIh
KqpRGqYdrfr9Sbvp0aHhnRZmqF7Q6GzAHrzYS5alsh1FiVwyyaRRbxg2O1Wc1YYrmwNH/5XC12Dv
0NklcJ1qrTZ2I8uTv2FkAYN9q7jHiMj8h7ADAFFIeoJv+5z7FwZXCt7CYvWHnTVSVs2nl/aF0fc6
Tttxx5gHLiIZc1S75prOdej4QP53Ar1LXhsYwuj2zGu4Q8uYqY0WRwFcMhGUEwCYdB53kzcRx03w
+aqgNrgnWcVz8Knfm7pl64asCbT5TtChk5aBkD9IreAezOn1pBHfs9qEoapwGs6twkwKoWdrLaLp
kn/AlpYQ1f7xIwl7Qq7wK1iV1pYWlVgPjXyl0czYFuVcmRQTqTHrQTyA2KslHvCUBI6/GjIEGeLu
p1641DJerVhWohBtX5QZJaU1b4Uhztart8QWSxjXnPlBCq/U97g5EITc9NubMMf+hM/a4k2g3pwB
uNBda13vONKbOZ/SfYHf3C2gEqsDtjnCC5JDnm67lnqcPwBBuG/Pwi/K8ZP6BzwerOGOOJM9uGy8
bK3rB9AOSsFiNWThYpo6YaZrbdm1ry08y2djQk4gs3HYZvfAGTRIBzsYVO5599ZXdWu0cgJyUebo
USEWttJ0KkhQHNMnW8Wk4zwtN0V3UdfAMUwjyHDArKDewK+HdKl2EPbbnDpBlhmU6T+LkE2/7VbQ
hL18DFVHmoR3yE8fWuyVUK2mKdIAdtD8d8QmVTdHOKfnzwyDTtB4fDQGhYxJ2ydiaUfaL9Ti0YMq
Zk3hO2z1bxSLM7d2swo1wyEZyix8DHAenImrxhKHwR/XjkQmGEASk3Jk7NwCvDNktrgXA9ge1SwT
c2UvTtA2VaXY/sJvGAmGqv6+2VPk0Uax8FeNlDljM4iItktYBEGoAoMgkDxa8bZJCKVZrgYDbYg1
/hvhfJngHJTENy4cUZfRd3NVzFHkXDZ7QFhyBOjuXr47ZGWAlFf4LXxizvuQSGRnE9e88d7XfN/L
9xFsYleGrHX/Qwb/UlZy5GvVg50bOg1+lA77t60hr5gPCh1EA5vRCnY7qSAJPZ6GxolD7Y+6XgC6
NtfMii+1/JctNQXTbOOcZUapZphAfJXvXNtmLn/aDk7S1Sd276996I9O2w9Rvb6D3ZJRACrs5czG
BkTyv2rglCcaEaga24nlL+2fNywJK6NWJhseL9zaaqgcA/DmNHeylbnBzIanfFfVm4aFH3p5Kre4
svd2XLbwZTOwWNS33rucsPm4dLTeyZAbRCmESwUCgSDYo9MxsqvvjIm9YoDBmJ42AmYWISx6OJo7
l/4jzx1Aai65VBBEEO1MtDz4CkDVEoflM72/W7GPEEj7p1DnnjQkVKuWmK5nvsE0zNeEYpuy1iZD
2iQ4QalNyXIInhKKxznEIrXGFynpdpIJSbl74k766oVGG0M1RvdhMJoxJN/FU+WM3YE6EIwWvAyS
IJkW9kx9x+Lp2ZNpREmH5gmKhaj/6bPhp5INtaKGmbqdsqM2pLDTlRPgi25DY1ugcE07ejjTPHlK
yBHPqFzlzGi66PPBJGMjUqVHC71Uuue1Kl3x3rosWMWFbQeWezUQn68T1+p5Eucy7D5aNgt9UQuo
HjE+AQEpdFyfW3qfpyUYhIYE4JIMWeJjRUupd9Ceb/6HM8nvLoug6bQYJan3unx6/xUApjntleIX
TG42SdG/HDub1Ce0QFsilBh2GMjpUgamMiq6/yzykCjpzOAywbv0mtZRhcGnp5eYs2cpyovlpXSD
Rtt2B4p8wjBiEZ0+o2wtQyd0SCOVdFUCnOqBKEKwD018HyU7a8EcMT48Hq5Qa78MdFEKZfltmRVA
5UdZJxf296nviOXrudYF3574d3gvlsr4kdI+Oojh1wMwnuWpj72TBjhspZ5G3X/YusgpvlG4OZRC
wfzieksW8gySS2CK2vxHee4b0ZLpg33qmTxXrbaYuhMfcgCDcGxcbubzJmicmA/OnDihyRk6XSwe
m5+u4WvhKoyKZ3ykkD3aFG3hzIMk0r5NVs95TTRYFipUfbGYU17j10d0LU6hjsXTB721q5sceM4W
pCGq3jz1aoljPRnNJIYIx35cOUibO2l29hLtsxgVmYa/XEC/GkqngmFNzkphsiJ8Zd2x1ZV6ETTA
RR8h3rPx2dPPsAuFedKPxx+8GZDckzAZuXjp5nA/XYIsXjPfIK4KMIGH/LojPfDhy5veTHs9KZaw
C3uDHB4oFiVZShgBBCfa3+5dG0g8QlkxlETeWlqPmUbo0OkNQNakMQhktvn7CN422sBYdvFyx6sp
Q+pw0qkiM246J9eRVzk0AuFlcZz2LmthYJoy5P9BrnX/0t//IzMFfXtsv4hGChLKGlm/yFaVP4MY
+vExcbljLwa04EhbBe5hUS2QMI6wTrcPT12+5MnbcvG1vjVRTC8+eSQ8L2/19JJS4vlP1YCrjTyM
Vupr/purlHrxgq8kMYrWWwL3Vr73JbtE8a9kA7Du1vpsdY7AOM7/0UcOqFukdlAfxjdy5ItBvInb
CkU/ZGF1TLXarV0PQws+itLlySdxW7oBpdFOI+jTNlqmuuELBKB+AF+8z73JSpYX0tKRhUxh5+y7
9V88fA/qrqM5pLGB4bHDNK3ryjwx84ct+zWwZSMLeE5MdbFY6dte7PpnPT+y9Ya8csJVqGNS0E9l
hq5qlKzZEiZVLzMyv5xPSIdGhQol6lD2WsuH5eT3ywd2/yAhBRqFDNAbSppT+/m2dYfi/xp8kD61
8OPqJ8uqP9Y131UsE0NhSrn9HAVroTOE8DVQd31TyH4igk+teVEIRwkmiBsDzxKoZw6tl2pQLti5
KBrf+9npehC1/EDKbnMTrx1y3uKyJ1/ddkzBwIuWE62h/v+gb5qEoQ4pQw91e4fPLDM40yynlnp2
6ulnzEKdJ3PPIJxuqHsGJzom2lOFzErdbapP/QayiDWfXrtWlPOs5OvL01SKyit2IuTHXzCzbzL6
kkFWAfjyIKdHuflYRLtzrmY+wU5Kbcx7uTKvWotgachqXQhUEENwXDeUR+gmhSRPHZ6v6hOf9sEw
NWTmOk2WE1bXOThMkipKzzGWtUDvhQxHEXT7UyF1sxhSt3tj9JIaXf2VcUqyQhuiJ03ED2nljrRD
Dea6Z6HHiybTHZllU0RkJUwH1QT4p/V4A7jHST2cxLZaH2yS5JSM+4QE2BZH/ub64ywEOBoI9Xiw
Aqqdw8snzTKNj7PJR3jnZ3rpBaCg50FKH3OnQymCoNZxSVjzM1VwvT+WFYE3NimQfNxSTmaAj7lS
+/u2kbnKrss3FX/hbHAxddFuh3Klek0Dx6/tl9e4+7JUXoxAa0YkzlfRTGzdAQiwQY3MPz6k74cM
f0QPwvN+RWpONHjxXVdT4O8AxAZFa7V265wDckFaVR/Y4jbppEoN2/8hVHANxTkYhFUnFBtzs8M+
fBK3PBkFDmAqYeqhRGaqDMDpP0jCpr4j/oeWimac4nlLRgB2auoVBGhY8G6nQ+UrL7pPk+4YRkln
oDiDdZxfyXJL149GJaPiaSDBRNyM2d5pR2/j6gqZ5e1p/i9AR4ktYtcABhzO9LfBSbf9xssjLhjF
ZGWZWGyw2JItNNbtIiGLAu16u9sHWbxRFQ3GvCyubMNpJUn3xaQ016aa5yiCJO51oKfLcUQR/dC4
O3LePW9Lg2Sg32n4HRTv+oee6rt9FzEdhErM/2zB0UPXlwqMIfKwwt62tUWIqjGRtIFV25SaDiEj
kPEuZwpPGHjn/5451EOGSQuRAcRkSNj/i78XbhGyPLGMd2fIDoaqPmyfaUWDJGFABL9pNLzWFNF5
6OS9lmAFNl0YSPLoESIZ0xUdbZoYaANQGBGhxzhn8P+r9giOWf7Ljb7nfXjaQHH1pWjdaW5Aj1S4
hN99HrlGAf47BkmHrgVyoGhB0QLVtSrt9nRpF/T1htxUlIt8GwfaLwdiSTAUqWnrKz2WP1k/svWW
bHRMcYSJXbZuXjaU0c5mX10SI1Oh5hb2wKn7ht9n5sWej9Fa5efZlSLBoSN3+js5HJ80fbvqO/fG
XgwyWtRvqKOEF98s34LxiXtyFvlASyXlCiP3K3fge+Lr3NlLHG2psvbPa2vXEi+4F5/ko3Qiqyqe
m90XNhsd2X2Z6D/ICxsHF67OvtA3vcQ0taM9fdkKf3s+CUMYyHa4rn7dKJU1KQ8ffY056G4LLlI7
Zrsso3BO6aETloThPjs+sJIV4b7ec19xuyxzBzypu+EKRH6uYh02mKPtpPOOdIp6qTaZyv41mCBN
mXhpSGBUgUKNa8j1tII5vY0gL4Zz3kX7FB3JAUafEwrDAmR+IPfEttdfrULRDrfBnjqG4DoYe1Pv
Cs81pt1vOLrgk7iXuY7Hu5GOpKUqHn7Yk0ULZzGLHogk4oWWEZ1oOyeD3SNf72eQq9yl0+jklgLX
12+lQNWyrcNyoMg9z5nM9PDSrYmfDE0dT8PJxN/TZxmr91r+MtZ0IvRbIqvIkJmy4ec7YrGwv67A
dUstlfgsJCCHASEzeP4VdJKWwhpO2V0FU3qdBdoETYfoLwDxfdlsI3yPbfvYTLWKQ6QNUTEq6hAE
WzLS/23ebcEqxeB0/wDWv/zbA0q/qc5TtvPoIJ5j/++Ag5oQTb4S27r2uq3qGu09YfIDz3Fh0Do5
NeOr94TtbzGl60zhrUXeWf8uVacAS3h4OrjSlU9QllEZt31CLZF2OezwUWEdkfSb003LNvVIIsXM
HKFzQurE769HiryB9wY4ig9FiF2jMuGPWEaAsONvEKA+xjJbdG8EffUYWYMb93cO3xYq5KGO7Equ
Rw64b+BEDcx0bYRWTeKPnCKpSPRmYUHd1rmjbS7frkns7NnJO2YuNtjfEY650I7S92KyGhFNbI/i
v+/QokNOHUOmGpp4P5NDS/z2X7R49Ho2H/HWibfsGVnPbNLtKarCTah6OZG4/l5ViI/gcAXUkGow
gvfNyTMZGaWYAeUy2I1waaD4+pFTWjYB3Hh8GGFHetSP2WcA2N8THtkZmyw2quit140I2xRX3z+s
9p8XPX3JRYiHx0Dy44G3HwV/UNtYva4hrZcy1mnPbA6JPAc/Ceze2ynGw4u5due/uujFSuVZMRgw
IxFsrukfr2g4zib1My7zD4B7Hxdsx5CXv/FfV5kVHw5wf5MwYXjaphXqNlkbpzuboUCUrYlUbxub
qtXgv8ikIxXjdHG3gB5KCBk9mxvPEY4AAcGN33UnNce3O6dqdVnSkuSDt57UxQeAaTl1KGxpZMsG
BC+H2SfXzIOFeK4r7Yvwy66w39VviC3h2E243jK5Qy+ROcPQ3HdSroXasZ6P2R1tupme8baIpGyD
W1YalVU9r9rqX+ii6pFBJeuwL5TxjW80THBd1NrDv+giplQ9220Fevih88Io9/7tIjUVy+0v7Jch
MBPc911QKvOaSIL4+39g6aZw6FNwrYJLgyxMlnU1ZWkU5gK2emapvT++Z2H8p9dBnUuKmrT3sRcI
c8E94XqDacnf89iVptCri4pQrmzU4MFsZ4J8/Us95SQtXP/7rj2cIegy8StNt424u6UJZkwINnp7
JIUJon0i3gnzUHYSohIKsJAZkUgEWppBxkE4Sad+zrEKQO+PNqfqNqfMh/gdNv8jFQ4xkWcNjn+8
NikIQI+ljxG4fo9dSdkFdqMkTN0PH3SUsZVPkBccdMaLiVVHBDaXH6dcxnI9jpD4ZJq19AcRjSpO
85d8E1zhG9lIgbr682+XrUTofYJnDPPGKWYFYGmZ1Dl9zW5tZu5GM1YXlwdUOT3HupHNYvTS9CRr
abuE87IYWnJiZKknhP3Y76F12Iw5axhs91KPmI0vv60ST4klNRhtS9EOzh+PC+b4DOHrTbY0kTnq
Axajyws2epFWspxJUdj1slykYRRZsA8fvyexdyX8q3HZL+AKtPLEYLvmMAY/r6W3p5RaMImttfCl
zUwnDTosUImy0gFrhXS4JW1JPUjMIpnYKaum7b/9Dx8LMoNHNXHdeCcrSlTUAj5zCrTgc3wAP8SY
sB/9GD1Drj/7xohozr3WYUae3HZydW/mSmdlwsmcTrQlSx/XnIGn+V/n1dpGUzwDRN3OFpQc7c+v
7PXQJG+i6gsnmwJZ6A1y/mmXwvNeein72qWHgAbsQU67jxi7cN1d3CS6wvU9yTKZEXEoLzEL0JxQ
h1CQjJKEyyYS5s90iyV/MiWMR6y0jJeH7Z3fBILs3NI75xLJnV9Xi7ve5QWNTwhaRuJvQ4aWJhji
U/ybkmPl9CR7NtnbS7k8x8wg+rFk/XsXr50YaLP1Lsis4HDDv9moJOB+8ToixWXi0YPXWBf6+2ft
5yKS7EPQ9cWzPUqTpibyr5KWk1nCSpOnwT3eJyq/Q37LQZgqFNa0qOlHn/pgwZOLwfFbUXxj6Bag
EMdnDWMZ3aphhPrViecsnHBQf2nA4+SQB05sv/e0cne94Kj99gBHHiVaZzFLPFpoc8XxvQQQb9U8
WP1BqH7spHOmc3r+wx+idcW4Govg6x96garXvKAX9eoeA8ZhtaYvjoMxi8Rr+l2wshEJBra5IDH9
+qvnGsTHngi0FZLfzSHL+YHHdIhdLql8iYvqcwgwBNggUlOdc9CNzFZbg7dENnArdgyKbwx8K4Or
y57PEov2WBMwHVhh10l/sJMawRCERWvVqYucisJw9PBV/CTvLQZY+ST32z8ktJj7DPIWi8TGaN0t
TKVawEf7w1qgGz8nuDhYjfLhT/IzImU8NzG+mCT0CNuYpEIqjiHPmNNXeq1cSAi3FONQdjQBEaNx
BALwRDZP3si6g5ymHLuOpMXiS+KDMzd4uJH8bxRcqKXHtzQip5NkBV0NOkvNCAZSUvq9cHc/7Zps
TwzDydgW2jGhVJAqgCVzYVxdNrDqAcQHzAeTxGObcOyOfmgeIU9xN95Nn2uhqqhJF4rxUa6SWULq
jVmZkhsBoF2Hyc1a3gG903TbQnejJ7A20NRvGYNIoSqRNH2s/wrWsdFN6Zm/5Dj3oFyVYTQYGsNd
ji0X/euJdCnHEIjrML3Uv2OqV5yhbL+6J8AtF4e1FlZeGKdzoFzL2Gerrly+rW1ubO11M5bUpfWt
6ZjdNaP83o/J+pwvNxJcpK78i0GZmsCM5BMiO/L8Cx6uuqczq1ff0xXdvS05cMlwVF2qyJayMjsr
OQ/RgARt/qDB94BXelxL4b8+IfZXogdEmxzYXG6+10sasW0RrzRHB2qwos44kAXB29zSzu5srVWm
qU60LEKCTr+mTVevlfoOMZeeayp74c2tCzVXelPjAjPIXk5UNgOTdjN9/iB4BF94kNFXh2HlV5Ld
xh37mxmt/oGIkYDhptPpYbg/bC8e6BFA8dZWxFUJyIdn0wNt0u9xZp/tY6EzLt9ORlKlNEvQGeeY
F/G+zfKLOhbKBCc8UWLbUgs99xSYaB41qe0gMn/4+Nxhsss6Ao2AHr0a5bcf2xO6JmQGLN/HsxyA
u5PRb/oEfEECV6ERVFKE3cL2sx956Kj7kCECOXxxQqDLIUfMVSiRh6NudYN65W5jo3/tpc7QqJq3
4co+0MhdYUOO/NwCCdNnBz1DtulyX6SZhyeRQVbcxb/dZv+0u4JO2Mwi6wdN1ZF8Y6nO5XeNXQPZ
+P8WKOieOPBh/D1AZa0pQq99qJm8Jr80dGi20t+r5OdXDrB89D04hzhe7fGfcTfx4ojZb0aiz9rh
8CVA2kRXnpblj9+9ceAHAJxRfAK7FLUTpqtzrf5evf4kIKGQC/zWvNSXnBdVG2CJg5rrBEhIzrmy
12y+SawIQ4y5NbJv/wLg/HO55D97G2y8AzenT0YQaQlkr1EDcxp/kULxVcs3MwRnQixqXSVDm9eu
mDepKaQwoRxnvaDKaIuIJj0dah4rHVpCoJj8AT7bGUB8mt2TUZceXifxwveQoN5XWHmGBqz5tah0
HhlzhcrQXc8y7yqI4qTFbg0GT9lanB9WavhsqhAeSojBgzBw824Z0kEmE74MRQaXF8/0b+FoGX5D
27WsHT6VhrGlgkZF82hnjOYN5kfocDfgW4UVnztexw5osToYWLq2eC5zu1b+ekZBTWcKWm5MF1EP
utzbM+3WQ8RW6tVKs0nJDM8mGteOkEa7EWo+FuYoubMLjlP4mWPBrXcgRap6pCgxbClagLBkeoA/
Pel1dLj8qNAQygjaQjG4ZDgfohm0Hp78NFbWUkS7auYeUzZ9oevhxPptKjcHP8LjEHbfrRoSW0vL
2VAIP5MGGWN8zyS23adMaqnoyJn99YswkwHkMjNitZWUioepPyY77cv4chGwYPTuJWV3qewNq/qR
AWs7iDH+Qj2AW+QtooorhkU15iRtmdf1Rpu8hQOXmYq/Wh1lyYEI47guB0uZKGp+kCroZ38RyOUM
tryJe28ElcH7h0V/d97IcmLqupHNx3cb4lnBCiY+PtiVUdAgFBxQJfo3LRK4SqLWHAt7FHkiNRzj
ypvG5s5LeaKiCaYfdkNurW6jYq3qRH5fOztdh087s533H29LkHg1vjhoj4WvDtM/Ua3iWyyGsdYP
RGGAHmhZB3VNENzBwT3rnEuiBmiL8Z3t1ILfPJ9amp5zaG+zOatSeKX+CQlvwavheDXzYupbiVEg
lkaYf3m231UuFaVnhzwvJrW6WBko5a2D0JSnEtbm4e3GTXXjRsbCiYF6dqx8QYTAr173FPsGCaWI
RcVfTmpvS2juFqyd7Ms+ie0ye3UC9D6zSjjW2lCzCnBb9USiY+GvZBU47m+Fu7vRFnOfMfGgQWZe
JZwgf+HqbuOUSYI6VYytOX7mLampbko1ChbEiwyoWINc77cUrTUXgHvBsNVl3IxuzGXclg4CdpJG
eHDkqFDDkYaKLEO2xjAPqTgbWgEQIiC8GsFJyMYDFAzDdN6QXw4lRm/NAfu+6sl1849Qp16tUx9z
PsWkkRhY0/jLiTEwqD9VZb9DY9kQVzIWrNL/+1R5u3LddwX78ZRrcpTv4dmnONyQP7yggpQZsVIw
RKA/s+TUCEdzY6PIW0d+MwV7Est8fnCnET0OwUo1y0rvsIL9eUeQyLWMy7Lzcw/PD/HtKjLwTRUM
leVvcFbQERQvPLgh1W1DO44qz3fkVfuxkTSX4R5H7L3S67CVi3aRzR+hAj9eJdHTfu34Vk2tYR68
prpNht5RC1YQCAZNi21nz1h0KyrPVvS5M9VvRxdos8QfUa/glRBE0kR3W4FmtdWzvCgRyHQKvUZ4
mPJ+05H2G2B2dyKxdCz2CCZ3trar7SwJmzFiIntOIbNks3UIdabP0/TWlqsv2b6iGtaapn9WKCul
WsT+0NZYMTO6+2J9ACM7pcmy36NFS9t5lfsKw6isqvdrrpbGVQ9C2/Z+nB3vDu6DQs2EOnILz6Jt
4NfsctCdhvgulYKXsv80iUB6DeJd7BSsyaEMidQ19Dz3ext5nXYKqwx9k3jufIHuhjbGFaV4YGdw
HsweKJoa1cshha0a9VGwobBN0+7AaT+PRUeq0nYskXJjVkYdBxjJx9yHbPyvR9lPVNuAEof6cyEX
ay6ZFY4Sl3wHpDvoat12CVZo4p5Zp9IEzaZhlzDg6GUq+jlftz6zF8EFUdnAlJh61h0ropLigBZ0
EImULWXie4xcPS4f7fX7X7qSn3zNad0qq+GSFvdI2Lit12ROdlhaZDAMQCiBf/Uk0RrcfJQGCRfr
/GVv4CZCgNJw3Uc7nEiKSM7Z+VCEKVsi5YS1+ZPw8zjFfmV1GyiFrlF0Gzq2MzM7xiV+pvCcHjPV
dUoUU2PDP+NwKhJBYkiSw/iILHdHTGtRlQ/YnudhwonWhqbDBE+nPc1JIhYLPKl7F4OV2XSZALdX
Tgwz6ixxzFKPcqB09n7FWJKJBo3Vu5xLdF+BbqX1G/x6HAhtnIz4SJGeMNfh+J/Djx/T9zUlNd41
kdCc+IJxKohcvSkq/wcRUpDOQQl0xW0NFams8XjIV1tT+Tp7zGFSFDMMtXC1xk7Y1hyDznZc3bYP
RwuZEF4CKhOKiOGW/0JzJ3vR2A8jSkiOTfoDAo/8KKEb0Lfp5f6kCat6wmuaSoXxGXFTd6DjXOYg
nRgy4R4OCpf5nHpAQipMLoec4fW86XBHq2lpT67p39FpaLFB3uhyYgv+5TFeOy7uJ2OMfg8wwi3n
o4yoJyigtqa8n/oVSDayWLMWGSx0gsCj0bF9nKYVZbmOgbvuPhjxdGDwelX7S+q05P+d3XuRpALS
dgAbF/NSo91f11HXeOLHAHYMhF5B8G/ohn67+e5pu4Kk3Qk+Ox3kej7ZcMcX4ntCw/1LcGafr0rG
JVKY5SWj4W+voiDoLihahn6cBEu1BoJUV90NMCO91oTDTCHD64CRqq/GoScqP8b3D2rj7/NDoQ9U
rUaQU3taGpduzPaQ69QktCBmYvpH99PKC0Fa611osQnMjTSifosg7b8lzhkORKCkPrdeBPQ5g0f9
SBwC9reZopOxstRNBEQrGjfEZHqNmTFRNdDK6wUfdnM0kO2YoQIcm2q4ZTuJLfr7qG5XKmzDNtfw
JY5Jib4zqgZm8TQ1A5oltw26yZ37xpnEqEbnmHtKSCVwq6n4wcR38sYCs4d8s6EDiLA50HZnvge4
/2Fn//7b6fdbsR3a1tb3/GLOOtvGMnb92cSQXCSe9vIem7Z4SKflj1i9JY8pxV02zioO8vOJEe4Q
X8l9peFJ6fKhlUY2gvTPPc2Dy+K2ctGDC/23ga5MZM5mCAIJlngY96s9ev9dbKUrA5TOEzNQS31j
kil/Jv3A/mjLSTjddQJ+1zfSs1ffVhpOMAKCMe6D0IZAhPpK7HxHh2mELOQNbyb+0dTfwArRtRbK
F+2Z5DdW6wUZF5lGQYKiG25NrWuhomxIibOs1BuHTdWR6lZTwTsedHZLQCOkz4fxrZL7c5cdevnH
LCLLKkWbALj/eukxnRGfCbrtA05ZxHu/gWub7E2yMgg4lXnFJrGCFs/ZFNlrBAqqkvLM9UD8Cs8G
JTiRu4c4GZSSHWIzz8v0xEhDeuO0PP4NXjHlDCsGN6s0gYJy5gM2t3Hr1T++SwNVX6k9tT6Uv9kv
lHfd+3b9OZmlHpFfMyOfQMDDuPMvwzMiASkd1iK5K3QEp0brfJ7ROb2lwvEF2ciA8kHgkCGkKpzz
nsI5EhI/ok+pr0gKz3OQmgKG0THtvazCNnNsSUbdzmTVLpsfCc6s1KYWzWdgroj6CdL038/56gW1
KfUDZNVB8GzpTNP3XnWLu3fZ58q7VADLu+DvSG6YLhBxI9Pby/f60yCxFC+OOKF5UGlU2yEtVReH
0UNQLXK00opC0FAE75VSJb0VhQ0I2rgF6Lk+d+vTAm0nHoqmwqxNjL5iv9zNDgUqxl6EACMvFC7/
PpRg5+KA3MoZgfSFIwTpB92SLNvM7nlVx4NDMVgaISwIQUJqoCOA4hBUiJvW8XiRD419aNTjd3v3
lnbC2OiPsP2CRzEqvGa8ANiTOzgORehdXIXaqJFr/cXsBLqt1jrfkOpkMwNIHdUcHNQcXVd1BkbD
22uegjUG6bToSYc4aCxnNYyeab0Jigz7njnSMgyrfALdOlRFnt/xHQWsplLfgSAY3WzUwvG+AXIq
johc0mc1tlf4obvXkaiiZW33dSee/8+tBw7VkSFDBQZCYk02BhtxEdgib4IVBjRPGO4XzoCksbfn
CAq996CClw7u0hyL0HaSbSUznK6rs9ZqW1rIRhiVSml2GKyyq8GMjYp+KeLSGvZ+0M+IW1yiUbVy
TLHG+hOoieSTc0PjIfxCASeyN45X3HcxwMd3usBy2yJxnEIJ+pZ/6sJw9wLKmM7CexeGVC2ctp7H
SKL//YG2l5X4XZrK7tOib9+PdcLkacSt86W5CoCsn7ck7Hi6FEp/a6eHQ62cQOKCBK2tU3RzjTlc
TZ8M/xVcWn8U3OdD9C3oRXj0qkKo/m/AQwrL9OSgku+kmBo6OT6fPHAotTq0wRgdLzIK30gdvf42
7XVvg6GDgi5voIA1sPDR4rW/CxzP+a9c3m36IiuS1dFvobCcoxK39xBDMHTgLAwzE7QsrmEw64KR
LjEE5Bt2QdHgvw3B4l96ahP+WMRsb5YC5+FtIJegv0AkNnai6PkZ3qRf4lubI3iEgKSdPDY58FFC
04dvydEkFnSLTuMN5w4cDm6BIzgIS407XuhaG+BbZStCqJTNcKAm7JE4hfOgKG/eYG5v5skcZApJ
OEoSNELiGSEkkw3FJ/ZStNSrgYqlDoqV7gnEYWUJKNl9FU5EUJqIyOWurNjW6DgnezBXUUwSwHx1
RfUxnTelsLb9flEth13GmVpg1PHvit+Hte1/mzwfVUyAAEs6WFPwNFzVu372tCS7UA4Wc0bClq1M
eCm0PVF2LJXE6miBCiCwXb1URVpqwLT8WvSRVjJteF8b0GFwZeK7Ck/xeas+mqFw2Y4swpUbhsuB
+fOzKr6caMXgVEPl+d9BQK+yH1sjv3Lpt5bAdBQvIEjNpSRTsBoxRRddTGT00CanQCuIfju/6Txx
ZCEp6QJiBb7bpZVa9AXhtundEvivifQa3icxZ99bEHooIVDC6C3SmUErWUaoOKV8RL43Azq0eSAn
YFibuBSqKkhYh1z4YFqvow4nHsCxsbsLy1IFlhm48Qb4UBuDVWITgfxcWwfD99ozN6yki+CkjyKq
GD8/LqprfOaUSUZhoj4ldA3lgS51Elfz2um/r67uAMZ+WSEziQ5DmQ3+uakX+JdkvrarVKMIGNjl
jvrJZdRmACc6UCKFfA81cTIzCjv9jI1MKkqnzUzUOIHjYxn9n7R3L5TBYoDPqoSJCsZ8dowannXN
W1GzmpbjNbXyihdE/1stwFRrLFTGSqJk0eWl6D5xWzDqg5HeLIzeD9mKl4C5u7kFbd2inBojI8CP
mWUKU565QWRrca3opqrdJlT7L00p1g1JoQmJEYzTrbkTZu3uLIT3TR+3MCabpLk7IOaMax6y6ZNe
VI6PSMJ2EJkI/Bo5whkNpdj4+0eg46PWSoOwvLYqovImHuZ5YRWZ4xb9uAREKUmjJOqhQYg95BNO
LlnA+Qb7q9Dhq5I6DFKcFpq9PsSbSLpwfKhoFFcyYm0pFqmUtYgyhA+XZOluH5icqmfBWoDt0daT
BJJwBGEpQQfpek2e8BshjQfzSrlMBE0Mv3PlXwmG3uzKrgGD886zV25eqfuqzOZhUUPPD5aV+qgd
LmnJcYCnaz0RyzFy5j+rahgoDVrVt24n6WSpKbjTUjwZpj2m7Ol7RQgCwTHMh/y1mhftZFzKwbyy
j9+OCfBA0KCQYT7pEIPB/83aMO2G1rGXF5jYutCBD4bODmx92kddOi5jFvEoZsEoIZbXbJYcBDTW
ThtqCfr4XIy7xjao8B1MYba4gBFI4C7xsBclaf0KgUORcBaSZ0HQGPhjkB8CjpOkmrIgLtxv91PY
BLtSkbWuH1nLYqrNqSIBCVdSMx6WL1lOnIyy5HuNg1dfWG4eNUtbtRJnKkxligS8VZkcK26etj/Z
nDl71iRTU4Ry8eSvf9tQ/sl8TcxXzUXC13TQvO5QzMv8i9vo3ddsVlbdTMQdEqhgMRyKx1T/9wal
6xC7caGj/BCosnlW3VMTN4LzPX1XROj+vxiBSFjHp7Z6K54JKQosQosEQRdyIWmN9ZBHWam9pvqw
mmHP8VwTMpkkV0hc8T3O8C9qVRVrbA0tun26MBScoCwY7rQz7qRbLA0IoiLP7IIsp6IquEowDjiR
ubcXujI8zi5HDvTZwNzTMlMYedbet37uJuUgr4PwWV315nCvCLkqoDNpcJYkx4TtDwjLVgX85Nex
dZPK/QwQBfgI9eyaMvewMHh0X1RWBYLRtOWPfkPg+GHTom0X1EJeglVOqMGmhmmow9HjCJ62mKP6
G6JuoXWmnqa4TGXJLbRjP++ST394RYnJR5prSnPY3hhlAMPC861jF9pprJQdk28hs6ZnuYUpqdb3
XpXK9XiNgY4VZa+qPo83HdSVkyUKf7l4G3Lzx2NKbmCDvrfqyuinOpflVuFHvoaEJFTu7kcQasR1
ky5K1Kx3DTUK7PUtTO7BgwqQRpFEnPBMPw8APFWdiyRmxwGUE6ohna4vo7HzSnEc40FpltfpZ1fm
mB13CosNBlOJXPnWbwW+muF6tCvmByYwijz1+kIX5HlYbFWz6tf3+srbH2XvfEXcbMYytU3ePa65
EMGvgQPPvE/0J158/ghawO1YrGGzMfHB3qY9uihTOsegIqY9jadM4RUv0XRJvatvh5Jf4F+2YCzJ
I8sbxOQhgK4qHG55zgEh1DumqCoAeavhTwcq7H4CoZt8lb51md6knSLLnvqE1qIxIEGsdhwI4Apu
BLcUl5+U+jHci10/+8r4xfk0LCfkfNm3sCHpBb2MBByFvmsuvvTqXUt4iILacFgwF5EbQ2a3nyHH
3GPeMJzVoRps3pIbIiXyOp6JTL2yQCm8F37NhGqbrn6hKQB+vJ3fLqiHyXDVDNikJkWHuW57vQvm
H0iPxetz5wvVTji9hfj8cBF+hn7XxwELDss1qqM6v7nZCoaacwCW1395McCJmaB32WtI0pELYltc
zrXYmQ53CyB9KC2HiSToAG2TZliqm4dDnum0ulPVtSDiYwp/cm9i3qs1w14ufDO52qY8GrZvjgm8
ZKOFeHxGHpkw/HgVLu0gaDrZFwL1v6ooiGVT0hQ7pwnhnyAchYMeykGV46AOEYTVcpQ6KmKfE82k
ERX53PWrPDCko2J+TneUPh/m8BCDexIhc9gcQPG07KmjQJTQ0FcA9huLPYqR0jXwCXEJjS5NlWZ5
0wGPutNYlDgL7wPdK4OoCECOhDaXm61CDu7rF50LEv14zV6S9kJVm2SNuCnIWnmghx6SEnTUJU3a
kD52ggajAOco6s8+XdYNOEAJ/u6Xz1PwvEmb/OQry/R/fr/eJyWVlVOn0BPGzkIG7/QMMZTDGSr9
nicIz7hHV/AfSpKPcIvcueOSuHSIQp3DAggScnYdEOYNIy4HwwUfwV+5vg9yUgwzk1Ti4ILX86UC
gp2Rb0QlSEAsCVk6k8mzX94lh50FpmawRFFFCOkwbUh+fgsuzOiNjHqYAXV08bhO6QWf0ELdoEBK
QEnl3/x1tG43IKCSJBExeLnfg49d2wM7H/P0xogHWtfgKTKRtVJZRKCplZhoh8OUI64e5LwgjYp7
YjQ/XyiLs7ZmgOBPcrQxv7hD8G3XlRnT4vCTt6xD5rS8G1oNeXq7kuem2uA5Qqj1yfDg6GTJp/lw
Xl4xx5iJZ2KYxB1/pNKSlt6Ud7VadWKCeg0fgKycUpzc9nCRk/hPfE+Sr0sj5mH2+V4j4BwmGPTV
02Q4Lor8SNWedA7EoFvAvWxE/MbSUdgjREPyw7NnZ3U0j+2PWYOC6wKDWAGlz/qGNnBe2DL6Wofs
2F1PNnry0c5k3lodgOIAs/ztiCJFgFuiRt+fEFn+m87jbB239PmEr/cPrQ+D24SUJPNEzRSVMZoT
8dRWjnUtKK/Ardc2VLT3GjvTUlGPId3A1DlVlt8BcnKl5v0uDFS1DgCz6ReX6XEMhe20Wd1JvqYM
JkdUW7POvbwfL8UkvnHBrVa4xi5xXDofrCXGs/tClJADFwx0tywk/tZdSmimStxaVFDTdE1fflAL
XzJSofCLU0+f23glCCzCckILXwpP4U/sRAR/hbw+4kfx5hxJ9o6QezO+MJcIMQT/ivlNFCjLKOju
TiF9wGim/Utjx2DOMQ08J8J+r8SCQ7lyht6mKx0/wEZi/wXbAZzBlh6SLFrKj4pETHWP1W9e4UJn
w1dm0ZqI2lB8vMtEzjSOg6Af2RV6ODnm49+Vm9CAlqNB/5gv57XylAV43BqOnEkCgJNEKUvKMInZ
abopPjWhQExw0so1itWjT5vY/q5wkkxTdLoeWjAdhcqVgPT9ycw//OsQ0dzSpTe3oafRMwlVwT1J
XD9NUiUtrpqTO6XkbFR0ESp1GLjV9lo+EE8TjYPrLsA/Rh6dh+wMDpXptbKLAAEQnd+mKWFWmJmB
lKwVTbTCaMWsmcpWOG5a1DYIZHVIExqmd/LRPUbS2TOx/f7oMzDTr+3Exs+qr+wZH+IzUZ3Ph2hx
CEm3nhSN2ewTlyqE4X0R1NHeRnz69ROT5p5vbxmEdFwGLLm3vjX6J19WKn6nAXK2zs9mYldkKVam
ZZqSW02Bm9PI1urlXvo6kMml4fh9CZwTlOEz/wsEGgABOxqfWupmgSv0rhnKKIL/I2lbE9bd1bEk
aBNWFqnmcCUEkIHMRM8iocwdq2CM0KTLJ54GWmwCVg626IUoWc/Go29GcHy0Eyi04MdDvzkXpx/2
inVxtMiVo40FzyrI5mK72/ieq5q+tMiQdhvEjmFW0ltfWKlbfN2QFSooTfTklgDKrX2yMDy7tqye
Hfgm0oD7HhDnjZISOefgSVasH6fsxaCFv9cKQM3Su8DusNfOIXm3Kf4jIK52AcnTCS9gfFJKMpsS
kc26S6wm4a3e34mLZ/ubk7WSQcyrz2aGHLuMQUJaNDEqyoSZF9bTSLw+FlC8oqkk+BvHc5qx5hVY
tyqI7xYa3VoNPXaZ4CwTArROrRqioo2Yo84grpPWYVZahzhjfROwDywTwrC2qt5lOtPZ/vbXLAY5
QbFOMzVrLJLu+Rr7ydm4HWaVK4DErLrrdAos8g2FwSrml+Viht25z0/pk7lijgHBGkkjWxvNCGkp
wX+09dj/ajz+YZ9f0muvnJzddPV1xilgNj7Rx2mHsiLAV0Skeba1qtcUH2iKfgXC1qW3uDB/lUtI
splSu+tzfXS2ZZUKqfx4Q8kcTvNEILgRbPBstQDPA/KBBOJFTkNPjvoauDJbuUBkm79AC2wdmA5c
32yMHCO78A8Jv/WyXjfdjAJfJ/lIccCsaIJq2b7AVnf40+GaZ4fJ/jpl+UpqwJwJi0JhT3L1rVH+
qf/zA5Lnpxrgois1J6gB/aj+wTg5AWh+lpMfptjhzZrx1yVQCIKiLmjPSNiEpzsmZord5mZZPUCR
tVhTZoAMBaVTlXTKYPNjKHDK3TNhTVu8XETDxNx4rBPDXorwkHtleTS12vxuGffDUlGj9KMpPuXw
0sG+qJmeMLNIbWY+End+Of/YAf5uGHTj/t0McBlA+s1iGDUrS57Uxid6RQUsYTp7p+WuHY5eOL5l
YlNSEf4NgTiAiIxnOafEv0WIakCaU+SHqy2QVvwkItKO6Jf4vHTIeuwRxt2H6tvm6unlboHpZX+l
JqON+Gv0iTUVVwZ0vWxpXyEWk5jmJZhATPbS22BQPY5QUj8iDqN2fkmRzLC++LlxdaJi0hczutVW
KOck/wKk9oBvlFfE27x3pNuf1qpF7L8TD4N5eVnmjxgw5FRX3CZNurMVc+A4iyeT+/g6oI/2m9JJ
TdMzlmRlvSbqNtu2P61noFKMsZIeU1HHdXDcSOiR7RAXmUoFMDAaPlsJEz4BnshrBajV6S5S4OjA
xfsHG0vWUo9MG/7fb87EyvdjO+zmoz28R6PR7vYCYNUjH57j0/MH+xvVcJxhfD28MmLr10GyPrAn
77gD7j+UHd97AesGzK83pWlPh+0m4tLKNo6V4uMADTxCdUSjpvrVdSPWB3c6j+pU44z+8ty1jXoM
OMUCIZSPG4H8QVr+gJlBNzWSo1qcVrtJOXvWdt/nuhqc6scY9MK9MFvg1UP7xF2miCfCbJ2dTRoW
/0wawNZTu++ZsCUpPPw/akH0LaAEPD+XxPW5ReF1hpe0k/lEjpnxFLvXX5t1VYpA2ogPdBH+Q4Yy
xzPoosCVngZJutmHvj/Txw6iV7YR7Fx/0aGDtbH1QR+K7IOFpeXG4Ql9zVWgOt/I4ktQTMf5U9tu
fHymffktonjgDc7ya6tHOV6LtAdwDkZvm0uNmzPGZwqkldINotdzAMGYvsbgwHxg32Mkc13MLa7d
Xo+faj0CN8T81fFRoXHoCexNsbo73AltVIN3xwwDLTHAxKiunVC9byA0bzWQ1KaDoyJAkL4lKK/Q
puC+n6p5vuKz+ZccEcPfClk5vKt6+c9k4GVj7mnSfwCure+/OngoMrcT/4XYe+Wpk85DC1WPDXdF
dNx4MSVjifQZd3kIXZsg7Y4Ui/88FsXSyhYvuk+Edp+OwCnaBe7jfxnG3gpGo2mC8jeRyUwu1ZY7
6PC/VYzT+zeiWEXBnUAbUbnq9c+QEXnun20VH7GYiK14Norwv7/Ec2As2jdFR1o2gHiI6NWwwLtg
R3t7ukHhh0fQDd0cVN/Kz0NdvJFXfHL6ULQjgeDBTe5478MWM7FE2OAddh4vmNPB0NhfA5aMeAiQ
7akMhxBPvKQ+Ak6m1eA+JGWKcynSsdJcDdhng21v/Whzcohk1YjKtajSLN0oYlkNv9OKQP0roLsu
SncAO2Er9/p5CRCXbjvZQ1cxxiZnzpdTh6OleZLNB78/1mPtXDpaw4uSFgu/DgYfL0K9Ma34qN/q
PJiaENzvIchZY21/cP2I3D/SyNV+qCseChAl2ckJccA3OAgnLPQg22FV3egNM275PYvM0ZcpPyR3
+JSrhmLgBgcO6Vl/DiM10kwxVnyuFYO1HujqlT5J2mueQRhdMvMtp1YrzTylR5F//HiEu+t1yj2V
4lbm0nMnc2kYbuVNON1N7uwmYtJSxDyY2PHuoVAsox6PW+1gFPrLKhvQTbexK2wn36dstF4erpMM
6E4L1hohHFu11omLZ5X0LmggtgEYBGw9M2ztv88NxB52BCkrkFlROqm/IGeaqE8Z09o96EMiogy4
q1iO4NKQ1RK3HVe7pIrwqGHxkUa/iJm2+zJYscH63FFzj72NAovbeasWv0zNQgorlnR4ixyMS32g
OHuO23M4+KqgvT3r2/EsTWWxk/lkzB4O6qaepKtucnXGjW1BroPJ87H150Iflwa4ahvCAvFUnXWJ
Fu/rZS6RvN/fknFyc20dNod4K4+IxX/8fmzHHAwzxT5W5htgNc49nvisKLlx2ORPxraQ1qGfeDUx
/hMQD2TdS+vQyWkkWXsmn65rPvKFlMkmjFzmHrVzQAR1uSSj8J64oHO8OuGLAJjeVKxZVVv3vgLN
8aDvOVJXRKjLCZna54+U2Z4WOiH6fP807UUBIK030PioJ/Cwq3zpKXUi79hlg4FGpsATf338bG5B
224VpKpnstdUxrcS0iEQK64JgLdbw2LL/QyDbrxeI3uzHrwFQ+GVUXOtc6nIrYOhfRQHufiu+YRO
C55wTc4t5D+wIfkAu7tGE4WDApvoJS/vJTmIPoLE/xx3hvLxndmUGnkJkXfnMiFr8LdJbjONoiUF
zT9cuoWM2eitE6QNsnn7t6XA/4FX/Wp3skbymplM/Wlxe7eNeIS+HYSReS02NNXgi78IP6kaMeFJ
s7sWlrM9GzU7ZCKLfVf5c9rGalI0LiVl9bQT03jbduFues4VbrH2cqpy+C/efHYTlSJ6dm5XctwB
4XQ9P745FBLsaU+XwPMw4LD1bBlA2FwiJnRwobMRZtDXk3cnpKhikzUHsgFd2y6WWws82VNSfm4N
JlpTZKVGm9Og762arwzECWeW/qG9U3IqU1W2yjKonHBoSGVQdiRMO1lNE+l24qXv6Lrh2lEICwsK
42UvLFN7bwOKLoqNfTTBR9Y6q9GEY/T15YcQABE6blH9anrLJFk1dI7eau/hJXRD6DMRB80KrbWS
ldPuEqOl14eFwjBriqV6SEh7veTTbYEKXXPVwrA0iNQue5b0zPZXh/wOc8yawHUrW29jwIk3nWaR
rmlk61+OCit/i8KL1VZe8qN1C2/0VMvGUBCE53XukkZ9RnWTv3VQZUhWpRyDNNVjVeKAvufmtXB7
+ZVCWqUGggJP6eue6C1vD/RKZKr/jrp5PK6I4fy7Ts8AfoE9TH/wgg1UfC0zbkk79b4qMGaIAsyN
QKwvZvZFClaTPoGXsCeZJWgdPxOqhh2+ELpXp88m9sMU7rnXfgUBLi1aKLe5I2gLdtiBKzdpWKyT
NUbIyoTFwfjJ2YqyhP4klt+XPa6FHZwu7RqwZrLWoyP8rYNSO3shF4M/8b0DP+Y3SE+a5tqt3uqI
2yiG7uBMR9JAgHTjeuTQ+O3hWR+wTxTIzdQGHCKC/DXSi4pZuNRgE5vakklYA9lhItNADIH9rLgc
uCCQMXQDFgUXBL4Wfc+UlKo/Q70iUL9mtjnGUZmtlSwvGDoWDwzTCY3ZrzqPLxFRcUyz9y045bAx
o+W7inMTzqbZW3ZMw766RCocYNg+P+vwnnDd0jK98TDHXWv15IVksDYOfqmCy5GxHli25CRns9y+
KsCd8Uv4SFfuBCr/6gbHQrmRL2hbjcbR0Gqmw9+L/Hihc8jobw4UFJ6N9n5s6hsK2aX1QLHblNgu
adjLQK0PIR+Y75/MCpARBrgxyqOlWx9uzGCpVi9mwDgAay8Q2C3P+tog9QauAGF4CeKFEIXQgYcG
w8uaULxDrLMhrdx5Kd2FhAOz61YY9+ygAwk4YzbCHtNT02GJkobJKcbzFqCEWW7MuqW7AD4o3f2Z
Hn7gbSmGgZtZnwD6r+XfyYC9c3bBaSUsMkZoaQ13C7PtLE5MVyFgN5wuLz4nknB76MVfQG+cDq+O
Lce3jH9DjAG+O71/9kxvgwBlE8OsvUgBfPXBdio1PvfeIj4pngraH4bamT/YKabYxujVJfjr6QFt
wcrjhtP0Jvi4HhWGHEZf8BmDIY3uUpqiCovOBRpsKvAKwJi7enm1IEfr+jal9uwFwUxXceccacEU
uVYQrYuvrhX8nOvLo9q7pbC5GmQmMSVl5rig6OJGOmgJIK9vsArZ399QRI+N8TbWolzQpN79oiR+
sVPfPN3mxpNxrw3CBkplRhhFmPEe48B3dke2e3ynfgNsq9R7HO9uwKxPjT/O65nD/PvN6omYOYuN
sMU6BOl1l6v5tti9OFOKrd015jgu6JFzL60KugMXDcr8oNYF+/0Wgcs64gLxCxqiCYG3fKVcrcFp
Oa9XsijqdSlsWV9OFlq/Pf6GBCgs6CEDhXGvjhEH0l7+/66hVA35OSPl98DWojnaH0K6OdIzMgnq
hgq3dpe6NrZG8EvplCwAlKOvQCi+QVJde1f/I+JH33S9S3e4l+H0prteDczYzNYzHljRKmzPHV1Z
jP4Mj7aEv1HMQ63HgFWgNxFrv4uwkBLaPdG1f6ajW34zDzZAtowjlmVKoukZzv3MYkkuarvD/bFl
OT9DZu/V5OjoCE21nrxV2949sxrwDiCgVAcb/zxHXCeQWWOUvtdC1MWM8m+R/vvWqASyshXV1kss
gq50I9zLUT5wTR8aJcje7/GDCJgPa9TIIhxxBvx9SSdIhagIOyPMYunhurdLtjteTenbQsioc6Bj
ybQgLSZDZyqoi0K0rAETk+YJznyyDXsAJvlF95iJacB7kOgMenoonPaZZH6SSZxyQKhRCI3jpMEL
nfvIRC9NEQAFuSup8LM34Hrwkm/bgREnr5Nt97Ha6/gkKDxWoDfqy/cXsDONDbf8+aarWTq6X/t9
A2zRyCu9LXdT3c7miTggA17Ngabm5bgyQqb+VqUYCQUdJjDwQP6eo7UT/WJM9M9FxcJlatKp85eg
0Yr0137vVnfxbegTZ/ZaNN3Ml2cR3tV/Q5Ny6ZpVUXbzImN8hAd/pNCm2mcvMJesUOIP0CzTg8N2
K+cWmIgzMFRLC3G7WheKCK/tZ4oIzq13Q+JQpMA2TGE+4GsUPU7cgH352bvTQHqMU9IJvxs/e6wJ
iD6WzvPKHcc3Kb+mp669tSn21JEIGC+tX+4yRwGCVPihCr+bZwxsm/0Ehx9B+bm8nCEEIxp8iRZz
mmzWLSczZKiSU5kd6lVOyb4nS89v1ygKBEHehBvP9OcPPtSYcGKm8Q3iueHKckRxeLxrbv2I9uWF
1zabVGmlrEis+AwdbFzvmv1AQmvT/3M0yOLJNO1zQmpHDJhiw0PgfoS0kLMIculJe4brwDZBucnT
P1N8eh4oloM7gOAPL16DOWgO2MDCzIK2lR4yCCcj1iPi496KvuXGWLiO/YeevFlnU2iAZNFsBQcj
4aEswz/wraBJkqoWnQvJQ1ADMIjOSs0ww8MiL+a3esHEG7Mf/UBp+ksdXE+6HW68xHI3p0L8sJrL
1hzNhgvJJRCE2qK30q0MPMj+ktUn1YyRAvdPgMygIe8GME4hpZYcckzQRzlhO12SZU2k1xKhnJCR
tflfX2I1vbTEImCmQYdg5DdsE5wh4QKbTLY4F/bRA5hkCKaRARIrJBegmYQnpS/ft6MY8TM+w5UJ
l6fMoUvyx7fOJEPg3TM0bntj0eUlUZX9CakLkmYrmruUH5gi1M8E30+e8HSswFDWVRWQkwFNpniG
2MNt8GLvjN1uO+mPgJYkk1cy512lGEb6jzdCWC6T/RxahbeRcGzb0oYMn8zGab4bDLCpjrw44V6V
MbN4KEgnW6W4FWL8wSTmRG1YQfW1n5B/TFm0Oj54zrnpRRpUwFD2MT/+TlNmrRV0JsQNEqUYK40F
L+DRt2FL/5maINLTMPMbKH5+Mhn95yecl3l3tJLHVNzuiyvuhtpSgQAXOLwExQ8akU9GNZ7z0Twh
Epbgk47XS5uDyoQIJLhoelC/pkqiuMHN0gHJLNCWVoPIkxeYbl74TrPqzX/CsT4gw95/HJ2raFJl
1f3L1CIumoYvYUMKFfj3fRIs/II+I9pB5U1ZbzlsHGGHzf2zvlC3Q421NFZsPtQBlFfoP4SrSPqD
/+cYj1INDZInzTy4rS8GI3U7AXz8r8rNtKKa669lfSckQ1gT+liFSNVhhqBcKwGiC/EgMleOsuij
a5VAO4TuFGI+wKClEsYTNHrIljUluSGYKaOpsrzlRTEU4E3HSKvowvyGzB77p+qoe4jPce16ytsc
ZDKxo8fkbXv9PgcVZyOT8z2X6tDBTVKP/ZIYYECyQLcnTfJELbDpxlSn4rDOAzlyqDWNidutD4Sp
9zL97oFbCw3Gx5PwBKz7jaQZcR69LS89gvWpVCaEEuNBue3d9M5cfuTYJvih8RUYvSFdWBOHDpUX
86cxaMxXWHxZg3wTD5sXyN5sQtjk0kM2N9y4nKBx272pb54u0XD9zE5eM7jFGnBIZwjYCLqZxieJ
sZwJkIrK1IFDVAFpv7LmhqD+9S2qHdLdTz0f3M5gk4v97SxEAMAW7640q9v2snvuOQuHJuYCaewd
HJqIRe093qdqv/4GKDh18YVIihdDU7lR0ZFjiM1ttQO5gy03nw24n13cjNsM8HOqbokXR1QpdSJ5
ounml4UFJf14oMorMqim+2KGpqGCgdefeE0o+yeaJ3KDzGO6AOWdBBsDltwU1R0yE+jKdRAw6Uo2
XmUQl6rqwFwhNCpkME/lZRqlAeRKz8VYelVxf97DZjLdMaeKpzQSxYk8tc0B01xaNqAaoShNZDPu
OsE8m6S9gabr2DmrdNClLn70tGd85DX4hvu8E1cKC8NVb5HeqGpbLJmY5r35aNslW8VqHc2rtjIj
VqAZjW1i4on96kXkumPkMdPyFMqsAO5U4xQORhwzVUeCgt5AqE1siG7q7n11UXofGYQi6BLQb8EE
EYBzYoElmsrGtOVA4A3wncRthdBVEGnPN5oQ6Jghcv7C9wstrfMFMfCFRiZQdCMi6BkzpbdZOaR4
j/OXN3sKG8voM/2rfCH9bVTp76jxXH7HEXX9H7UpVl7UjvEzhrA6pLOEwOXu1a+pKwMM6klE4RY3
s6ex4Cqvh91OBoM7eauAQGeRfI7/7siJylrLIB4Lan5JQfTmh7vi3XgdufgNb0StcAoLNbkLV/Tw
KhOIMM0OCJfRaaj+VZzC2NmX21UGVHpzXZNxw7UKEqK+w6a6gnor0nkKv4qt6t3c7kkDhJKyQXjb
5IdDljR34UOHFMo9ud8CURy8gRYY/k0/9+IiF8+yBS1jAyzc89VsjIIlAh5NhIC1d0FXX3uz9Z9F
OK3zjUb3hUIvje2BOq+ReQO07V9PVn8ZnoGP3BB87bRANyRgz6HCv82wH1NsDnb3HHRBolsH+v7u
yRgXK4LMfvekZ1uJkEDSWdlPqUZt1LWnXrYT2BQa3ahPS4akfuOoYN6wa0YPLLzst1kSjEMI4Ize
iaXdgm400mdZ4DEk5JnKwv0/P7WaR5XV8/xlClYlQf3/ixU28VzeZ4G5ahDM+OGAjri9dBmw66U6
p7BSQHVPawlXd11emQJniCw7wOiVoeDQnmVRBiOFN9WSL6Pe4O0Fzq+fy86ekkGl8ovZyz0JIiD8
iIUSyXbf5DVoZDAmbSCkSER1RatgxGSeEoibTvqg/O0J2322bRi1yBgcgdZg53KwiJ1e90tmyupf
CjtuUToSqfclRp3MwZmp7Xx7FZuqfCuVwvWo7EHNxNrK3DW/HL715k8uWeZhuXaFLUri2tNIUGcw
7SSkO0gxmLt7jtg5Wfh5cuCbwUY2ztO1saer4ooWCrVI2+p8Sp18XL7KhcUygz3WFKHj1XuhpZyI
fwpHok1TK5SvfdWhWDut9yMBAlNz7VrPgRfmDlqcxOjSEBEV+icHvkRgSq7q4TJikDaq+9y9rWB9
rUnC11O0eiWZ/3Sjcl+B3FtBYoG3wRVlVl/YUK2dvtWxP79zbCDFFOz9mWW7fW3rVuaCw+gUTGWD
aO90kwqJunZ9O+bDKAadHlZraXo2W+u/PAWDk6x7KKxq5xbyaAf3EkAiOs0IGqBEf/PARNR4aimY
6LdAd21byPt8Hu1+tVWyXTGdeX8fyr9aYalDBO44Y2iR+5j1nmxwa8axlhfKdQLePqSC/bnPZgVt
JVBZaKnCDneGGuyVWU35krMjlnlXs44Gg0eblGO8xn1QMJHQDwFP/DlBKBJMsqMUWXxMVQ7fcO23
vzL5GnXvQThFq09XcEQmDhdIih4LqZt9ymdRt+zxrwVNBkUvWGhCspZiZb1cNQfFlphZvQbBw9ts
62Zhbq7SvdET9pSWGwPhffDzd8KM4udRN6TfKJehj4+tKW93stHzFU/JQ1DaJfmRr6H26YUh8rA+
XTXfAiF0Q7lCTPMn3Ltr4tMZNi11u42aru1WH2e95jdsiLCrOgS4nMWAds6zQcSxfJg16IL+iiej
A+/4YAq6Qqh1kkoIsVpe75TvzzEAQQL0tvxo5FaAAHazMwIukO0POLYlU+EiiYjmEZQ6noACaamy
oYc8+4y3pHt8yjWtBNCxADU5nqeT+ERQeF7uWJoMU7uISZsU5NI8i9HrNGQ/sGKAz0mZcp+ZcRFJ
qvahaxst3/kWaU7WfdPKHI9tI4wlFVhCCdU0F3UnUdj1/ilXyLs1p5C6YLyo3tD8Kb86O5232L/U
qVj4XD1hCyTmBpB5BTds/1q8DtOilvE9pc/iNnEYms6uI8OeKZgFbLLFFENN1ONyORL/bIt0bsYA
ZhWWkgzN8O/enLKKXeQFeYBr0sRED3R2NhOZvu+dmO83CfWqhBQILo047wyIuVIwpgywoO4M1eoa
G5wsbPeH858gNG+hjw8OKx3ApqIqk7vT8hfJtC9hEDa+GcXLAMOSPr/8e94cwMtS7zUrvc+mtHDk
EWS6W5gYXkco9qBFAWsZMFRaXkyKxfmtNNI3oIJHBcNutXPtkRbzFAVWlwzA9OIDpQztTbQW5KB8
4iA3qPcOveNP1p0zbYSsVIAgpAmmCnWoDim/S23BrgYevdnAxe5VfVwdoWA/wMGxfdA6e4gFjT0d
VUzznjWGf5b1/indjwDXBkBvHPWHDw7dI/UZUM5dOkOisNTnHRKKxR1GzxBgU4W5wvncSoP5g9fx
TrbXhRexr18NZa1zH0HZr9XizOvZ/3w7nYShcLBEc2mcSvh8yUTfdBA3pMLh46ULsk8EeGKkiUI0
UVqCXsxa22nV0xksI0H4nMwfaLXoI04v8tEZ99GxgQVDrRs9aqbUXJczNKSwkar4gKkQ7lOGJpAb
/PysqVUYekpDIasXbFMO9Xv0L8nFyHM8K+We0/BVHRlmBvSBxIIH7Qk5S5XYctbM8+BdbucAeSiK
u6/+Tj5eKwvUH/gNModBccV0V6ZWUJtvX6le5tZ9dwNL1q/qETcfXuj1X1xXD5IhVsDfRztGomiE
tGKEr1bO539aP5vWVqC/aFcNh/u7Xyzw+2MuwyrSGs9LKfizGOew16ijnrA+1Mmu9hQFU63kCs+X
n6lCSagR0IEKtMObhUX2P2vI4iL2ii7+DNhqdJBi3qcu6DBHps+rpkRk3qiAAxzXdodLAS6e4szf
c2Eut1nAW7g+jYWqWu+8BC5f7/ncS+aJXb4jLsMRJqxCuMu4Hb7Q9TXy2CKyyVSf5K3WyP0BANEl
iN6Tme6OpGtuF4NP1Ss7SsVsZaft5g07mKA1YgUKds6VbSS6rSXdOF1ZOjH4SVhDi9HEtW90MPaf
P6rkyViLjayVbN82HvMeb24khDiH3GWhfQAkee376vLmFkrDVf6f0l7qHaGrafGZnJHVSmugTYn8
0iD7CpZ5Jt6H7oYTv6mM99r/Y/LquYIcjSokb1SYTS8UttVQ5sypMklMhuZ807Tu+24H8tWuoCX1
TQxHwYXDPsulFBG5ihAmAsdB9P8sTK8VyOYe8kbV09izvuNVDGs8nk1SwF7xZYPKZEniQmHE52i0
9kEtp4rATgx2vE/bXKjvzL5JR7FSqoPbpJrG/5+wqYf64vKCbzMTsgZV6mwSKPFZVqqEGojTIfOp
EJkC+YGfriQGTO1FYYia3HHg3KG0UAzSZ1KB1f21zgrhd6NqX1a4wXM814XWpMxz6fPBF+Vl5ICS
OwEZR96rr/jlg4cxpJyyEmqWcNb8///kzioUb+wwF2z4ZBzPGERyJRVUUMWRP17rtAjvbc7ShSiH
mwNBLcg7yiib0tj722jwDIeuSrfbhtSObhPqP0dMJhUXL7SDwaFYTPzlGW4uAUegslWNjuWC6yDb
uor/Xfm1I51MgETasRUJu7CD2Q5JxG9/ugcSc8ev1dAoicA5wjKHgzK9Ocil5Bg/7cg5TpIl6nA1
LiO5kbaKQOKierOmeRLlF2uVwiuaahPXFWNRKRjwwSHwNNcBNgFXCPgKps80W8KM4CgpKWUEBdJM
knVVewyTo2q1Vr2aawlNvlcxQohZd8vk4bTU/yRUdtX2umbEPeWY4WONuHq7aoFwdzDDpJAnZtAy
AF4Lk4tcKMtzvBLVBOwKX4wi6VHLxxLAyvKButKs27ADYdFrwfaA/yfAuARue1ojIlhyEAj7C5F9
Kgb+UEnAOgFqTl64HV+kPOVLPGR/aiENf4DnqJwgnOGSvv3oPEW1+wb+ZyzDnOGjEmrcWSxR2cm6
o7zJylnBv77RLiCH0Y0s32+SvhdW4nYFyQqxowSL4oQ2njQghYOEtbOVAic4TAb6+aVCBghhm8kk
RLtADuBomewnNdKNgY49JQZTHDlGpcrwvGUPXsIeIKKQUlE/1tVqC9fQxjb/ix9fBXpba6yE7byN
RtEgPe4A80auLlgE/t5YhlBg3E2CzFVhViz7MmvpRws3xqmyCx5sufwdD9F1Wlk88WjKPuv/vcts
oAL3gNdjTwBApgyHgsJ+yTZeMFjpZncl4MuEXjulQHTz16qINJaEavCDyfNKmpQRCp2myuo8aTWR
ThVsqaCqCyauFFHJC9RQLVMoKXtTF2eS1SCtimVyo8zeXNJ0SUTA+wpnDQ3ox5YBqDROREhtSPxE
rfWPZBVIw5bc9rRsGXsqZPjnmmWzztVyR9Rq5lX/MBHm46V5Qdf8QUvLOiohKSfSI4vCXSjyfsto
pqo1rJe4hIw1W/TN8BJ+psu3/dN5qy/hd0B8GI9pNecrtoOFuuy/pZ2gG8xFj3W08bp/kMXN4oRW
FsIW1IT8c/d9/gML5ASmv+IH51oDq9iG8DO2Rar/Q1ByWcLzbzjTQFpU8HXyyOwWx6klnpkBoT/A
p6uU3PMVT6uK+3YtjVHM2gqPQpiJpDi4k1R6KJ8rTkjZq5u/rCJZMnsrnh8M3sPeuBoRlC11Kybl
HFSM/z4kI/WlJsVHVcXTgpLyJZF9jyRnLKXfsF4GcimFc/CPDdu5d6EBhNU9arV2tRU4J0zNssuP
B0M7INRlpdR2ZvbbiAGqRArswFZem3q9adEonkR3LCNVXTItsykcqGQQo3UjQUngaln1/LFbC4bO
VkxVNvztvx/gOakq2VBkUOIjmYqkbzlM+EeubdeAQeTcceLdkBo7+ZOcnVzN/bqBG3Wj4ljlQnik
v4RaTOHBXgjM6aTVkHpZu30RWMFoTlvchOoFmedpPfaA947uHleFnQt+J37UutaveNYD2uNtsYMB
okdF/WHmV+UIFVWaau0UWh0v0mJWW2o9eW4JdXdSbL78TXo7ovh5RZq7fwppHULfPhjTpYURtz9a
8kI3g72wsrcbMzwg+Lf74qScKe2EiniOzjIDASXFfym+vLbsKGmbEplRtlChEoErp6IhWEYdnsKi
2wGzcivPm/IMsQTdle5Ayp7m8OqaiOeE6VRgtffEbyL5V+WfPd+DUQNtkRogOFzHjR5duM+goJDK
R99ylT4/Vse8MYsNXu8DJK/pn3g8gIRJob9fS6XTD86pvcm98CWg5UaZt05sXr76FcDrZuTJ51Mo
GG3obMPpCS9kZv/kolVEXuD9FoKnBfUCcFtXnNcsLdqVpXG8LWwZI7yNciXpEGOueuDFO9qTJJ7r
EROrkFUBnuzWRh0dIrsBFu6EfooTAPx40Xptg/Q3IJ/4AYgV+v5QMbTjcjxHQzpCqF1C7KFZvYEm
kWEFjp76pTI/914weBCUfyKjCVOqmFae3dylBKctvDTFCpP9O+sHgOUDOpJbND/rkzTAwfiYBRjU
f81s52dCtzbhEJijBQrvhcg4KFbbg8wKajPlpAS1Oh7GYNywhG+Wyt6hRof5CE6Vd6v7lBQmbRlu
9E6+OOpG0TYlOYSQJ3KYTW+6dli82htqs1mGmG83kr/z9YBvjIlKJtXtfptKp49E399wRX0s+3sj
TWSabworw4yQOAxAAZ6cNrJHaXRc6LtLOJlMOtVo0fvb9HU4jOX/IGL3UUXXs4+6kTIdRgvcnyZh
6ygGgw4nubSp2fptz11VQ3k1wShuauGH6HlH2VWmjxdxKXWERKlKHNzL6hNCMxalraQ8dd7NGAb+
n6kh48J2dsZSuzCTxXdRJNuy/gs/+RhwvHeYHLmlC12CrbfOGgJ3Bdfr/5IGxJB5rlucxgQXGAKn
5kwmIr1oofVi1Y7RzzKKTm4QH0mlqQmkmu2azXL3tb4GhppU61o/eJNfgcq0LME7SpqjSFDQZHqH
cN8zBO1fIsFqWI7dLFMk3odsAhsqDkCjQUTgiD7qtsHUNWLjkI/gSF57LMqJZyGmHQm2QwGB/6JP
RVZ49tQt1T8LtBIR2Y9BBJL00gJpQo9jZWFr9x2AcS0XC8GQ865yLNVyM11l+A5x7u1tMMjIUsjR
CyHOLUnng0K4jsLPKb2PfX/rtd48fVzb6QejDQ9AIXa50d8Msg/dHwzb9Q4fGEFxhLBycDF9/Nzg
TLNEddTngGfYUmpEgj69Aupmk5dhdOz0BAoEEOCxOazA9mnzoJ+ZQkGMrebTTcy35r9Ix7YXOnLZ
NfW/5JNDgpT/qeoxRYMBJEIW7nMnDhYwxfPQFH7VSJ+yfugIoBB3isG4QfACryBvF+MJVTBlZozC
3mSLJSpZTS24aS4QmqJLoEsX2NdUfTwLUYzr7y+3RC2bjOTGQr3eivIG6BAHHDnIyHu3LuC/vaXd
tmURzoU5p8cdC4F3Fxno5LCD8vbOPQQfq9qT/cQkP45bYiEYHeCmHhd0D9801npX2a0zH1ozhRIO
CdcHZwVNZmgcczEoWMJ0LFMAL5r9YnxsY6WqY/ojgenur6vXdbvbiNOgXqFsNPI0dKP+rBtWkBUc
ICGKPtu9QJLPMuZiPi83nvj9C/j2F7ra3Y7DkxHXwyj5nQglcY9a86A4VbJ94ZGR3DCH/6OBxWBB
1eSeyY0kZ+imKhiru8DTsLgV2b/VUcJnxTzYCENPCXYHaY/c31vVeuPl+z6rF+3oGmIanE1ZDC+8
rNK27aqr/msvJGOmMUahLDL7UD6WsXqP1siJt31Qj68ELzQtmAkieFxOchVtNFHOhZ/0fCAbLpOA
GLBcQaTwUdhDD0tnL0SapoO2S71VSQkNv1muv3QaLpDIAHPxBOEAw+CxLlIs1Ql00tfLfx8m3VTN
Q9xCT1KhgpNO2Qdu4lCIp/PCfpoQQkRlI4yBEADtDtRjAvnSps6MhewFVXmYLIQXCuVUv6tErsQx
79rWb0TZemlV8Hd7mKymumXnn7ZFkaGecuh5upOZ3UN2/DsUOrIhyRAQBucL2suD6L65NZfYwRe9
QZUqe+vjsVX/tDLiZVphcwpR9lF53IoWX7bsfPa6WmSXY8ZU58mtj4w02mI38kTsmvEegQ9O2Egz
HC7Hl4apBesbFocwUO22TXaK6SSB++r9CgGI2Q1MtmcGRLMmhI297Mr+6+Nh9hbdzP0pJQPNx/VV
btvQdwKGlPb9ffy7Mu2A5LaAMpcYszZe1xHjWcLy/HUFkPAe/p3rhTDNljOp05fFyPdEx2tGM67J
NlccMyDsWVQd4t8RYKJaVx6J3aNoIRUt2YJq9HO2BZkOM6STobqR6T3cGQwuHeUyzZ5rwbHVjk0W
/RUb+0LhPv4tHKoR1+N6mG9hRX0kMMBJQ5i5dAQqW0Zsr7njPq20L3ln+1835hJGmujTlqG9PCqy
nznSolczBpO4NmR5hgF1OzZHe/0fafkPVJg3CM1qK1tq4xRLN6DPAidrOEGXyrPZvGLFQMktJ5aL
4GwEDYIFtTGq+BIW8DkWy2MnVB+bsrv+ZRcWOn72x8R6w5siBZJEQpvPkzoNMunKeFTUatOd1NjG
DrtQO98Va3GDIW4JbQggWk1XS0Lmz58FI4bp2VD3FJEtvFllRKJOm7Z1vOK4VKfxrDTgrF2+uL+0
4m1utAbS45InAcDlyNGt357+EedVmhjs0gfXFb1yGmdvMWL0J9Epdl5Wy/S53mtcy2Vhw5m0S0+p
QLlaHV4IASfEyCj7bpwXmhnT+Nvf1CRky5hny3V0Eq7CFK/b1+RzYfPN1Kz2sGDswQCt3X+vZIXe
mLriWMR0S73Nt18FKqS7WJ9TcCx1MDaaN1xdZamx5oFmuNAXtQaFOSb3pnaMk6o9qR5i6fhKk/c4
3BPGpQd+SrBFgQnQkGiD0zaYFqGCvQAVr+WsQC1fS14PN/2s/lT9l9vjW6cJI88JXrcg3wHM3PNd
vy3uThFgqviCwfXw4t8JbLOzHZWzxbqwyHJEnHNIsshsi2G8teGKyn84CVJhmqUdkQtdaqIPMoh9
QP2r+kNdQGS+aJOuVWZEIKVvG2bP9ANp4K0TtsysMfMvpD28DGwbyW14A/OWJtKaXHcMpeaKGmfl
H1D2Ein3XMoGBdYZuYK+2/wqnK67uPBQLROe0pUPZzc3muhnKY1/cOG5llwJSPkiGFqWeAd3/ySA
43eu+ABvLQ4bEY2AXfbZeIuje1LDZ1RkuLAfpB5+hsueYUH+wcBjy4pYllcEabWdhSYGXtG4J250
f1OAN+EOubaqY0E1a8xtGjP/Mj+TQSNX3ieK+gYvLh9dAdzNtuPc3eqOosX9mAHvTLMBw2WO9CKR
1z6UPtz/q+cynL3noTlOEQTh76HRCbiKuGRpioVAwi77KTD/fJuLA8HnRgxj/26+MkuPA8P/G3qq
H+zlMvHEDe6gYBFaNQMRcN7UKT4TyR/cJjbK8XKZtsWFiME9DC32i8n4ECk1fw2hKZWWrjXwdIKR
0X9ah4bIIN87/U8KelE4Yj3InDwfvYxY+d2LABVAoDnsB4x0DIbkzLlAk/CI+WpvLw+3XOcQhkEL
7+UGTKbk7JrSTvKZ3eG5vyNro5ut5F+VjeF8pCKBB0UwAWuPmuZNqNx8P96qbtQbxzV6nq/WrSoM
PmrgxjM2xs9vpyxl/CocVqC4k6yghm1rUeTRQioXEkttWgLEvPkfeRazge/uPy0Jm7gR/QBkNuDw
IxdhGBnqLkUWbQqVTZcmkO35ck3bq8oASdQpca2a3x7YfAJba2MCVkg0SdsP3y+fu4yPC7YSgrnj
LIjxu8mMRNsc+lqJqW3iptMg8nwq8qImL/FDMFt9j3tTOYvVWKNDtj5q8HpjbH5YoQT7hQqaPY+8
WuyxxBXYbWUFcIy7TQZsr6rH9u7tHabyTB9Zi59iWenR8bHuQf7IdS/xst8djUFSsKA9UfLn3m2A
BZn21c6eZqdUfqgDOVCOuOjSqrwHHDcsgO/7eqBAtbh7oIzfaCE/YRPVJL6PtaJSz452UKXLRnPr
1QQ2fw7jl+dolbeY14yT/s5PxpBJjoVk5m87VGEAHx7Ups1ZdOWxYQpPoQKZ/yOsa+Ou9hw0m8bf
FWlZFScWsWT2W6widUfYuHGQIzgTuHV2zjdixCQHCHQPtFpLCYnKNvUIIOsegbE5lKOLOln2XKFs
9TDuOSzcCFXgBwK8tBnhsr1nTXgQOFLQPQJ19ig5glLqZsDZVX9SQT9KYM0x0fUokawwePo9CTjZ
p1tH7OVxWB+U4POzUKGlrzB5IMFITVhRlSlkP+4BS1OJ72IsquT2dWKvydnmbRwW1MosSCcR9Nlv
gC/vybOWoAUn4oRgAN7AiMmd7BRjNDGe90ubsRnAUVcPpunpwdllTUnR7kv6ERhxQ+5a4fYpiuIB
1QCs9HTYYL2z3WJdURYq4NZkCgZ7fxORviudV2OmE9l2wq13TYm7CCDGzP9AJNxy6rfHneK8aBE0
TCCKco833birO9cE+448jX6oxfMeWWl+xEZVwiQs0uhYc6j8/8p1X+CPzU9r5evt0QVbufDuuZRt
7JFJNAJORrbXjVyKwZoyLAVC7T9CTJAJgr9HffxvyDpGV5D6zO8/5sD1geAjHvyCt9sKv57pM0EV
Wi2gUIA00oV6wVz5SiBImNlAazw6Jv8TzFlTUyjj/W4QDjWMBrEMot8AGWFXjjDyDfFr6YY3FTwm
lvJtQUm99DdKVLa1Zw3ZW3RmFdiM8pO/xApS9klLCrH/3qDiBWU0HHXo10lDvBxnUgDg5S5ZA4AQ
ST7FYolx/nKXvkCD0CGFmJD1DoWDiChW2XJm09dL/rlpMH90togXAYYqVisiZ8Ol7amOSNR8hzVJ
F9wogZWWU9sw6+kVzXhqNIXTNsFbif6DakFpBKcWJoLzBO/ZawjrgZUBmiVehgioGbasao1hKNpE
qXaIChyGOYQ61vCKMFaezLtkK4KbVlJWpDXl0Bg8yvqUuQb94VqceTEQ6WTVFalaRzAl4IusvPHm
pgf2VCCDIunMFu5pt74pHTgM7xFnHFgx75WSgCtNn7C0OS7jIATxh0xArgGeM+iwTSl5iF2EKzlK
rTC3fDMlO2OXxVWBNC0mPHrbEC7lpvto4So5mAjcEcoh7RugLfllvidqk1I9Gy8OHLHXgxkxPvun
5kC27sKjUgO81As9fUF1NBSYfh4mFuFS271yH1O2/Q7dyrmswH36Sv2QcUNAn93CYjswcitPF+xu
HrNQ/bQQol2cIkfSGfAMZW8i/ZTHlnHHT5LnGJSjN7UM+OJNMHMVKyeFtKDZAM35i9o8maLOOuQ4
bt3onOJwQplbsQqdI/3eAehI1KN/bXeBBwExDmWUFU8RDO7uJ9/icCMD7jdgT+N6XRkesLyvUASi
9Avaqja4WhG/CUi06XXrg/P0++ClFepSmPiEg2xCuDbUKUbfhCVTOVXsvwrSc6meQXK2XMgkkHyG
l7V9oWEh2ad8XcgKM3UWIcy1T4FmvNqgEN7TGCglGWWSiBJwIAlzcZQHvpRsDXdGq27quwsEb+b9
Ggd8uAAiH+9A1io4hMplPjrGY9wNjeTOmHT40iiQHqowdiOhMcZ42BDYniOk/yB0/bZKiKEhymfr
cGMy2wFPTHOmu8Vp9rVyv2vQFXYIGJpraxsYtt0+hRUPSxfgMT9aZ7F+8Vk/a2HlfK/ztYDxAl0O
KeUqVkVyAGGbFxgEtpadNDNJOptiqMhGIFBf0ssq9ojDED8+57ulQWS7QoAbD6w3cDtLIK49ziJ/
lDhdj0B+OrheAdSPbvsurl1nIF4sW/FzvqTKJyIC4zPF2Y3qSG6GpsHgPKXm5vjgxCG53gj5egcx
bCvzF3befHba7OxWcrHYvH9LiV21FBzt8/hZKOkeTS/NBugP5OyXm88SuV0YM4s9iXXpV5+a/Mk9
sWK83FKmhZM6vILAcPTQnlkLkrdzLTEXDtYcTmesT+TIBEJOhE2hCRpy9i/jFMb3fX/uyKmN10lD
IlQ5+jnS8TbcFnFnpZqjRDsKFlGaMqK30kJmp8oTWcF2CO/k1iEypUFGJ6k1ruTZe+7RiycZYuCy
dxTAyNKdRzMOja6bsA6q26mQg43RMncFKeypTS2PykVEzbb6BLu8qpjSdxYdq7DxUj/34Fvvya06
itDK5DeOUc8OZ6iTf1Larc4QOBd5/TPZASPUIRQBKeqMLdI7KJCFyksNtei03sUyEoZUOf2rHMjp
mivtnxPc+ZxDp6kjGxKjOy7Bv3E8oLTRCcMB+rzshTyDd2XDtZcaKNruziEM2Xxoy7iCQ5FyhQ7J
3Mm6ekRiaHYkIMBYeNIOM971SNzynRUSU5EbQF3FKq5sJpu5vfOZ3K8GHhpXV23wpv1y1Hh9uLt3
NhI0Asj2W0LEoYr9ROBMTit0KoSUpCnXzStt0cz6P/V7gv8B3JH0S07icpc1oT0V5ovKaV2oKxCC
/8GOrSl0ac2DbKgvALmsk5FPVc63ePuV7oy6cw+Li28kRXGsAYtp4BgoKnwVBDG0r6dLRpnJQvCi
BK2tjI26ltd1KpbPrk2BtxZ0tn8O/k+98CDoPtH0S3vZy69YknVQdudVyZ8osz49DGudWvA9bt7U
zwj3bb7lnxDktf2CNMtVeTYsbFzLlvC+XSRllMP5MccsGMWzd+r4VTnP+ks0HKPzlAqecKw3kZwB
32F8xl/IzrIDXYDijjQ/H8meXcR8N6T5Ss8IIQ80ClWuCyvyKEAi5ux/kYQ7ORN5GvdCrWMBD5Bt
9DeYTmOyF+3SdF87N+6QZtY1cnNkGONb3wJadcGrSE6DU8SVhBDLj95E0JZFFg/vSooXNlkieZjA
CZfkEuacK6Ubz0VZndHBBdY7370HZnkg7IuGn25IMEZURH6I8YF2OKBICTF/1D+zPUSIkBkMe4k/
m/O8XKlmTgiDAu0E5II5UB1N3hYmClOkI+dlcK6LfPS4RZOT935/9iOk++BfhZlypqU9J7I1N+PY
AAJjhFwcUGCR9tHWfx++CaOokEDV4XwWNTTZhHixOc0yibgWZQuolSVK2gHEAbQxj8Zk9VShTMQq
K0O9AstZGDUPy41Gi0dHe3x5BY65PqwIVUKFdFowIdEM3cZeHOm1Bj97KkpKXLlCAbPMqQYOeffG
K4/f/Xx6CnqvBV8CQxQawdJyQ/ujhem7ufNddgLUEuehBrhvijicXTEv2hfiHlPhQWZxz1YMaHjX
YU6OptYq2tKVfkD4f+4515iPOFXQ73EhXFhiXQOYrGGtSmDQmCe02zB+mRuQ+GtLjG/SVuA8oDZD
wDrVdoIZcpJMAKQbHwUtZTGlUOwax6Otcvz+SyYQMWUmKMYTumT04Deler2Rw9WFTLzlc1453HbV
+vnQqgMsuhlpm8lpMQH3f3ZWWMjTgdTqsMIgAbbVyjXYlWhZePEJwuFhqXUFdO+pkG80Rqiyq9Qv
BIMPJHQZa1RCbKnD5SHn+5n9UjRo6nNc08zNr9EuBT6GtX3805Dp7o2vb6I+IhAaVGV59LAG9Kz0
HPfphm/H1Pb8TmWwdFj9FXBZo0HjRSXHfxCGFhyWISY9HlutQ1Gp56mvlSIgT9/ZyZBWX4kmIESY
AitQC5myZy0sYcHR5rV7uZOUR1OLKwXKgdldKJIQNJQN+U5XFx0NQp81ot/qx3H/sY5YkjuHBNZE
OTYY10oQz5sVrV7/NjS5Baz9cnd/dY4yyPqL6rN2qPScfQXEBH6IbDGVzJvuGW36LEtV54QHllYV
ZLuiWMjZsh2hRtcOK9WrEk0RJ37GF1+3E/H9ENf0938WvI1tXEVeHwbY2+BMSqc2y9mxedN3af2i
Z9D7BZlKc685zjh41o3UHeXVgVmAUVfszs/TYbicRpp/CHyJxm8C7OfoFzHL4piNglTuPMBl7bEx
Uyaft5Mzi+4Ih5KYNqC/Zov/f8xqZTbi9jOPG+XnUydlpMY9OzFYIsh3su3y6JA7jqQbZvjRZFQV
Q6AgSvOLXQuVVnzwQaYY4tn3CxlWSo0+oMd1kA0TcRScLSEQzHxgMzalzHapFE++PZ+URuM/mE4B
9Hn8Z53eEXwAsfG6E0eJngsNCGJEL9B1vTtH9Cb65sPv6RpWxYWVoUW1Lm+BZGR+eimW2FyhAzxR
c7be4hKyg8OHGm1XBJr+PPpvVEfQbbcaI98Yav/v3OODokP+h2PCMDQIMb1ReFb5s5UmtmkWxLbs
BpxKHrbKfhn5d4AR1gRYpQMun9mRgI4O3Yh6FPxuqfKYhxl4LFwGFXpHJNXTu5WWbBV6E1xAKYvp
qq792fBS1Q8I1WOkcRED6xohjeJC+Clq8xLe6xQaRLdWG2TZZjaT1Ek9lgmdEdn8btO6p+Cp3cbo
0NbgP/o9XwYHLAvD8gwzmRiPisI3Lc9tgxQozCpvdyCvZXacwacWnqO4duao1Jd49SMhAtFKShym
jCjgHiBVXlhAYGVloN+hJjgu+kKcCnrZH4/GYpDBOx98E8bQ9/b2b5Z3h5+VMRyP/HRBNRyAV1QU
IzHPGs19df2VVFOqQ5QmWh+EwXz+fjLpkrcyG9o/a2Ix117K09KtsGWEbsfzG2ERMzLn+7Il5kws
WOJK5E3P82wtRJGo51wy0oPlC3WlNK7nhUqTK/FkAT1mKvXcLlGUl7zrT3uvIhLyu15GmaO4xJqe
ifQaodpYjGQyUfZU9/p6dQ2i3KD+Qmj+NCT2TsoT9UJI7/wn/qy/WhenJKjuDr466IZ8bm1TvxGr
8cwoQpke7jQQ2fkpLVDhxiILwzWQRwkEnGBTCPfiKthBEnlyhf3dzZmVRXn+3WzCVXw+TUmCCcB1
ypKj+maphlzHdFpVOwYOe9UhosEkXR4ggzTY8P9w7xpWi5gVk7WQnCxU4gFhRGeDVv/oOPxdquza
NN5EEwaWlPq2lbuUSC+C36il7DqIPCVIWFOxodcjFjtryCjMG7uTqzzved443pGR4LTBpeLw4Rmb
DmyOmxYDMWqrar42IlmCusvpHe8EVuLtnXWSX3CovjDQSkopt9C95/po4iUjwa3R5dJK49gxOh9e
F7gK0Ji6ODS41D6kH9W5sDDyc1qxVYPM7PzfNjm6iTdQHv3H7KeuXw2JbKWm520ECQekLTFc4z4m
bufNKBXUMANb5Qmtw3UG46J4+bsa647IV05DVe6EjdRtGsmbRyKp13BJ8J/20trblnjR2wmPaFA5
AZzwhCctSHuP3o0vQJOi3etUN1OvznEyTCNQawpNA38GUO14MHCzFEab1rcPEdw9KImoxWrGc0m6
lcEx7fzGxnWrE3XkYMuejWUTe+9FBm5Jq0xc6Fh4gN4352Q78H1i5CGsiul8Rw6Z1wAFdrvtudxF
e35Mgdt4I+hjsUJoeFkEkElu6WVxkMCuPHf6FEuOyNISCLrWsbOUqc536PDx1UK8p33QRnXMfIV6
LVO2rQQd6EkpTsS/P0KujMmK60fkSLr3H/HR1xawCdLWCZt3Q0DHzWQp9t9lNa2X94PEDuMgEeQ/
6aEEAg9TkXHcwQ6+xqshiblKyjozLconXvHNGX2Mue+Yc/GJsnNSxCpnST4P9rHO386jQElBv6Si
HCaxj1ULsrIV2dDlR7ELFCwCApr7akbBaTdLTUhmQPVCE3wUk4mrqhQdY8tvqutnuST+M0lmVmLw
6fRzepkUollZ8yJ1UdaRdYDfNDoqNKomihFcEyIyDtr+jjy9Q6LjRt0sa4MURsFu8UFaZ+jUQ+6m
xgOQkYsiboi9B7coYr7hfD5XOYoRKD6R82Wcv+UJ+AG8OlKy9IxAP47FJUQFMxbJhpmVMFyYQqgr
am8I0HoqMdJk730jF+19GA2FCsICy/jV7Gv89Sb8wdvk/vaIRAld3PFp1YAh6MzHi2tb48kZmf9E
3kK058W7Jyv621din8zhDBDkffmK74ADvX55TD2OXd5Vv5eamc3B90ZsJkewuO6U67ZwnETuXeI4
OcCfmzR0V2QOPuxIgOVCZAysTED4njKSMI93iYptajharnvmvOFu8ZGaYFb8lZjqNiFTYmeRe0iD
yx3Hp4FNvGgBKTT6x39Ka+K2UKgQgy8WFkAun+kc57alyeri22vb45zpe1qMM7PiOfXZbyM1mM3z
xiMN+rKIyTjAxjj4mnNIFzt2oiAEp/WypptZBvzWSkYwHjVsyAZfUbr2NpSqE9TQOdPFZpXenT82
4i7/s0VDiJPLXP/sRAoBzNL03LqMfLo4V0jCsMgl2AjrkO7vT++tJE1r3ZsOLbPD3kVCj7wFb5eH
hy7fedxqGbWsSCE4LkM1tK9GhKoWuehuu7gC3T0m6jYRUFJCWoIeL5Qxms6q2OyLN3lm+csn4vyz
hg5+1fhfCDJhBqDX92C6putHl1iWgELZ1S1QWUd+VF8oW8PcUb7XMYJ94JBFwTACnBKubF1l04lv
944cFvtNHLwTzFzUi2PoLgzkbO3WlGgF7xRtcF/a8RZYKvAD9mWsi5uBUqGvvyrJ8QX/Rhleyu8Z
/BtA+A3ILSBeNRhROnuTaQYaJeA5gJgZizIS2FBaEWW11Lsi8apyfVZkSQeuBALfV2AOXTSSUusx
jKaOdqypoqH4rew9VJUbmSEkuV7/uXSUh14AJtl/tET4tEB1CTVvpIeC1cUnY1sD73Dv8O5eyEro
sjwlwfQHLiIBUT06cM21Enyu6+DbkU9my4fbAkn65U/DtpJ8V4YzJRifZ/o4LEmw69L0BcQE1W+D
PQ99c5yYDfTicJpZQCsc0tYFTDdrFg7Dfj4dfmFEn+Hc7xNVgcP446iuwpnDGhuMBiYCPVjKE32X
uyY1gyAlU3KNiAijfQ8czaO97cL2985SVDLrjrA51JEzxjC8jq7jnBioPEJpAYcwMsi/Khh6WuAn
9IHkGnhAlMk6QaayvofIaTVqr4kGCHCpDgUM+JSYy8h34yEqGWQ2k90q7bFYeh7OtW9Ii3Qejm6V
fixKYMf9Ca+quk1fhlVhGtAGLJm0qQZGbACDlNdU0ZFV8IwXJoh3kwnTNg6WCzM6oFl30K/sqMLB
1N1mVNtQYbiajZIS6D7VSPO5xSpmX9bB68MwbXIgaaUlpmc2plIO0xR8Mz891bvpI4Z+pgsGpTNa
WYVd7QwsAwfwuH11lyN61YCaDjheEBktUIKoryyaLF9v9f/4DaU7nozOisprTYrWirBQsJdKpgCZ
GkUV/d4AOT/aO/2rzqMmWSnKZnWXOOOVlsTXMSWunlXwXKhmMCtjUbASdKGuFtKuCn1jnno5+nEm
UXXuoz83rEWhcEGHcT+wclnqbcEvjzTKdESZvcIPfhJA3OwUEnWmpp0cQUmJX/Hj6GPX3+MO1V11
7BGGbQLNGMW3zqp2EMIPc27TBaLS54vA0/tHwq/0VYGcuJW6De5OmOoS07DGLo2CBSFJSQKhdaGW
53tXlmVpxgllQ9Zlqd+SoVhqiB8HYs4N4G8bgJkyWTwtPob5GxNYbrnELKK+GZuI4/bNv8aLJN6w
2zKcI4pAPFazaMtWqyn0qDD5Yo2+3qwn4XrmFeU7gBIeoZ3BA9JPkN5ZNCy5rIZ0sI+aVPxI4cju
GQ7kd/17/Sgjoh0msaUurs0sOHKbHW9cWaEH5prYlVd84HfbjnXTAH3GxHpZpwAlrcX1OIYj9G5k
OSJZZxJb+XuDgiu8tr4wxFPmyQwI4TxBMcjSl4CDTF9ZxZu3YZJhmaM2+6fvkTrHcmt78PdErHqr
p+Wr3wwTEn/5+ysb8rrkHaMlaMb7TrrdTzg0qjCaIlZK3knY9wLsVdJstMJ0dhlbnO9Suksw38dk
9yNgSKfaW4d+4L38upBTB40tig6wUY0Pqf/mXa33Ys+bT9q6QslwqgnzG5WoyTBvH/4pajdfMBW3
iWW0AKEBdUzZ9iEMON86ep8uymlyM/1qxlib3jHmKgBX2Q1krwdajyq4jbFTN4X9CzjF1e6zI4ND
CKOrixcDGkizlbODDoPrwnMf3EWt5FEQWvx+C5T6yi9I3pxeRrb14BQPsfRfEYHrO6RrwkZZ22O3
FbboMAqpza/PvHpCdsRO8bfUaU6hQCFrkdBxM9yPdX47li2CXnaSRjvrfJRjxB6nx51c2Cha+dIk
q/PoRaH9JXBnhbdZK6rdugAGg97X/TsWZUTDNOVJVZ4hmpP65fLF/AVCgqSOpl0pJHPofzksdVZf
W2y5M7TnFs4VKE+9RarylJp1Q0uRk1RAPD9zXCtSAVQozcvQ3VoL0q0YlHkqdJLslPVjnOFAufxR
9G/hnFZ+r2O3SNwJdx4DgjKIAoyuTSNgEp41WauG4RdsZDgk09qgGi9pz9ScLXn0dcMpl9DC5ApT
H6jc86aAuE7nHQicxVpmIory50vBwqwwfzwKEDhr1Y7ht+Bx06I/vMbLwFeqMSOkOSw8obvQC564
30qN+wGZJUSHIp49pXkRjbrMakM+fOY44/QXefnAmCJpISFppngMMVJiGcgxK7+yswqqoyb4nQ40
P2ikKYpVhVpJ81ItjyrtRY2DTbLF5/pBMaFXGrgapglcswUohfq7tpyXtmJi2Alg28BvIFAKWfep
jl1ZQ6IAqvd5vdEXH4ip6dmyaz2ThcaYYBFvzq32l3ZABxKdxteaXyj4NfxJ/j6+FmdzW/tHgiVY
cNS3aeSxOOJMcY6MEDwMSKZe9hmie+tcIUIPz7+sAQsHQSWMwCuUehR2WoaV8Q349OekXStthHft
EJkyJhzoW7tQ1UX7XJ451WLjk+KMZhm7C0beh21Xq9Fgt0ai+CCOhSsjg12oiOQXnSq0reLfTcYl
HhxkG6ok38UskdE+S0UBXiX4UmU60eEzWXNb7zn9Iwta/hBwYFhRHTRmUFWpeLkgsdb3r5Jgjxfa
ZTzVSq2AEifm/eCRNQWD9jG96ed5D3pUjroOdgEFJm7Nfiw3zrs7M+BhoWmI/kke+I5kgU1GcwAL
287RS8ukzYrvnZAo31yUewJBSegQBftfpjmWQ72gXvIMF5uhKT108+bqF+cIWGYh1tcWLRB7RYX1
Om2R1oYuylzeG/w/NSbJLBIN8XNwwjNe7bHFWKEu1+pBMzjSA25Mxk1jpdJ6t3ag30Wg+6Vwaza4
sQiVipeKyFF/SFJNx6wFvr1y9ZXDREWwyQuH4/kWUSP/cZ5Xjgl/62sz6ayOzL8yJ+MDO42vSKDx
WqX4Fy2W7aPS3JTSGrnTc4uKY9j7Kf7FWNU7nQtHu0c8Dfl7dry8o1GNqeUvQ07cDBHQQHIEws34
23cQXqm6CZV1OsaKyiqIp8MZW65Teb0VaNGq1aT3gYaLI2YVMPw+QudFgLWgxtrUU8sdHo7DVNPF
dSn37hY6/m85T2DhWJ1SJY3pk0u7jvkhuamFL3KjjRkgLnO7Y8rH4jZEXNVm1tVHnhEi7yjMx71D
0JcVWnwYgYSOpo7IS44+eNDzHRI1xKg++bAWFoy5w1bDUFS5VCTvPf38jEx+cmfCK1+JW6bW0eFA
82CcsZjM+dn9pZmyOuHcX2ICUgNpbysoDKtxnDL5gKKo511lT9pKH/LdHxU4qdIDZLOUhwQeraws
LsJwOnMZKKPXC34GCYuGFoi4VIHQQqxDyQLswix+/krUhUj1evHRhQ9LQTfkVqm0JgkF8TPkuxzh
6e0eADYYHrx6AAJAG9p3NSZDnNVu3OiSgTqeVhDxRsClQxNWfO8Fi88jFRP64Fq0xa98v1LrydbH
qfsl9k/vsN/Q4KTFmKvigajcyqcj8QPzMIGwjX3t6gAnB7/hK1jWZy7G9cql5raZnI1eXez3bKmo
rzb+GUskmUXjZWJD+1utD0gwVxRcujfnmLwn34znE839GMEisxYnsNGJc2Vr4F+sQJGUz5AS8NS0
G1RXrQPpGUQxWh+iqzmVnzjszlmXurFNdq9zlqFHEO29JpuI1/2HBlpXtYrH+/Ww7UojS87nFpcs
7FqKVbRakzk69v6EiJrhuVfRKxbAjlPKi3VKUtkDDkG9ZKuvQ9jehyggXP1JhvkUce+5tJBwt+lw
dKsZUBc2WeTvvU09hc2useJ7xqzdqXnnlceclDoM8qRrnC7R4+WX7lIZ6nCXtdMWQrVSnNVaqOAV
JPWr9lW9P3EexCXTexlyfOQOY+upxknKuOQB+ROq75UW9LwrJKATnm9PkEUbEzrqsMKHP/U61IG7
jD3l2W00cgfyRPTn3ZYTZcmAu/TdPz0t/1Lrhdcf9oBHR+JaExZszW95I3Dy07l3grP5WBqHeDTs
+gGCP12/8kqUU2PHnO3YeyvFLCZrqaEMvM0oe7/lYLH5HAt4U6oGs/NvoD+d4u3RJqbWTzbLvsKz
p1WsnUej7XOLvfaLED7RWtRzmXHKW+dw7TnYe8FBJy01/siAiNASwFX6yaNE9u0rNcOFBuS8jQ0n
ezpg3bjABYK6L1WjyZKnqCwY4yNwZc4OOT8uuNdmAG2DfETqYsICEIMfz3EFVJgflZ1O4GfnokXd
2qAPpX3AUaQTZ5oly9gFX5ruP4/R9oJGl074iH4Dbp2G5zNzs2/ZiJdoHkfKP0nMtrYJZ99+x/2t
iFlGRznmDuvIjFsZEvk63G4HW37u+P+QIaInbE0Kx7wXbETt5ElXdNYNTpU8qkogWVJgLxE7lmWI
SD2Ir+RQRxUD4vaE9x2hbdPxaFYaVxopsE6f3Gz7c1o9Sc3DGjGxfSDt5D11c1F4ElU9alUCwYFt
JQMh56VrhJqT2xdGTY0XtJM0TBtsaDryzUY5GQ9sq3L/XhKVHo95dEiVpMtW3tvg/pba4iCP2p+7
DIK16/cGC50RWlc9MZZlccYu1wy2PDpNCxYBd49Eoj/qI8pZAL7xY7eQw9+PGbYS9sK9WpFZ1Kqo
Ca4y1MLnhiY+ITFyalGjuRhJ8L10y2R39NHiWXOZ033cGZY05/sHjDDlwMoTvLGTjMllvMbccat4
RvVQim6iIteJQIuHK8R6zeIf4aigXBT8v6OuwoyR9dIG+ZLc7yHED7DIo8WjFIF2BBi5YBLVT99Z
lmHB34QkSw2e9BuMV3OL+AYjcWbqps/CtWE4d88E9x3t4cKSvSxbcrD1K0VVIe4T0Ei5K1F3+jQZ
1KptoLLaEEGl7jkYJ1bRQhPE9rnhrH8Zhd+AVF3lfliyyy1B6Us2qyFTr8ecLbc1iBqjd7qrk3hb
AVA8SOVrQ9Qu4lP+anrYTNQJn56dkNgNx/XuID8WRLKSvKSHBJ9+gLaT5MpO03TrH+rTC8g+LMVL
qHowxHd8MEnZ7PWU/oneXK/lH7+58NOJuZqXUxeSZjhl9pyItYRbbSJlC/7eW97XBVgf5/SsnBzS
cA1/GA+ycZOE1AKDmyEVZ1PupY2DexJNuc9Ks+YNRytmqTWk2Od1V1jt4wPyzhsqtDFpopYHy2AE
RwFDt395r7ZQND71Yn1MIfS5ep2h2z/jHfTgoCQaxj+g1LRiDqUessJjiELNe+E6VXmzKKAyjXhn
m6Sm9kcJjktooqrANCSCNPwvWOzad+LqiaOTXFu+tfKjsG3WCKs72sDdu3w6+ZoDnh9XmQaf6FE6
MpB6QfZOWMSViBcTZ2PTPjNYM2gyMSOSijHaQgDW2P6HIYku9loMy9Q469qCNPbnUxTYcCS/RPgx
BhK3pRddfAIg2oky6Tjw7F1J1QvPL+epjxfLz3tiQ4rCcG2X82dI8Wynt2BfDXoKF2VbPPR3W5eA
1LAPkd/PhcJXS93ra19f4TNc3cuan4l8PEEg3tJApePsTXnls7KAqdxzmEfSLBjhMpbbhtQpW9zR
Z2j3Ylqlp0O4BVwEqBDjsEEGSIGFtyNOwYHRk3AP8z9Oiw0eJB+1bvO9FPfHu2tAcKf7HVJ8cyb+
Lnurw8z0+7M/3vLh+FIHiAMj36RZ+A44PGqe3yKRnN9mGkTnF28he39pZOkq+plqbkB47yhSbZsu
m6nxwCCOclj5InqvBVXJufnVTWVuZLxdKeE4L+3zc8gT0x+wr8rm+CCSbBxBUI7ItKl5EY4ybHMb
A5Dc1dFqRnJhDcug2lAVjWDGJwmv13GZJ2uNz6rtGrpvt1wTAgvxKbcdRr/+W91imYAW9XTtBNMu
gQAcA45NOBDgIebyr5QSO5+7PmhWt7VCx8UNv2/BMOXJ+OyAQrVOhqTXf85SWZDkgc1fCkubaeRy
bbe30lmFjEsK3TlhuUjHL+8Z2uiDlLeEwU9H3motukToZ1PacK863cYK2aUAtn92PgJYwcNzErOo
Gp2ZodXh6QyKU6s3haiukTC8gLW9tYxW5Jbngps2TWqHTr0Nn6D35qbsuNspT+NEShjHE3Ssgeo/
xFDTk8o6YbjCuBekPJ3wgUH/wERUOAxz8KPfdM84k899Jb49eT1tfq4GVp/PYJ9fdWCwzOEiA1+H
CbW3vwNnrnwjsO8QSLGXmCJXCrowQyO8q7nAkzwk1arclluf8sC/0zlk6gFXGvJm6WqiTNfJ7eSW
iNmMry8wivL/VvIM/jbpg4feBbsEWA0eHhzret545yJKSRbx4qUc/jVlH5VMyw5Oyvz06ugT7tkO
TPHCJ4GUgrBUciVfCCfLyBK1wGLPY5t5GSaLFYGyIEC4TLExZKmzS/xVNW9fBT08Wlm10tL8NQqM
+iGYEIpPXXUegb1oct15ylXz5rz4MLCLhDzNXXDaEaJ/o16RFz0vGUTZkjl7+sIzGq/o85+tEgvQ
F2NsQsxy6Q5nimHufDAe8dQYECS7EXugxfhMBe1GbUzDK93M8t61iqv/N+37VUES9DCNATEUSN4/
Tak3qGHiKKELAAdieC41DefkqDKaKfgMlDGxJze4x2x5dtmWDR33Vq8amFWbWaKO627pt7powuvi
lu/jzNoHCx/wyKn3WBEumU0xl1dvDB4pOZY7SOEcb6kdNVcCSCfl4y4zhVX1C2EhHsyxexpFC4DA
G2IH5mngtD8jptSsP1b0SLAGXdUocKsSGQ3sWgt1ncF8YpXMelJrycy97ekZEscZNCvxujyDlh7F
zlw0pvijgEdobmsDjfN/Vm+cI+Sttehob+y1XRBPoJZOkaXG1TQDnHSoAL4vAV36CxtUGy8KQO2X
NnZWI+mHK6kgVZ5n7dXYrRlqfhachWhijVXLdg+yfGltRf9cyo6JPdWmWvihrU1zeRgn2pZ4NZlj
jGh/Y8WLVTR6/lZoREISp3PAMSQz/QH1PnBda9JwWwe7Dm39nsxz/CiflTqZK4Jxo6Jcp/xX4Qgb
OF3zMWtuTcTtugLD38TaRYI3xbAiZksUeP+EB0WJKmdn9fpGkvtKKNH9kKkjW573LFzuBa8cWMe1
L8A6h6g81hhcFzmCMvrwgQh3BQm6WtG9Wq/H2k3EBha6IvpT0nP7O6wVbPPnrrGc2Llmqd0BJRC3
gdwIbFmNN1I1AS/CRevbpuOGBwUcRgCOb++UJapgElZzXDKH4gO8TwTO6XIK/Z96gWzTE1wgr6Li
71Or7+oAiwsfGIM+AfK/Uo7UoQWk6ItyenTnai5IgzbsRpbh+LiPtBSfArHkbxTeAVc7QWGKMij1
veIcXY+zPAwbVzVhydeA9801wxEV2egvSnYmngk8MQgdSfPwOadkWNRFImwOtnMk1Uy1mWndx+hf
eVAJV+SaCE67jX3/9WVM73UygR2bsvAwbqv8G6rQS88/pdTISaZQBRMZ1KXGPco6wNu7zHwZMk1y
6jHr9ngpZs/2sNPKUWLOzVpzYU48pYTCImzzGJAswVeJGdCUxvclFYi/njjZeVu7bhvw3sO7Body
q4SxrvZyFyzLx0RbZ4IMH3/JLuJGWT5Os4EUSahluBOZioSEl0xvVw9ra/sSwdb0ZonCofFfkjxK
APEXZ0ZKAQ3IlFcjfWnA7JZ5U8t3B15rxJpfeUW9VugEm9/GELmNWs6EszoM0OEWsyNEb5SFanpz
oZkeEn6tEDhIg5rc7yq8Qv6Tok/MvHORIQxKKlFjZ/EY8zskKip/mosW57+Wlo9f/0E3auxKduiG
mLm/hpPlsixiAHVYg2J4UQ9TVBLts2E4gKVerJebcoC7dA+2R8Bwufuzq8XCgaGNvWesgZefBMJQ
SM8/LR1YZEQ6fy72bzpyW0xeHDTjewQhLX3kzY27bs033GYNuoIx+f8B++OFjP7fVTGjuDfzIr3Z
P5EM1C6EeWabcUJXdL/5XPMRBONKB5kdzVVM5fQNb5gY/uIcYNM/OidDU33L3WpRPI5iYxsxkOpq
kGz8+84ITUau0XfrUOofEyGKMa0xIlYFmjZHDf8u7VMmqv5Qg9Paz7FeIs7P/MvvZoqfTrwpiHBx
CGsr3asJg75Ej+pDtiCUjnUUvmypmamjujYhcD88SG6WZRdTS3GK0OvEYSeM10fQvSmx/+Nlbgjx
maBBbe53jFXIA+zvyVYWbJJWM6T/kUUCePQ1/mEnsAte0Y/kMS6WoUqaJR9txrhYOHzUUYQhWeuz
BREnQxlUfrNxsWef5LKC1FQfu/d3UL133Xt60m9ao3c973W1HVIY8pDeKY5O7y+TSkoeoKmXIhXg
UmcWOqBBJ42OB+LCW3Y2ox2+4l73pc2gpPbwXbhePAdfifQivXBnsbaTOKTlHR8mIMj0mUhOsY/N
XQs9tD11Jh9EvTCHshGhjt15o8weCbjgfCUWzLpZ6VrdbjUi5dePvbUSGNyaPDAqFpkv6XvCRn9f
Waj87pmdOY19HQ2SNaglB37BBmOzqKcaYGETJPn3yisrIa0QJlJmoK/mikHjWRZpLAK26neCapX2
0LbmGt2+bVppVAR1ck/VmifRhm16Mf3LGUS3zpwAs4dLffPriODZsfBg5+8lB3m0gbg2VpdZM9Xq
bTbHsfnvs5fwIaov3N7n6NLWS1tnYpUTC+gCDeNRx1ZVz2xIn6YL5hvbwuadfM75NmjsLwGxU3Q0
t7z8gYt2BAR4puX5yWpqTZs1Qy2fZAnkcMxrS+60U3mPfRVWO/vEucBJ4a7lNFdfxPNkMfZh568S
M91uKQ+42pldFYF6VumGfg/xqcfaJ6diqDjT2CsznaB/N4oHsY2p7ypLTTVQfAJTCV3bZt9/9fkk
K265ST71iuFCRziGy40M1+EoIj2F844TsS18wH5woCZuO445wH3r3M48nvjA6QGroHbaXD79T45T
uyYmWXXd+7BX0BW/Og4p1SGVijAk+VZc9+e/H4sA/O1MQWfIFbS0ZXiXU9R8ZZfVF0cS05ZSrIy4
Ag75GBeHCAcHkevfM7mF4u2gISQDcyuIaUO51opI9tq1waFRlnPM4nRCuyIvLVf66Ez3UFOgIDJJ
pDNmjSFA6KnrPu2KBAfnUPtTXOwHPk/ZM5Lkj1n8gHkQst/pyi1Bku7rZpKMLneBDJOvN35xHqMJ
NEAJGvQsX/GQ+ibRThyLN7t7x1iSGizGMjUVthrttzXCGpdHx504yewpHWdSLb+9PacrQmsLXb1B
v7voGLJBV+tuqP9vOzPPyilBkIXIDXWdzdK00TY9SRHkbTUQdki1YjTMjuBUFXVdlTWBPVIEYIXw
BwDP57KOS8wFhvQP7tDluiL1CqdiYgszFGXnmwBOR5jxl7AtLjTNwV/pmdxrAiCicYnB6naARwZ7
bRz5b3ovxdJ1GITRcumFLD3YXDewAyF85biJRnfRryLrx/X/90Xu7x4tfKBXd4CKKcO8tXii1G6l
k94bf5v09K8g1A6MyeGqs0+c75UaYzBVZiqybpaYqcbCcZKzHsVHG8Mju0qAuxiZPj+T2obobmwK
q2wDoIPvdqp5qV9ctp/yGEfZVaBRO0oggLLPMNijodrZb6ArGJoH5w1qjV5d36ZUU4vwOS8ToFqb
GnpOjhxj55BaROUf+KyDT9vxIem0BeTiD9UemIWDchGhDedRCrgJcTrJyHcW2YbGuK+c98gmCIYe
+T3EjQjDrBGipKuEu8MYEjOihrc8yw/wSFu2cj6nV8+Bm12eyuhcJcRXHEOWgHyIrqFgrOcBgaVS
iymH9qGZIfPPP/TNNiVFP3cst/erw3IuPi32Y37wm7TbifQzh3sWzRJoaH9H5LVGXAwtWscQW6XY
x03sQfebY0dDUhVC/vuf62s9zylYnCzxEfsOG5DaJCaI1F0r4DLkotbPshfabVOy4z5dxxWkblDG
v2Lx7eI4obeh+V/DUFWzxXna2a112z33VlOGVTEDrkMEloGXtQlOsVYHCnmSSlK4w/Kt8edyBSDo
j3Yx1rvdle71+3N+2o2z7fV9ppTw01uQhqwoHyeQlTuxVKEqqIHp3Pfspe8ZPWP3ZQt/QMxRH6ga
uCe5SkGRmOFvLMQoHsqwDic4gdQXUnLuNPOxPu/AV0cuINmI/vnJlP3x+N39FDcggFDtJqp4VG+8
zAzTVwm792VFY5Zpe474mWYXvA6MnfzFl4C7OJgtvegEpICBrBi9CZYVS0ANiPnyv76mwg88OmOS
5P0iJ4o59qj//xt7sC0B5vWv+NlP4Uk9ce1b95MLVyvx4cyWmsrjOpUfXgbqRm0/XsdLn9hRxTPG
3jTSYQuAHlgjw/wN0TiofzZznNhOMZkPL2O7tXyhOHHVe+eGGudhFlbDgxinBCRShRmn+Khqtch/
RWRC8mN0UU1ZBoRcVd186M7VbW7rKsVSKjX9nCO0jXYT69GgWwb1K4hnCbqMDz38I6IUFcRItKmM
imFUNashkSOuLQwtq+8TJ3bIJDe4UNFEsXOo2n0kqMEjvdWSVbtQamFinTuilVBErm3XBBXN9keE
ZEhYg/nYNV76haAqb5gHzElM02Y+FXHuaDuGoPKOmnq6ajYDqPSxqew6G/haj7rCN2STun8x3kA1
v7k3IlB0ocgfNc+mQXtOcU1IYydVV6AhXLz1/lEfHjQTEtOZyUBSlcmF15pZwIlaKBlVkgjlcXtM
2Km9YQVWgHZsNFN4NchNexoWWAuf6Z0s+qyjSAvn2rGSExlTi6mRGkoNvch3CmmwPVl7udtgQr0I
Lbaxv1B+VtD6aeYGjK+eqjZ6W18ZMgM4RzomchvcwsZRnH5jm71CjBZ1TKbEsgxt946sgSWNn9mq
FTmQSDxi0/LpltUm0hx7GN+a1Vqxhx4JX9WQC4zIwT7hYt5ig2SoUU9RDfPpVBP4N3ZtRZnq59Q3
HjonUad23WLaUUua+v/mNzhGDKWWbw7JSsxUTJuOBz17E58gidyxtrjH9zNWuqCn5O0Y17r2jhz5
4i7OwTWE/FhIKoc3VQKHegLL+COPdXFWE5yS15Ok0s4csSbetKSQw+jeZ4JL8JuPtDjjPTkDim1l
g7V109Qc3B/PLFFAxa3xNhvTBIoH5+VHmaSUgd6roTfCKp3Lj5ZDFI8zU2Dt0/sT+roNPnOs9GMM
GiYF/dOj7qyV9c5jq/2GEtzE1kU+CWMEGtxi8cEvxuUz0pXGtBfCpAeQnR/id7YAh3m9upfAdYYt
fkUmRVhF0VLFB4bOj60AAVnc1P0SxvnJVyXl78xVCQeOgCC23NIfzaLrx3OV1XQ62uu9ilgqbeei
aanaxqo7ZF0uF9/adi8QdR+tzTF8e2fFkbE8JInMT4eDPXvLtchxQGd+1gw94fF8ZmP4TjLwzkks
zcyPtsDb0jGmQWxr1d/I7vugLWJIeBqLzebjS8/NtnFwc03v/ByaCZjMTb5n6kuWTQPMIYTx+K7i
uFB8sgBHvLeFOpY0B8/G5/6hpTkf3VUtDt18Mqxpews1QAJYQ4CCFKr00yYt4PcYUZTumPe/Fzbe
+1D9tbR5i/bE6gypJeYdbqSjYlEhj0BwuBo1b/yFQzVbbNnwnjThN2JB0uk5BFE+yxbvx1naGXOJ
vJltWqt1413FnnEP+Phn2t+KlAQ1z3FNBbhzvTjCQAXXcNGr2/t2LgTxjwC2EqW+0/smLS6Ku4uJ
rY6/lukZC1mGE85rP59R5RaKrFlMl6jhD0MMtOwNCsN0/XBnouuevUwJekyvpIADCMyUcMrcBiKm
2jafIf9pYOZKBqjaOfJy7NuJc8ZCnR8AfE2y9OwyRn7fbrhFjv6cCrW2yDLQcdEUFOM+baCwXdte
H6a/3hbfrW1YhVTyv8LVnzw4of1mz7myMRqqYyXO0BO/Yhwv2IqJKWN0NxUXO/IPypylMkEEKmq2
AvDidqm9HxWMXeU2Dobo+GUobr0uKHLTHbWzGwi83Xvl7OBgdzSUwFNY2ffbum5WBnZtjQ2wfiSj
vquQ1nTJnkcxauMS4plo/VmF3a2iWxdro3NnMLskIb6OCxj3xfjrnKw1MmHpYZVoxvTIEfsg5m/8
mNY24io9v/hRwMTLsKG/Za9ls8LEbsECxNwCy/OrvUJYbSo9kMt60TiD2n3PiW+qkpjWcju+A1nI
Kx+lrFZEVHb4dWnUl37CPDsleREJoADQokRaFTlyexiYfRoQWwRGNTEjJbrE1xnFV6QdDhOpIcEN
8LaNQYOMjO69ugoFs6ywv1qcoSRJT4SebaYMLzemSNSVg7IofrP5mt32Em30N2L+rNv8DjA3XxO6
nE5avk4rh57jBgbA/pXYV1wjJccfC2rdJ2vQTMQJ8yS6oa4Cv/CKSFjQpGWVGx2BgJm7+0ZQ1YhF
S/llb4xEuvEvIEiBoyaLV9eoHQpvzNuRGm1lVdIuMHIBB6n/5H8Yb/TcpN6YigZoDxoJgmdftDuU
HihqEMz5BCTtO3X73Tn/LIpFFwH9bwjKDtHDLjfA9zAawE1t98nTP3dPkxJsBxE/S1e41p3srVH6
YD17VTWfhC+5lWIzkmrWPpuGIA00gYwbnfQ4f7DpPsTNDlhoExpaKHDtNrqW9WEQlPviKMcEZ+U3
mNyL5QGNxlbeFbV+q0nAoEOzY+b8z6uR5D9p2yzr+vSeaE0BDZMNX//egSED3IJaPw0R8dTXNC+H
vHCxPbUWAt8YSj8d1/NttqJTS6e8+FbgvpgaZNH1S9jBPPBcrqUu59DXDA0xV/hIFQfAcMqZL3dU
MZx+P8/N2yVYaLm0YkR6pnRSfHmjy/H9CwQV/DBmeY6oX+JF+PjIIcceT6DAcBZuAGiqX7E/mUe2
tL1p8r7UDk4raufNdkz4MryspX547tqSaJg7YbTSQAkE7F5yhVAviKzzmoDwLYucMNMWNjyjHzme
3sn3BsHEgZC/b/N/PqFphZkogxxbQuriDL/teQkWlJ4qB5RXwePl608EfmpUUVnJJa8OcnwB6Ii6
I0qV7gHR8UxSo+81Afyf1/tmncyNBlho06w37Z/9x69739i9rqqPyziq4Kx03sjjJBSRYaWkdHIa
ZrNLxH5GpLkcFly7Y44ZN7Zq/Km62NCsjKlwqIOHpRbRYaJGkHFzRuyCJH+FFdbPKPGAyqzU1qMZ
UsOWsdJ/q55rvm6V4wo+QvnsOwiVQB3/O/xTuwxCMYiarPzyQSpIv3GZoJ5B4Zt3es0T5UAu/SvM
SPP3W3gSv0m5a3A9k/lQ2ycKfDhZOrhlrakalDoYQmomYYGAPB5c/pJI2eQj1dqObpKqHxrPVFlH
gKC9onm6ffWEHTJa/VOVW7vspjNr2E/5RDKIKpaZkq8vJnB4CVxcISQwfEdAxisdkbeumOtAgNdj
oDduicWjPoU8+nCGNU21DtTksp7uHVwcROc+53oJrcnG4pvuj9HSpK3b/5CS6MdRy2rvPMy/rKFe
OTCUT/9HSHZBmXIjO77Xv8bG+NoGjXcTJeqgHnqBFGSuYyqIFYoks83q33ive9rgp+ec1E8BYsiA
yKcFmLJzl9I7KVD3AoQoywOy8Uo/jrBuwCYujHOlEAU8B4KEYhGyrMAcoGKM8zqD63BS9Kq5h/72
RJCGTIxHLOhik9fkDxYvUrfhy/rYalDb1HbefUDqu/sWP/IZm7lYKlwiTcuhd2c4UiP5bs2iZmOQ
CcGYgSFbSwrIEBfJ/2Jy21SR1VPYweoaPTnfeSA1pFnWPmEP4ZdXONpHWaZw1KJWBeMk/CK5S2Y9
sAHnrUCDVyRbff2QGG6FBg+dNPBllhbUW6WPHIdkPmYjB1XZkpmQ3s2JAJ9LE/6NFP8Ng4L686MU
ptBOhfo71fRQmTDR9DWF5v623+6Gua/Rf9BHR2AiC17Xj+jq2/IrbkwLaHCJjw/ELUFBLgXysfpY
Fvo2+PAJNYtLYhGraCzFFi26Kh6lv2wSBztqV33D96cFnNbism7kFCThCW/wE0HF7/XGA0bLRJkS
PJQ5JXlzktnQ4rNke3hmH/Etm9ZVfDoATR/cUvts0hKRMh1VyQPpMryIPxD3ny4FbB5X/NHZaIcG
28dpkumqF65X7W6Uwrf8a20NO151Ei929vB2cCAhZL7MmwdG3MUL4pERpr6dwj8Po2fDQqMixtJC
zY1yA6posOQKYXd+NlYVWVTOf0u9Zuerp+3HHUJfWurkfZ9cHZ3opii+3aEhbP9f2Mlo3xTW019H
cVX/mJK170ulYBzN+5d47SYIupJz/3dMBpgPiqYLM1NPCEhIfFpETNj7olpKOgZRj2lqxmH1JQT8
KLlrQ/vCdmTGDv8B7mu8KAMlOS2i9ZtPnJms97buXiPdE/+iPKdklOx/7OZ/zscKeYMDqjcX2IO+
YZJbk02ZgVmEc+vtGODJFHwFu9wmsuuh1UVEzt+Msm94DsytRhFdalLBYP6gtzmi+keYClJCG5F8
ijg8EZ0uBOyejfEkBNeaHru4nXnBBvtURSfo1q0NZYp4+fh9DuZFwjPbSWdzc6CfPHLmFGvUHxIH
NZ9Jstve5G20fMzmnIa5vsyJtLMbC+mxjaD8JjtZ8XGmC2jWJABhy3kJrUmxj8EpfiO3OLmSqjF2
07EVac7vrp2bIdb1TUYUbzToacoGzNyVNMmw56+n7pvYfKyCSt3XgG+aV6dyECSOezx+pi/NsQHU
DkG4dqLFMk+cXk5phN7lLzRICtErFIYI85/RtuDNk4Zzt0VvI8s1lx64wvSuR/B2PZzrf+r3xqMw
AdokQ2wquGfFHVM9j5kZqfR0oaEF+ykjQdt1Tb45qegGMMZG1HHEpRBPlPgZlfHvwJkwSw6K7k/m
ET4rUbQFtyars0vpdS183Clyfc5+mBzvm+GeQwIZDd2Ww1x8QHU1xaSRQ4BNZdb035Awi1L3RgXs
McNEKEXHQWaiXn1YQ4hbi3K5roUTEjk6SS9Fvb+H5Tihsa8oaS/VyDlEg/ZjzV2kQf582OLfooRp
pADNzIIde6KOyEiG9mHYg2CDo+8Y+4ElbqYVuAGgkPGIlv6BqlNn7twbkRlr7KxhwT0tWO2Uq1rA
WMGJd0dzxefGP6a4snH2kuVISx2aKgi2cUzfomnUuI6HE/VA58k/wZdjnLaLhLFGlRyBvd+Bc3it
WJy9L5k43oS1PJlJL/G1/4yWkOsXGGoB591IbWiPZTqLq2QxfCpTnF8DPzW2nBgPg2vc7GRFSTVQ
PIQGsypr1AOSO+C7b4W1VdaiWCkknc3/zmlbAmPfQWDbX0kcl0aJz/TdrXaiDenPzlbnhedrRF3j
594eaXXINBnF2kAM1vbMBLE9taHGs27wR+HtjoDXixrTp3CFB57aGQRs/+ZcrI88MBK6YrepHMIv
g5OFAptxrIDDPTyCaJD93t1RNMH3/cUYgaRyB7NdL44ihqzPgmtlByeNLaGswhBbdY4jKde2167j
gmyGMVhzhwrQexKLpCx4vVGS4WH1fONd0DYIzzvKmCn+ockh0y8NtiDey3vTsn1QxnAu+UUJmeNK
vWiggHMShiDW1fj9FBTZHbEsoZ+gW/Nyo3BS5bzP5IzWg6pzs8+VqRNQArfrbelz/JU1h3C1WNIA
JuRCiAJFnCuaN48b2XPAE1rjg61S9pYJU41ibAai3jYl9ciQyInzzaRNp/iWAfkwzUsbBfSRPAQT
dUg3AAD3sCx1e94cqZKGo2pftMJ+BCiQkXxlqQpcNNOXrG6CAO4Yp1kOdhyPZ5QWI/lQmYYfHffV
ShnI/Bz9VzyzkiU7IwGhzmoH3tTbJypdq4UUYJm06GiEhN6nldxf1Ifq4+nzxCQrgLgK/QPHlYzd
ZVBfvrj7ztJc/TQ3ItzG7ioTk5RGyyma+woHV1jRbrz4s4t13EwgRKikvCtpCw8qrTntEOW90JaG
TyoYWHnhUCOb56YMROCW5mvnEMng1/kRIwsyVlYsjcm9GcavWl4NgcVJRtnWJ/TdRVr0CT2ukOZO
QRnSZBlvRNQMxjHCImQctgpheluMLlGudTXSjpMg3QyJTKxZjgrwIhQbX/P1q58C2TC1UjeoE4kX
heDqbZGIs0f5jCkyYy3FcheTx0stJL2y79QhHgcHhm0xJxS6HrSrZUPpJT6pbaxSDfpdwxW4K8J1
Vvy3slO/psUnlogASHbw74CmbI2KLUS0L1ZUcaxbGHwKeYVZz6IjDbw94CzhIgeb55tc60eirIWG
Zpgamv1gYqxUDaFlUawRM+lvbSBlqYmulXwfgZECjkiNFB0cWSuJDWe5nO4s44DD1GtNFpV1clVC
7DH2hafiQhzjotA8JLWOBJ+ambEHcyrtdcXqvBl/zV1fu6jZEexXuPn/IHbBFFCKQqoFV2oOaE76
zRK1N/nSA3Kscpe9YihhY4FPPrTvzXrcRP87pGWV0iTRo05llgPOEK6YKeaPBZHqOrQu6U8Xb1Tc
U9m7h8FaLzmpqMN0m0ELHriGLvOGGh2t0uEUE/5WGSvlhWWAYFhX7GgnbhzBxIE22y8BaWMfvbGc
JNrJCizegPzMxEuDKXopEDPlMw8z9c8ecQTu/Vng3Dowf9LVLtWwtqhGMX82FFQNE1oxYCsEoFq8
219VYAh6XNNSvVLdog18RlHPitZx8yYKM+j4gAOoacOtoYGslkNUcSMqWQACbNaDrCoa7WC9P+ZJ
HqBoTOSlUb2/o0131Jumt3+Fe3aYoXFHOm7YsuXHa7N9ZNQlckPpkyFgQ07GmkFaPIumfRsvaX0l
Tw/pATn2zlvIAbtqWLNAKZ+R6ATg4zkG/Htq3cMmAs5WC8eEUjE5SASUM4ivq5wftUkupCXUwn92
Mr5EM5T2WzukyaXxphr3bPRsK7NQP0dL9FacwJKdvMFvAyilXK2qwiI/j8HOpDR+WeDvhUiHJufA
5asvLP453t6x2FbHNJShNYtQdhLIjtpjTQ2TVdZwsSqDxmba72+lAZGB8rF1IQv4Jfjcg4HaPs+h
Lx8oMClKjdRWxI6eYGgijs3fJM/x3cpJpNiD8SVjs+QZ2S+sS8KDqc/H/foCaczN/J4kvW7mcn0g
Z8CZyBzcYKKnFEyXWAjNIiZxZ7thfRaRfIXswU7QfRuNT+O6P+8akS7Suw31K7xw+UMWg30f29t+
XpKgEJFyXqsNKYir3PdTQWGsqlG2U4cibRM2lVPvlx5iC1WgDI3S2ndvgFGIT4YXK3P+iynWW3Wy
RlVAHlQyMGWwRFE2D75OcNGYhuyx6faYdHdKa1vas9NUBBVOH7OYQI7/PJUzKpAa5uLdjFf9TuZZ
8BSdPcHEjMzhDxRTCUCRlRxUXYD422n48qIMJfAj8y8VH11MGJQX09RGA5f8orG2iAYBQAgfr9Yu
Rzf98kcnEDFv+ScG5jVsQ9ygY5d39qesCNUt2pkzZI+WK7+vf8CGmUjL62elJTaLS1y3mcMzYzlF
6HdMjEU/UkG+op1NzbJOOhQYCYMRBwomELtoA9wVPHg4je2tjkqvNVbGDR8PHL9WTEeVlthSyrGG
1AyhfU0Ddi9qD+fuNppOAVqH+TgwuY2JrdjIy3KWLFqr3L8dq1mA0x4fO0PIUxv8ECYj3AINgBvR
k3B1b0m/XsAdG8KtwflJcBwPWMiWj50bQFwcwYOqpyqAhrKLssj0WRyCpjFhIDAyBW+nAfoxVTQI
624VF42idd6SnCxVeBAzQBE0x8b7sqV7kXFzxWI1CapH+CVP0W8cWE7khCVr1Fokh+97cWyq8Mui
j3ooloOPmBCYmAle2s0Cp2lH+E5UQtAWIh7qf1pf94O/y0X73UOC3IK02x+4pxONIztA7o50FcCU
OfIfLxSGEhvrBYDMlKemXEIdEx94SZjlxUM4FEyzNQerMFSGDjEo9teqCj5TuybFijsSYqklY+Lc
xd7oCqCHqNKKu6EcSJ3GDSQ+M0ZFSedRHpht7UYORQQfllUUoD8Ykd9LWqhV0/eTrPwrE7Osnygk
uwX+fal46+Ln80r8HWSQDpbrF2hQk4JZGHapJvbV+YPtfgbQPCW4Ojn9mtVNNMnabZSBMvwntlQE
nCdQbRyZxqPUBThm5IcyPcvC/cO8Y7uBuGJUHBDX/eWx6tAq6EEHVetXIuGrvFVbjbutOT58kt9u
GklOErofixgRoR88NrOwOeqIyqbezxjAgN3LmNZUUhOI3EZEgWE0ygNhU7uyZljWV5uCzyNFbEde
Ba1uMZ+4rKXL+XBI7HK5MlsvgdIcEk6u+fg6uYbcfV5NsflsndKQNZuz2VX5uu96409hXz6N5dGN
BpI387Y/UAg9ooUHuWu9jSeeZxvPejmyG5T54fbpdHegm/voB145ZcQBlK6pbXRZHl0ZNUsEWhgc
7A+KnFeMrzWMeKjcWocqYoCp3acweGgq2i7+I74+bdwLuYLA+RWUNEQveo762RliJMTjLuKQOVYo
66pZy0sx8AwfgdYI8WEC6aeqF/XdvNM5mfgOBWbgl11Eb9TndmPqexI74qf5GoCBXr17OHJIFuVM
DsnWrKt/xwRqucT77eggF2Z4RNL6LmeqY3sdSLsm62ucvd9RHOGMIdfW4YdISin5iqGSrFVe1mcZ
OP7ceplwLoaNLSbnbaMRzHICk9PK9fjgCzsOp9uc7+3QzrC+x0rq9bUqQW6Wy+PA05svh/lujKME
uS8zl1DAtut1Bo9wk6+zlCsO2K4W/xZEnY3pl0WdDLxB4tHEnalziNPOvpR+enj+/oan+/h29MLS
L/zktBpPWRCgXowqR/9SMh+XYsnIaZI+NWAF7aevYmYjYc1sqNMlV4EOY+ZK+6Lk1R3vN86j7Ctu
tnDoHmOeVhHZoCaq45K4MAqCeenvoq2fLtaid8XHzDIFa7YlfGY/5B+JecInf8yUguyAm+9291YC
OstFonulgiiYThq8XmUTBQwXOyutLj/QdeJktEPPgP0U0YGx+SosVDVzE+ZRuAKr+K6XZapHgtqK
b8KxBgNdgtgmJnKkXgn1dZq2yqE3VBgQzz5luQl9whbZHTttZA4KKr8ffkTX+O1YGtG7EDRG8QMb
riPQ8CK3EAww6a9jduw7OIcVLgq3XRpQNESHY198bDVXd/rUpt0T88yn5EbCmLOOR1p/wk96ds3j
wKj4LNuiLxj/ejHbte3Idwbra7H0ANj1xmsqHdKiRTrfa1zbsIN0GFWfHIW/DbLr4ztcGPNiXsUv
yYgi/cecR2VO8niI9ouKsEbba31Z6A2QhOfEfZOuMWcQ12sHEk+U9y9NhmuqepHNcgKY6bSyp/rh
yF0/FIICghyk2KeWydoSss1CFepRNcyiKQ4ZUprZulT86zGPBM6qtzPZ/WocmFW4DavPK0NXa2U7
DVWnhcnLrdjvrbgtsb9kdvGCg43o17lsN2ubxQQs7WvH7j+WTTRqxjZiF/FbE3NLL+81GgsmjkDM
aoVnh2ysQ3O7Me7Ff1XhEeD5Z24/zZaZ/6Ghr3PqumJbqP+Jw5SV8FbglkXOUbUFCYuTqobAnZse
O/dk079d25AkPdIw0Wq+yeMYFtAMXYNM99uvNoOOPCvHAJ184YYyfr1MpFAR6Oe9kZs2BEik0uKA
vA4/Y11LlMWkK6VFSC+ZLP1E6+dj8sQ2+AcrgvLvYw+yPY0ExT4Pfta1l97Rs+mfWgCcDzeTvsuf
hfeIRRGcoFUBgnSSqvApf77AprGowobFBw//PUF3vIolPGcDEXJ1XyGWppaV2HqpkF/HRE8IIb5O
/33iXOFKsZdrddgf/tYF1AvVmV3ncqNufQilRkAnFP+tOxSrzeSLIh1fsy88YAn7Le+4ArJhc0N2
u1Fg1xsx9wbUJ47e0Ry8y5AFNEAHp0omA+F0sr7SMu6LwhG/d+IP/MNTNuzx9TfY8EXSrU4fPzLw
e1/1LlvJtd6ZeTjq3hM0J8jEssDjwFVyxlkXqxJbGS0PCC2VTUQc8g9vcJ53VJK10ZZIcJxFq0xp
rkgNj5qIJ68fDxKIj26nXMbF7LHSK+/zNWyhkAtYoE9W0/fz7wLc5wCjIQfGD976O+Pn1rLHlDfp
9e9xLGCyKuKlizdXs6T5Mmy5jhQZWIKi8wbcxNMR/2YflipuCNmlbb68nYLlBeqtlSHhmXQ6lj14
FE3tUI0D5vMlCu7whzQ6650SUpTpO8w2fXNC79sHLG3QhnCvjNaiPUUHmx+tITiWytoiKtG4jw4Z
2268LqPbLzr1VdCgIi1J3SHu6Lgauo3B5BgekBW/Cs9JQUz7HoOzoPckkDG0bbt6W8nKwmsaR+sa
NzRdjqVfFNtBonoFUSK68GrmfstwIq1w9FWIugGJ2OAPJYiyOpGIl/ovRXDYiRuVOoEa5stP+Au7
3MHllI0GR/LqgPDT/DrGiLfRvj+oymrL9A6Q/6rIbFEVTzu1IsDxF4QkyDWmBDKvvJgG2FZQiS4A
TlNFoAkqY8JIhgDKXz5ucMB7Ta/c2wc4vTyJjk8boAFLH8u+V3OlYBqKpOl/sbmQG4HPxYfT/NV7
08uiykgl1fU2FqtiDYjA6GPHfYY1UxkGST6XhoQTzvEcO9+cyhuwJKAr46rFmedWwDDyUtZeniz5
g6dY7n0ca6FkYnpq3LEfmzixijZjVjdU6euyFPOebO+tyDvP9ZJgfm7AnBoOjABtJpqpq16YATdd
bwxmdKM2W1lBuB7jKnMV0wVGYmTNA67SnvhKDloAa1cQ5eYv2KGBIoCt6MkkbYBkGAhhIM0NGZ1i
RqYhAuNbs+kjI/+6k5rp30elpA37yQt6Xg9k+hd+9gJvrXkfFxtRkQRWpyB0ilWpgrTX+0988tTu
2m9+H53Dcztzz9frxGKZVQkZTc046oN9ox4UwlxA26nlyrx1O3VuFmdqKLTbAiDdS7fuHpqL6NLW
ZOMLx9EOxIAq8PGaQl8ynzF+Ucx9pOfgQZUHoU7lLabrUR0oh9B+kcWdU3oDx17xs/38RRh2z9LT
a8FjbhwAd/SGFnLv1odrk/jt5SxAQLz1b8OnM8DK0LMAK56KTKQQWp3DBhSqeMDDOGYyhBMU+as+
zKCbHxE+D/5WsORZ+f+xoggebtjiIlUogb3OatdmK+Lo9xWxVQzHrJZFKgid4mSGsW5xQ+/YAUdi
7mcZGVmfikYuoQozXSa+okt9fbKMp0tZj3ay6DugmMQrloTWchMV6gMGmrB5xyNb9FvqzJqp45AI
yfCr0Z287mNPiDIb1oNxehB4impERQ1VLRZxC/PgbKUsL6ipT5jWaZnyKzReeu2KI46OMnXbaO4N
AN0490393plqXfgxUI9lhbJredoONFTp/0muaTOKVL9iVjKVuRaDaA9fasiuuTDRt1lkaM4O2E0J
JLoKXrgvDX6eaRmolnxIsJ0htSPtQ8auQ1QpibKzmM0ZhKjZT7wfY9Evbk5jrrdqyNNtE16OSBCc
paSQXumDYDCA50l3StepQa8j6ptxmU3IBXOws0N/yMVYVT2C9qVs9PYUq5nYT95ny8S++tAvHaLf
p3KgEkH/4BNcrS6G5TxzQmjTZCDG5yYH34imwYFNS6wc9SRZ+iDxp61pd3Rp1uIN7bZ2mFaiF8Gu
AWMh5RR2PTkx75NSH9TBUY44W2YgFHoiYgX16VIUKB+gnYmeAjr/e9Y19Lx6Vso96X3PdxY1CBOi
m1J0fHyTiV4XoRyaqRNz3QKQUbCPw97CqDIoyNL/SpIauhcjqnw4staybjSwX2sSYFk2Y2dp0xXF
yjdVRd5RF4NfQ+TbxfcQgj2Znq66sZVdYePtFraPXq/UwoXKzj4LHy63S+i2TAObnbDXWSADVRL8
3e4z+mBbhEK27/d1hPFduPIZWXWpa/BWHGu9z/7K5GkGnVaFaoOkhIBVFeP8DgiwUy67bYHo66o/
5Xzb5okey8u+KeunhqZsfzsv7cfMpsUMT4RuzIys4b6qX6R+XspP1HZpZ9KFI3Te0AVRTtbqkx5U
8WLcjNGPZAJr514qrSV6G7ZsuWx4LhAzbW+XswQHc1v009OtqmRPvBIsgB/ze9HNs+hodLbmCsqk
tHvZRr+IHJVQ0IcxXiO7If08mLP9IdIs0kXNLFIycoSStRYH9VBfHiePerv2Yw9kKzxbTpL50CN0
TzWkoyKlgVNAeR6LzC2Uj2IEamB545tD3XaBZ//885wjdxK3T/A7RRyT+8sGIpXV8+Zu4XEPIMSL
ErGF+IYO48bpuhl6XuuMt2N9svB0IqSp9+GSf/xYdyjSbWNIu+SwwFaw3fb2kCuWxWkRxdAIPRy8
S8y7tgphiZUyadNX0gudmE9Oh9iZbit5mxTRF3j3LBZlGKfGCCyRtwd/Gko9VOJCDCYKR48WIybX
ITB7kY0bmbJRo8pQ4xHQ4LKN3gxEWlX46ydyE6qnkgzu/uucJ0mpavk3iTB3dAoF7VzYCZGt5bGv
fXsTbK5YYEA9cnC5PKMUzuwXrwgDJuFRX1Fkzv78WQOF9ACwBfH2Q57iaXnAS5v952whraB5sClZ
+LE2NFjRn/UPCzAB+at7N0gbI2D2oeoptiGAs/AmWA3ELiD0PatpzKnT9iL8K8pc0rTWlQghkH9i
PeunnYNRmbMfFzG1xVzn3Kk3MnBvX/qzdq72IrJOleW8bQ2/RXhyvOd5w3gFhsMYqEJn3m8C+c5r
oU4vIQkklTmmNZb5Jhd4CJAl5HQ9cw+E62C9fIxGQQ+NGnzjB6Ddq5uSZbru4w284RNaXHp6naXO
lK8fpe5siApCTf6KE6f5ZiL1fHAv/AAHmWYZkRv8/RKPHObrPf6XOlxvJ+oLD5Rt8e2k9d6im88f
S1EeSeDo1jjhPF8MY9AWf+l/hf+SWyHYy4YsqjM3PKtSS8yzJSvUbldfRVounl6UApVTp3Md2j9i
Xl2urG/S3/70f3tXZuQbRypBGMcf2SH4hnl2NsA1+sId0XHnurww63pFL20dKf+004JCXHoYcNQp
JmLucVG9twW/sN6vEhuYeMWF9maE0JHaS+Lv5eSNkpJrrmxC8t6OK6ErPtbiZAo5OLpKetsZN80+
uo9wDypHfDR+aA4HkYV7S7WlKjB63+gl/2UejUXAKhimc+c6SS5H1LHeEfDGedReF4hLClJozleR
N8l30zofcAOIIGFVK1krX0u4GWmpQyaulHxRi6fbeehCZ6BLi6sinv9Ka7tv3pH5a/BCzNP23s2Z
Xt9byhsGXPaeTPqDOh3TR81cNcUw9oZ15B0wEXNA+IqV5KtQLb79Ig1K7y7/VNit+0Q7dkLpNgmr
30yjM43IINDpCDOIXVla863cqmLblm/un7ZJ3Nd9Da+tjMxoXM1neaZCSVQ/q1Vr8rUmVliQIGHC
/p+XHj4bg0f/Gcm73/lO5lhwamyyiLyu9g52oIH92Gd5e7GoMHYJa4ib4KgGtpAuJULSW/dmo6Nw
PI2RDF0UsCOgKX7k9zKiEKo1SXILVA+XZhz5ZYtb82vOGScRdPcMlRChZwF4wLhigKCwOobFHhOd
l3iqlMHAq7YKOrXS0+EtuMV7v+wXSxk6vsECV9L6+JOoJ+Qvh4W0LT6mrJXDp04EL/E/4KoByoYY
oJipvjgITaRFp3d7O/HXk3wrBGzdEliPV9HhR59S/G/kVeP8PdGtaAfnW2zqAmclVpu1V5kLQTEn
swnETyLrSfKwjiYKjA2FjTzG6RbSEmRw+OO/VXootD9bRrN/9cCsKoXjKRWBpPj/bQPoUCOZg2Re
dtevRRIj3D8161PFXwNxWbLzEU1+nrwXjHlElvpI12LAQBkWlQxhasHsI52pyq0+s9xNRFdR66rm
sUh2s+ezE4K3rmyMi2BHkSvSSlkmDufupmETiuPKmFOFMe3uzG7Ql2NmgSwz66t8nEcAEFb+d9Mr
gg5KJdjsSrjteMAVg3xl2vToBY7c9XbJDYeAZyIxB+Np9UxhRfVB/OAuB/xUOAB+biGxBhG4webS
zjU9TIZ9Eet2WAo0+9UGit3EnUghJGbhpEFWXnXkN5VHWvK7gtahx4SCdo8yNMD/kBnJUqsfd4Ph
0c5uBU228aaaUvynK7yAvTdjsG0qnq0M+HcGf9opGCXe2XEqsNvfIm1e3hJJG1dm8HasLRhsTrA2
OgJ3fXHRpAT7G2yanDRAg/OSHEDbyWaseSs7yfuZkujV3svyJ6QrVGarBX5pqNIo7Y/zEoPyPz3F
1Hq/gTscrhQITIvBypHIZ31yWByiEAyF/tnc8xTRAMx1lut3ZO+f54prFI+nqdfUnAB+jZVA/Dn6
8g5JhME1KwgC5GPNnKyLUkMWlJjwPTf1cXxb4Lt0ozrVCZaACIfxAQ96J17qBElL+DUxsp3pmXNh
dssNc9myBAmA/m06e+rwLjwMxMeMsmVhNuqjXZ2wyVKAZJvdBHhejyD95Wr76x84OU+7OAgmFWe3
Qh72FE0je9DXuN0PVbYn6plIWUMd1soH+Db4/k7+X1l2NO14JQhGGEHym8VoSnvV94c6DiYXz8lT
5jDDADawaA8CkiGRflQVpntRNFBaswy3/9KHc82zW/aPb2Qm/7STuPM7NVOeaXbt3sVOjaehbe/3
ZJ3UXu0JXx/GIq3iXFnOy3BYnEEoodelS0B5D7zvhAi+W6j9wFrf1lNkFOZ3DS/I5k2nMn7wUrco
OPRwpTKylPlSqfAtnOYWTTbv4T6FpVH7UoR+1bkfF93OqdJPwKh/khhQ+SS2/gTFn8tnSLsAfknk
B4Jx8PcihERZyq9e/s/fnDwgPtFS3VYJboGP0i84RvMRGaY3xH0qpYsgXtxPUcbZYPd4myE8IA9E
VJ+NiCXpAtDgVL7g6moDlxh6GHzwo4yHa7x+UMsYxY/2/MSElKmJLsaU6zfga7qGzmMJ8bBq4MiZ
uLJcNMld7NvtfTYIiLsUx4Z/ZRelDcHHDwe6JUwA0o96fubRghn5F4210H1z8/bKpe8LNbQEm/Cf
MSgutjo0NlTqcToZhCJ9Te7o06/ZSzsudfUwlxYUMW+VRydvF6ORcH1Z/6QgSzwisOK7neiLLqBd
nDIAPi6RZaea95OuDmDH+s0OgVvAchSoPQYlfNGxlw1WO0PSZzkxsRTy2fHkDzFRgk8nBn3Enfkc
5uP/iVbsnMHx0+5qQc5BkjmYhTJant6EQ9Erd55Elj2LFe5KBRz0Ihg9/xd+apHdE8edExriGD9Z
gmrvhai0mb4rnJA4ybeKhXxf4OOpTk395Tf8Sp4pPgi9p00DO6vg8lN7OTEKwmFj2oLT1HQVLBpZ
3ntUAHAMerxMwhmMAx/XigbpkpXNvv4rf7i/YNH7imDMGtUBqpz2edWUjZV0HKUnUGvD9MiMWWot
bUU9E4tMcQOIdcbtRwU9Bj6PVg7vqLg6NYeq8L7PiKWgBe+s84goWOe86DXX4YvSH/ojepJQJVO2
+ihLv3+Hw3yRggjO4SqBQ3YcyNJ+qm7q1LFDEwnXNI0rnHfv1mKs7gnyqPOi4xd84Itx2WcTulEN
ZLIDmYRICR1wnGFBMaO3HMgiXgm5f4px1qNE/Io7KgV/SyiXaeOr62LbXbRcsHn0w6V7FjfvGV0Z
1o5DQjgbpfU4YQl3c+GDEz9fPtLASiI0oXhYuvJDas68FgpN2fxuJLtQ6bgcZ935DUS6tHRBEXiD
Pzzkd5XNFCAsFP4s19bOxNF5MxAgvVp4OYvpg5C36oDLCuV5ulSYoas4XOyYqMpnnDLG9la2uVjD
n0w/NVT8OiFYf/U2CAyzxALB7tymEUtc4IQMnpo9q/014cUm53Stm1ALJCSqmnRhWLGkhFk0F/OI
j6/xj5PQ529XtQ4+HmZmN+jY/cTNQ+IgLFLBJkZZ9JDz9tE2OCAwG5aTm/Ah8TR9wTzM0GBE/aUL
EExq+66uuEfkgxFFItuonXXoAi/aq5nL6g8JbeXVWmTyUA+5AxVxS+37TmmXSQJqmR/gZsqclUU5
gpvzyTzK01V8fnoUglQKVKvwN/uVZ3AYg1t16qIYd7sDjZcyCf9LpGnE2tU3Am5sUjhi5LyeeEu6
v/9o1Ghvm21hOAr299aGYnNGtC3bDVMqhPf5zm29t00zt1a9zFLmMUNlVXN0+5UIeY9hdYNYqmBT
G2xAWvMM85gzuX1zDpIIbjU5A0RkSvOV77Uccfg/ccdZxFmgsmi8IjbeqcWzHKrZGqxtqFx70f40
fKduOSMlNLYa6zDnbu6Lo19BRFLderWoYiSZNV1JGlehlIHCPN2/xBT5MMqP6IVcsWqf9EIUFpBB
nP43qtdeL1thAb7NLB9siEJboioIU/Z1rktxgh/50+nbavgwjDVreYg2B84uiB3dN3lAfCC4be22
cYOF4rfClSTS/Gf7pKkMPDJxQERYvgMU4o3wHSE1ctbP0Cjg+kLmfS/KVgbcQMdSUUMVxxdphu3z
0wdUriLjmEDv4/6y06JCUGTDN0Gi+KlnKFMKo4DJAqoGBZloJ6t8hHt4uFWfqTDqh5EocMHmga27
6xJb79+juVr4ITMREkLwScyni++82XNO+HK2pCdnlTbqlgMmXeXH6dAlkaE7hd9eiYgaYdBC3oEM
2WFRVdDAWHsK39kGiw+DOPyjBSSLjdUP8kWzoVjUPg1I+DmJ599pTuG8wfMR4SL8zkkspZaon9/w
6/FvoGktKXeW9oYT+1LqZoq+PyBpLIyWL7m32CdjsqsRYzQLPcEz+DmPJeWnIQMn891qakcK7sOi
oN3cSBOEEdbq/akJzR7metjCAMAskqRSGFQfYPtTkhDiu4YnALoajy5Sn2R8z7QY45TjKhnOh1Zc
69QqySnfQ6UbC8YNmPwbxONItp4FJ/RsrOIq70PvtjgjTv3xMw2qmmi21d76C4HxKNo67t4T8osd
VsLPGQrdPGpLiG6btWzVdNIxtKINbNzMumbDYa0E3sdUjMYALMZsIWp1ikaEpGMHb/NbjvZWA1Y6
z1U3DZ6jD1fDatSnEPmqcfy0dpMrE/0Mc4WgKkeQfjIhj1uNsCq7dbAaXu7P1OtOLaXJuvHrIxhf
rlCPdFscczmYicBurm78UlZoxICo08KSXdSOlF9t/dodL/c5hQyJEiBg6cKHwMSKO0isJtzUt0w2
8iCzQoKQtiIiEzXxQcEyTmkruyMYcLQOduXaZBVbmhX7SBOFuj8qacm0fUNhvCEwZo9DJW+16M+C
7ZmNbUpx6fFGmL2zicCCekWcFNjOtYzBDgBoNOuALuO+tsbwYVzKhrlpIhrmaenq/Q7S95QEIkw9
3JKCGHHryvQnjRWSEu8DUnRwQrjf+vRMN7nR4dJQWssLieshAwfDLm7nX+dw6sCyK0s6IkesXLer
Oepw/6iZsl2hC3shsJCoGgRzP2L/b4wGAqgnpPHJlwP58SSACcXkYOieqVsBOZO/1pPoUsSYuHNB
XK5fP6eH9OqOvM41u7mr1e2uFm6PMAQGxQebeM48hDqtt9uOTm6YueTC1TNbqPMZz35iBqe5JppZ
RTcyuP/DTngYAHGqBkeRTI8F5dXuKKOd89B1PhuiSlGk7caHfLsY+TCxWXSAokXRaWvpLKvqvlh/
c9UQ2zTRFhGgoxo6f75N5W+24FJ3pc6xzeGWafy3qKG7dr2/HuVgafVyoq2n+E4z00qhaLmrlud4
S2DkawVUDFn7UXPWzie4W0Ip3V6LQ8HCmHpmtuwVqJhpc2/alTNBu3ajy/VWRbcREt/j/PNy0BnR
8xXlfNd4eB+eFaniQa2uKUQwDgaHBAQME6bVUMf4PF4rH5ovatvYXRmvlhA9/+3bQBr3jOcxfZoI
D0MGqOruOtvC9Gq/V8zspmfe1YJrGuQHEsKX/xDTXYZ9PDmXU4LEXkZj6e/yMA6a/lg2st1eT4UV
G+qV4O0SWdyiadNjfsNs57zjkXV3f3pxW+Kuuzfapkwj5doVRSyhajuRi5Mmc4+UQNTFwsAGJjpk
WLKadUr+No2j7UqMgy+C31PbJKLEdevExATAP1MbnBwzQ9ayEUeJNMcKArdh4uQO7/lPoqCuzUr5
oO2JbWlO4NhZkMZCMNT8sCwNHggg0QiwJGLAEC1kMbyxoT0BLGiuiYTFJleRyXrJu64EmiNAT20h
yclhKvDYgUfc927NmuEPdMZ2RUiNVZMlNtMZyJWpP/9rGhzmHUoCcY0VZKErbX2FBA3P3eJCQg6x
MlBZZ3Zwuq0k1bNXvRNc1FL1W7ySstiy7ZtTVXjyyibQ2h1pw3oqtijT5dzEP5bU30oXbRoxNSI+
HBbteA62sog+dBRbExtuPVf9vHcAVrCVKKLlqIm0BsDw68pPMtYcaiR/Gly8fHpHWZ9z6HXwLlGY
Kex330Ra1UKVLPdX5crom5Tc/zcETWbloxcLiiDaEUf32ReUV0RYQI+9o1NLsdS5L0bjklntYZl4
DheaRb6QcQ4EuqFDfrhFbJNoENY0+raT0iWeHwRZ+z4g4dRUjfgQ68xToAdMFyZMUfbHF9MjF7P8
W5JCDS8Kzn5VTi0Bov7Q6VAvy1HNZN/iCk1lPp+4uQU2JEzSGEEsQOmx9e+P1MFdo4WEN5z76eZd
VW75VDyx+zyqscRdV6CI95uXJ5j47em5gNcuLEQ9V+dQo+GGBMaqB/DT+gjOeNgmXwSfpD85AWxG
CKVE+VR/9pjT4opaRbeTGpFo9d5w4+0r61jyRUyGgkfaMSdcK6TlLYOoH1Wgvdx1UEqKsIvP+T9l
cl8rUn8FRkC84eBoKw/SM7vEoGU8b1doup3WQzUrXpw6M6o2rwVEpzmBhZh7nXycyftkVr90fvR1
oMTM7wPs6URWI7rbbjUanhpC7SQU1g89ox+D5SqftCKZ0LhApQHXPM31ZJgM8H59eL3xfvfrTKfa
dxIiaMJ5AmPFsAY6HLixjGQm67+DTb8+P07AsW0kBI/5cVjwTks3mJpmPlSqmxBUpGOtiIR9W4Jd
kiHKVFmgPCMoGVaw2dTJwmBGn7g3Av3WDTiACsRCM8wQ7YoSMRM37W8CYbVgCGdLOw35fijpAHxv
noDUoPEpuGpp4rKTr1++aF0ilRRUeIxUua9iG3ZWcoPOG3IeOmHzKg7rcqWCkc7z1ah1zNLE5wVz
lKzTlH+By+PZhZO1nqx3DOLF36XwBecjOez59T53siLwXLYwk8vExBG93MOyXLfNpLHnn98myDix
RHNkNDylSPWE8CGs3xGiM/9FjLrA7Ig7QrCTEmnmsXGigia3NJX7RQLGi0DkfZTLnC2CZYSsktmB
KZL3Nu67p37QsIzCAPRnmLAZvWP/9UuhhiiOf0bAO5vF+Jo0iz0NDtPudofbOb9BMiGyAILex6Nk
vTWvVkQShohMPlBzQrfcbURY+A6xvbZwN5IBja6mJzdvlwPtQjwGricXJb1rZ68RvsxRJ9bbfUYV
NqQudymC3PuPeR6U7ysauLo3faeT24b6wm1EeX7MG6LYOAQJzLfE7ZaNsSaz1aCSy0AhxRaPR1vv
PJItswFeOvEG1PB9/BiBaSmbLDHEfooqupavyUId85nF8gkK6tBmZzQmWvlmtdz02BqCnWupelLU
yhhJEq9CHDEOeSeOA5fz+1xzE/+B5U9aaU3fn7Bd3OTWhelILKcm7z8AzyMKjZM1A5rYbETjV9Xa
LqAi9UlzuZFsP7w4R3kjaOFVbqsKWUjHQqfhzv1V7i7vLDllMDe8Sf4QBb+4n7I09RUipAR/KyvY
UjW9I7uL/5GB8tyzv6XAFMe4gFahDgwjDSbmEd5JcwoHUBV1FgPnTOsQNG7oK0BzCCh15mitI+CX
6KGBbtNl22YpszJvXmc2lS4qcYG8ixSDVb09JOlOeRa00z1VDhy45BHkK1ft0sEgWKbt0KZ0ZuTc
zUX8U6Sg+0fXuQ9inEzpDgfIKd1giMhvhUvghMJRDJfWV5UAR8Lfnmh6iikV+ZGgXiYqnS/mHw1s
6luVPOm9d36awDaS5eGqjJ0a/sFSGLxesi/RP+oT5+NfWnkqHkI8kBhWNzs7X576mM6cipWWXHVt
je4spNoWzIgRveQ3Xo6v+dXMRVybWTtLljJ2aXc2N/OPynXhCoJ3IHYcGN6cuD8pqVQmlQPBRkfl
SYM+dO5cJ42Q2fjzMT7lz0kf4zgjhd6tMGp6wYmxzQIT2U3k8Nx/OPYn7tlQZGQt6OCx8ZtkS1I8
Ergc/HdyrHyRjlJH1h8jZOmE4Iep7tx9+HrEzQLWZOXUp2it0QKnDkXR3R7dI5CTMb05oTZCOsyy
l5rdiwOLicdpNLRFHa4A5apjx0Ox4PkWZCtimxGQvrs2jn4d1tH4DaHKl1mTS1iaudk/v2WHj1Qs
Ahel/JYlaTzv3lQRPyWz4HwKjhVD5UxUUhypdry5ZDNpJpotgGjAfReWJJNg2iHqvxeywY1wn9sd
W3xNljydP/8bpiIxRl4VpflJ9IGMOq3AOoDJDdVCJgSdFQ8sMF5tZj45AzUhoXDpeP7RGRNkLlze
+pcSKWhcC3ExokTTrEIf1ccDEZFmzc6uq9udy6pg6pv4ifhhIDnxu3A3hMJzr3eZHvqZzU7K/l4D
1wzN1dwarKznwBzu1JiIXe9/RJA8zA9huHkDRGaVbtSIH55NhFn9YpY+wcAEdaeub6TPmfoVZylR
/Q2fCxOLl1zfyngiOvJ2vp3and+oVbkjfOL7Iej0W5UzehNqMl12Z0daQXxp/nF7yrIHVbIfvJl/
cEZrM90AmT2ivsX7UCWRdipH/mGPB09IA7P7uHOmg1/iPo9aTzM3lkkN+2wSXI6flmzZrTnaDcBG
tPYlAb6TkgPHBub525g7H9chZJaPBBOPDXxyohEAiEC7PmJ0fu9bueqoMca7sb/f2MGhF2Z3D2PL
x7dUQdyIsa/2CQ5Dxjv0JBZD1yG/H+Gvn5jc1BJTysUaQRhNrdZLmRuP5id9ZAt/fZ0nL+hIQsGg
mbtvKeQGiPCGTEuot+QVGvdEJEW8Tahbt1F0Mswj9SihlyyyOB1N6jKcKN0m5+i5ITib3bkUJMn9
YK1OGTBp9Uewdm4MDcO467tP92EGyoYzjiHHCZXdkEP+3kCtMlc8XXiz09cQ/3BRHXnJwjQIZmKN
lhkCMBKVpCEIpVrn+ksllQwwBYqfudgTv0WVSCzoufj4oiZXIsRKUE1CvBC38KjuxrT0DQWgHTYQ
TydT07CeSR4V+NNuSbzYZTCGD/jvWPa36jnHL5C0SheIkEBIp7IisPZ/yank+myikJHAgjsTc+w3
hPPzXt1KeEtBv9tAlrqR5PNr7OdERL8pnGpXMK5uUH87oS8gGJEkXrtdM+2C6oSQ+RRMtLFkcgjM
+OcrfLf4Xtwp7xRnPb3ew2Ql+sDlGUFy5d9Ra9LGIMu/5BC+PVhveg+ywVWJpCdyVq5lkNAM/yjl
ArztpGR3nR7NhLzkdvd+jonq2WTxrAOTIYdOhM78nECxwDKvT0ODvRguPiqRrmRcPMm54259Pn5A
x6t9kMAwuzrs/Pe2dI64X+e9m8NfqMOJny/8iXgCximfGq6FjPOaynd7avLLqfsEz4uLAjlAbme4
/xmcK0SG6kDYRMrkdDjS2EymJQhjr7NC9c/aLTyEmS8/FOwFjQEc/DOwW8/RXfXulZqxrkCRtiHY
eDIn6tsABrDIZdDvyOAQoujPLH6cZZcWLtZiob9guspRKs+gXQMe0A6QNcgnnflizNREMRAZo0zR
q+khqa36NNpnh8gaGOXwDLgSyHT0ykh/orCDxBBF/sXndGPbbhBjKjhqOqt5VLXFDmk5XGN1il5o
ihpA+6lfu4YGPPYF030rqfS66LVmjlM85h0/njM8mBrSuIujzt3ucKOMMOs5JZTVoO594l3UGlmm
+QWt19xUV3QuxVga+dpI6M4NooOSHPBFjRMgquYgwBTap6SVGSLk+915w3b+JD+R8rReTYFArPm4
wVANv7Ps9xxB3v7TSJtpsDiNbVnmKPJ9TM1+skPcArcc6UubJMRA19po567tRgNvGud7YZvfrXCJ
TxlCegUbJc92Sub9cAB1uDS8xneMiDKYqYFkpP0BRlO0AzdHZnvdVZfkm13uzIXC7R8Sa2BOvpWw
reNH9Bfv1asZFmfO662m5lP4SbWKOhmYlt7t+LEtJYDP1ocFXJ4uoIDjU07OybR8kPJRtAXRXnJw
Ap0Tf8VVtbzBY4F2ysZAkNoBZQoJ3JxhJtykJiMld1Dh0TeLhEkE3wNC7aGjQ1tGAePBpNxL3uUq
Ipa6J5ixcC8PkpCBgEtJY6JeiNPNa4NrNOhSBgR8G6lUSoRrI+gytiKHgimJxfdoRpRtkL3b/tf7
tJBo+fX5SKIQo2+fCFcWxSnEMefVSV6/xwic0l7AfrxWzjaU28nw2SfVx7a7wznOOpD04ig6W/rr
Z+K6QfJr9K7o56STGV11t5Uvia4/drF7+u81LUh3pAJ84E9Z9w0zUnNusijAqveAnarae74/IpA1
6tqPTwyZ+6PkJajSfynm5FLqmsY3fZVc+WdyNNk2Weabxb//VSnfHHESmJbYz55KAg192fwbSRmk
x6GoClBoVFrkvjZt4Qhe+ftaOXor9X+MyqxqqPq8HbIGeBqdLMSKPwQuLFl5wnlzVBONsXShHmJT
Ho3DutFlTpN5Gp6beQJLMuqMyIU9x0Q/SLRR7i+yyZTKrbaGVic8BErfC85+CJadCcd+R8YzkuV/
wuio+YFxQOzALXs8U/8X+z0v1ryLsRU7Fon32PZjuZBSts37vzjj8aOeJy2WA/LLeYEBjRsKHJsI
N8l09wau1B90+vr/xRLJts3o35Si0z6T+zWBDeKaz/WvVFdtvfw0ibM/OyCiY3DvU4JM8ye9PzEI
FK3D9eXMmnQDHEqH4e8BoTfVGN3pl8qnjVhrwkjUJY06VoX/xh/nqfjIel74W4uTst0qbhNPQ06U
WXtjKHSylCLciPcEYm0cCBoyE9sqGRjdaalVPp/mmpwIaRxwdEci/6+jfk0WngvLBDXoyn3gIPyy
MQRYhXunBY2M3kfOtHjJ+Yj1mgf6jEB2crQlz2CYxxsSPtWr6nlL0OFq1YxmY7nLhmL9Fjv8IgCG
MhGr++qv9+NzbPBCZcK5062CBo/JeWHbeEM4EVicvy8t6pLXnQKHV+foKYcnH83qnLeL5Owx81vE
FRlpdYGOQHKcICXJxzvdNQAhl9sYBI0HfeeIKK+WNS3M+uUNzaaPFrZtqoNfhyDAQMoqEn36WMgM
wTZEYRjovCQch6RxL6ne6IY6EkI4b5l0UlJi+oeBRg1M4WbcDzoADqrhThEZqZdEsjkQ+MWzEtm7
4QZi6qP3q2+gT3d4fBZtmXb2xmQZD1mTMNuwynmkWIJFJT5dQ5o4whJs/bn9AoipoIFAd2uwPGq0
1tHHTeLvUfFOFKHTKpmPEftHL8fpFUlAl9Lr8pHP258aWvmi/anv5DWF6iIM/Uu0cUqhA2RlJN01
SpM0cbD1qB1PTZlNnDD9ZMDrTx1c2BHMByiFrjY/lreN3DkGm0gDwSj6FbQCX1GpZYNa9eaEk90I
PJJ0/jhtnAOMqwUOYUuRbjlkd4rlhx5LRlLX9Pb8w1SZnKiIr3l5Mk37yZ0iWzqSxAIUjKyiEIvD
WKyNnUIzikAI9Ot+EV86GbRe5JNyV9Fo8FcRN7LcXIb3TX5OMec6qi4D7VeFyYoKYBgKs7mQdpj2
itF+TL2Xpn5IG6Jy52UixQywmeaPjhY7IudoD3em5DUvUyHsfGeeav4Mvbg85AeECG+zaFvFtZX3
Krk+/xHE24aJgMA9ACSTh4P4uBgcPT2PHRb9zICJ5XGUTNHDJD96+CnMcyWS3jVd8bggWMtD7hCe
nJX1uoGev73fy3KG1VwWnbSJjaHdFQH6bjEBywGKW4wEGPVBgYjQI2FrGzlZ56TIssYmLeTAJ3u9
b7JF7yZMsGQZsFH4P6L9o7uXUDriyw3B5lMWo+1tEuoh/dY5EKGXnuBCC4Kv8DN7FiciofCtk9YK
Le8dxYUeC6hfVzfNy89HwPcgOxbBp0Ti+KfGokr4dKc4bTzGRVBYpVzMs0X3LqWCKyX5JWmhFUXP
FLB6xjG9Wcs2HZWM8zIrNFUBYdf2W5gNxifEeoTEqgOe36Hu3ZtZ5IDy+J8rvzw7U3fAY4jbdsdN
11R3s0/iUMe3mIbJ308jkC+itFTjS3oJPt+F0Pj+2E8Z58FutIWMoi7hpWEu6faSaDbUHK9Mkzzz
0QHYb7mkKzdAaNTIYTQAUYY0qsQxAbE6X6HHs3WVEZuRvOwGDhfjhvMbWnbpOcqml3s2YwMbgnOa
E6SS71L2Hj8pU5nYZXWjkdDALGU0Ca0rUHoFcKVBngTxzEYz/GSUgafXAHdemJcX6aV9PAsWUhOQ
a+PMUekD0ImLgRxicg4LQja5uAj4ymcL9LOrxho4CaI2hJJWlS/kv1O96lP7N4xVm4XlC/I24MEj
6/ZsGkyHwfPKzyH2UbLySIw+zXwOBTYSMtArP9+8P+KZzhTj7gjSvU3gmIx2U8e3ZOu0Np/H/tSb
QuDP6yq3zrzusE3yGT9X+JnwmhopYcYhDwoeB6hjfEVa9AG0OKgIEh064evkQ0hxwsBa4sp8f6Pm
24ILUjd67HLKa1WyhkH0VwIpSzDTKYoSyvJLa7ztei0ALHhy0KqUmAkwmx3dKPyA5wmuJNPAJJWB
Q3CeIvVtg+jcCECC3J+VZm/rJyS3DsSY2Oyh98RjgJV25LsBewwYdbG9V3RvGEtMTTQtQnMREbFc
ef8AjsbuWpouuPFBip0KyQy4qXDFQJCbUS8UwA1Gzgf4Lxpnx2oSAj1AshEARmlbgbrv+/YymIx9
Sv7563c3QF3o+yigBDXaCjsp+IUwWOGbsv5x2TV7m+B2dLRXJCsrF+K/gc/JUkl1wm8rlX9Wy/Ql
OC2yN6NmiCpG1qJIg6KafTqhWXio9YMlcpFFZCAtyNpHTkBU1ZXfJ2BUMaWLPj+1IbkC78/soafT
fdM+grGLz9ZGmeGJrXjCjSeLqCYYUJ/eoMSnCl9ad8EJkM5tgyteFO3yCpJn9uyKyaJoOWrVS99o
m4i0H4mmYJOzYJ3w6T1tRcyxdIJh+wfvBHc/qrfLDZsCa4NQeOumxCHXioDuKMtGcsvCl6MmGnim
H635Q2drmLcUK58NTKG+kXCIrXlc0hUlkIX7mwoXpKZnFt3tZ2dR6fP/Z1jDib6HE9QrtKzVYal7
uOWbK/7NTtTmvD7Q61d9MSjYd1mGLDK25cY8kMHRHkBVnLsEZNW+15qyXl5bQfd8y4SgW1kQsrT/
Rd8p2g22iOhb1AqYLGOafsUZhkBNlG5zeKsyYxBBjsNS5U1A93P5VRgQVmOt40dEv5C0RPJRcjgS
MaNS20bDPfeVWI6az9VizA1tFKrOjRdmXg65K9+sVlly4fwyMr8RD+uZfN70JJzlDsE14oGrHTdY
hzIljfdJ3k3TSCA/saAARtir+sGWFXfchQNqL0RYXspsRtNnnD7cWeQaHx2mkkLHFrZJf/ncmnQG
UhhtGDQfK2ZWdY8nREn1tiVZhgdxx/Xc28v6J/ZhV2yAqUyeQO2Nni5EBnAhyj/6tpOfQjSpOGd7
ccti2rjCaSuPm5/BaT2vJnXUaG0q12kSqptMmiR625BaqhX0fF0nLOevVGCdxUUYxzBimJlet70p
VV/HK4Ecb/2no+mSJvoaPxTaf7g9C32cZdgP77ijjsyRqFSCGA1PUFT4THc24MjwGIg1SZ3Ppaod
E0pIkIh+JDfzNO/SZGXX3WKZJNcBM4gjlodN/8GsUi3FDZoH2KdqJVLxFgZpTH++L+FRCcEEsex3
OHy6tSJ2wnm7yCmVFYlHPq33ia8H2Ww87hDzRA3c4UeS05VGKvDMFT3++pFFSyuguRHC3YYw3Ue3
qy8h/XjsS83iYMaG1nBWPAuiiUuoc9UWUENyWLCIt+1AWkDgdySVE8DBljFqVrNEQy0XvNBEXhAR
oGQRyD89pbGkxJD93TNs+ieIhaznWKdyRWqhGJNahhtEhaE92EP+lK+mGPBJ/qFOejedtMgqRN0x
KSKyIy9cIAIK6w7NEZLq8KXaO/hX8kQbOEAm9II3275lpOftRG1gmHt5PVf//d4SIJKWysppj7rG
iJR0PN7VL12E4lOaWoip95riFenMzoutYVbuZQBuZhP1veu+QocZ/MzIp9rLCq7RW4z9dKoxhx3z
0JFmYe9e8lXO2wcBfqMQYdmxC/Pf16Bis0NhdD5jw3TJ3/m3md3UqiB6F+EGoLrgifF83CO1NL/I
gnLUihKAKXyZN9/XGNj8mJ3ZKcVO48FAWfPyqYcb6aF4mFv6APxpJFLb51P81tqK8IHi22kYTdyM
xcOKMV0wuuqrjgdfOUiyIfkHmDXivAIF0gyELf2Q2DGZJ2/iuBwJ2inRIBKrVNxPLbdMqM5YYR3r
GPugb/0mEbOMPkolbUYef+VKV7zGQPNxnDyESvbupR1W5G0E5706WhxqUn0wXCBnuJ/OuN+bSXU6
xHmb0WUxIOwUE4rlvPVsOV6vAS9mepC7mpUY4zGjr0VXFpLhul5zj1W8KqWLqMUBa/nxC3wXLZGd
2GWBeRB/w+FUvq4Eex9ydem+5Sit4W6uTEsCRtUr6/+Hviiec1tjRHrSlCC5QED6xoZL2sox2+zx
WOLT0oyj3oGUFFAjQk5dLO+IZZd8G/6dM5hzjdvd0AsUu+LfTYKAbGABMAVg9V0RHHI3VLGVmz+J
dcIhLnzQjCRTKkcRRrEosPGse0hvTcmsY1EvviNLXpirnPKMp1QSZiCmp+67jDD9pvGIwQhrQfwt
V6EUeDfkKsJfTeyDXnXRC21wwjw8vXojd9HMR2Si0Oq4V+GvFeiAYj21opALXqR99S9sLC+pGj7F
1YZDkPVLhJVUbu1njYl+yQCjSplVdiL/QxVkuhl4/+RESfN7y1KB4N6q7R1Iqjd6C2qXhqTIeF9W
F/QsLuP7Qhm1L3p3ord04fU/f5c4h1JmvShbjDukQNfuekPg7TpavE+/GCD8Tj6Z9zi2C8GhnQAc
C8o19P0F4La5am8bTTnYbBN+GMdLFLlIKTlbgQKy0rdJUVK6LO5LAmR8z9yXFflwVtCVCbrmgOei
BJLa9AL91usDVfUQVfs10V6OE3g/afeSgVG8FW8nIBjRhXBplLpRo3YSpPGBzyaXjP1F6MYdFx29
h5UFXJUCxF0K6OLz0srKlq9Jxn+CYzN14fVDOog6X0Yu12tRR+DnSPHzyIAXtDbfSK9MAxUyuV3t
ZgtMyPgduDhfL893jVguaAjHp9SJctXabmklYAxjc+4XYgQ7IlB5TwfmYGe7d9TtS28vneqGMUF+
2x/p4hPN/glDIieGajY2gUjt5bwaaABce01MiqZ0zMQUSKPamPHouukIz6cvi1n4q/qsQwGYK3gv
EWgIfq8cPA6mGHYYiD5Zpg2IAHujOMQptyfVw4Ma2sC+H9yUWAsGffbDlY/nD0J6nCKm0Nkv8QCl
e0uhTN5QwqiQN0rH4I/GMjiBBG09q2v1/WsiK0s3BszW0QD4iF1J8Z01uBnV23KloIaUSMZOKKtD
68IfQSpUR9Qy1f5q4vEGLuJWaucBEO1/XtsrbimtGbRRYexFLK2bNA/CD0fRKf6kOYOD5fGQPM/t
IrjeaUm9HVs6B5lgFWvWVV4JimUP8xeYIObcEBTP4YHULY/IbsLHbA5hicda7oIHHzYlpgLYoUsj
GF5CgdtJFzaw4Z7wzVfl2ZxZyKP1b1lbhwqlu/6YrjkWr8uPzy9UZVoj5dKsGNlW+ErlCcF0mcL/
ahc4nkZGj8xlOUvkxADRxXVNueNvjXnzJF2i91fXXuYBaR26KW+g0yBTzJ7R9MqIDTffGqlj5C8o
+11hzK/7IJ1VqXpWdOVrq1AioFENK8yldB2PIpwFZlpKc1jT74vKs/0cUtvQOSi8HUwzevDZw8Fb
9vLCM6QRnewRRO1LInXDE5O9Ar7boXh7ewscGldvZCH5CdxfM1eZARf/vpcH6/EdDV4GKLPoyJAq
9wbQix9maVL3wZsq0pn4/3RuD4rRtPhbOfOZvHd+d7x1KTmEfbsftcPNl0WyH4kAF9YjIWA7XorK
jlRGlWT6N26Izzx2pQ+JP1Bcr4P8gdpwbOWjyL0W9jd9XMec+r3krjT2YrknJZ4VYm4Vec24Ht8c
+U7QpddREgWNKskBYiQT0Ack7WuGHwQkLnp/3MDTV22AAUaJWZyY8Ok+gVNtmUxO0llN/+poi/jP
asWHpzq6rdzChGsEawm8/oz8paGiOKBKpBk35PxiuwEu4q3H26q4NgReRnRKIrlXzvLgHvnjRuAe
Ge9pYsy+Ypw53mbWEMHNoucGgHGmGbEwzJ+EFcDY0aL+treth6jrIMyzBdaqJklPapvlLzJ7pK7i
DHxBGFe6adlxoRMc06hQYFH3Fk/ybhDrRfn/tWG1Qm1gOa9Bzg7KmP3y65a9zapSstDiZsBlGaRB
MmXY4L6o+O/oqYiD5QLJKP0E+2ksuTGC3EamhDvdZnHijeI8bkfp8V3V4XGiMzuAkrcoQCKQjPzl
LWtXwja2HEnf7YUwLkU+i+Qge4qi3mK8VpwaJXB/SRqnYxdkZPAGdLoq9gjC+pHXNfCqn+cX+rtJ
o1IuHeBgtMNUCTHf7I8jAauW3cTpeo+80GAeOqf2rBxKHRwbwo5ErJ2xYmeDmzT3BNl+3SvnPH0d
6k5TVAxs28F/mLX+1EEmLZc50GncnN/eRFZDjLnoJXs79LKdfzOCAhLd+LapJDk66m7yZptU4bTw
SInZVLELRZFbSE6IDNjT/KRFovbGJHn33VGH3LijALsZbRcacVuIPomO2hKznF9DyS+1woC1qWwc
zXkc1pBP3ep/fc/5FutLJkXs/grtDpY6JeUPoi0VIx2dPSsyb4PV6uM0AFJ+O/eHa6ek91MWSUVC
5Z8flbsxSqeZhnzVbGOQ3e2DHNsTam2GhNvePl57AHPiVArIaSbvvvj1T3D0pA+SLajw/9qWqOnb
Cio03cGz20CnKXoobkKl1Ue4RGb+aIXP1UGKJzGMjTABPKFI1CUFiAP2Uiooierh51skvogBNAtI
ACQi4KQTfK5J4Q7CoBH8w0YkUhiyftV51RxZw+OKQ/0msN+cVmiQseXPbortEyW3nhV2idRDzdE0
lfhH9P1QTz9+TkXTju2S10Rx66cQyk+wmXA3zSZSKyMEk5ZqHF+qylzQ41DJFIoxIQVVT7LSXKk/
SFyHFhpjUEwO1aBKXROqt2Avqb2X1strAoM+1r5hZddrvd3Iu+BNhAY+qgZU0bSd1OqP/Q3bRFc1
qgK/ZbeOffn/gZhdFFrRDi1ZMsaeTudb+aqY8jWmtqSfu+DeWFVlNf/IYe5qYlHR0i2kFxCQFRaz
7MVhxYqCXC/qLpOoUgKzwJIMBhv/YLlMuzanGF+sJtLolp+84fhBG4RIBElL0JdpMcKNh+pCJ8vO
1vYl8RzfQpWYm26682YjvXDIxu6VJvkokoo/mQ5UkJj8/DJoDDTBjiowlk5B7kCTMKMvFZ54NB4L
gp7ohdXxTocsPjEalwaI/YOcA9CXewNrNTe+L7mwguiaToRAz8B9DGNGzyFlzDRRyWetcswVNqBF
dTB10KVHYqgLFr59TYdtytmuMENVAJEuSu0Ofw72TGI1OWM5osBeDMq+XreowqXw711oAF3+36uL
cuFiDyvQNBWe3huuy9wA+C26J49VjPRH2NDqLqYRksUHo1sErvZrJqvvmTZ+KVcKS3Rt/2prncwA
1+4JxPkybJyeBy1GrnaIZkjVDOvS4h8Vs2BEUcr3UnVPiH69bg7Discheth4AmqjEtsIKz7IXZRR
R2n0SmWp5x5s0P9rU313M+dCFIPsHVXDxfjdfxsQMCjdDypQWLNk7lvBP0WaVOSn3UeDysDJFDVs
QLduiyIhsHU71RONwzLvAoSn9VxCjKR8gYjvNZJKIo/D87/jsi1mNsMPGvhy935YnzYqvrq3Q5Gm
dRHSeIbrxemtAKB17V1Imet0Ekp6rI63O9kSWzvsUj4Gz/UNmGIh2ClciPIULnSRIHfll8Kl0XGg
Bp7hXM9J8CbV9dFFXFOkTyeKySS/6hKf7OjRtjyYTPn28eRQeNDtDYptRjkaVh+e3K9TGZfJil0S
ANQlDbSdltiYme/0/DCGJFQ7iCXl+zqdlbdmyIlIow89uqEvr4Z+ADPDcaxVzXFxEwPXJmiIruiJ
CUAtY1EXsMgsFqQYJCxltrNaPbfwcfIbxgZ7/HYl96pfNRQcyu4t9Saj1n5z0udz16ZrfZTtlpLd
3nWz+Si5jI31Ov1oyq+NWV9T2gySpyNOkp+y3rUdoeibUSrtHh8Vf0iVTtcVMFiH/ggZR57Av2tq
6pye/gJ5o1LoMmQczm6uSmIDleSmOxe5VPwEOEtrZlcK486Atm+JR8VLLY+ha/fTMqnMPW6pRnF0
O3HTKrEIP8GrowUAl7bDzj7pVj4WONOlzE4rj5cqbItTMl0g1RSdgsclVjPO4l+Y1L0IaPAo06vT
5n9Pt1XakBrjhwhI/1Ts5EbU5IoCexyx9LHDUd0b5TEloHAeas4WIIZx2KhLmzauvlbso22emJfP
OUoSHGg3tpD2c7UkKglykihZxs6UJQESzMtBfmBjXUbxlJt/thHRass5YKl/gvHPYx2U/Of21Wzv
Mdq17xF0Me5jgqNMptRDXoa2tnFUG3rSGxwB1MjvWGcRCYjbpxJt/8iPToz8+3zBkypTwFPj2L5T
prvOWH6uz04VukgRHx1M4E+XFnNTPGoF/c1I3bb6peiliTsP/cy87RughY4Y6Tk6IhCMjBWB5piI
X/CUD4inSOqObp695gxploKZNk1gc/Wcq9UEDArdI1oCG4zR7+SQpsSEJa34D3oVzYhpRyX1KIQr
j/57eLlYv2st2ijqrToCRvaiRy99LTttb3r/rIKhaDIFcg6NgZehxfAWBNl0IYeVGWP08NuKQw2l
y5ivPzDfsZ/MKSgFBCArGArv6/jwjfFbo6qHnKo+b7Kt173TdzwkC/+qMMPd54WF4jRIxJ3QzDFF
DegQJ/1/2BhTCHNGNtCnx+u6HmJMQj6eHvRjECWOnnVfwIvQ3hSmOAVy//zmmgyVxQQx9UVgZayU
QvnNxYGzd1xp1rdVyyGMotwk1axENdHlZ2CfP/V06JwHdMBAzUIhU4QLOy2WhS+puYpAgxsin0gM
cy+q/lZ9KQmAoUUbokUQn5+gAHeklS8ZXYD7XHkUHRZhvWWxH5GSDcp+IMMQOQDQo4AdEIoL3rKm
mKiOSXpb9Fi7VFIzgGdkXv7raLMkF4UVbybzI4T6VkyaqAkbay80MYCjxXmUIR/2i02UXxPe1w2Q
dEaObn/fSbCLdubKdJsQsmvv0sbcUZElFaQL36jH2K5PqpTdiCDYYj/IWBKpWnx2fEn4slGubBa6
FJNIuzjvBtCtzOM13vpJCo68lcsSO/rkyo522jL9p60cxJ258OW1/qRj8tBZ7ThvoRvEjxV91zf9
aQJIewFYB4ugEiaWE8aFCmFWeFrToY/8oaihZ/6dcr9pCHRGBOX96HTD6vrjrKIjm1UeEdOZOZ3l
yTbdLU+cdmHfwGnD40lddPL98xkgbwSPOrCpttnhVEenxRz7lL3kbazaZHHu1rdFgYmMau9Qle/t
vHVkOnVhnRh2cw1BkAQx7o9SREVRz+Ky/jhsa21qFCeLWz06lbRegrKwmfprNXyyVB/7MAQfvNzU
y1faZZKBqG9NbBIEIqFQ4ZpvTkn0j+Bq/ggIG5kyMhwooOKpkpLGoR5BGyT8/Jz7IFzX5MPjJjJB
cE+XpqH1FaQ6qWb2/7z9tPuSv/BjpMAJhaGOKA8f/sILyUl9/AbNFPoSGynKF2zCdaq88bYE8OTQ
2SeCx3lZpdFTbbsNltCbR8J0hzadWHpAYIswcp2NRnvRhfrzSF8i/9+Q6QsNsEoRnZOACSRBYdhy
7GhfA2RQut0RYqqxGw9jYNC/wOYGi10XtyIw7KlxGgrCypeXZnZPMFzxuYNaUMOw2Ynhcb38pzsE
27eeJHqP33j1DGXd59yc++0mEvUsUrJFi1iHJ3HcUp42ODXiBuiIrrPRCrWAkr0oXM/kS1oqTsBe
H/CwQR2/745FgUd/tH5jfUyrJgjbeeZ0ufl+WI3fWVq1zGpU85F59A2f1cA3tNOFwRTR6VoQ0egB
l16NNGMcFr3boZifGdXrH2BKcsve6ZO9jw4BfNbPsXZwrKFin++TZddyVEejGlpvngarfaW84SgK
Ho3I8PjBqcLDLcWkSFHM3xZdVaxKs6FJ70KBIFT7EwQT0ZPfI9vZ29ovlajBPYyVUlfJe5NvpxBO
FMp90aKqYyDtbc+pO6drlXvBLFbMUGg2+70sYsPHOLL3jPcWSGtZ9FcPBpjWpk2bmLVS1qGQyCpY
SMF+PGgL99C2XgIT8k028kisbMn7aqDcmHVJgFSU5lo4ZiI8L31WrO3sZ2NRg7nWaEKCCQVfCZ0A
vKgc9PqlW/jr1UWGGzTcXvNQBNacM5MGWJZCQ91HGwa5tnas4Stm+5qOE1z4Gq3mW4S22m0ROW2w
9BfvP86aSmTuVbOlHjwqjOazYzBjTgRHMV00OoH6b68oZCCQBoeIq+euX/ZbSeTvVjnkq7QZDUqF
d/HXrD8Rswu9KPeFQzaniOlfe9eY/EZ1y5UQ4eCeu4djLwX65KwiKs9laBGVwxyp9qTmIfILR6ab
ZTnagsFMhgX9yERlVK5ldfN0fbQBYKpTIrrx0uuU+rEIuoAqAKeAGiBdJeUDk+W/tS8lgJ3IKRjb
qPgGnPJan7t+WoWI3ds/1PuXzMTqje44NQTIo/2wj7r5+7Pdr9Khl4t3kxGnkS+6afKQBWk6GSui
6MtxFXCylBZ00ZtEN3xgcD8b9hSdJhZqWwlXCCTyqdFbs+1Nn8IGGYWwP8c+pBOdILfuk3QAg8/I
UXEREbswYKHgZBqwfsmYhHRN30iFOLRdHbErCU/O0fk43OcOl4ZeJzIvrHN9AEKKkWtyT190U9z9
aWYimx6HRQ++AOEjk4uu0IA3Nll0OXAES85aaX3Kt5ROuquQHRXoeyz8eNPeu4/vyhJCu2U3MCaS
RdTvkVI99i85WmXiIjD72YTzwL8C4EWH9tmbq3Oed3ETt7S82EI4EoSRnwXwrRS7jECkOD9k1CVl
I6isZuhI+n+UX0pkWK/rxhHrMZJsswaoVxEUsk1VFULcowEkoeLfYJe9H8/y1rSReWA+6stfkeuj
lbnTgSPsll5lK02tHa2TCLQAVaxJtDus6XuWJ8AVR8WmGQyqEyGH/UiNClE2PY47T7nzkB+Qiu6Q
LRfg8s+8CjjjUiyvwwFq+p7TK2zq18Mfsbz+OTyLIYoaj/9wQ/7Q9/F+wDNooxP4dgqJOH16DSi+
GYCPY5qpU5B/ot7usThQIajXJdScpNdFCFuwBVWcgyLtrloYr9bzhGpmzaM0cl2BnJ/mtG6WnDcK
AvlAdIwZ4HJmBWM2UjmPAloEWdymyPQkGSrHBEttO6JqcJH1lbFfVBSx/MrL1UyNaf2GPINlNcLl
86mJmsF6kmY9Us3jrE88AndR/gMgr3l1XlYAsAZ3GpL1XGWLGX/nlHDdSM34zNVXCzu3ppmKSI54
DyeQ+9HTgngDfwr7Zbz6bs35plUb3BrLhSmygq9XTX6i5JCjsQY56fTzH1K73eQXq1P1shcMwL6z
WCcwA3NjThn2iv3DRVYfhHAiJFPafiHBPggVrve+xcjGmfm5GsUXek0jVhYmz2IZ3SKE4iqyJFjK
eRsbJHCpWI11Yg1L1rJTfMZLI44pqy/ogAukbb5xqWskiHPtPYlxRdIhlHMtHY1CEqFKc4kPioE3
4iQwZ3LnWA2D7ZVzab8w1QuCGUMcphflI9t4IPb/11rAJ0M1VfEkuFeu4JJop4VMXAidvUVKlCq6
wtRHEFzOJLINjAxWYPaLRLfcHMX6jxZLLu4/YrO0pyHI54jZjo4goI1y/F+SlNWBSH4DV+sdtpW5
ZXcsqRhzgIGDiuFCL7UA9Vc2ty9zyGMFgxfQpqWFSdNXu1bVPJ0Snh3mlIvQyJ9OAtwGLtxl/ND8
yP/rvqMC1e8OAEnoJPSfo2l8rvPNOZGpXWP+ADGLIZ6Cd9dGnk2S7joYV/SRjYzjJzGifAEdBphi
cDtUanifJqwqiCj7wGXe2JYK21CTtBJ1mZaMvP9yMpxnpq8fq9bNz7f0On5rFxwBKMXjLeFTMl4a
io84DYjLNJt+E89I2tj9Psaf2z5i8JIaau+MDVOuowiO6v+6lfEeVVYf9Y/58sbIEd9sD/pNE3sP
Te3lfDPUsXDImUH6Y4bbveKo0LNoIoLiPITukxQ0cD7QzK6wtoS8J7XTlpIB4N82BnFa77oHPBi2
zl2nblFabqnsLlv+3MgIgR4N7AhSBBqgjbTKVr15SDtc1UiqRkKDmwv5PYVe/CT29a7CtoAq0U1S
dN4iHMcqHWgO2LxfxuAmMbepJvdN8YxCCAOc5A6mbcaCHKSqjvG+XfDE4Cksm1qpTJz0AlquxsGy
XAPYsDpTN2yMOp7QDlymW6pcYdUghYDEwDgmIWzx3g0fTPpxxVARPhprdBHlJTos/jHHobhNwZUA
wrTmUjE/8LdfZcE+h/1a2LO9/vCP8ogyBazc6dqcnaoRjOd58hUJAHLMn2qkXKbU2DEGkQYww1Cu
ybYtxxNW9PWgBoa8Id25e0Ovcu9ZQbt+7Q+UrifpdDDgyDvOzPMWmp5qEkRsiBJ7NwfBKMy/FO5w
0fHlvgoRzXRX4O0GLA3DzdzXSUJEA0Hm1wy7ZDebd3unTngZppgi9WE5MJmmHNvYvd/hKUrLqQeJ
r7SiyCDHbpWAnIz8dKHnt30ZLS0Ax3tgRNt0ZgMFAuBmM9MNwSsWpo86+C4IREYukxExCUda4EVK
4BelHRGj4fXG/Od2mtI/jK6w/2AAtzio614CpzN7+zoSnh71BwPMuNS5ZTk9PNAMKTT5AEDvw3Er
H8Dk8LE6OS/0OoN+Dc4An4VnT80m8dt2fpQ6Fn7YdfICdE7yyfLchLL/LTEThmOx8Fc+8NpBWknl
qpYyHHslbt/cxJPOu30Vq7E0XOn8jQxXFHBFiZ8GVp37zunE3i96gecx/ijh4ibPyIkutyOn1Vw5
QixSrK4+DtOOcQzpJ+plgqXYsO5O7WkDg4onop1G+qA54lPjE+p/I3rkv3EyCJNYNIzprv9QC+2w
VBGKUEKq8ANmdXhU5P/ww/KO/B8uZF+ACM7Q/YbBtkTps9b4yGpYOb0Xckkj8rNWXG6jYkSO0Set
AlW5T5NCFSG/5rBtH455JrbjKjmfPUrd31jFGVM+rHQM5CG3L0RqTdMBKdMh3uk3TSE4bRlUMZjd
ueextwi0Gi+5fprAND61dj/jegETcj3EF7kXFx30yk5FqQO9+VIJBu/+P6YpIb2i3kxG51oWtfwM
KEKlGzhxospSFs4DItijeC1ImDELyr9RCs9wwxHaZGHQea9I4VnxA83CaLEzdZUeyTEX2zJ1qRZW
/4ENu5repwE3z2OJwciTnQcg6+OvWkQNLMigLvq/pk+6sjMuZPvkgQOgj8xQdjLVpyw/6GCW+S+e
i3Wl8sOsZbTFe8i2gntSNdQ+zskE9zoJHKYnjvAj/CQ3VCKk391W+HalYg9kS9ppbh/nWnt5cSFE
C0D7JGA5GINoQm4To72fL/HhzpHqKHhfIA+KFW07MGOJf8VEyf2jfjA4OysXh1ONSoRU/H4tZR9L
HH5JhV1H3+CfagjX2pM5p494qcfnxKR5SqEn7A+9s9/2tEyAgqmkit89cjbyGa/2LqjMPW+2T0vw
y0fEKVZ1Zh19IIOMtDb3T3fT/H63QhYg24tKZgjB4uB6U77+qOo0WxaMuIG/zWSAgYpMtj9lLrZq
eZOktd/Wlxz00uesKC+2FtZqGdtlaIRt8v12okVg64ec7pXEnh8/yG/rsJaADabZJSqkmkICDTBa
kfJON3uvoirIuVfbmGiayZejq/JfZFX4iNpnwg7Yt8yN2IbGVOi8UYpowJJTo2v0rLGMmv1W47cK
I9cxkiVgjpHSsCm5NCYfNAPLerQ7oHV+e08aGpm+QycOsw2H1sHifV0jRBzJ0+O1mWkortAi5rm+
+Q8T88IoMyUyYNkj2scdZYFUVSTUr+M7rr9evjMB6lJ8nGH+lSXskKcG/rF/2cQlhfLDhvxGuiWi
ZURuKJ7IpdCQWbVTiXrM8s0o/DC/O3BRfwCiR182rsoObVEIsgZ34YhnhCCgB9OGvq60ZApZlZ3q
vSK/Vmsxwapz/cnt6M1xVw7eUMVFG+dAAx0V3oxQD6mRIeocvZ0JX3tXjdeE9yrmXkrxBPgahNCQ
+ogyIQeJSoRE6tMJlLSAQbQLvHKNtV6fEqj/2PshUpE9UfVOqXeq9tZI5JVPJ1M7cnShrqE7JLaW
31gx15tDwgcCQdGOiwTLM9tosBZHxxNR3e0aWStc3H+xYw2z85ax+dYfUOSIuGtAXO+fOH4/dM5B
Nkh1gLTHWTWFscmCLfAoiPmAGVKIUTfi1dzylvOVED/2cbxwrn0jJRvPLhWf18Z8c7t8bzsKQPm4
9Kmg7FrGjOWEr0xCL339qWInucICSdhkEfETxeDWnUHzLw0GB/jY8fzs4oRWl/OTbBUKv/p2CF0o
Hb6HIko4L+Fn/uvBluS/ZzoYTqy+7TavaJWoEfltcleA1oowGxwfAR8sqgvStt9fdWOE12AnCaVt
5aB8/5Gpb+oh/rmiZz6YKdxR/hgwXRrHsv5FQd9QkueUpB54RjXkyXNkm4xEBbqnlW9Cny8cA4ZE
k9RHiBGuyc5lHs6lPiGqFIBkI1g3OjL1aWovefc7/W2o1N5F1ez4ovTtds00C37NsW9wmag4Vu8y
/B8QDTBWbquQlhS69lWW02uWGu8RY4jIisAZc8F/QH7mlHSbeNeudExafQaYX9m57ya5mGsLEktr
WqipbqEVMwvw+kyoVatTS61Kw15Mjx8vt1HyKGHFM4ARh/qCzMvAQ6LbLCwra5jUucpO6NTQdSNd
Dd+15UXW5x00L0JLjmDmASEkJSI+ZNIrVl6BwhNcdPTlg4EXSns2+lxDpShEfhJyHK6Tuv6jPgDx
KSAB6pXtL4blgFpaKadm9Axl8BJCnUM9zHmrwq8sPynZRNeqin5PTi31vHqn/NeT6f3lRtmFKOfE
kG9aV8lccB68gf8uRrxn+zEZqquCrwNLCDqh3naRcAh0pFzWh3AvIEyMecWNW0q7nFxLKtP1Rw2G
rvpqwdrA9OxJ2VyQD9Ek5fqFwPL4yALBGjv+CP9aJXJyFH0rg9HAFjd6T7ODY9IBsF+T0V8J8pSI
ocDHwvEnt/f08NxoeURH+cpO0eZ4BuiIHXPs/I9wgVBF/oGBpQi56F1w421hyUFWJGJ2hCuh5XVt
w/pr/QobVhPAHnCl5hF5swUbWuZ8gED1jfd9Be6SiopPoKfpEJgTHfmmt3cnGuO1CKw/uE9VCRvg
4EtVitpjqz0HTT5NjtPzB/7+dIRXHMIUkc8HO2XTEbNbPQdfw7LZv5ADQBvC4XaGC73cIKm5AtWH
r+MvxvjdoMrDa4hwlvsh8xQ9ZVB3Re8U20+8Z6h7PFtM5krWAkgn+f+Xim7d4yjBOFrpGOBrHDgO
yQmHbzc55HzI62V9lOO76NgQIJUy8e7yLgJR7lQHVOvuI29FaMMpoCS+gLaaiPv4jxhNNL2jW6f1
RJY+nTwAleZLCxMkgqyPt85tnirTw/oOMLCNh7DZhzVmN9jtuknEoyukqMi57iOpnKdvhHfzopBi
FDTFqrDlvSU19IoQ/cQc6YQ7ciBZnrUzbbrPMmgwB+IpH39Vpx/fqmTnXB302xZHeCRYS28OZdhZ
f8nISFFgpZAQC6s1oyosRlU8FSIIuMm+gVhlqB0dPP9o9xsTmHR8MnkaUtNpYbGHH2vtCQbFSWu5
LoRsvyCrPN0PF/UMrrW6RFoZov1R1700Uh6BurdbINPx2lfGwRC9AXfI6YXY+oCSpN0p/uAgKSzg
+KECdgYnEW/cWttnsOIRlQlz23a0qggu1SJZcecnEJRnapgRrTtZOoifpepWswpVjihrLriuYs9R
vHHH6EgEcrI5MdE85XULgGlo4DwolQiW0cbkW5Fd8qmAbWlg+YU9KmI7PY5VyR4OD42GpJdVuyIt
hlOmIahW1dPZt+OSK7hCeSYglHpB0GnBxsEt18M93PKY0o5kb5Lk9LMv/hsKdaQUE9gs61bObU9n
fyR36ABI/P04cP1GfxnQIyRAgeet4wo3KTfXoSkcejODhFR9FX7M8fFIKSejTPanwAcJG8XPPuB2
XlCB5JC3cJxgCzZEik3TZz2Q5KpHzBdalfBkLGno2VSquLFu5vzIQfIsc9+0rxkbZF5vbNeIYq/+
QuxH5z75Sgzd7rLJBVTD534en7rbJwpyzrW/eRRVUjVUpL1Chbo9bHgWpFllKuMzhvyptPsz1iht
1+Aj8mkVe3Ug8r2Cnffkhn4dsQY0ZxI602mwT9sV3xtBPhbH22zL5NTEMuqtFEtCKl0sZilWyNJU
XDQdmAeuPNtX2kpZwO5SeIFx92ib4XfPcZhsQvH+3wg/p6WDw55xTLekWoZpVOld4lQ4EguCMPrR
ff5lH3kSpU+OjokPBwB1CwOgy6Uec0xRBBIwwjiiCi19skOI05ac+EmaX59aX4qA9Yx4G+oEGNJe
66ErnqYjEjKvfNS1qCEOS7chQ4KPwHdhveZjVo/HufpJC4eOMe4Kihyk1dyGkHJ+Tyz5lsw+4Ols
Oa1X7vJs4bQAka/Y/a6jJ2RBwWwOCh2gMTeeEdhigkH5yyMh9rPSCuDZFd2yQHFEQZWq3QxJXaqS
clNcE4YOnqxNnH72djEpzA5HVMdHNNDi/5QsCL0Q9DN2EuehsMfAjpaCypLhxNSroASFcnIdb05Q
UgoGUMHHFs7uvtaBwvN3fM3YoTPEc75UYGSsTaKbP3RXNfY8xZQgm2XbXlX5a3HGBC56ZhY6LKyT
in3Af5OxUb28dKQ9Ala9o0Dq8s3cD9IMeiDW9wp8aeCUcgdDFkx9coHIuvB9QT0zr+QxtPzYuuPn
rcdMxqJq3w/THZHqoeyMjTQ/UKVBijKLxS6apQElmd2c/pkfpq1DzR53nWL7HH+K2QPc39A+O4d8
VLwaDtwts66DTM54G5ZL5K7HE+6XHHJ2AaO/pjiT6x/HfmrYIAFkTaAHvCPPsRtuc7oS2KvqZa3p
7QY5gRGXp2AG0Os+ZDAkTu7M8OrRQQl8FJjMc4r2LDyI9V2PMkK6zV6uOPcNKL8JeSlX/bvXlnFZ
b2fWadSrr3lfmQOxnCBO174YfxxbF9pQbNVZLiE/ZrZJkkKBD1Vi2zH478PtxFQMACx5iqsHQXlY
HCpz5843P46/ZTox9gIxmZvAMMwQ6eHQhLJFwFZBmM2iLDikbIPKPxzGl2aSQq83L9m27lloqXA4
Gn9fgyHv+i9Vwc9zD6P6YiUnzoLmcQm+K56a+4xYP5BZRmeWvQ8ZHlE3UIy5qFoM1aIWDxgun017
yZH4wtTJaih0Zx4HC7Et5HtHlaP/Cf7pBlmE8S+DrNlSGebSg0bu7gRv1YOREBFu2/uow1XP61xu
wOk8qG67oIWeoiEt1Ki/RKpmml81uDJf0QhEkV8lWTkCTRKHkDlWqt+FcLxmLmTlG1Rt6NZbBb+S
SPO+ZHQgCsBFwGMcKawhLcYH6ZjhUTARg8O01wBkHGOgodCeDMgJnfwriQyDKYtaoP+qyqSFdArp
v3+7r1DpyN8EpoRSr8b8chzSUWXd7cnDad0BnSH59NX0GMGBMBit2pcRZ9R612qod6+AZdmJP+zm
kO0RpupU9SVVGWvO/cgs/IqzjVs7BW3+6NJSeMQW7bBIsrcl3obw5ylTyGcbmjtNtK+6QJl3H124
22f/ZcVosomuATZm8b+vIiirCirccawGt6Q0ls17MkohOCcNTWA2p356d1+e8WlMOHyMvXiboOuY
TidojC/5dvwAd6NvwZQSI9eOsXiEts/oSMBPjLOVO63piAOUAYvFSc5xxtXS6cuATZX1XOfwcNoE
3poAGaEim+Hrrv9Ww3OEecmf3VscAOnAFWCCkwtJl6XpgE6dXLNgEgti7z1wlLPEiSr66DPlrBWa
TOg3WFjC14YKgILo1kI4/+ZYjvVHdYwqTZAB1xq710JWoHS4WQL1pMgOKWQ8eeWbQq3cVxLJx5UM
Q+atl4vOPmb5K6Zs40N1v1ig367ZOjN+L8aHTfXKHuXNUQw6ykDL1liWQ1QILNoASFAjrqXh44Fu
rvm5U45LE94Fx/5Qk//UIl/KmZOnu0pIv4g4P2OsnrDQ5Paq9mJ7Xf0JMY+yeMIjiINWp5eu2EmP
RKsqlubRT9Ngulqrg9GYgbFqC2MnKxJo8Vb2xa/m+BaqGz5l/VUWdEbUr3DnmAtOv/nUO/RwaTzu
Gi2JPzMOmm9HkXMYa/eyvIRGcLLbydBnTL+zkn6G67dltBukEq8iuSVi2uMAVuHZ4gQOw3Gpvq7G
5nW+OnwKjGfvyPnOCBIxQQRVY8P/WpV9y2KfT6SAtX8ylI7u1DBD8PnQMnKwg+TgKczwwTScvIIL
/ofudWZA55BhVpycgyEoseX9nsX8D0oYkkOwq9S3LNRJLOrEbuOTmfSfaqWC49eAmREn9vjG63Yp
17QjdE3NJSKWX0YCBFgBQPngCs6A2+tQkuzg2Ol6oqr44d2ZsCam6phjpXY8CgipagWsg6iSlYVN
OS/SN9LQ0v4W0hpi8b5ZR7SoWcjmlkT2NbHe8RTc8c66xGlwVCtu4Ayu4vSF3L+fAeF3UXn+QaZy
DK/FzLw/DhtYvT8vg4VeovM+S01JuCl0g7zGp0klZurWtlNu+I4PVPh33LMTQIkH+XbRJoL+7Xai
b6cBq4WzzA7cBEx000uSH62WnaycbXLi6IRze+Pnz3x9NLtD92yty+h9fbDrN2Src+GQvmJMKTv8
n2/DvaVWCTBAmCgbyV1Rp0szlMo+O4F/bI/HIwPLLyR4DRLBEWZf0ZF0EYm96cawaMuBSsBULTBt
Lspofv9FdY3JwlUOrundQQ97TJOGPlKkCgPnQEJxESUUArU3wagPqx8udJy+yq45lj1DwxdsnTbE
wumI2jpCtUh8krj4szsYAKkIkBWHGZ2YpzipLGlkilaYESdhfjPn/qCPW46WWAmx8ckBZzsgAHNq
nq9SJAZU65R1ACAOVVvIt2YTXnDLtVrzNMS1MWCgW4EFw1DNXUgb8VBrZ1r1zUPB9l2blssjnsiP
tvdj2Pt1PwCrdVUfnhLBpr/i6uA3LcNgN6TIIvAeP38apBYYjWtUTpW31WeNBXkaRUHadwZ+RqyA
LEdzP3Bdg2wmUY2XRowoV+6R2MXkk2ZtkOcKPgiLoFKFtt1oaBh4yXMpor7r2PZS+buKm8tIz8ob
GhiMMRRC99oeDd5C4/ohBDxkj2KlQSEX3VLcbJ0qIPGVtICh2/uhgYC9T4aSOqsMjydSrOJ65q23
JyhRElODxkUUjNBAGtj62yZKeA2HTigz6GL790X3JsRGtJRlvBQwMzvmgth91y2pkd9pKo2emcGO
QSFKUK/rYXepAlsGV60s2W0Q4fG0LvNscWCBla4vNysxge3lkNmo2AsASdcXzvCtVX2LIvYd9mVX
nl8umK0mEXbJwq3uFlsYED1HpLKdeAZdYmWZY38FChmbZCuOOZdHNW7FYq+htnwg4qpBW1LaVKQn
V/yD7qs5HYgMKwC5Z93eAB19/pGLY3Ix03otvwV+a6HCnoB66yq3OaXwNXQZP6g5kA4IjmU4U/Kv
H9tRY6hTI+24RIM6s+YdNOWjZHoxslpq294wnpcLbRenZImj9kzjRZTrBDNyhmXxlEmf8eh7JutF
m9AVe4UI8PpPAEi9iSBfJXWiRhEL3gHzGjltTllGJERMEkS5jxurKYGn7o1R9JOEk9qhpOy9QXZN
nsRTSLOfWb2cjstumY3cRMyRjQ6fdVqkaO1nFf/00izqu358XIzC1PKxGFJV3QYDb/nkFWaIXvyv
rG0MydF1+gb3MNAbo6EC6d5MVboU6ugLJ0y4KWCWfTBjOh0EBIoeEihXmgN3SX/lIXDRbdEQk/hy
GUqKytqb02picsKBUiDLUdf2EkXvnET1jH9z14SRmdlslDe/umWYrfllvZsn0oU+PYYrxaylgdmC
c7f2NLuge60U1sBs6Lu8Tb0YTILtz1XdonpybolCpFFZJfVByvzH3mpGOB+SsNGaTgMH0ywbfOko
dnXr1u4A4zRNHNeWEtlwypkhWq6zWg4qMtvqeAXb3Pvswer0VhChW7yfF+Qazy+3c3xNjY+Wjb6z
8ucJjwffN16k6nrqQifKY9TqgMpaBVuM6yf+GfG7Ewp+YZZTFkwgnMmGVIUyYagGjOT9mMP6D/hy
fWNaPOZUPPPi384VQIcBw0GS6gt06G3aLdSOx7GIlq4fmtRyUdPVRrftWhqDXOkgAilfELbD6MkL
gLWpM5VDan2h082Hrlh8HN+Dqjf8nOUX5bx+aUcK55+n3/TiiX5PgnnSZiBGQylBpzDM9piEz8MO
z+y5PR/HaO4CKjPoAmLlTXbsWkZ0pTgg8CpACcDQIx9OplqZ8SL/yOKU9J8CCbv/JalUlcs9clqr
kkiiIuRW7/pXXO0zINoDsIcWvv2RBBUZRVTsXmttn9ybMoPeBGPijYQTkebItGV0UEN/8x2mu1U9
4ePRecEhU8Dmymnq6KFp2mbjdR3rY3zHa/aLCVewcO+HLQfQRhcDTH/EYqLy8p+GlmmfufC7GEHW
L0D/TQmw0oWYB/xo/2R6k2SvIBfKsvuFqX3C0xC8qdZ00LdxZ8KE9rKx8/x7cglDqyF9XUoSXTFF
jRvjcu8zxsWg43MOBkLu7g4hXZWJwxtoNzjF2ptkW3lyGhMV1bITLQpNtru3DlJW/SpyGKGJi89E
7ax/ChuNIzSY5hQT0GGBZJhShwIwV9yALupIjM8e+1NoXUsudK8QoADcTvD33AMmBBfEz2hgxWoi
X1QF56ixc3SCI3fy6T/+YB5hDXWfjejXc86Jpc+9Chue8ITa9BTwK1+PD3zV1VEffVuLoJhGczm2
tBoJwsI9BrKdsr0h5xWP7jj5ASeZOOTP4gA77L/sTXdd6HRqA/yoMGr1EUP0btS+ryjFxEc+hgRM
tL4DdJgwO1pvPeAEfCSH6kdTiqZsjXYF1RIWxLSMGP2L4Q20LPyI6/84gwL6s9KgeXTiyumPahyG
zH9ovOMLDHN8YUecBA+PSSAXlF9SXYpPQRnUIQh3P4ILk7Z5qpSIPJmtBootkDsa776ewvFVdF8H
KOPsA3oFdPKv08Stpls+cJXcdSCW3MjZp/bp8sPyRsZKvC0IBbFdh5BmOa8dgSYJe2+b2LPTS1bP
2sGpPNEASqwdtNzScwzAMeGCEnCnFQsCi+ivV7SNaA+pAKgVE/4cq7JlBOUKCwQ2KmY2ap9EP4PL
kmfUUbpkVoKbK48dsKITa46MR0TLOiKM3qGBM20uTXO5AqLc5K/JzKxqEO953yW3wPJ3vELhI4XA
56X/+cYqWcvwItzjBMQS/yxxrlv2YXz9emkqhgT0G6f8DmZi7NqDXvCH+WP0+TQfmqUvF/1XI0Bb
YJLJym8393LYVrl12DFB1KpM9rSU45Vp5GSd8UW/a07QF+ucfwSUf7FA31AxVw33RBNfWSIiRep5
DjX1Aid9B68p2HaptGrmYJzGlV4HZWXksS5fTg5RflpB+mfEaQZz2O8dpBFP950ecCNxDUbpsr35
zs+eS1oY90R2krjQV+wHVUpGrqViEf7AErN3cQjgAY5pUrII2NpBUe+nkISDyLiNH3lhzfA/8NIt
yZsgPJ915BGo0Jy/l5qQa24kTNH2nOQMiD4Z8o4ZO7le0m8SpgeamIwi9NGj6DAYxFe+DoPwT6FR
afltqItaHQsJ1cBEIgIlYGwyCc3JWodg2kInu3iZllCYWo1uGLHii/jYXlvzYHy/FMuHxMHxEqfA
vue+jaiiLy8vljfAY1BxUKmgUPDB45IXUznXo9BUFNfKTPzs7k1+Ww1muCw0fs0rBh+bZlVfAI2G
uK1V/RfbEW04B0Bd7pQG7OYbRH7McdaLM3+jAq0dXfLAlHoskD/P4Nd1iQVQwBNMKBnFkALSc7C2
jeM2m7USx62G0PMUkMI0P5L+crdpUZlsBAZZwYIfjtM7EzUicM4c1/cw/oaZqORZxsFkJ+JipzeD
dX74in4EQ6v1QGiUX7tD2qBN030NZbJg1CS6Kv7/1JLPQHlqXbFO9fgCs7gpG1hMw+2dg0DbQdYE
DX3rIOxJ+3mBxEfApi1LbOrBEmsO2ol1Z1N09bHrmB3hAurP61zxpfD2RmFxx7rL5IxICZ2G/N75
u49VoPlYWCOIcMM33idh93ZFZVrf8iNlkaRvR49/ymQN48G8mEbPWKEmxa0acxE/hRV9iyCnF/6j
gDRcGxeikMZxfRkP7FkAW1XeSjflazI4ANTRoSLNh7BY8Qv9dmla6O/nkcuEl0hso2X9Vhfwoic1
jFHyc+eFyA5uyfbZsnmWCtAhpXQWsUkQItr7wXg7e+Mw3UdFFE+ZG3Ih1zv/JS45jccYFHSbX+PV
bVyzVqglAE+NgIsCweeq3geR+r5FJKZl3aBz8vC6clSa0e/30E5qJOoGNC8zRJ2eQbqbK3TVO9he
sSBzwN2RJBbBkX2mk1f5rS8Dc9HAi2gfiPoiOPO4dg6W2kUNp1DrDBshM0AXQ12RNOy1DbufUEgD
Fh/F8AoT5qLkII23ZUVzyi6bpQKrbTvHqRl+MFY1SPsY3OoYQe8liQ/tt8ntp5tvSvZaw0zasJw/
gOKswe0YbuXu7OJxSiA6CJo+46eBkfAvnN+jWCWWmPlHk+e61FD8hWxsEWAif2aRSF9hKQnGTwjr
Y9s9LvSoCG977WWiLQaPXuwV0bbzZaiRRhKjB9JZT1AiT9p3MN1QXR6H57NXwvjnQrKu9wUBOaH+
L9cMmX1V2wBHbVHXgB5GWWhhM1vpNarb2GkgHLTyyFl5F9QtDvrZIPJOGO5EiCKaCPDQWqBzixLl
gdNhTwxyvFVRvg/eTpvv9LjizpZrHFoktrFmYYXoGf/T9tRafNKpxd1NlX+QgV15urLxINAzo4jM
umyinTQrR4HHkJwUH2WnQH8+cSyKzlnsnxzHZiE4HaHM0yOtTnUjx233WgqJnuOcWs8WSAWY1m4w
Fcmk3xYr9pgaXO1roxCiYqD/MrpIpI+fq1KMylsaB7so3UVarlba7qevXBKzUKts4iHxoXbdJxkw
5CqtiIMRKSl5wx9pDqfZdfPati7llDePdW0R+/TqWHrfrZvr9XkS8mIShur8Q82/+HCeW6ekjStR
q2FabQE+Iaph7r/rlmySP3qx/xAhecDiL+K7A5r9+/n3wUULoeOeHvgAlYLXQf1Oth1uvfDGU8VS
j+4RdVOym8SROIf9R+x0P92plNl/qyUwU/kZ4VvwmfiaTaJF8faO6AJqH8uq8ocn6wbbs3Sm7psQ
YbLZF17dWCO7Kuv2CDfiVYUvBTZO7QltooIswuRQf1FjKl+Q97H3Ba+7VvGNZwddR5Sg6Bui60qY
AQx+cBlljHmZXGGQhB4wQVIHYvNGCrAgd34KntaI/wHJ2Ljdvz4vHMvWAdED+Lvm1lr1herJfEp6
o6oTayriLu1FiwQVkImEu4vGzHfPNwNsyQGv5o1gAlpQB3jQCDmFke1b9kCtKIZNGf38F2+LqdGT
+5M2Vug74OHI/6lKB8giQteOSpewdWi2nR1tzEcprkxBm9kC+hwGoDNX+ggBuFuFN6DkdGWXrN6q
TUdonOd9KoeBhLplUbm4S9E1cEeuDUjcfzOshcv4nAkwXpaLh/2sgNuiTajQyYTK9I1AeI6fiiSC
Pm1gcagJ8fUwPceOlp5jg0RkryYqUIFMHgum3jA+M2Y/K54n9jC79Mqy2Q9imYx3FzyC7Bj+SW0+
7J1x0WGNuvMD5T0yFA7ElWPbfy1DFh/+aHJTWnzsTN9CqMfupcwOKVjgcfydN6bJG95NCV82GjKS
MyEm+8Tnjpki+RclQYZJGnlbWkLk6aGq1UhHGgVOdD1WFvWxQv84pGsH13F0EVYo+z4ulti+glry
J/PWjAb410oN/LOWD6nv3uijkjxCtmts+iPOKM8jaJgsdHUvTL4JULJYM3xX0vTgzJJa2jLrEMFJ
t0mdCEbHK22XaavpEEw+JPt/+qxZ4wxodlXDDQD3sDAEquYwS/RMaolzb+18zy6eNt03SrEgWRJI
G+nfiKS5EekF9R8VUfwQpfGTBUUuz7DIVU+rVgEAaKmm3pveUAXscN+7vForgQELk9PDED+pSJaD
tdPkIthlerboTHBouP3RXyT4wpC7enKHDyKY97qLn+PFi0nCfbrgCBiIjKnGPgdSEzAZa+fR8GP1
YFT1/LprTNL3nK4exL1nW6uhMY0ipFLX9X0i34pLvz0FJHpDYBuXoHTdft0BAj01EjxdC+S7/Nrj
rNbxPI0Alx9c3dD0yOWMchg77CdlG+OVCiSf1ClujOx4iurq92aP4bMVReMvsST3veSWEFBLNlNa
EisB5U7hLqHK4bBjOYt4rkscSuFxuBwrmMIsxjGfCTQC4yu3QNs1JYrb5RGgYzdNkP7QkuXTxz4v
J73776nXbF05jsw0R6cZR1nhiRsJoMZT1P/S5QuVTQ0s3EH0B1aR/0c/H4LbZGsT9XM2rRi3IBxE
2xgh9DGrJFhgJar5p8+kwEXjSzRsHNoGEB/OG7/E54f8H5Hz2+impeOv5cysKjMhO2/pzehjpAdO
2kH4q3rSt+sYNxehe5knC8AplmYZDF0nq3DtU/mvgzO/EhkDKfuQe9lUk1i709O8HoyyQQddDqw+
yfHK2O134zgK7zH62SMxXtzrNBWI7Q88m3L/1i+TwDynWuRQRqgYcuzLqGx75Y/PSFLJiMIut/+u
HA4XfDCAZ58IAd3LCyn1D9atuAHQOi0Aqs6ol1np8QfPcXvJXjWtcpDdEQUzXrV2mpeKfdpjOGOJ
n4W/FFOcP98F+itRka4Z2m62XPtiio29PXsyENAv805PUihgkjEA/Q++gWcM1/iKC8d2IvgfjrK3
Q/D6wAPDLpN2bLUwdK0mR6SygpODeddfPHjpwexaPtj4xAzcIlwNP4xxXHAT8/OAsd2kOczQk11O
59lrkPNePypU2QOgl0KO8UBGyV+XxQa1GT2xoUxGPnc40QnhyYyc1vulpCj5Tdrmhio9UM8qeFBb
D2PbNsC15I3N+WOzJ4l92w7peZN9aNsw0JFkP5X6EPg0rNXWtFjj7QnxdCQcvzbA/ex5vkKUnlgA
R1uJoIcMMncfMQ57LwMQMaTYfBvdAo/kj1fjAPQuiK1Dcyyosu3ozUUigduePPrjLZKsboOXxx7d
5KqBP9rs1U7UZXSVWfz7YYtCDXXt2W+dyC9qXhdQ6U9PwP3cGWxH8B8JjqK0DZPOCJ9DRG08uQMo
uCHArpnHjoJ895DBpeIx7NF8OUD4kgbZfrgHg0cUaXrsdAuYoGOml9HAt38XnnMmuT0r/ZGkHONC
ANKb7XqZF3ow3eCnTK3pewsNb0S5qmTPyEDdjBYNqJsA9E3NUcdx4TnMdf+5UtWD9LWIWxoQFkDW
dSNdxD7velRs+/uMSz2xUlyeLUZUOPbUFoH8AhUwVJX1AKtaAxurjQ7DaljBay7s2UnLpAJZTat1
OZeNxvECIpRD4UDF0qiMwfPVSlq47/WNJdcPqdPdInU7GmjCT+8E720e3BBZ9xQ7R5yCT1dsvPiJ
VC2Bcsh+cAgzWO+o0b5aiu2culxoAKkBz8v++0rsHJP8t422lMTDTeZtKW7D8j1cf2X9w58k11yy
cVRzGRuEIScgpHjYgP9FCDVNLZQiKfMJtQi7P6T6DSBf44n/OnXtuUsxe6swnzpHycyQYzJJ5Vma
ffG2Ee/lMtMKR7mWKIKLYinf2nuXyk1agS9mSSzyT+cL/GPkp9cutbLzahC26O9Lc6AWBqA/vXVh
kDeXuNjyFyPZMNSIxeK52U14UlEA5+XLFZ3fvgfts+WIMO+X2AKv4H5Zz3HuWMLWBx00+QdWYBc1
pGKE5rz1rRBqwplDymjY4MHebESsvOdPN785EBir1aqHzoP29Aodpkim8B44UvJk57grhVZ0YrvW
o6Acn/xHqvyuWROuUSjA5hIYscCSMWHh5JT6w5Zd+4D2Ni9nezGqRi8QBVYEkAzp20acMibuhTYf
a3zh1mSoyVD9R26DPKYO6MH6xL0suW0BgPlBiBO1MCXKQz9Y9C3fk1l2GNcET/Mx2DUe237wGSgd
XafHPkgd3YqLi6nyjZ2nD06B5F83s/a/wqCguw5+aZX+PRAeWz85t6fhLZs/DOxY6E0FrPayvJce
gaop5hCQl0qkDGTDI8WCUV+Y7luBsXsDMDrjBVVIbuINFMUfdnQbFGnCSzYF9A7QUmvnN/qDrDsm
WXMIe2qN7F4IKK9or4nHCqhzUj6ethcekOiBYnDo+6lQ3EW2L8KejCXENTctMb8/aTmkg7T11CQZ
HQMsPvMnbuibBNJ6MNBqnIPdXCRVKhE4oFoGdoLKmwEq9FqioNXpeNsQJE9eUyTjBGukfI+AWy1Q
cQsd+QJ/jQKKF3rkfyEAeCt9Ds0IJd+h06gDUi80kltTF+hDB7qUhxS1nyz1pVAaLIhtQYIUGizf
dB7j2bbSaViyF3HDGmfaz+o9IQas8MlGSAcZ7YZdPIZNG7MRuevpCdTN7aYhQr/qHwa9ZNkKkK7N
J7JbvWOqRdWaQxNTlSeMOg9vn7vI6BCORR58Vrn86bHlqDTfjhRJNunajnUvjguNcBqDAqBew/gm
I8Y8JGsjD9HTU1IKQGpA4mrkwBdK95IUsmHnllbIFvekn+lXR7N6R5h+98wUkF3ogGJ+UUkdjd9z
DX47LC1JZTmWraHc7Fg8tN4IhsnqM9ZK1D9G8sEs1pQg/kz0fYm0kxnQIM9SwREZGWIwWKX9Wlvo
1Q8b6fpbw4SEFdWpi6scMaYdInMUXMwxDb1dpGZS0RGKTauDRbBL0hdu+TNzT/x1oXCoCwJ362CR
m6qDPfD1YDzq5JhO8N489pZ0OvFf5XkVwo+AizCqSkZX8LUKkJv/zv8LPomfdzTvP4/hz5b4rsBH
cmCFmhPD5vUJ61yEZQaRA98ebkG6grC3XsyKF1w0jsDQ/3oOSP/vqC3lViFYiJd9e0FdCxobgrsv
wFGnvZgr6FwEUqxMUh+zUMqhQT6RsnwbYYhf+mirG1TI0NHdMM3xe3KDdC9of9kWpdimP5ssYPwp
IS6Z9zkQn5HJihQjqwRs7U84QDLoBeec016aXSleNKKMzzgyp4Ce1irGNw6rMKaOJnxXZvTrTwdw
8TH/BnW3n8bEVrJUimarIb8PPdyJHRU8FuQ9qqrQeb2qh96bhKTKPsPNvtY508WsQBNEgvSyXDe/
gzAh2Gz9iW8KggbFSu/oIAJMDF+0pdd48SRzvSfyoX92CSsLltVgxgacLM2hQoo2COnj8KYE3I28
xfTy+cBQMswXb70Sym3dDmtOHioMvzTWKqdF+oIVDVM+0TgtecB/QiEJOnGP4SBOJyvrvJCWhKgo
I6mlH7V6evp5MNPV7pD8AJ2JQf5x+Umwq/5aP8Ex1bV1FBHzzjxwiJUS9H0y5VpKVJBeDw33M2lj
4Op7GGmESTWJxfhg05y5L982MNBM8boXXh38xrLuLBzVNklrDw8nymodzQIdzYyh9pazOcOQBC8J
9mX4C3faLl/M5K6yZh1KJRd17+diZQjcE/cKwd6iuGW1NJKBT62AL7Hk1FCyyRYC/HOjyAkLgBy0
p63hofvJOHs+gB5ltmXsZvG7luJIRNAFRVHBQQGt3xiM0qpzrjR8H6gzNMzOyOcVqs8xCf+vTxch
C9Y+CVQ549UnSSPpkaxkB8LvS8lrwhRfcqPxz6p/5fWJjOyCVXwxotM5q8lVLbE3E7iiEWOKRykr
0MJwViTD1q8e+e3qttWKhX7ZSGtHsQjpWtrergxoLTQq/cW66i7GFGboW62k8e10cOl21iQWYdxt
csIOfhwmLfdCIKkT/du2/PNUaMLhXJUn+hdNaN+/DQ30Cee5XXFx4sCxAgX3YhXiyI5wRhh5zOe3
48Qtq3vC9yfxDOU/+NJ8vY0JBvWe3++wLf5XfVwvsiwJKDakbx69fdYeXRmGzqjrp4mYstNmMMxM
oTFqHM1Bjs2BCmjMYgpEc4CoqbZ6/xDsGRsKj/3fOAP43sqvTFvdi9rCYRlmnYBhxKXUlzgle/+Y
xKOgKPBerId9GZMDpI6blmGo0C4y77++WdC2XppJiWxeTjsRf/uf+vTPbSYUboTDt1D8EAwf2eKe
Ok4lE4hTXL7r2XeiLjYe52AIvrO4yUNN0Tj4yTRqlhE9QwvbcbQN7SnFdM7B3vLMPt9NTnoYDDdX
prKxLHMfu6ggzrTE07IxAUgC0dmRc/l5hLmkhDzeM2XYFviYAeqt0vNxiV4eD9llPI7CxxQVPl8H
TXvNElo06+k+erqJcbbA7SmLBaEVHffQp1FqF1Z5sRMyQ5lrzGCzZABqaAGYarfReuj/hpS7UjJl
cdP/mqDrwvIVye/V+7fBAEBH2VUlDiRGJFewsaXQQBxTQ5kXjRPSHlfjt0jFBpuEASJ3kvGvUTzQ
9oamx11aXfJ+Z/N4UYxhggWsKJOfopG0kuOq5JtGMEteyaV1c3qm7SVretVzakJ8HLUdVcKlfpeL
rfjyZlZwHFvn8mk+q+SiWL7Usvc8uU1I87nVkPUjZfPafNn+aZC4xWBIjcmeYg5cMryBQSbVbUGo
I+9WPxPQglOw0fvUNL8CVKXOILZOpVDtCc+6kO0XB34Uq1CWEd/bycV7+aCbKN/k66biI7C/4Nj9
WXyOfh0gqVB7Edb6eSe2Z3pGxeGeMJApmA8m5tmLsQCsxKc9sE9YrRWl6fgdRh3vfMXW6Hc0Q7CZ
sVhk3iRO9dwciyZL4QV0dTbgd0kYNXvb8fWzBRfaBbZgEtgrWY/4C+CZfDfaJEuKtES045/JobEZ
baEFCRfy44G7y5P15gk7xpcpYMtkxiAOKKsm+OnxcvheoNM7EBMSwVth65EeLX13qQKpON5kfm9N
fVMnVFyr4X6+wHd4oDxYcUmKzmqVVG0mKW9YHN/rvZkGmVJCbKPe/fdcwJBGgxWF0ZUmYRByJFtB
rTX8kuvUDvEwmgA9gIYo/pJcLOAB4/ElX4pJUTGNJJWR6SyN6XIE4E19Vuwl0QKujaCU0721xxbf
+IuRZ4jsm8D+cxyGUzXTHniRkOFoBdfFad0L0zRaIK0giqnxTojBUvLwvbYu6Rd0eHzfhdmzXxXJ
C3oMGQcFlx0dzkhugdZ4y+MrbK/V1sZSB81qtIuTSlGN1cbrk3WGiNfbwq3IP7YFKL976751YMR2
zlQU0OAu5w/QXdWndVGzGmN51T79x9Q1LfP5QmQNgMWohEy1TPLibaE1a3X6LUv4kBuGkjqP6lgK
Hi3MBQUzOVvEfSibUkaMsqXwVDgs3N5G+QdeQosoeTy7IIVhsX/A8B3lNQENhT+QGII++4+3Q4lV
kKHJY5AJ3xOCSj5dqO1BVtggA380Ia1OI/Nl8Icm7e3Wvy7xkOZXJ18wH//T8OHT1lfLWRoBo+7G
E40xdcZDNijFWoop+Eq75v2hzO0w7qKK8ACaNQRniWyI2m0xfph2bWAu+V1CbQ5PUsG0s9OstG1Y
K8Q8pyMysuguEGomzvupaRnNwAo9pKaENnQJ+wkqUpLP3uvYOzjSDDlMyXAF2xQUbgNZ4FVfEzZS
VpOLKcbFdjrxUr/wbvRNMMwOQItwXvdjn3TOgnGescY/ZZb1Dp3ZdztGias+snls0dDwJrN230tt
PwV2e306Bs2Q+R/K0gHcC4BrlPfUab0IaAvkA9Ic517vidTGsPhOmqqVmXf33XzsSpzp0ZT6wTbX
WRUus3VMlfzaJkFZKhPYHLRy/is7aK9/Tw83ojUdQmPflVPr1OyOCpPOhdzZPvYBUmjdDvFtDcHP
AE36NzlMQPQ9qfx9SePZXZ/S1Dn/Ec32PX8L7sGT5ZiBGFrFvakhTnum9zRA8JkZ8Kg7FyVpD2X3
xmZKFoRodnihxZD9HUtW+N5Wmi4XEvD0ptLVZWOW7O+M1YVZId7ETrGtdoMmpXMkg5eyjs/8bnku
VHrJh2ZxOWqTPYXNHKNY2GQyrDueNGW4krwPexAtsC9S/u4mkpFhBV10TiSUAxIDPUxTbaRopd49
v1NWwOjl3i/O9wCFW4QE4wiChKITjKXqtcT0jT2USxX89yYSOeL8cl/9Q2Zm9A6X/HJjsjetty7b
ehs31711e+qawwfJJeHzPj0ig30UeAs14mMjreIyUQMl7UYNgg1aUzF5hTH4HvqPoJmVfUkpTiTE
sGjbdHXpgoMIpNgMl4GrQX5k/hpdFo5rozmznobjPABbBCJCUMY5LL2URPweQp1sbV7YjnXoTiW1
JhK10BCx9iOu9k+89Eqdwa88GBVNdN+kfwGsLFsLgkK/h1aPnZIZcIoXzybbE3QgoP8i2Q28z/BK
efdXrOMvll8pCMfrXpxCyfNb5emLURBYHQCuTlYeD5iH7gAaZG/qs0SNMXcGFiDFL9l5+1pN0xmD
NUBw3me9CKxV4vBGM6C7/n8+KT0CQdvlTaMswZQbbLXkHFIGz4J3cyhq8mCRaPFoMpdgjUTtkHcc
3/Z/w83nWoyHCt9zAfBo+xevtA5ON4SUdmX6JLHyQho5fd9gQY9cqit1KfbLhKw7XMk+YJTbuoW2
AhUBIWYruve04CR3QmJ70vTZlY92g0TGzHrebDvWbMLA2lDIVRhvWPr9hP/i1uuMTv7Q8VEFbxxZ
1A0GhPXg9rctee7CYWQzeQyMsWNsEomjRG1hMvNzhy4SFA0XMai/Y8TBB8ifFV2F2PJW6UdV1gzu
/BmxlOjN3Vm+DiSXbm67owyT4W7n/6yGkB/gYB3fRalNWc2Dg/WtYdKCEpQxKNG4b84mPi4rQX8M
yfUCp5QZ+VySMJSS7yYN/kiGMTDScNTNrk5809VrFsSVk4jOHD225JWTbTDZPpqUi0mOM34Jl0It
GqTHPhSPqWZSmaeWeajrYPnwFNem/d6vAJc1ZjOA4kkGeBhdghcB4FMD69V4xZxXW3BqgW4OErzd
0ir9oiUPr74CYmni3fb4/VwFsZlKzbylx+nOPdtaMV9LVsfWhLUlcO3NJUBFk4DH2yvTCHAhdLgp
W0HMv/o/eqfk0w1/TAMkl5NdXZD1BgwcYIXnTxo5H2yMy5ilHvm/xzSoNMNXQE9hLuGSZhwnURcm
vrUht8S67Q5oIp1ei1+/1ZhOJj0E8cWqiFg4bv4njsTLLIlBSkvhKVypkronoMQ3e+Zq+3heD1vK
7Xx7Shjo7PSTTfmw+yO2+WLcoBwyu7L23UX5t/WVc+/LCtHWocXgGzjwPYbO/6Dd7GcYX64cvf9r
H71xbm5AK1J8hNFsMgw7I7x0I560MXw8M1RNaOhc1M0PqxiPaOQ98f8e7CQHZsIf23QFWoqedg2d
lDNsBRFYEGyHBk6CPnpNDUFfgBkwr8FUMgaoV3rmP3SVIM59KG/OLNrNqsLxtKmOSjsRacRut9G6
8FXcVLMJt1y5w09infEwIaVf8bcowniQBBRUKh8yIe0KIm79iCZiWxUH7m8jkwAli1kActdVXEOM
+i7C34tFATwZoH1wovq6x+kqGXrgg495i7ngsSpqt4rmB4BXGO+eUTbFJV32avWmf+1HbN08ZDs7
ftWcMKFQS9yfMPQbF9eyvRbypsuhDTTDovUXqB2GVTKehF8vFi0db5Wf4ZEVIndNaXyHHqvMWRM9
klWDNwNcnDl2J0YXQ5y/t5QcmtMZVTCWzrHlNwO/AI4PvhigQKw+jM8VgKYIcfMdGEIEVR8iJ86l
mr0tpchkMy8Gd/tALi+eczx7OVvaUVcZme0c+zit+Tl1h1bCnrom6LQ08fqXaGvOalCNCeIhnt0t
+Iqo04sxbkOsfZj+xF0dQbHa3Y1x08Z46GKq8+5O8JdaHjklZ/1wDzycRvW6ze8pf4Iq1xDY4Pb1
iYJzh2lJ2Xi7e/S0L85GjaYrBOSyxwHKtuAG1ZlgZm7SDG5+cN1YMryM4liKWRtAEB3/a1q8hQSK
CXIgXqwxU3HfRF5ZqwU3Z4n7+QMJmDVdFGoMndH+4aLDa3FSygYvb6Y8nW1hbzHUhwDn7lQTpG1n
cvB4ubEZ+n4DiD/+UQeN9VxRNwAz8t90VX3THDfl+KYHMaDyAC39MCXDPlIjPBcbtKO87ghf2EAk
CIb8tstqdX9wvv+rw1E5QDKfGFXlhzpoucyflw+hv1XRaS2EO8xjpN3DuP7VatME+admGF8cQfvx
PhT08vP6bO+5VxTc+A4OUJAPzI4d7xatGowSEH4CmGqLEjLZZKpMfjmBcHeeu7sKRP8679nfT6T3
DGpf0kfsVYitGNuux3Fcml/bLrvt7gWp4mqjFvC0/+VwaqkSTZ2ZmHHE1CwN7Y9O4QXEWQz4gI/v
M51rlXGzS6ORZ0ekLMmu0Pjp+H5qqHDD47RoOeqgypbAgwxame4NnRFhPH2UMG+5G27f4vVdUyF5
S0mXXlGO31qPYivbAiMqGeixg5pjbOTu/dl9NJDa4LKuCSvnMBbG7hnlRIIpID9Rd2ztC2yDiozh
UENGTGuE1HGOXdJlZYR/qXZ/FwYoki6LpQ9b7XRzb0LV/9mFt0CB8bgPy61F+fH96zY9O0wAis51
ZqfKJyx3X9VNExa8PYy81dkBWgIjOpqWUFU4JVas4wlqT3FS0qRnrSzO3axn/RiC1lSf0FV8/xfb
FTTnb08qF/GpFW9b75wai/8/m3ujh+8cgBfOKJvRtZeZQrYF0C5wJ/edhXuujiRIkN9Eet8nfAr7
/yGiv7VpSuIXJfLCNMJp9K86U/KI0BOqwXYM/3vbFhuss352zbpuy48XkxMujWxqX1PxFC5FX8b1
tNilTdZGLBRTXn6HRMNyR+d5J4xS7HbZlDZeLBHirzT8Gygn29jHIvoYv1sJhiCUY0kGRtUwK2qR
2dedOr46uTUafz7nIYirJEUn1UkZCwoB71mMMAGmRXUKAFV0Te+24xB7r35X/mGAzgRaQFzmbCcH
Q7+TInAKt7r/p3019htBQ987oRLT6djGYqXJnSBRCfvstqHNeJaYCdU1v2lWegJR4cKx5yRMhJ4o
sRHBldKt55J5bUL5cocWq4bJpGYzY7wc9d4ASks9T4z1eNXB2sIe5TabPEOdvZQKlNuak93Q91+i
8CfK3pt6aCP6szM2SBYyuqHTNjRcmTk955OaeLj9bUqQIQmVbX5DgQ4oY8woTKj1mx7l3zUQ5PfA
oe+bNVqMChm4lJ2akvNhbvFUWyT8IIXPdv/07q3M//JWFrdGCErMywHcNWRzDrgw2y01IWmiBADY
XuYyYK2N3dgs5zZegnb/uKWsSs7cj+WK2TbLJpKO4To+Gnk11MHCPTbNIcCzNhQCbcWiyzVmIAZ4
cFzUfsitWMdCp3czGLzjOW8tQA5UE1hXQQeinoJthKZcopPuM8RvmyKmldb93Ahh9jkVLORl8NNq
nNuC6qjzGFtShtmfTXq1pfLl1mXbdlm4p+vvfw7nDR7pCA6mqZga+/SahrUsYCnHFJ8yNpLNJyG8
UXhnUMhgeQk+2dwumedGGZNlhTmOrZafj47jYMhaOjVwCUBibmB8IbKDadtucXBvmCEfE03wXaGm
gZUGcvD1Zdt00KIz+z2Z4ntYmBstnSl2BcVD1werTRDNlONU2XR9mWN/62KvuDmPaXKWi0PDBHLF
ddKoGp+i4Z31BXyA9/jxACi8YvWe+qjI1j/Da9zSbSqdowOc96AmRdWMKd+R39OmOXEA+jeirr30
io+iSHjbPywbYm93MQ9fvC/QgV9NrQ8Dn6xv7xNZST+iH3vhGD4ZBmeEygsZLMrCg1/jxA9soW85
pn7OmgUpvrZFP9p2dLhgcvJqcrBnsWBKtGbMK3M3I9lF9fCCjPcKdf845sl1bIVQQsYx9ajcOLLa
Atthed3nA+v3lDjwoj2VCgZs5BFM8Z4Fu8RA7pqhLGqu2xfJhh7O0S8RJiK4SPRCYXu2CFc+owdV
yrGn8bXGs9r1JbYPRrsEdWo4OYm/E9aDABxVt5cWE5ITko8fD9nQTNu+tnfb9pTqQ35i5ltIU2rJ
kw5MbPxzWqhmiGdO4K0I21evqsr0OpsMrf4myLakbsrxR2n+Mvk1SfpiXXst+SsbO7djnnTaLlUk
v04u3YB9ErinnqTHSaLumJxpH7ajv2AaWXQm/j6+IFsx03pG56t8fTkhKrLAbmVU9N0nxTcYJeHY
e9+F6oFCi1q15ouxE8y8CmpVLnFbduwWAmRL07GVW4QQZcMblYei3CY/hGolp1G7EdwIAqd6LAeV
eSSotXyVtz8XGJ4OK1no894LaI3oOdOcBojau1RdoF7qQtuNW38f+NDYDGHC/lLBl4JV11nEfGOi
MgkHh9Yl6ChMCLW0JZOPNiEwv1qHPAnyjrJKdMTdjlZ+WI+ApUVE7PdbEFDqwZHcmpqcklSwN51e
izvgB5KxI/fQmuSJTJ5JX0Zq9DFggZhoW8g1dgu5+0vzMRbCSL13QqeAIEoGH1JEq8olOXq73+5v
40l6flr2ILI+w7Hbta110yHhCmgZhTFQgJnskOdswR3xYqKf83Bz2tlRKu6iwWWWFH+MjHLGH8MA
OCFHQHu1JjeCp9RHePP4vk9cwBLvBDoXzTux8rxyTdVkxBdqcWwQiZPmILyfqqgkmW/gHvnaYw7F
Qyc91Yp3agjLf9s1ED/zjoU1hkntMSWAoSSEA2jLto5aQ3eBQq5gjcw305ZmgMgYEZ0hAveCIwIB
9fW/EN8IYYR1zwwO1K/ooa5Sbvda4Y4l97bxUqL0FoVXx6BlZ3mqMMuTUcQguYQoE/do3wLQpDK2
0Xu+inf8rbag9hXtQz83SLmrBrbhr4gh07Kjc7JVm3M3F4saIQUx0WVgOgl0SK9nJiWDo1uB5yUc
bs18bcC4vDeoMsNSvMQTrfiSA2dIBkR/nJxI2ArpoECPuJ18pbabUjDiJ7xvSR+RrcklCN8oNRcw
vGM363bX48ZUZ2VY4XdxzssdZgAfpdJBSLlIcl+NqwYq2A8ejf6ZVw67INoB/HK4TcAmamqO7le8
lN0JU3h0ONt5aJeoBYk7MIPhOucHKw49jf7S+j9bCLbLOF7FdjALPPxeOCrGedW90JsBi5sd/J6a
igJFgV7O4QIBTY4QJZZrq44VT995YoZbZvvmI3+cy6yXXaK1OchsO98S8sKKfu7UoCipZy7YZtBI
44rHGhGiWg9FwC7QDFHQVs//b7yN4rRQxxyUeDDpLnbxpjhjg5WRm4G7wAdDl+eyqlJoyTCbFVwO
rmfn6Gye9TwqnNyJ5f3HzzyKVWoMKzUF3TQxq9UyC72T+ycEeLSdfFucvxyFfvI96/rZ7O8IRFRA
818qaPwdoTIygISja3BnpH8/OiZR7POdzjMmJaQQbSlNSICMeLHTf18Mt7FNjf/P6ke1LHSsd+8t
bhz26MrPOi4O6O/PIbG2Gy5iLNHXj/QN2vIZdWTedwO/R3THpraG5cUXmhHvcOWc8fnMEbvSVhSo
qMjR3pjDFRrBNzexDUjfnZaZl15v2GnwCq9UdBRLsmsi2ybLbOKIZwr+EwMD3VGong+pMKCsJKEd
6Lu5fmXu3NaPgT6TNZD1bqng38p9L7uPTztkhJzV7BUqFBBbRWP0xd/ZVttaWHD4ObFyqWjN4/9N
MF95rS4aV1YVKOjoUnWDtz8KD9owUD8ETMngoXIuPn85xgfAzBlQ6wzZsQM67JXx7li+PdG7i8ti
0fBorJU1uQpZQfc2kn2q89y63aZ8aAHXZOi3lEH4bRhD6tH9qLqazteygm6mGpRS+8v2y3SDCO8t
3ANRXQgkAEbt3o2u+7H5r36eSC9HRzQDsTdYDmHhJ6dlJ2zYGtKci6cl1b0Cmv7XnAAHVxL62oKr
QPoXedTDAXalSRLRbMyZqJ0398WsN+FkXAENQlynMX0QPN8UwrXOog6EESDQN7SmsKsGKeQ3m8Eh
FA9/3wt1YUnYpt4pdYNJWCqjx+oj2Jq/hZZk+Pg7SGjNQeFLPxmR9g0TrgF1qVyiIkBhS7UngSxp
qwV8zPkusLuly14EOccgANHkT7IBAyOeLMXyNxHjRE0hBemMGdD8RrucmqKRRxKrfQFZsDAMyCkH
6h/YunHWFZ9hbUFeMUnbkMlFKWWsbt3UqTCvO/EyQeEWF/+V2YlAIB9vM1oHUlBD5aTNmdE2H6Kj
QKRtbofwzVKDmuTQTyKY01MJD+NHFfxmdRNh1JazUPfq38jxPgvI7OciwzL5bGNu/h6uOAS4n2kZ
R4fE+a79n57aW7walZ1rPfNWTTnF4rujjmAnADXVkYAxF4ihQ50UUjB1NRqmWSTHEfqLu47IGUZR
cm6BNRjlW3NeZ38XEWWZ8vW5VqkKureFmcw+n08aPJXd696xSWGPzYzyvd3SaHllUFi4ac4Lb3sc
EKMbzfONaMgmfNGnFY6jsEqP5F3l/FmcS5cdo4KzkJMAjc6qTMSjzgrGdzxBLXfEmg9UKC6GZVaq
AXUUjdkxdl2HpjP4oeNfodgqG4GiE4LmgrwhMvd8JUwey1+yz29A+GI+hD4nEBUz1SkKi5OzOb8L
hftE9VsRXesbmUnsfsIarT+M4vRDnkxo7V5PrOs0stuEkzS14FW7Lbh4XmrsCXbrG3fJmyC6BSlz
9XeQ97kOWdyD+VjwRTlusk/G5ShUTEL4OvQEEAlsmEHYjgfr4vQz225TrQkKn6WLHDhsVmpqcKKn
rTt7Vf770qfnkj5OVpBrFKEfIID89nJoSiFTsjbKlJJ3wsuLtsH9hc26OPOlq5zTyfc7s0f7QIpa
u7Vui8e8nEgmblouNrzVLvJtPBbU2hAsbjFLrElI9wTcWzm3DiCHjWyAf9hhZhsIxUlNuiKp5zCw
UVkq+GJBFUaoT8r6Lvs7DcGse5Sd83f9dmkk34Do/C/soR8dZhP07Iob/i1SHD6zdNNU4XfD0zbH
lgbafOEvejrojCB640vYKpuoIRCdrfk0UaROso2IpzjqhzDbCB4YI7rqMZszCLKAgz0m4ggceE5I
/sRm+KEDpISwPDS25Zb5PC1M2GMlpTmhMhSUNPOead53s+h6ADnxfY02pko/UlL7Jq9Q5edxdzOf
0FlzTfl85+xSwfNDXcagTj8F2TQ61FMHJSM0Y/QGyOBHWhIt1nAXe/1Tm9R96Rr9Ifp/qp4JQCtL
G34HNYSITV0ayY1iA2Kk6lUDKxjAKaf9w6F9+9d4WyZxnID657AHyBdYlgL20fwOaMrulj+d/hj4
Edz2KoFGgqU94VaXEVy0e1v+jUZNWARDewrFxKdIIcfz0tqMKhidlDZ4/nEBAsoHczysHzqQR2Ew
/L3lw3IpefupKVhEy8P6cdhDBVU4XBzIsEqXE1NpC8Lkl1fJ1gui10Wa6DHuXZfVW5wQIWAhRH6I
AJ+9CKzxoPcnGF7pCFctKlfVE2k3nZCfmQcBuVA3OIbOu+A6AK+0Is6SgJXvpy/LHmmFQzdyt9Bj
X3zy3CMiFUNrPVD1bNvdWhblzrbqkMwhYko1k+Mxock7RhqTqMMYfyfkz3wlqNrxdpoBBnwf8Wa7
UENfbj+5wsfCCfOChX48b3f4UDdcCrV8JkivGX/I3eHn1J2xGpL6q4aMoPHNmB99y1TsEcJYCFn2
5p110gqyjPwSB38gtcB2Bn92ZDVJUJvARj4TLkQD+Da1GGIchmRxrbMtJhEmkhu8Drsk6L99Mb1j
iN3miLsKEWfOTC3xhmIgIQefYbZfs0GROvNRiFwz6DCRpkbrOyOlsuPIjoCBmABgKiFhAuV4aMUs
WjMni3WrG4Zo93OVrvyL/frQldYgLz2l1HptLty5eTI8YfK7h5xwmHFB6DCQz+RYsx76d5bPW6Hi
AZ7110Vmf6uAJ/vuPu7atM2vQpPJDDYwbfrWUzxk0vS2iuaWiJb+bQAHe0rmt2YBlKiDLzs3Eses
guUWpcsuXojgAX6Jycm8IGSgog5ulMdglIY/I0wqj/5U7mxM7SCaAjEVbDH9dZ6Vfh97wjey6E+P
xRu9KsTE8Rr8EsJPC+mTimOH+lg8jcdmYYp5j09+AAWp5piHz0objpMGB1pgjKRw6123DtY4So8L
07nD940GAY5GB5xPQAAADgm05sscGYZBBViURJPa/mqLfZ+ZFVt2WvNSkBWzvctu0FeF7hrHf/ye
yKZw0w5QcufjiDfPJCCTvy8npHAeUFXDjFJImEA88Ga70pi8yPOfzb6CgY7KWZu9WS+On5feIkms
lLk42uOYKrpAYDjkCPTlQr+w0uoUgL7yFcpgxDorBwbreBc+aa/evqyuxHCCGTNF1HbxQ8AjNCVP
r/y6h7AtbVbg4DcPFZXdbaVcWNiPyCgbkD/dQiURYE+c7jVeLMxYb/pwenJBA4czntK8kN2+IYlT
21CokL7inHlBf9+a8aFoZ7rsc0wZIeSSpyuBffCl+Ib+FZlyOPNCF/U7fzyIi1Vq06DjEsbYjuaa
D7/Q90TFrU1jFCL979KnAJOWS//cVhPuvsa8Vj1xlGM7d4MCi6018OEL2Va3NIvkNboFXFiPMWgp
ZIxRE1DNXoN0j//NNuxwigzwC71Rh82Sq55HJWGKyN0VNgQiZTFzsjZ6KZXMv/HmKhpcHt09dYMX
cAZ5pDhh71N05C/phdg8BCOZIojtNt6W9tHC9T5Dn2uy5+xTVCOpinWv2HTRM34z+Yg7X4xHBW+1
HR5ws4Jpyw+9kS6TCJTmKO4cwdYBZBQqg74v+V6dKQNUqFPrgQw/yBp1E0FdldCAevluE5lITBPH
uHzmf0RVKtqcqrI7PzPnCpuQB3g9R3EGB7mQ0pt22K46utyCAwXoBM0yIEe/iTNZQh+e/koZsFi1
QPLpBlD3D2dMiVbw4vRr075e1Wis1Om9eUUXeHC8XUs1t0ePf4Wu6zaxpB3380cQWp30BG/GMTgX
oRZa/K43kRPQIC07CwTvoudC1NuHH9HnWHXW2qFc7C7Owwbv5bFSv3Ux0VmZtD2NebEm/XFfk3GD
ereB6vzv34h7ojsC/IGiLzqcgU8w5QNHs6hX3f6yD+rAXYKijS1X4gQlfoDRpBCgRgPTPCdvePqA
XpvUdGmsQeDCYjePVR/CEfzpuMRs998hHVHRhHXz5vI07DRDVz1EAzXNZwGZ0Eh+Dl1xcXHjDqDA
hAL8TxQP+N7oF8+zEGD6t7OragU7nmb8mscgrMQrrHHm/Cp2vOme0W/x8uQszQHUJ4kHCZzgUrO1
yclHQ2dXU5x+tXUhBc5a4EmLQswmDheQx3vmdIjAsqDSfCd7OzdMDFKGM/X57vU03Ksq3LcnxWVQ
/Xe+EulCYQPIS8iqe73px2YTSV85SvNpiof++9slqUirMuFe01cF5OY+fEqYO67Pik6oPAEgKnjd
Vh4qpHVpx0P9tqjShdwAGk4w7P5aGC36pNtPpfmdZB64KkI1zCYn6zCCty9+zNOIZ8FEQgrq95ZS
02q5UwfQuh1V6suygCKdCYwHEv0oraBGfTwPVipeeggz4E9itl9iyqaDR8+n/JgFiv9m2WFxZ7/j
y/DWiay7JQRNxjPhzXT9fp9pfazfJmCFNBbx8DePBj3Tfhj9CzhBiiJv3iTsqhsB4rF0utifNNn2
oO+9izRXLvo320J/8whLAv5wyQOE5q5LBk6dLuYiABioPIXt1pSyydNWTh9Y+lUFUndK97ONgm6O
wnpnD0s05d4r8UFDcQb13Mjp1CTG+hzLKGQoE+GtvehE219hUWxYL6NiuHotAFYlJ9ozPuQMT0FN
ElGeunz6SqjT1yNQUojPNDDc/gXty/sCJ56m3Uqir7Q8SYyPoxgwL4I046ZC25ja0bKAFq6R+FIY
dsyKRHEmFuXVhWFqFicwymtvOf9d/IYS+5PA7h2Hbk4EhiYedO5bsatgnnCxon8zqR72Yq6vW8GL
nyli/g8mZ58VAMf0pRPROfg4a6o+3D00sroxKwtU1pXFy0O10oqDvAyXtazmE5uAIy1ks7SwuUhU
5q1FT1EQHSg85NY5YHJkp/5QHUD4bVofVNFyZq3bw8+S8YQvQ2EFND34JEAolRgkrr2bQU6EgR5T
aCmWZ5jgO9rzvJ27kDNm6ao20vdZep7sNOijmyBEn5GEbDuQb8oHVlNlvML80m5cI+w7ks7RLROG
swfe+mh2KUOccX1A9Z5WjxJkJlUpAtQ1EiftDjgIuMgVDPiojsxw2f2NkreQ8IUHzK00fqqDVvAh
VvU175nNAP6cCbr6+mH84mLHSgHPCLcuo4dY2wolKG57gk34O6G36tlQl3RueMz/FEFRgZ7KoGKh
U+bo5QafysHdGrgdvsbaXE7gMi3Sn1w635kgOz0q4Og8q+XN8lSo8SqSgRGwq07RR6X1zvRctoiE
Ww7oiiB/fRrEDf4/OSo0TSzR+mAY3G0qGt1y5LjUT9mWIwPGe3XxTTotkXkgH0sUc14+mhmp4aw5
Z9dQPOHhae3CaNlBHO9s6DY4D+jgUIflhyFoizGK7EtagaftAyBo9spMtOBOnBwgEp5FDWJAo/sy
sNiL6ZF/l1dxxQg1+7Eq57IIPIoZkkw1p5gYIYh0bZ85BmkCFwuG3AaUlSnAauD7R5sEYNXbXQ1E
Qpg3G/CMHc7wQkV4HFBKoZ1cAacu1UqzTx90xi8LsZPsnLc0ruPe5FSriaU6JngC6a4KpY7iPCLm
AtShJWdUbhqUHuKYCa0OeVwIzdDTjKTx7Thqz7859jlhwAOXjJeT3LbfPW/VpDF54mK/4xe134ga
+0tGRQeGCMaCifJg/QDBI7rjMXCUiUosogee4jQcK8uLD4mW+YCee7tXUHsJJ+t29yg2JdSivQQ3
Nx+F+iduJBAoOTN7xG09bue3EkNmoVAaBcHvAu7XvCSWwO4l1dKPUdm9wjQ81H/4KGSLplD05X71
2AVZZtlfmgsc0OsdLEJoXXXEIuxYJkFuhO1mq7K9luVcRqQfdztqa0Rog8gTy+xSgSPZbsJQ1fXd
IqcWoJ0+moh/3pjfofGrb4UxC9hGFNB2yGwpXtkpozUeKfEFfAMqgoDYEKV/xNyMiiSfMEoN4VL4
G1meVdMlqjcuMiHNFXZxEc7/OVTA2pKJa3AMPwBLSnK5DU81KOLwNLMST/EdA5UyZ1IXERyzGJ4x
B5/NDun3Yce9JOk3ARKCcvOa9/0fyEC7HzKq/um0kracCnW4pcqEGe0++6scsoCLX+76JY4lJs9p
ZEAB8vI90jJs+Z5oT1e0XOUztDIhPPh1PDkWWLRT/S3bTEEackgevSPDIGbZ0HFOzGxq40/gmbqL
avzWJr10l/LJN6wDOr1CYHWyuSFjT/pzMT5jExe6iz9Qcui8PiGTlNvc9O+KxrRRIakoe6WQ77Sv
NNrokHghJT6uOaP5YEgs0LXBpo2jH8SAKvjz9LBm3k7uKNPCmZzEgPlvxl4LMNA3WfvkoJcY5oV0
oszSsHg/pmGD41Y+sc/QcR8UaV4QSXl8fDvr5HwRvJOg0JTcw/54Ui8t+1xcQzif3/MSaMr/aDhw
BcmYdaa5HFXXKPRkqMDkLe3M8lpGt+OUwKOWeCvRt2V600Lkla+NzoYgkTcLbPodkdOuynZBiTLB
TfI82o2GAbBH3d9mKdq64FcAGK9zQmACPigoXXt7UC8YlubLm0ZVTNy6+DmTKIGZ7IoQsRf0vOBD
lKw+jwfsBcT5BG6yuXRNyaiUonaFc2LxjVMlRfTukSXZHdZpN1Z8zn262vl7BgZRaITyfnCgXaUT
HfFvRTeU7by/2cPbpnmKQLz//lG+M2S40+mpxX0epfWAE5NZgIzwDz+bmSARK4dOL6eJKviUe4D0
muo88y/fuvs2emYngk7bBqM/+QcFlY83YgfByfpNyKJtfaJBk4RkoUnnvaT3aXzhqsPURsgnbkVF
Sy97Vzg6wxwNziuJBGY9EV64MQM50P9FYTtJLPV+oFtSehPoVsYy2TgBVKfLwARz9J7QqoJt8F+A
JNbP6As1HHuZzpqDTeEjx6+EgpoVSFozUMq6XBoGaAqPFBV45wvsY4xuVwGe7t5HOnaFQifH9mqs
BwYZVST9UZKQ5IA48ZOtaquRwifXPubneMUbe3NPvAO5CXDyBSYF24aHPKZUdDSTNBCOztTFGXxQ
iSFw5TK/r/0kQU7upli1t0M5X8qg+vIoaejwoPbnVDdnlBO5JmGLItF2BGpIGRw3ck40EfUCwmMJ
G/g8wg3LLtIZ45beHfbNdhnlcziIzYDzGx32TT0hj8VjywDchoujqfWMMYHhLKGCtEWKsVUHwSsH
Ljcn8VYErrEkAlnEEaJq0PXc+ZmPiUEeTxOvWQRgexHCLTSlnauywI688U/ZOtx3ijCxbf9roHW7
VZe59dw/tcp9XXQ/tOoOY+I/TA9D7TxZ+8Yx35KIqqHMAFBOx+CNg9jFexnwHghBqGd0+fShu1Pn
qP3xWeA2JyQVoO7zuFhbkR3Yfqo/js27jKdgIPrmIG99D0WOHQtfTuTmKuCAvsj5nVtqzgazq7Xw
vc0aE1dMW1ZNi/g6xZ9ykeMgpf2UAe2/tu/jCDLkktdw8VoAaNVYq37geWGI7Z/d3D6GwlNbSHYP
KeanKTYiXbZf7hDhJbtPxVGR40xTtPeADGonUwpVoTQl4gDFy3KGCVb/Z3aSep97oiG9mLX7ZhWa
RjmCctYFgwdRaXX1MsrvbkyGKI9LGop7zjZ2y21CFI2aFXjzR3udDVoNpMoiOwHVRz7ONocHvGxI
N09s7Y+I8Al4L8FKty3ycIaj8EmBxKntmeWM0DiI3fCOHC+566bbY8CWRwKbQkwAfE6QWInXKwt5
mVIyj9TYQi0MyLjL/mh60+uAFoMGZkcnEAZSYNasvlVRP3p5v6MxmqktusrdWdxfKuUmzdnCs4Mc
TQSmpPu2foxfMgv+Hz9V89BcdocCWpikZrMZoBKB5208jjvXKaX8/3v0oHUW6f31GmeapQ87y8X4
9p4brhnMyfd4CGQ6KUns1kaDeEzh2u2U17YVeuGjOON7D3s/Il67j/2OBFkaIDM4m/FSW3L3uaba
rtZCtv9kOsVaRyWn2Oknp06AdGguDm5f+l8nhtZ+neYhbxBYvhZh6SPYbQ4M8DkwSvjVwy6W7rG5
mNov9zkmhaNmBQm39qwoeZO3DXsbgPXuaRKZKqqDEhtr+2wl/U+yD74Cf+OnCjRhQp1d962KNk3Q
1ZhGIACRC61q8INpDaikPFJAPTxAnn6fHqK9qtNBCRRt6i2+BZGyRbEblUn7m9gKgh4+g2ST/8ZJ
kO8GRWkdJgOYcL08sj6bzL16NKgIlXFfFn8JH9c5qeDUsaFj4EgaMfxxbXnNLT/Bgr3ICfeMEM9e
PBSXrvGrt94kYTnBbpIaTyzpLls+oyp8ZSJW81eu6veubFNIn5eEmvyvYTl+5FTzBbEfezbxcrkP
o6bdSvHTUhs9SyQJd+hAfS5fMzylWJb2gTMOO4YuFzFlZGA5QYE3pz+PMjXInY9ofj8V0wnpPIUz
toyponrKXhAyDKiNLbkgrxLt9N9FcEu2Usd3IaHhEaMvB122vpqkjlQJYfp4usNI6FLF1chjaQfp
6ksAtY8Uo/0mr1zQPDWhGSePAKiH3tJN+PtCnGv8eZvsgg3yjyBKw2a1TuCfGGBrbAzJ/cjMb2gU
162+uGTndXFDb8EkoEkcTGLeZ1ULZSoDxa/3OVum720wO/+irMQS729pxXgzxUYxZ0ls3VHQrDCW
ekrDdjzBALDsz+RXpBPuHI30+jEUnvE0Oj9h/dGMElK2GrcpU2qU7a5kk9B8Wc3/lO4LlWy0Ld6v
KB593eWfTLZSMcF7wA5eAy7CWfTKzwkmsdp2vbsKQZvudugf7rdjkEIcgpB1Z4Rtz++AhYGrwLix
UZaBkViruTGsnsmN4mFSAkrVNOoAUOa1mjAWjmUuRHBJTT/c5kwkUE6v7zUMqNGkX655ZgP2ev1Y
mJ9Qdqmom0d47a+nYrZ1SxdmgYbo1HUKU9PZloCjpWXRJk/xa5++w278EHHvkdXT/l7B+StrMsqY
JhRRpkP1K0nMDZchEMSy4Di641i7h0ekDeODHTZnibmA93F87CmgH6pUZfnM7+Nn3cKMph4OMphB
gATsg6bdF8AiqVtINLJQHxBzKfXHh0xf76sk4kJYhD6F8C6fpvqyO9I/hqPffHY5Z8hr7ttvt4ce
BEb8dkOzu01TCs7Yifil18F65NLTiusP+R1wVx+lI1uMwZwsugeFLAgzg6pbDW0cC1WS6/rBqD+J
pS6rNG0rCRJjFaC3LjkyviShhfXsKf/HuJj2AmKQEHth2MHYfOn7iu8lTxNT1jm14uzAwoubuu5d
+MpSnGLO49H+8Klw96+aP2/JN2jIKhKMik6GmpqGGnuod4gzYk7D+0C/yI6otWb31DbcGItuonTw
+6aOPR9OlAl4b2Js42Clkup+avlIJLzofb2NS7MFD6lo0Rzi4uE53HdA4xKsyPvJVHOkW9yzUedH
DQMgh84ooY/64cvsf3yRqA0RYe30CRvSdio1Xuwfe5ToKcx8oXLBNmqCSIBlCL5vEkvQCd7tkbyW
OSLWYZFuF+OF5cfyKmweeIYVbkIJpmPk6XKT9ewWT9C6MRKnELWL7EbPwx+u2onH1U8Yh/FtSdbK
oox/1JQHgOyKC338L2l/mXvf3UQyASCoTzhYx+sjVgp1x5Q3+/FzIO7NoDjfVAI40mmgKYNVIIOa
D94/XRFjtOjlfEAxGe4nwO1Rw19Q9sXpFkuJfMcZH2bCEstu6IsBo5fGwpTEBGBbHY1NoAxhTw9y
yddBGLBFob2JVzJ3afjazdan8W3+lFYOiPlqTO/kkMxGh/GfujSLp9Bm4KOCR8Vgzhf3rMYw8RIS
PHw3m3RiwjNyITL/PIniieFdb1Zi2DVFU8HJ+JS5VLML6n2c+TFnfx1TQR0uK1EXXUH9sHlCI6Sb
WRg30bvhnjsZzFq0nrCvgU3gSdvEicX4jkj9/ytBKErU8xh1F67A7V38d67blc7qwcaPSB5NyYUI
3LfCf/EmOueKkLoglZQAiISFHy9rUean1ZwrAKvxL0c6R2/uZL7vJtFN6Pk+ftB90Mky60UlLiNL
qhdGa46MCKS7zjeykGs2btEpaaLEw3jthFwsOhRez7G8Q3mPJ1VQL1yplf26LKH5DHd/wQTdnjLs
6jSj5rW4SGMEwboiAyXr5e9/3DHhpt4svmfnAEP3XEuQdnYteOu8g9qenSNv+NKIuG/6uecCpVZM
UFRGBmT+ZZ74jWnAWiAArUCeghwQXB3OxKUOP2jnkR2CPYbjh2uMdyVADmM0pT7sDX9Sf6RQmLnF
EVPZIYavIdZAQbANckQHe04SGIF1bUyRpsatWHa6/TWOA6cfyFIufTKD8Zx+huVtFHvwrYKdGpiO
O1UbwUKWAUOjPkdiM6tbzRnQfSecNFgzjx/GrEXx52yVZjww0oZAkHPgdZ38UWtYpVmGH4dSNr2t
4TFQUsMRqMIvIod+bsD1Zus7qQ1DVIdWzO8g9mwTxSMJ1prEdOewW/UkZRS66Y8YiALtOdMQ2kVT
KnKXJv2NtT3Y5xqqh08CL9UaT7dzZsxvui2++PHI206mNbN6C/Ao27D21mep7PKi9sMOSpxpycuL
ub9cFcVMomzdI+2ih6pIRa9D4OedvCiLwmz8AxfgB+X7oGbFN/DcZ80/QPyfE/O7906ECWtA7DCA
CWAgF17gd40u1UtFGOmnavyNpTezejsVdptzLObrGIyTNjrPZb+p+je6L4CsuDkvWwNq/AzVTN0T
QzHwXtkNDgOXO1MFERV2qCl9wKCy7aJbFCXOFzV816JK0W23XoF8y5BnN8hSeLnBvEgpyt7bSjeE
iN74KvkRviWp2/kYvMUAQeMengvsSVdkMDFUpDiTErwWVJjjPHX8IH8hwsXOi9marvr0lpU8bstR
ziXRrzbusCZaftMZNxSvf21r1GgKXplP4Viw0fV2UWssWFSL0HEHRCk8DZ9TWEsivcYiHhVhLhc7
8ynois0/WUTxiH6uCIwcQWxT8iXvw9TeZnaVRM14UVR9UOG/Ih7YWTgIqlIUcwi20eafwhlEUQu3
kR++lQxwM38GWm4uyUhe+LJdhLTN+rJ9yyV7+HFcdMVhixQW+MBa1s7AZRAZioDudTO8nsUbeQfI
Tmy0YGDmHaXx8fPnQ90nKzCdubQ/vS5g40RTMFsTp/UWhOW/Emirt77PIpxqzp+KAUbOpxBgW7Vr
35fEGq0rHux4p9m1r3XIBrtWPt571VUfswAOsm1KVq4zOsH7jb+TSQnL4NfUF8QRvttCMqcJ1/Uw
9MZKQCKWjBGVSSriiFBFmfxUZB2PPLdXSq8RnfKe87mRRZkeIlLJWCvs2n/0/maH6fCCPSb8ObzL
Uuu06dFOrTK7B9r9E3LeBQVSRG9S+zaHtUF8PtZWGjlERUo3sG7ALznOZmcxPwhAbLTNq0HjOTIS
CguObSVeuLCuDRosourveZZFG73pd5u7uRGBF4dOsnrSocNnwGljuS3U+j8I6Nf2fIw7wbADlMvN
PcTBSoDkhAYbZ2OmanVb5n5U4jh/F5RUZ12SVw/Rwcr7brbecSV9ZsBOWhG74HK5pCjJ+gixX3uC
iyKEoqcSllJYI5k0NohyFuS3J3Kwycvx9eNO+/PP1W7Zc0V1Vv1eC7HamdWtOohc74Uav4/9mqEf
bXoj2BqFK5JVkIpydTstzwhoZ4Yu4vfHuZcV2/voiS41wvZKz342cWXz99fLiORfojzaSgBUmTlJ
Ggd9s4NnEuoB077STIh35jbgGO51i3FJUroGxa5Neyu54s/K/YfepfvNkCVI0R6K9SmmpakAwZvd
M54knuUrgasC51+tQv53YT4yTZmPwatAg8222jjNw7OqFQ9vrBTDPHgy2brJPIu4t6zv2es5y7cf
eYsuFsZ//cEJDN4n5osKgrsFhqTUiV4NjxWsGFmvfrzXvR3x3WH7OOrVyWHAQuY1RgJ32f5K6Xn8
hVOLE8PJB9eavVGnmr9TNIp2dheEpGbiQbqXhgFMum3SKG/GCxuDfeQEMEhu1gNpAz6C1j5HO9R9
7w0CpFoNBi0wDmLFn2cQNN2v9UZDhA0wUw7Q2JeWJylxKxVOYi4RhTp6QAJ2u0pwKEzeI86z1dbV
9QeyhFSZV6hfWofeydbiUEreeJY3UZieHMPF5NPSAzrbu7iYk9unYd23slrIR1CsyLT1ZSiHVC5T
A1dM6aU7Vx/R9pTslR4B/HRzxiLlCwptCO3iLHSE8904uGR9YxNjzbWRIE0eSjJgahm7kvVym4lc
qZcQufg9ttNlW1XIzDPVTmVM/rsDzjQhlNtX9XraUJhkhcqezxrcOgJ0KqupBiRu3frsHlP2O9y2
KU8Efwb3/kl4mjQWVnFmE3gVtlN1vPQ4s9FAjpeGXMb1baiKfTTsfnfEpVyayYDSREb6aYalTKzM
rgWIoHdBhLd8O2u1u7OTDLjyXGO32UiccEgwkyAvZwWOIPRLvIChOHeA5wAvFopjU1ZTOBx58i3E
rJpUnwaCUAIWeykvUv68X1/sTLa6oAhJGd9YlJOQjTXEqJaAbuYtJPgL+ttiC+P0+1jnAQosCt/O
BqbOjbAKwApT8glIOSoA0Lg3ett4O0yN3OAAhLOQy9LbsKZkn/wjuPhc79grWCqPoTWTCgXoqHHg
gEg6fSQtH+Iw5ZMhI37NhombCIt/fXYhMwWlJrO5LXO6F3x+zGjMd4CQMGJ3yZx54UIQYpHnf4D+
NYm6wgv6qztekwQEuO6FFmu5bmXLP/Y+wvha3MTV3VXxybMsdVaM0QohW2IMrDC/Ol7Aw2QLt5q+
p3S9AKOgZ8NsRpWOvZvEQTkeecp60QGwmxYL2Q01CN4ZmHrUdYHvs6Y1jy894tCAwZrxNcWnWX4Q
Ej/M5gX3Harg+Q7j9zpzq2gDa0u+E+XS78/2W1UCGYXNvkGPUfWFJwpbycwF+57t2Rinb5Y8zlVm
pRFR2QfBC9/we6oKBPGOBzn3DMjbboX8XR16VHo4UVAesjlk7gM6CUUUX5FKKpxm8vgzGDy483pM
O31ZSJ8Sxm6HtyHw5N9sKUSgsBQv9yOmYfXkznIzcRSYQfLHaPOanecjdgk3slnfNppmEaBuoUHr
qzR8G6TN2NicSMYkBDP3ctaQMjZxBmMduQ7XZCKyyPY4gojdt5ZKGNl5LOQzt4xfskygZuI/O+h2
NRBI+kC7uQMomz2nwJRodsJh4IUDDv5AwruK0ahnZEX1Fi7McQBjLYk0qFoBM00AG5D3zQ1Ioy4o
XDb3e7415zGiRZyWtu9fuHCK1czzdIrN1ZD5K3pP/cpZgfmD58gCWfN/y1BjblT6Aj8giezcOvhy
1Nid8+ksE2VeA40iiE1133jKPieloe8VVtt/59q4NrGpJC5I/AqNhZe97xijddAMZrFsUTVaB3XE
q+084l0jSwhwaXs6THBgQkZW9PT61hjvUxy+oQ2Jsg+EnnpdUz2XlrA2DsC496kOly1/JUwc+KbS
sK1Nhx46fYli/y6C6Q+nYAqrMlw2/RBAtkdCPrKJTjAn7h0F+p5K2SBWggEiWobSb+lKpcsMiwwW
xc4fONSz8iLd0ufA+VXP/jt6GWWS7Og5eBhjwqhkdLMTj3/vkxbOnCHCEQtRycUs7A/qbatSc0y5
BxOHW5AsAwgjSk0jUyct9szh5uLwKJsKC40TUjzTwex0tG4pQ6cVlhWnqkaSGrFKxf6AT13eFoyo
88FC6y+aYdfyu8YCMz8kNbOeVo8UT6KbShBl6/KiYYA1dhcJQoONolQ/Ow68Wcwt/jlWckalm2PZ
w66vGo28m74Wyn1hNaGlHviqmQK0fk4DxvF9FA9qaGWZ5/KZcycUnon97Vfvf/zLA486Rl60opej
XzfZPikMq9QHFz9cGGosxVpE/GWbu4HZhsdFjqzpVnfog7ljPK6qcxehO8FywEtAEHeeSMMbFk8m
qVJL8iqHuZxPKTIuJ7eGKBT1rRC8GxgJwlxnfbNM2XWe8gUXeMvFsU/DBGyJ1UXkPnM2CVO8BbbG
rsrB0kzuUI6mhweUCkOqIM3WcriB6830BNzPUFzyY1oU81keuehWsRJiiUMKCXop1eQ0KXyPFg2e
uXu3hT5zWQpLq7RmwU3a6ne7/0bPZMgQwC49n23DV6CeRMnbN+bQL94Caxgz0chGpvB9W5sIGBEC
xd69v065zkp4zqyOfcJFhxGHx7NZPmuCul2dx5vXk9eFjPUKM+svX67dzsyLnnW6PsKPH/G2w/ba
VqBPkgMT8FwWP/8+YR9XKm6jHv5HDd+wIq43MB6fwX82if9yn3HslYs+7pU81ITc0ZIIEZNmAgbw
x6e7jM7S28sfxdUbSpQSonlqIAdnBikEUHN93+UAGCppkdg9+ox7+QyOJVpCZfTch8xchd0ZkCns
UcRchp5x0IQzk7eNDVFaggDHUzSa7s/4AIE55dbWB/FAKIFyUWv+pB+ybhIXB1v4djshf8v0j6rP
YBUVe9uYOymduANmkDGmnvtk8nFHDzd92Vf+RYPTaIKSih5cM0H07M7dLHfbHcW4JyB4GNZpBNZQ
KvTUWHJCTkzumlVeOmcJX4yaVcw1O3ZhrgCgeKEfxrmfMBeyWkzR3crIsEpDVnZ0VvjAN9m14hXB
ccNF399jN47OVLM7goxngPoANsYrOx5aOc1oiV4s3LUo23Yyc75mSflnHqQ67HWRSeEMLU58d8Wp
8vQ4use9XtbjL+/KG9SYvT9FD/kDG9MZ7ZrValwhOzkSrWKlsvR7dpzj5o63jNFDU1vO1nu3phg9
wMiSE08letMb4m3RI7hpClWgaBgf59EvffVWGpngGqRQuuItLJO0Dh/Ktbe+5rJtIKTm8dgKXDYn
+OkG0yg3bjhqsKhhVh/E+uVBSBBZjt/swzcm0Vdq7dZVbPr7iULUbkNg1EF1YwSOUVxD5Vd5bkmI
352r0vxKPtsJsJsiwtsmepd5C+0kJb4xoC6kurI0uXGn8gPzBlZ4MySE0p+yuNd8sz/4NsRakwey
VzoyOEYZp2KEqy8muVjBIHtCPtx8VK9xmjwruWdgHiBEpC8H8mlu8PTsiylCJGiN7FVaPqBQgvLy
rDzzUINA/Ti70JWinMRjgunmkdqtMazPNgOZFMfHjS0rBD913kJZQYDrEhCyvBfvn3n73GOt3p88
279rfMrxfV4O0D45TVfWN6Rl0HS9qZzhlFYybiqRZp2f0tKSyjKEpbw6RU3PvsoWcOpEuybApaQG
9sB8T4HVVM73AFW46W4KUz2UIovRRqvQyxbLdTWD2wvc7Sou5u6i5k4BzYKW3ryeq5wN6by/WZP7
wROu05oC4uwV9muKWkuVBAbn8kylq3e5SspMw1B0zvUvY3H6N/boHjhvWN2JoP00O95rKMJ3PB5L
PvMzGQwRnMhCxdXjgbi1JkwTxNGGxE6HzuLX4Voy2DlkqNY5vOAawgtUPDGnoa3+gznjP9LOI04X
6g1MIFQ1l+SnHMu+Kn/brPyz140gW8puPs0YLc+BSFhSSNYJpQklmctwJL9FMkDnxJc+o9/ptQlB
vvpH1bfR97Me94zx5SISkn8VgwoWBx8P+CZAxbxCSaB5Lf+QbqNksoHC8aZebRKBaFf5s2z6yKXP
/Q56TKAV2YzqivexkUA2GdObacXZZIlwdqAMsi3iBlFWzt7uMXvvXhjh2/363RLe1rNCeWK22+hq
IVa16zpvSklOa1oyLO6vDEwJtf3YJjgXW1V8d4a7qg6tlBsNRj3tRHh+Inx6fQY0jue6Hc4gJBIP
mAqgBS3PVPQWXi4FAGvkUp3KLZ0D61Nb2wZ+l1GA4OhsCHuJRliUlfBm7v63v8h0dRyw5IQs7M/8
smFiwDhOgp7UqHs/3fuK2AtyrOQsNkNRIq/ZPfxh/G7/WXBubUTn5h/23JJkus3KrAbzkotXTOeI
ZruKfIQr0Zeb0rNWpnT67zf15XVohpFy3RopTScvJRuSIX0K0vHNyOU/aMaECkI/yJxqhyRCCn3b
nSSvnbFQNSvovbyvfBcZlfJ1rsvAsVpPVwVu5upaVbNUbDfT7FJkAf5OH8SGZWwPQVrCyMAVyvmV
K3OLkru1RT/HAWhWU0MR9SLEnjmve/6wzAu2dLrAz8ViuJiFRinbzTUPNOLoBolvvbOu4XyZDZ+l
izz9QIW3x/wNxPo3TBorTN/Pcp0c8qIqlRz7O8K4excramAcA+qJy/jcEfdLYUXkIzFiB35McTIz
dwKN75nPpPBnenXq6NIkdvCE5Kf9x+jy1qGyOsAdYsnOuWbFpnQfhLJ9Eyt8l41rRAaK6LRjeV5o
GU0feIJ5KXs+ZDxVm3MulrSxJwDzZgZc4/KjdYT+Re6+Uzdk63lR+CS6hYFVHuGguxjVWCCd1rdW
rZeiGoTB5qbkVYoQuRACxFY98DcDsdgjEe4oMj40UGXf7/W/MphrzSv5IB2A3WbuVlOP3jLod862
RGhlUAobWPHmyD8O2qj84nKyIlvWnbC/rUKk3r/sRtDWSLTTMRpTxQvef4gb8q/Fjy7qik4UJjad
yQcWw3dTEq75EapWNk2vUqadrRk9RCzKT0nwuVA8gdu3ULLjyawB+WWmVO8M/I4SGXoZiNTxn0lU
nlJRUcuEV9rqOJG5NSxhMrFFOOPFo5+3qNahAOMDLFCLytZ+p+ORloWCUbX+QpEk2ytUNq+8pmo4
p4DHQTEDQBrkZtKIuvNB1zEzCMWmuaJQZspOM8y86xu/qBZCTZ91x5lxg6R9uB9cXV9gw26XM13p
w8VJKQQr7mc8H8sVGb9cdwuFBUQxGynEeGN12BU9qr845KAtb9MlueXc82kaWY/BKmGjBho+MTMi
5BDv9ejdQ6K96gpbqM5N8kjWm8Gqd3R/4bUlr9v2pii4zHv+4YzcWBTl0IvVEymHFWFmNI9jGqGA
xozdM4G7RHTQnDF1kuN484VwQBlMfRPbI4MwRrYOwSgrM/PfR4bHK5wvox+CZZ7dycS//znqlSQi
B/dmIUxG3eYdSHQWKGBWY/H/49YTE4yFnb/zMMFz3JAZXTYWqn8l+q/to9fpgfmX7Ns9/OXv0Zll
Czc0xkYuYb2ixptFFgnnuEOOui7j/guOtsPUPzLI4myjQjs1kcUBDfUaFj44UYnOxjGDfQKDQSwk
ILbaz2AuaQYygPuHqeIZMjxB1b9LbFoueMLcRGXYRgHfKXxIn3ekbD+L1/UlIqHxDbBb0TbBt05R
K0NRQshGpUWzODIWY8I+1qIniKniGNCmXif+WFCcRmLN8hsrCfcAOGBKGceAfXJU7SYMFy/ufh4s
nh1twPGK176YxI7wGfnAB+GRUxYIX5si+AJI8k786FR/80553VBW6/48RVEQpxEb4ANEzhJm51Co
YqoD7rN2lACzUEgowDLXMOoH6OWzBfQq3Cp4JpMAoTB5hhO+YXwiWUeCHSxJNxDUY4AhEu6sBcM2
nWGwKI2U59F+4WA4edX+mALa+ZApe65xva5/6oTh8jLCkPWDOqsl15tiinSL66oEZY7GNirba/7b
aiB47+RJ0ivJ9EoJp977WZeMo20eTx7sbM6CkAo2bY0bWSOUgrECEkrtJLSXOIQKPEfPx0QSi8Fe
swEY7G5hoxWafk13jYDibuX1438TY/YpmO8XO5CuABvOIvr4Akdfr+fiKNwI7Y/3KaIi7tInwmly
cvI0l2SJDsCB6kGEyiJ19cmxHTVjwD/dauvCJpabH4tdEne6IHkqt3w2faebmpy0zhFjt4C0JMP9
zlPj5ZZk/cgLrc6IyK/TT3+NjtCepe2yVUwF/GNmGozJVcZ22jEGDFZOmtKtzrG2Up9MKrtKlB9I
SCPFSFgyWZ5FC6kvC5ShCWD5N7dzAVbOM0xi/gc4ZvFL1TmsFETUTV4rOr/Lf3CvaZUwefOy9Udd
75IQZjzeu/CNEnkuS9OPjs7PD85nKhwYdWXgYgTHZqCl+BmnV4tY6ExqkZn6RcKm/ehtTExBrbR9
f1Gb66L9dPw039G/IEGfiCYZ8dMmQpNrBWvVf2lXYVCyaDAhEgLJQ9HekxsDSIL7Kj+/Mk9MBk1C
TSefTK//MSxNYpLMBnYsNl6DMLsK7F2qCwqYAS5Lb7Cobqq5rMKCtZIVBzqND7y7Yz18FXNZLA5k
aFvd2qwWgl1owUiXUXYAMfia6+5hIemA4thvdSbELFvH9iT1kma9Km20fdrfD9eh9x9o/Zo0H/dt
IHmeVeKKQlLnugCFtuejaUr8j7J6wwRTYoBlpD+OFppU9IjcsvfDFJMBUllS6RPSfai+NDNn0KxV
+nUiPpHYV1xgMph/hQEA6LevEC7slGhrALGljEALK0bGW6Fkk8WOHLuoC5Dh6K+VjWQlFbs/ron2
/FJgnfdinlRjj3BkAj9pGzlVPMK8DKmplpVyCIaf/tIn2Opb8+7Js8+h5izTlpEd3C1o2XzAE/rp
7cQgscvr8rDqX3D2rcLU5Vs2sLm3V1fH6PI6KGh6+4TKJSi+/hLUo0XQUIYgJTMuMNEiF5x2QcMb
OKvaPagUN3m6YfTLm62xjpHaC0+ofNQS265Mxfffd/wzNgKZeJsrz18kBH7KHDcf3qw7nyWFm4zM
11lYCh0gea5N6f/bo9bIFioBjjexDoW8LMJymxzbVgZWtVNZtoemy33tBWdCDEKM1YJHtizsTwtN
HBRxVUZf7EVLUIKQGlUkhSuMAcO04gOiwxuUFca/waXTjNOFPazjNau2eCKbd+1yGacevD9us+J9
r6jNh8/271gofmcj52kk+KR3nzSddgn+iBwFh5/AtP6xlr+r4tuhEMQWKf1pka1xgraCw/hXyUhw
xhavbNco50+iR3bzsN8ATnZJAYbt9YUCEqMjcJhaRHVmMoUriZE3mmLCCHjLLbd7nX8LmD/vXGXe
WlVA/51s5HH1jbUcngOE77Z6iFUBY3z5XkleNH/QMXDdb8zU2fJVjRt2D9LHvZRO19E3my8CLslK
5E4XyhAjwCLC12ON4rlQAPAMVXPbWlfk6mV0hLiQucUMzbps1IOgzRiol3MMym/qK2QWn+LorG6C
PGMH0UBLkT7h8A8q+eHVd4ywuJqdAgRbk8yzw7u5MiLE8z5it8xBsMJZrZq1AdutS2mGVhhvyWTw
dLpSgS1SEO7KC+OKSNdJ2DLUq/4nN40/VyqR9mxBjurvWG/rvhtz3iDwO6lGg5sm+g4VaX14hFZV
EUPPiSwguJgpZGwiMhxV7Fj2nZIKNDmuj+atbQoETkwi1gPKoJQJKLXrp5iMWdAuoXtY5eSnMnUQ
oCDf4xyWb/tbIaukOxZ843hJKwjrf23Wmx30/1eC36CUZzSqPHByacVxNtccuNp55ANq0avJnwcw
RuUvsYEX8fB74tiCFaF8YWfqreFx6yjMFeOYgizMLVoK7LHWHufMG8byV2iy1bZsZ4F2w1AMofWx
WO+k+8Ya4/DD07rilTYkfQO3G8oksiCUSpO4FPLqdx3zpkZeircGCrgCj5X6pmdPUFA0yVbRUhDs
FghSTl8jfOhONGTA4xx4usoGlSWfgEmzG+xb5yQ1auDq3DHuE4EZ+4OKl9yjeYyLD+cJ6PBegy+1
7i+KljJefJ2rS3GpCF+TCvsUnHMs4/mssTNNE9zEqG1fyFZyj2avsxvo86+1rdMp1VvaXU2beuZk
GqtvsTCVVdf3og+x1AqzDXHVSPzZoSG547U/L2jeQ1zaxD1iXcr/rHxjqUL07mDeUEjdvi9s8Ign
xqMqCIzAz4zzUeW18BD1eO0jFSl1hKnIzKNzdKUqdE/HtojR5M6D86uC0C1MyAej+gever+MCC/n
UBLp/zM8neqaadAZMczgTe03icLNeyIzRjFCVCbE4wvbInQ8R/nfYELYQOREIe5HziWtl45B75ho
QulP+kDcLWFlr78D99DsVHa8LSbEAZIqdIqbsvNOoaqYC1ZaA5KHbuLzDJx/YO3JmaO2hLJPLZSU
WVuYXbeHQOtRxIyCGI/MdeSoV25eW8Be3GIIVbnpNQ0WsKEAKvgBRUybU59vzj5IbFb9go8MIGPc
LhOdJ54dn6WAgmearZ4SVutMYz9h3rvuAicsnL9BCBk+yjgYpXnMY6TwMEdvRPsA5p5Pr1ulI5Nb
0kPQte+1rUObiYhirge1kgnSf6FAEvJSv2BKezKR5f//hT5MEQr78qTelo4x+59HbyqNvFUfQDM3
kGDnnpNKOf5VcxL+vWOFyJ+r6lstYu1A+IqNdLBGnaPdJ83HFUIIUh6S8e8dVrVo42xGkTrXnmjo
5OxrIJ2FEqFfUW7JPrqYl9IyTPTSToI4ZzFWz8NdLxLsFkD2WBUynM9ZTqMe/VU2UEHH/knRBkGv
MdnSpahTs+jsjwpT7RzemWtkeHZnEC4ZafaJ5k/wb8wU0kt1XsZdydlqbSAkdF1UW4JrMbyHFsX2
2N9li9K0gcHBuLR+HQPphW6mVEsdKsRNJgta/mtHN9x3tdBxfiXNakX16wy/u5nZ2+gFqsIlvaC0
1HAZkx8pPEirN5gybZ4xR6m320MMlNb/42OUfh2RIwlS3zMy0PHD38LU8omM5jlbL2XMc9L4nyZu
tXZRkO6rc+q2ugJuEV0N+Ny+4W/fMmEgA+blpDg451woLFeLEBGvjbc36zdXpgV9SQ8r/dwbldv8
icMcvh9xJT/Aqb4tGbCvZGS90eO53gCgkGDw4JBs0fW9wwdAbA2V81E8kpnTWAxWN5Pdt/Z2EfvP
c1mNs9LjWDE09qZb3Tb43UOgGKDK646WnXJHK8C8QdazmCFmd26FT9SDJ2IfARKVFgnqYVnHs73m
DEJpe/AseUF++pSboJFTLcQiguhYzW80gN1n/7I6GzWwnjsZeRgVuJooGFSFfA4d/wHaaxVp7Xg8
LbE3Sk2ffbZe0hMP/CuCM1qD2+cYB8qkJWnqtWMNK3A+V+vB+ovpyYBL/oh+zhDRNPXCzrYoxgyq
J5AQsvqz/uTRyfDD6N5SbkSV4EVJjcew8ilM8kfp4gcteK86sd2q09q3/m0vbtBY/IC/69R1SHqK
HjBjtlFUT1q6scmi4v4YTDKdUio+1318L7jF3SMNVGfc/X6duIZ6WahcctmAscAWR2ya5SqOz3Qj
WUm8ppeM18/CGHEuL+aty7eQy7AsVrWzNy8RqAqTIflax+MImKkpnn563bQJT4juXVwf0ruuFgE4
YI/luSI6pSeloE1bg/Zenf4tkoPbwQMiGbAlbS2j46YMcpFwu77C1JvByRqQUoXcPPspHGUdBIlz
LjEL8iPoqXzhP+I5DFV5WhK+QmEZwIAv0Y5OFZfc2tlckZ52WR6anqVKB1yVuI56bd/WPKIqi+zn
1NErd3HVKTYd6KsA+cYqb2y9/BnFqG3fFRMUlUBoBTiP2FtiqEHYPNS6RJCGNPy3LAn8FEzvrunZ
XSfm8EPidIHA7rIPWQrLVfdmwwF+fuvRBKR1sAMyPe2n1/MHvpq31FpeDPjSqVjc2jcOD7lnyyt9
7WOgYFlxOr+KjNZJb7ehByLhQHuGdpu5ZV+ZbuIpdHNj94qBDs6Pv28OZ7YL42CRWlUChgtl3vSG
sNRC8zh2b/7uRADKlvecuFfwT0fRN70/JRpdFE+WWbigXuyzcgVEU5ohs2Jlken5SI0g0vZpxlSQ
pcoIabgAI/bINE84UfjCmY0HK12Yxty/OttGUboWmqmuO8als7GPjE1unqsbQQ5KqUvW9QCQm+bm
xUu5Tub8b3b6O0vRulQ75L0REj67H2A1idncZstYO+vYRofY0h/E2Gv8fAeN/G/JdDMzoPlQKokj
r6b5bcRAvQi8QAfy/tT498Q6cGnLr46Z4nAV9lWMRrx1oiVenHpMedQVrP0iuf2Jw2P14p+wuq6G
s5oN4xcD1YJ+Jo7lJMsDMeTu3mimUTq7QYZKv6YMhcsihAxfoLB9mk4jqf/Zc2FI6y0xHSWHpB9f
FTmbo3mXuRuBJwfQIvzo37ZBVbwIe+xcqZgMttFt3RuYnrlIwhYAiHdtMLlGPk29RyN+vnHCpZtx
LVUC9NQU8ZAgj+I/vm4D8rTaWPK4vdaHvByrrsuvIE4hw0GO3WrGw89GZLTqPvDdApYm+1cNFDYM
6KtH5N99xfgNG4+nfP1Ct/HVKTwoUYL+ypK+pFrkpb1ivhcwDstb4fq/o+TAYRJsqUArOEl73gfy
X5fCxw4B5A85b4YzeXVPrhc2yMiXgBHJb0YW0JiXlPlwKffJ6Cf6xJpvVpYiUE3og7VSwe4zBhtf
okmprcoeLQWBw3EGs0bvd00n3XttDnhTkWgIJ6cVvsN8qq1woAw0KdToPZgxedKvI22MD1LPlOO2
+etC3RPSk3yEW3jgcpkO9NDs+R+xkZKIcST/SBOI2i2qmn1Ia85+SsrE+46BTRnpPLpQMe/QxMPk
ZQ9i//9s2TGAe8hjdsdLXeyX5j5qsZYm0qnlc3rlo5oHLNVzyNQpySeWbLQWEQvY11se/t2bPYmY
2LZrJXTqwIbMQZKq9AqgbVaLUJhSZyKENJuvSzEXqre+f51iT2E+1Qt4UehYa4bZEzYHboTP4XbT
tF8tsgCK6rcacZERwHUfnVxvIb0JzH5RX5ZEFxB7YPBibFntT/eLuG1NsGMA84OZZQQTjFp8/KOW
1qYS5Oec2wLsEzCDxM10qtdNu/fk03Shie4uIdvq3gaYXynT9CdwRNx2zVPP8LA1KdekwKkbD79/
72/mTYzIIemKV16HNGppiIDxK+i0HMiO8kZ+8PqL8v1AlnroUH0OAUtJNkNwj7BQcTK4a5E5X9hw
Do7W4XgKDyx7MBQ6pzE2r34YBz8uZizfdggkNrbFbIpoPRZ0ngJ3URYmMTG62VphjorwPJJMKNrj
ibkXHbXhO5BACUNVlEs/FyDP/2SSv1taXxJ0E0rgql1Jyf8qmTRrysMkyohVn/RlFZy02HgvrcCh
wc4FTcRJeRQEAcynHAHlf7ifO1eeC2pcxnR5/NoAIS8RQJiVVp+AEOj4sgdKpX5wEBv58Qlpegqt
PYm2AYmg5P9U47ylZK/fUtVcrTpuDx1FV4rPnKxMrXF3I11qmy77IQRWvIKYU/1+7+z17O8xaxu7
0+bwfQeQbTrkpukC+s4JUMZqIQQrKBtlHf9n/ULpEshMDpRA6IyMcxPy/Qm2b22bPFNjxdOBMdtu
lMY2R79XGXyeqx6bCcQ8jfsGmsYqblJnKCQh0Zlqezf3uVmPyWo5XfYQ/gz6ntPoCBXV0PucGU54
WvWUPYIH5CrsyqfqmFx+lEyFplWx4ZGUM1ou1NIFCbwdUQsiBhofpKwz7DSyUDoVz9C2S/f77QHE
GZ4FnY1Wzkj7PAFW+gqJh315FaNHt1h3d1Qord7Nev1+oKp78TX/bTrSIvhWkszo0ki85J0qjeLq
C7FG8sha3Om4I2ifBNaOUnbSmYiL4ogIL6FPZTJ8Dz7L4m/8M1vc7sIBu0qr+6UUN5EIJ2euEEsW
Lck69DCvolpRB5t/bUVf9taItRb0HoAHo+iCiyqrIbkpUNhtMWjNYnleLIjrSLRbwXU3508IvtIF
uZyQmelOkeLXiSxfNXtTyXk9N2rqh2yGCT4kgYoJ9UubAo14GzTSvBxkQZtNXUcX165otS0lNCEp
kK2ivWlyRGeLilkU1yOEDPorQswNGrKi3KZC8NKYEUGBnMvVmpTL1/Qd+C+ikoLNezcJufAB/mIP
NbfbhVSaNP82mLl2R15nRLAMX8XvAfdv2ttRDf6a667RV8L9Eujm73udefTHbJ89ZTDk54kazdFy
QbYgATjKd6xKnhbYOfhTFyUhAlfFpO0q1VL5FZaH0ibaQBF1O9L75uAqvMHEkRt9fm0BxWh7HHVK
y9rXzjeAeWD1vFA6x9k6OWyY0RuG0jic+Wf/eMFmjnKMnym33j/WS51DrlrdwCtgYvTMc1eJoadr
t3Fh7ypzC3pdrkHn5Laa+4qD4l2xwIIjBUTloJrbN/Zg2eHCpqgoVQcM1UxjZ64MKpqaRj+0UWO5
49gSmWiCWXNd3lOyZp6JzW15pdTqPkEMRBZZGiCLMarv4LQNy2fQ788SNagB1zMq/sKs0HUrrRcJ
j8t5NOqwvbzRO6QY7ChcK0FB+0c6z0DTZCUqgezORWS3EXqpQJmJMtRp6LXjZlW2mFaZSiyBnoui
ZSZeIk15eUYTo0kWEPKR5LcGZxL+T5RKo/zYhM5pRa+1q2GXJYxbzDkzDcebJ9ulMAV5H2o5Zm8F
wBhL9w9iI47H7Umms65hn8dQtZsTHKVx/iqmDB/IcJlIWV+ypNn2eBk+OjWaGmbNcB8GryJaKab+
WrR8lz5scrU/7YB8Ve9bwigK57/B/kdYXQNPhOi/u9kseZM47f9PQjpeqTxT0wc77wp80/D9r9Ky
V4kT0vXlQGyB/ufUVM2W66CrLDiNmoE+nT2SRzpSCsWA+9Qe1hvFBcjD3nzX3mF1uWsF/UaWH73O
tBOtbiMC19DbMm9HFzkoSAMTiA/grStYwhqAZ6N/YjcmNmHmFr4XNjmo07hJAQk64YRmA8DqfXJS
oW7LgUMGJ2s47IOlv0WV54FycIEQ8KcOQdN30+xvmU42KisSEenM0Tx2GWTUcmhgQNcCeecn2SJ2
iOX7swE1H0A6k3w9eNYnp1n85FJpbhEmG6jGhAQWI4/+HmUZxPoEC554o+KSITGv0lAabaN/4CSD
zA0+lS3CCqVqQZswZFgRXOtSdJgPzVyCvVyvH3kw4oZBDp8MIQQlxvoxeVfblIE8A//CMcKWw9nr
RNVMC2uYC85r2LF/s4qj11EBq4XMUftxFcZoEV6tKJbg/5C9O5B+yDI5sTBtNvHVnG/dF4Byxioh
P7W30SRHVOtdE+N51++2oNJM2DJFnrbixwM2HwSUfENeqo3ukXBsjOLvho4JoVgxRoB1ucecP+g8
o7lJ/DyroUN97SsIKZT5XFSC8xxHoh2fbzGy5h8dxSkeTkvJ3I3Vw4lsSMM+1hvdgQczJLka8eCw
1XYAD11Ank9/fKZJT3TY2JMnnW7ZPceyACE3/69U6qhCDIzbwU109FuKTnWHAoVTr8KGNxA5DFvt
Q3CNT+ICzZWz0Xurnmo6wyWMZZqVfftnkf7VEDx4w+T4I/E4DcnyeI189/Js8a46qSc/b1F5odcc
kWRnd9yq9nWuGlPqObdOp9UsO6qbbnQZm6/Y/61xJrkYNnS8c8zsLe2oVR/YFyjph3hDjWaDDDjb
Sul3DID4To1FFzvZGuxCNIGNNfYI6H/3l1E+12P7pING25YpB+Ufl+9H2lFcWH2TK5myZHhmcvI2
54UNd2mTF5ucH1LE5FHQkK8/57SRXxVLfrdTq/vQos3U/rA2/BpkFLFpY7XWck6gDHcbw9t1hHN7
o/mlnvCmyg44MFJ3aYNUwTFiv5EBEldOAtOcZ6rEF7le4MRAmgvUeiIvBra2sxljPXClcZcRUfSe
7VqsRSd36fxwU+bxKdfQQ3ZTd8T73OpIkx9cdYj9XiIbBTpgB2q3QAH7+zix+eXSo+Z8XZRMRqZ/
YCNAaCxgNZb6PkShpmUzRn1vzI6N1+Xa79PomjM95rj1DfmdCHeoS7wTWKm/ouWd1Tq2NSrdnOtN
5PaEPViQDDD7KpnVIg6RJVqp2yuZtrjZxJ6V2koi4LonLFp8hZqsBPhBSTboEC3DXuicxaLeJ/DW
a8+/mtBiKR4kzkgHFE8CJ59LraSc6zraEG8MI7rbEMsbwqtXt4rY2aH5ncrwklr3rHExgsZFB/Is
rYuZ1W0MLgwGGkv+HGz9aD4NPxSVm3oAsEyCycv82VDXL0qt1BbWC7WzkEuDdaG3pEZnA7k/JfEO
Jv92oI6IU5/++7+CfuWDnIkngR+Dcf3nnCKvyAG3bK1sRQ5rO0q3IHhwCqAjj9McuFYwp+ri+O16
0gxh6Rsh2y2uoN6s4yZd8cqoKNJRDETLO6ItbxkEj5RxKqAR6fvzWdEfKn878l5KUYC9Zsx4DFew
/uyG2M/cSZ77KRCou/Z7DgTQuE/AGQ3JmC0E61Dm4FUT1SCFPY+vqgMKU5TW/3kSY+G82p1MdGYb
q54k8H4jOl92kz8KU+tqQ6J8q+4Uarr8sgI4qGtM4tsx5c6mjQBWGlOSnf/NYsBD+Gk47jsm0T/U
L2FeBjjs2be5Jd8p1lUZzhXn0TGztdvitQa2LpkfxitJnGcBiyOibWtTTiKzYAc0RPJAZ7/bJygP
Dp3pMdEQaWaylubN9amHWANWH7xQCh0bJd9nFZSvZScHkpbWY6kN8+ANbegqWlNPEYNOYeHziP3D
cJXxF6CNsBP4cJvCER5vEUPaQQe3izslPE8HoPKmyBdmJB6st4Im+1hqT562GAhUNnK8CLUKCoeb
3YZnjkO89OmsoyRBiM/d8KPyIDFUwHCafI4jNZhZlPt9rCZXScoWHWCoRdgbU3vwMWUdbe8MWe63
ZawtvfNNxi2ROzZL6lAP08GLMvXLfg3CO/4v+iimB0aWZm3UZOC73gVFqbN35Dzp3k94GNZ2SBsa
/uVaZhuMsxINtKo1S0KppSbesLKk6LJqyd7biMk1lMrsH9uVqCtx/6y0pWpywJzJxbAiPcKzqUs4
4Lr/SeRdHbXajBOY/hxdSx7PaOvq9QhOn/5ZMyQWtpsnGNCz7qs0YY4zoaW4c4kbRP5Mdw+NI8rv
HL7Kv30Sod0GrilQ9drGtPVStufUKQdkBsIAtWTWuHvK43rEVab3wRQqETojAZwzofVoztXesLgP
Rpyajmvd8ONv4jA03MmUgAIp7gs+T6NsbMC/aMgjn5kQD0W76DzwWYF6viWiae7Ez4o2TMhEJ2Kf
Rhq2ncYbaxhY4ce3DrsFbKE5KN7WRVEu2U2JPvB0XxODVvymm+GnolELvcsM92XzFcqWJUf++CUr
cBsHvtECd2bkNAdTYq4xv0R77dBubaIx3jEp0Dhks2HyQzCjsNdMh9l6QUF73JCSQjmQsY3mECWJ
T/TYCtKbcg5U0nMAU0jg+5Xqv0i2ZjqQ5ybDTrO3cWR2s2vEFONh2IstNO2cXR7mO9pvfVXaPN+L
xRNiySGKDg+wXxlqBQHzdI6wMCYW4IMf+MGWmKcbXZ2Mbsqn2QSXwNLS8GhzfHlk/hCvkry2at6u
eqZWttVpZPn8Zhj1KgeJGqSSIDkc5+QaHz5CBKki30TQXQ2Emr3j3gHVuM+jQIqBuuAFSLNVdbgc
dA7nIss3oE0vpGUZgMRZUeurX1/5JN5UoFULD0mBU1J7LBsmUk0JHmRE2NEz6hAzv/z11c8kZp3n
yZ6bSFm/Jm2tAiq/fyVHY28LV9Ms2q1HWVVcQGfahpuiZh4xPOTZ1n52SQ8a0T4j9V+m1tItGMld
0Y4AFcGyeKdNK4jBpBZEke1WDPdE26lr3FiKeYy4jevnQolqHKgOnKpzdjb+7D/W5VOQ3Gbem7gl
CGwsIEKmoeUJSLu3HrODknKUEUB8oL4g6JJ4ZiXN8T812WdFoJ3AlXaaX2odUetGMMPvHxfA8B6U
/7ebpR157VDpjEnNFInv4tPcGxmXrpsWUr/8QCpE98Shj6Gr7QluRj3oS3JFVih24dTcoNaVjso+
AqC/+tFJh/LXa9euwuGsmXav/QMWERz2a5I5nmoFMxFq52/yd+1m25y2jHVLLk7IYhx8WT2mLLki
HS9QIqWYS4F/rkBa/El9fOrpQEv8UKqrk3LNJKHnzqP8kX9UFNxboLWCNMLodls6VKPtE905zrYa
8kwmvzP2bGyUZryylPTkO4FdvgOe9+vCvw3Lus/rYk1hrDldvy4ZDR4fNel05DMJ/9EnNIAFTMmh
wL74SsfygtvLWfje/rsp3aBvPulZzUoYyArTX6VzwhxfLcN0S5OGdAb6X9WYDZAogg4ZJepp7K2e
x5OoiY23bRsUVPTBiV5kBNVu99leKxiYIebpXVsNV/a4Sehg9QX7AgtPm7FFE6rsm2Js8OFj2SB+
rwQTGm4o2BKlyP5oyQPTwmsfm8kGQRJsUADNRuAB0+ahy52HPPf00UTtopfSO7sDEt7RK0Yud/3u
T6s+eedyd10doNj5KoyrUTiH4kWFgSdgjj2LgSZzsVqPYNR8ecIWOcofMEXtNnN+NCi0Y//41JGf
hL3+yZyRb7/BUbDbfrzzZH9HxwvYDQCSRIhjvMwKaPkQFH9LIxXyGeZsLL8Tawi5+GGPqgVafvFp
j8RLxabTCEHtfwUwoWkiX9BwZ5uJQsgxKg5Jvt9QFxj/WxOnb5NXbYpaNhErkzg0r/pfvVAicTq2
FuYgoIW4LbjwBnVBMLisUzq5OC4L8+lzxvJR7dfc1SuEL76yQE6MIfF5v17MVoPfvNIVn7Xcd+6Q
uy++5m1p/oY7TUxdI0hJfvsTQ61pvR/QT8mvjXoQ4sr/nFFp6P4iNjw/QEkNYW1AoNteHJIxjPQs
m9VzTpYXM1hS7/EXwL4zAhMo6PsSfBYHALlOvbFBIKJvxtxYlptOmSnIXdI0m9xzNhMHdF/hw2tO
wFGrBYcX7soCIu9yeKjaLl3Ka0A9z0zZar+gXixHVML8R8uRms3gweggiLl3M4SeenfGXwHX05rs
eVC+Sw8bc0N10hVN2oQt1DMWBiphZOVhIdY6FipkNP+cNqZrx7BTzZqhj1QxQHBsvVXaq74b1PcA
quVEXAahCfCvWiBPFlZKXV4NVjLA8lXHuSOzDkvYZ2eNHRECiB3ooNmpbf8t06+yuTOhEkkjQ3cL
KN8LB2IukjQul86WpVlQdEjfuNlAFPgJTa0JBc4KpGJ7EZ8SopOxqNkJ87EiITaP4e0KU7eTpQKR
3Hab/tsdrsxWkbdfWr/tXi93nInS5sqBfrJeCxo4aNhSJCtUsJvydloT5b6rV7C1b7oL+BNizhO9
nJYhB6n5ZCz3+loETT46yMl754AqF1W2buwSuOysrQXuPoR08wXT3LaM/TtoMdpbxwhFydQh/PWZ
gmqRAd45inPtsw7Ezh7qRP4K2KCzTSsD91emQjrtizxOka9S6zCgt4159+e+LcxSd3TpTNGrVOrj
ek43Z6VTdVH6fP05d001+rfn/mHv5hoCt2tADg9GtSAhh53H8ki/sYxxMBuBrEFLDm627mg4zGyW
Xb20RtwfYkXLcKGzsqYyIEh/nzfygNrG9axEqWfez3jWd1L+RrepVqY/J0tQmSqFqUdz/ShnPodf
3kWezOsyijHzFiYYmmYNiAIFeJosphS6TnBbuA0uzacYQnlxmyvZGrGuVyAUkjrhLaQM0yagGsvq
tcRgYn+3ExmKgCa1uIwAu5TqBmM6N+PLa8QKx7WhkgBewMx1pLt5yg3oWST7tgH2/8xHJ83ZHXoU
HhgwLqyY+JMprV31vDdvcHmE6lTH3ARzHRdOB7AgLMobLL/FyBtC5J3pTI1YQZ0dgbOEMlwdL0xk
/sY6gD9wtsZVF5kkS+y/UemOz6dB4OlJwpUvrkjQqWuEo7ERLd6QXVWIVxZlqIO3sV3S9Z6OfEmd
tSiQzVSfVGBkSB3/KkUdSfZl3oNKaq7lMRUG7aoYg1mwovJ+dNdjBeZgV8mkPsZN5tXgIUOZ84RK
ubuUTpBgZOSVFjWUB6C5aisbe5+WnEY05ni7dFWrFZIqdEIn2JF9WS6cMGY/BaPcmqQBBFyETPW1
fv5TZcGv9+bifI5a373w5ltwrXjhlBOdU8UUR6D/7jVlsNPElx8kIOKMqXRNQt9rYsDgHtEQWJg5
Ces7V67EHGE2/r8ruUri6yw0G1w+ki79Wuqrj01qYZiuKTwRr+f/jYHYugNpALGZzMT2CVXvd4Pg
HBh7kCpPyq5VOC4xYNEyE+v6JuXHLFQ3zUMblJZJxgyuMRQ8KD1yXslqnT6OJaSlDmvf5aRWCy/N
RVejqKmI2GZXf0OeVnIAn5FjUNAGb5LQ+Y/yWvbJ5DyPiK5SCqsh6hUbTgdkldc2t1lVRD9/GDQ0
Mrq7gErOL81sKcyxziq+DQQUrm1zbxl+5ASuJ4DGMrSHinYneVxj7CADC0lGikl9jo/oZf+S8BRR
ke7PExKp8K67RQFvfQGzZL1/F7FRwyaLnPQTmQq/SpGqinZNYVNMdB+3r1blY7Hd+cazPWqoFZ0Z
102+R3fihomzJCOtvOf3VKaSTupcb/HL8lnTUb+VGTZWpXtcQZx8M2npIafTByxtq7UIc75QD9UQ
Kx2uBZGaoiZStMZhJKU/M+aqwEKJkN2fvw8Uhmr/yOzI+77bebCXBv8tdc5JGGWxTLS0C+iomHaD
dAS7BSrQK/GjFZ+J0Xl9JLkWZ4G4USrTxtBXSjrbGjE+e5k0eeftCGof3t7Uyj3AFIq/0asukFvR
tOQHMfannKZt3n6imAFpg3A14QdrV70cpY0548ngSoscTLyFbQs7UjWCECmsY1/GoHMbz9YdIupl
ZF/OGscgHTRfyPe4nwgqVwzGySx5bawtICJJ7O4my+kNRfnBGN/brlLEbKrvG+npRl3CdrxhMa40
Ip6kAmnlrZaJMc+xS+13wl11T0oWQI1Cbt+uv6ZmNbH1rz8cjUjM7rPEkJwNx+dsglFxrubT+pP+
qcZY3PiTPqaVb+L23UY3kmySzrw0W9gdwahRat7qDYtmQyjU0wbnpZx0Ilz0LsO6DGtZZAb7yf+4
jQjpJIY6eVxbJpXxs17tN7FCP/WVnbFDu3vPvky3jxdssKprcBPIb9nHboXIUHwB9si1tIvW1VSk
uTWCDauz0fHmfghiSkDPwBbvUcF+y9gyxnu1aftbCX7BeO572TAhxt/6gscPVoLe6Nc6IrpPKsS9
cXaNPHXd7tDqftSqYcY1VXUK3JWZsO2vnu9PtjRyA/kmdsOjvnN8Z0wgperbdwh8z7vncoxPlZ+n
3kcBopmVjT1g/oJLFdvXZssaIkPnWo8SFvux4t8T8CYcAdhZ7MVz6lH5AB65AOdfu5g9OCDgNjx7
b46aocRWDjrkeu6JUl4KlrJpD0VtFLu2YFa9+W1Do1UJLohRQ+i477GiVq4yQpbNBX5/LPzPi+zU
3os43xkah/aGsmMcxxO/GvCz/2Ql2BjRO4w+H9K5LpG3KRwj5W5lot/Qxz6cGCBPtcHdvy0j7uO6
E53zpC/ZRjhsKYHLJ6fNzfQK/1ZjqxBRmywK8s/R8lwArpmae2VXX5D8Gts6biaHuvaVjJyPZDtE
HCatfhAQyde3O6HCPAEegMla3XLUPjQ2Ajh8ztxT8GichJ7+91LRR4TjIQknXJFcym4MSwZ0bkud
QY7e6xpjKIH7VllFedyRewE7vcv3mt0PE77k8qyEJzwRjvwpsXMZrYptuHsl4ppvIZq11pD9GHXr
wI8epN8KExuFwhgMemlI//ykSvagWvfXs9xGJyveoMy7QIqfJ6vzghhr5qCTBnMZVHl31Emf96qN
GId69pSHFejXMux8sGjtZI3qyVvw52B4S4xsr3ju7PzMaCrbf+6ksbj3aROlAis67SObIqlfE3v9
IY+JRUIRSjgzCfuaiq1rJftZYWpYtWqpX7wga25seYP5z0D1oVm3IdVNeoZ7T/zj+rB+P4NrQTh2
X7PhxCa1yK86XlnimVmqhVzpg0/l+PwcNBSJa3Hceh2NglHvINMk7ms5skNBuGvFq3ELHP4EqSx0
bDPIGxZbg0bThg/fP+PpTis9ifVH4a5TZiZTaFdwv3yBKF4T5QAa6ZLWvQsh6zo1M6igL7xJei2K
6hlVwl/LoRI6nzz9GR5rcIA4mxGJ4chLeRlgbvoUIbyyPo4tNCslgu5p+6A6eUctjhnhF+DrPl6o
X7OC8UjpjGJW14HGBmiBpBqvKrgep2AVjifeU3AKfIa+8L1pB5m+2CxejFq1N2UaP/S8IgbtLEYi
dh0g3loxGfa0T1SNdlv2pQ+GYqX5lWqw+gKCi9t03bTOlZ5oY2hTJwP5ED4c5h606kA1UNuv1DS9
MXpzgRzAns9ak2zmYnWsWT98uKLUuLYzqIOkCouc7kE/luA2iRjvaSfuHjVSVDMlUkXPodXwz1aM
fRHfyYaCjix/Kcq2I+cq03RNtrf3HC3c0TR/xcOcmzIFNKVkFo2PDnLT3qfEfaiQJTBoEZNPdDZc
cVEete2dUt94lv9vIm2j3FOT/hr5PohwQP+IinZqOCmlQ8qfGs+fN91GZA3NBhl6nOZw0gytuFYv
bHeo7eO7DagzBOBCU3SNv0OabLhbuUXkzFo3pQ6QcbpiZhHG7skCQequee9YCCfOb4csNff2Xqaq
MniFRFCKx9u+UxJ8m+X6cKouYOKx0mQy3WSbstCPWsbNdAwn8VwijJL49yqSVxrEcp28SjwzPBjJ
ujPPzTp2WQW/RuSjhoIZrae1IbDea3TZrCuYt/sK3eImBaS5U7Tj4db2rbKSUQQ4vH8o7skKsefL
kVzc9iHikcK3LMBLwjiyC/m8iIl9oDdfQqjZRbaN6feLZe4ZnteciwMB9ZU4ttu0ACkVkgGjuCoJ
7M5uMnKi0U1J8mxIV2Vt6bkGPs5wYFcXF5S3qeBrT5HaFt4oRBvodM3cwrFmtEvpDtbFFfBCXt5K
AmRb/ANwiN2cJVAQI4gcImbXePtv5s3d+gFusSgLU+kvycXNYqyiLB6BfuoNWBetqY1/swhg6wAM
OotaDeWDB0BshhCAKdOafw7js58OvXomqUA6NEbvgFlPJrE7TxWPByEet4TK21exWk112Qf+dF/k
ZQnDLlcXKY66L3wKLRHS77xJ2f880inpBtCupxlyaA4UbejV0pYHr4HsL0Rv6XVr6RzHJPaY8gCS
IziKIKoerOZWAIFLK0f1H0vfes48C1iyMfsQiBuqsY293Cbh1p1tioXKNDBDnvS52AlCr/A4Bab+
MgOqSqjo7LHpPlFn4XMru1wjp4Bc8fyboaQRqgJZgocsJaIx7KZ4+MzeH6HM2UPsShQ1PhHIrqIl
TquAG67hEb5/09Teitun5oXZYkC2rp6XTzfcF20z4MsHVZMKE5BgiokJn2hJAtBBESvjFw3nMxD5
AVS7JNt18yMuq4OK6ANhEGoBibWCL81d0pY33pVOtFLxe/T/0EROk5M8iXRODAnOk3ckAJwRV/xi
69zWQ/on7fKJ7ZXcRPx2W+AcypV20ip62lijF/n3OgzofecBQBQSpzjdEhSQmrkcFSwb7PR97SRj
9zI42xWqlaa7PvuMTL0p2+UJcnCkmND5S22Bj26KGySloKZ+aCAE9xWbtUoUtFijnPZClC7g1oUT
N9rxMuyHXZzWnVHj/efZ2Lfo4LUhDc5xZ05X4q8D0TqJ9IeDXpszAl0Udj+dJl1ReTzjJyikM7KR
rBwyeW2e1eFQzIdN+K1XWbG++phWSTs1vijXWWM7/Hccbg5lyvhrqMnE4Crj4Q1ZYy8i5H3LnMWK
YUWqwgJk5qC0pmxT2tr2HaC9H2VL7d6yLSOLSmSC5MdOUhKvm36dv8VFAHzdOIgnph3xENHwuiMq
qe3oFtvzFjDNwm1YLy7KvIDmRQJlkU8Td1FKWIoL/qDv2qoYd2To4cra3m1CCbgFM2sDibLNiQcm
vwkYKIo+rCGUYoIqAxihZ2XEZOkcDEhQCcHZQU+yEk0K62Yfwo3hnSoR6I+B2V+Kgsr6W+0drcOc
mAaHSDNnnZODj6kZUyoRJKU74h06ZbrsEB6aCzdb2crb6DBZpcExwHvebyAZXswZ/x2wrMLHH5v0
QVah7cd7jB4ky+2V3CeCbw64yTGMfOUowoFrGMeLNDTVAjmru/w+KpxWvWca1ixCmi9GbaQvn/0q
GClou75tb0YdfFKcRzxlmJhqlvn+FMLvtR6RAQVex3QPhF5wFrB7iBRvrYV28w+Ds2/thZpsq+qJ
bE6/OSD9t5iJ6AQUy6G5eXSGahdJsz5v6WtoraDVPI8Vk7QiJJ+T6qVzN4mtPogHrU5U1vWFtHj2
q8Uv81I7+Y2eBY0TC+yhrTRUFLEf5tse8fbkgxBBiQJqygrUBATZAaEZPIHf5GN/OPnfyixFXHKb
7PRVa/6zXQS9e/Ej4L4UUzvfWunQxzyBMoIc0EI4mwvdydyI1ZSrnpbQo3pcRXdQOuJr/TgY9S8A
KkF0QKmutYPcoqctqnrW1G13MAxplurNV+3BqZauPHhbnpmEAR+OYmp1ag1ac+e9S5KShheRlo2O
gtAm3NK+pocE/FQ5mrpgX/VUeXOMFcjovxqRE15GGY4V3AZEbvgUJ7/Aii96Wk4H3Jy/7A/q4e7k
yhBVW7FwZucqJebfE7/WxMkfyoOpJh0o4ScOm09ubvParJTdol/PwOjk4c+6CzEn3eLGQ6ERTw+Q
Xyk8moBaC4M+MztVTcS0swVXnfsbob1SzQqSzxSB1Nb8wekHNDpQH7SXHiK4N3HncjbnPn2MjC0o
Aq7QBFLmOWkCRsUcLxg3rPbiFUPJwQyHnBt6Vi7Jtx18+DCGgbKK/eyAi4AtaZn29luPeuWA73dm
7Mbeom2s12jcxNI2EHBenVRPApt2oHASrfeczyhTc9eDjo1pIuMMOjqB2CIvXJJBsOvW9c0KJwml
odQJ4LBFJiHeFGIJZwOXodgC6gAHiuTRf/I1b4xBsOhgeEoILPm/NZkWnUsKsqxTorLbDbOULAJw
Er4oiys396s1Kgh/hco2YsXTg2zK7f8Fkf1t9xi0gYUkwg4G8qJxu36zFdbwOV9qsuUcQKc//5RV
qYomPAKmGo7YHwJpuGq9tBCoqcYEdWVAjwBrNoGIXnJamkJAEU0mSpqRsLRD6Vu8awKnCqCjgKDN
KLCptyn1M/1ElZ+bq8SY1v7+rI4b1vmqvNK6nTSr8kyMQN/5wTTNk7EfyQg/Ffd2xI3DfdgANYaA
68QcpSBuHQMXQURphR/JUX6iaZNQIHPCJhSU1btH2cDPtW1evCwqG0gsE9zPnBcdnS3h/rBl3Z10
MTf2RGA4fCXwomdxNM8RWnUsth32SVmw63FVKyN+27NsIZHtBRunY3J7lwBUhpNomdLOEg5Id8AM
OwddwsuQxtQaRr0bECdepT0/Lnd0uMjR+awLd3mnmkHYTBXZj80lb5BGOcfGebbW0GogaSNa364R
t8pkcH2+s9a5vWaovlO0Wn7+optcHKzo+6J2BE7/TxFkP7duoaaKP4YGAyskix2BfAN+FGrGg2u8
gbdh4ExItVTj4hHjaNfGk+R65brpnn+M1VVa81SlBAUHvNsMoGFr9QBmRcnJmgIitWuwOCatY2hS
Inr0ZD/9QPUIkQbDT1t8BBHxIraoNysVV900Tz2alIBkjKqIOEFNPQ61ruIyzIjG5jiaNeDXxwir
izBpRkxRYHkvUwDNFwX4h6Erlt4DVoKVorf89SiuzV4UUddPtuqYVWqSxPBJwrKvCJv76wXWvS3G
4/qLxnICo4c0VBIuMHEWqT7fBIlWa10mMh13QGjyMLF6nnIMp8A/NZ9TGE78Bp8k5yr2jRACorQw
Hlz+kDgWD2UebGwM0tZqDAKzXC8CHb1uIB8P0tzqiy/W80Nsm1V5pj4AOkUZDoHfNakVdWiVleWb
Bro3hup60QNz7iHBW5J/Y3Wu3JBiDcbnXbI/zJSvBgDNpX6yBNgoGj6GhQBhiae5f4/yo5j/EtqG
SotZBSOPzMl1zk4ess/xWkIyfvhf0iqjtJgp/+wTzu0zRPf2Ro4ismP1GIhANpVcZEcpuUt2PJVr
fy3b0Ft/TjLKwvSUyBX0CYGEKhyBVFuFXP4HgRxiDDBdqjrO3N6CGZ1PaLCe6yrWxcdEJKKi+GKj
s/RUM8kjxD37UY497MLNRWQOXKHl0wZc7AeADloKgh0q5RvKOlvvfiQ1ulMqCf17qvduylaDeQx5
VdsuR0mT2Nmxikw12PnjFNWfhUxXl2WlnU45n0QbmuZp9LCh+zfnNrSFaASTLbml2Dvqo+g8pHSU
R6/7c2ZpyMiC7Q4fVXXGHcyIsUJxTjazVqPGwynfP9hjbX8ItP+nVZQ6SSVDUxVCsWQ4+Uae/7rW
1NYNM+NkWheK+E1p2cvodqdISxRmZofIHwQ4T7R5stUky6Pimzz+WIqiqo2YXs+UvvMLrhPi58La
dW/TOVlhR9rUhtQIN0ODwzqP5vFJtHWQIQfQpfa3Ao/xtuA0UJz9DNnSoFzhR+l/nodtW8Z+QvUD
WjW6qYpcqvycp748Yub/Y4Y3SF2Ps4HOvKCVgVFRxHJ1RUJlBPsCUC+9zPsdWoBG9wRnsJIpZbVn
WVCFXNL6V9R/MfABfIfHVrVa2VMmWo8B4m5GSNZmgSa4aTMpMEuSZZBpi8GRB5oY+pmDfV09vQNO
7uJlnras1BMnez7bEws6GSnvTAKu6nfdprPCsbgxMbt+QnIVVA+1rd4qe0lhta+z3OMXxsN7/Y4Y
eEopDGW0z5hEgmgv3FF13AyjaV8qUelfIrQbReJR4HKxHIo3tmWvIhgzC4fRAtQtDeJvAiYG+D6t
pknhVgKkbe6Nbpv7bBMjnmBRaj0J0Q1yrI+3Ov+uqu8kyj2pvoeaoIG6iJ0NUzMT675C4T3WExOf
U3vS6mlKjbcF/mWJ+Kh0lsONbQyX6HKYTjDWq3ZPpH0bcoDD80uRWQ8xX1v/jSBZim/9aDcvAl00
oKin4o2xIG3x4mn3NoNNapnKscCM/lYFVKeevwpeaz1LG2qey+A2poTxCfo5Z11pU+ag9i4ePA7e
kcc5PZZS1u7hx4ZUppdFw0PiK5v+rj0ahyh3VkjMVlgLfN3WzbH5Mjph6fSMPPmvr6XBMBpPKXRy
vSHZDN2gSEoIDcJLoRosoqgIzc57ft0aRglnhPK7ULxoO8rrD6K3kggyn2qTYc+53cB4sp8bUbmJ
6pVWX2wSujUgoP1oB+uz/DNSRFkHVreTlk0qkmbCzYXNZNgdt2u05KgXYI69jNIquYaK3GNCYHkC
WQRA3jAti+5axhHpBTswHFutYGgyZVFoz3LIoCKvKVrddAPE5ITm4WfnUXtTWF0OUkc2xfSkQpl/
2ajebxlvMqMNuEG6St8OlLLTbsYYpPXUvfpdA5Rbjl+UaSxRI1+UTA8SSPiKxppNAm/Q8a/M/yPc
sIfDJXVUFrPC+jFNY51tDdBZDUNVkigSp5wbS1kSR0wTI/ljz13RiOZZdw1Mq9rnD6zCfREq3viG
hQCCWKLNjsxUcmmmzNBI+djYPXsyBK7+/Ne602YLVIUQUPpJBuY9MvowM0NrgY3AcffGGtPRHirj
gbHClmWsV4BTemNaNc5Jrs+2UrO2OV47MV3vNKfYH17SRKMZThj9sBbU4XjvWv0RLFdNSIoTsFBo
fVAn3s5CiLZuHYG1dqFMAb+gDP/Y0Yd7XpmBkadvqUuc6hQwdiM+EXuu5GiKZnruODG/327L6X8n
VSDUuAUkXMF57zvXe0Udm+mfy4Zgxnn9+/VrOuLopbCoLKhE34QQ9BE8bLN2ORqIRH2s70Flcjyl
L7MCCIUCfwx70U/xgrQl3F/OsC/yfhskanpibVYdXwWlPrYhTYq9ssu121722RqRji6NRlMT0DEv
rZTWKZTkxBQgW0zMVC5ZlQ8e7K+wvYdAGsI4zzU231XYd+urB+G6wETDk5C8H8qMGQnHmVYFgIJB
it9Alp74KEJXcVQqoSrBsm223EGT/r5xlYXromyBpXYHge/x4v+ubF0RLPOyfgSz3+9djisl/MF8
zzz6iiFjcuI7ChSRDOeCi8JpdM3bOBMyC/yLDL83DlZbRM8iujtnL+SdCICfq41xdR5TwztGtGdY
tyqZoDpszJSuP+QsjkH+0fDP9eVlGMEg8VcdaBERgYfcO8rXAbaM5acYQCd3QEGM4rqEw/7zcjD+
XbM5beAL/QnlXeaaWAsS1bxWWFs7+iZfLHBAvdmN+6cWRdhPr2qZOvic1fqKgcWGTeKep3/f+vyk
rc/hbqCAUjOy6qD3Wo+YuJNCcKgu7BRhT3eWlC6L0ruHmfPe0lWMyB3TaJC3EYoyFpw2/liqyQBV
nHKOAOWBFKclWvEejXgscjmiXMvnbmW2ZwMzPVleppyAOJ5kPpKVzSGp0zaPidbDqJeG9yGqwDcs
RnY82I+B3ohVOBFgA0kpI1QvQWSSw0kxRUvJkxsuW9OIl/X8371GlbTCCyF7QZp8bLGCIAGebk4e
E5dZPEXTjXQcBm1QAux2QnNSvAschIOzmYP1PlCgfVgXmg2hsunkDeyQ10is7bRM3dDpbi+FRaBu
lhdUJPhICIBIPJUaPv7P8VRRjLAd/l+ch9LbK6EX16Mv6+vRfsh6iQtP6Sljq3TScnBmy7YtB+C8
tj0SL77vEulTU9qg4qTQi4vyvzSxH0S6pU5Tii1PdMw2AQaayVFpmDSAg4Ol6J191LX8mLWMVKI4
L1UkZ64fzT7XLoI1pHhI24gpMkHVuvrrWSOfWYM2/0co3PDUWJqJeG/qrwDm1nZj5doNSEDDjsJn
rjBVDBfZDOnAx3dw2h5eVNBmFg0AV2AMaCrQbpO8bhFxInGKsDyxIaZI+Ql/6X0TeubMr7Gg2kNf
qRgGgAtuTxqXP3IGbnu6YMrVU90kBBowHDyRl56HsbvbWkmHHuNUNKuS2ihN73eFg40Wk76j2uvt
qQVmstCbF+4w4QPEMxlcfpCMKwIX+HIjlLnqIjtIKqeDrXXKdCCMWX73qFs1ck2yKvXnrO/qZX0c
I+rVTswy2bZEBeKzti7Xbfc9XFkSuhLBsjcpdVJ6ux+hNE3uLRpBJkJ2NrKNzESN2A/Vuix4MYFa
5u4fvSwW3KMudHaBPNGME4SqxPj/9r0REkfNdMFSF0n6dGiHqRaE6GJ02yPcPDcaQ06TnY9yl1Ke
lfHlxKwPruijUPQvu9hWbBXoKIuPuJxsuGvrF9hnvXbtf2ui4pzb60F5TON7s923+fSU9e2z0tIq
xCC+nvNtVijIh5GQnFFPEnPJCb2Uo/1ePElutxSu90fSVDpJ/1KF9j5dlOr8m+BoYxrF4YpvxiHt
g0u5zdccaxt2d7YEzCADm3SE61sXOfawvyS0RjezCD+wGspfv995lHIkntUI/GBc3lqgWOwk5WD3
wylB2/gjON4Y+KbuBi3CY4maUkQp4OnnzPGxnZ6WXj7me51306F+8nWycJXfCg2azNQUFKoSMXST
7eyNQ9REgJVPLYj7bpsIb0M68dpyix0ODibwvlaHSQOdNv95jpjlQHDS6IY0Hoeds6ecZwpZz50O
ds8k2z8VjXe8CM41pKN1hRnhZwVw4JUMEqOcyxJRAUAQVQ0RMG9mrc+llNQlskAHC6gVQ6QeYKTq
48JbwVQFPi4MQXyw1YHa/l3ceJEntijSIVhZT9RwuQiDRJboHwhTPBd/DAfa5JF04Ecy6CrK7vOf
Anzr8Ni6+dzHVbDz4NQ632On81VHPZtPiejTcVvodLuMrEZFz/3hS/bZwY/5HSgKMZRAoLmGYvZ+
UDGzLgguSp1ZZ5dJp2k4t2FKx1fJ8ypixPTg7V1YxjKwVAPKSn98nPoGl0BNht3CG24mwc1XGfDu
hU3RKxwDBJMejyf4FfPWBaqcuMAu1VDiDvMWrRhb09yLfvxroeiJA0kUQNwJWfaowd5ZgGKn+6lM
wEEG9wHGFPk0dcwNmDpubM7Z/EwMFQJ/Bl+eHgBT956CY2k0F7QvBXO8dwbKfQRS0QhaEcpcmtMO
oTXOI2KS3UO8Ufw6joJrvAK6cP2ddXmerNGOxjf1yd8yhxY8G8yF8goXu8H9LXIgAqg178hu2o9o
T2ryMUoB29Pn3YCB+DjGmqe/vLkKTcJJogipZn9K0se9HKYN4eIX/Wd0RVxfZgZPZt4kFkrhaGu7
JbWhLlsGaUsStHFvsthHLDinCtbzrDTALFucyNxGSXysdGkKoqqhtgI87OijMhK4HCyrqdNubY7E
qcEhyf+bcO2UyYnMjT8gZBbnMpV4ZnRpzfTwUXXYrn0OukqApT8fatPrjWniybUFcA0LVzi5tEMY
kdApVKm9uH9wxj9JgUP+QidvmSOsMkCMFXhSYKljqIfTT3UvkrIKo8Vp9XzSc7NqkQxGfQjYoErF
3lwWQ3bnmSaVrV5XGszfIMBhm2sTGZTxmtr/jDlBoZvmHZ5klzGKlomrx9XshIn/+W4Mf6sqKpXL
7FWPTrkHUdxH37/YXCLSdUrvenfb3lpe7gnScefZBtZSlwYVJDGzIg7w6IzNwl/2SN14yMc7Zf9R
zMZGMj++yFg+d4EGvkJM9/+wtTdeHGuOjqQpj0LvFzuIbn39m4DOA4OyZ9F5V505L44h10QQ8Knk
+DbR+CwP5hUxb7kQb7Xfd+Gehjxe4jnkfsfr6kK6wRAofqwW4YsZpJWovgbYJ5qfgBk+HpuHgMfg
I7SlpIZsoOQhOvccEo4mld5wDPaqIzMbo8QzuYDD6xumvjhAjrwD9ZsPPZa1YXZt1A1WXFVOpaoz
isajy25imOfzcfpVe9rcoUR7jU3xjQpnBdCyH5ApOkvmPZEud51I3pRdrkVE/IigO2AaQgnYBny0
I9gUUGlAtTGvXNE8yCOtnASS6JS1zCkv4mkv9/NUNAJCmKHCLenBLllp46//fwVpzzMnqjnkZiHz
p2lWefsUjpSJEO/7s+oS6PFTmsmsToN5H7DaxqKQYRVmyhPSWwctCG9Bo0SlCd/eDcYcCbzqR3oc
wz+DZObYP+CaAW3SgBRN4uDolomT6kdqWUth2c8+tHb5kA0j83FoXd/ryTs5cR9hXmnmANfaCbRA
0elhvxEZ/KSsImtm3XCDxZLBG8nEj/3EQ9K5mgBs2QNTcTrmw09X+oW4MwVBVrLPenktgt3pXuJ2
5rD8VvqP7vzFJXeVVy37D4+8Kahl/MnNCVsKCSs49bAkLDd1EWlOi8RAO+URzdG+6MOQsUSsFGHI
7/ZqORIY+TcgxwBiv5dnf39y69q+MVMltXKYyB3PiD4DHj/+Kzu6toZFVmieBOaix9yU5M/bQvYc
X8WlXrbsNG3fIFcTcnKgupXn1EEvDXgDqW5y6rIomKm3y+3IuhEIeWD/C+mvIP6myR7vr/zf85S2
ZaYGx7Raz8g58gxp//0gzYj7znbFyyDMFM5KNMVWTN8oBKOuG9Ne5JlE5KFOqOdVMAiuEnjkip0m
c/3OUEJbv1HGo6zKNKUz8g0xy7W7CejLlXpcSZMGhqHsMv+lhEmEmRoHfKUsvF8GUeOZwbvTF+r+
abnQDtWRE/s0aANFOI5JpFU7ysH2TCtrE5eTBVYRFdJRvwPAbuQ5bwuk7rrzbyl2Wo8vVaneTW1U
b4SDnUpPydcfyXpjT4/l204GcY2GJXekpex8LICfMJkpQRpQxSBnVJn494Emn/5II6R1vq+7robM
+jmZW6yUJ/k2hWU9yyDcVylLVzGEv10QqtZQ7F1pXjgQxtxXrBXPZEiD6xJVeW88Naquh9RpYccH
mG+4HdG7FhfsLBwZwdUYZM9+GoVaFzMmTGU7FeAz02WMgMPmRSKpm4s3ioVY/5mBExlsJucVBUok
PESMEJu4CU7G2n4FS2W2MbbPCohG8vNCjcpGcgqm0k7FYFcDhPslv+QwBG1K5tjVwW8WPz+J3Qbl
iFmUfIv7ZRau/DeT/s104QDXg27OhwIEvbUYz2eQIYFMsmz3IXT71DxufnlVWfu5Kd5PkM2QO2Ya
O3NhJv6jYFRYdMpf8lKPxTQ+zybWyLc6sqO8bx8+mcJwXJHJ1fI5k38sTVYIvISlMjDVKDmVEPF1
EsSnsDbasFk9YKJ70Dta+nkOv59Tb0dpI0k0nJQ6VvUYUbVAev5ur5FOjykx0S8mgBzwx4iwoR0A
YHGhehADu0ilN8aUMnw/5GDz6K+mxRDky6J/2brHJ5GlIi12JR6dG5eOkteKv8dSns8bvkEDb999
4r9no7zyR4/1ricd9UVcGxr20Il1j736rEamgEvgsazTnr3AEcPKHKBkRVZGZlwzyENg858N6dEY
jR9xWn5yt+gXOl0blYdzyE1+rM5RKPWmKiku/9km/Uq4SoRZxuHmYk4JlO61xWPN4uZZiweLjLlf
J0dYd4+Y1BxUoDHka+D8NUcbD1HbKaCXKQ1njWmKNtZYDqTVHoDNOuOwtOxE3c+mf2y/w9NWkMW4
tTZyECon/2uqcvPjRDnzIILEvJehgeheX30GZh8rf/yR0dzj4phH1FiDWtUKh1ZG/jM6XLJzLwus
n8Hu4734KrSeIY2u4y8CulW3iB7IPnpjKQxHoDGKh+OfAUt8jqWoTkAOHGGJcijiUK4/Yl3YYQ5b
f396gL7257CNwpp86uLuK5OB6teKn0IhWgXQrPaSTSxHB0cd9cWQPNz6MfTGxtFmcJI/eZW9IiO7
Bd8zOBSoREApuIC9GXfO/pUEZOzPSsh/rR7G2W2kdFBeYi9ujnAixx2YZmTTjVW0D1et1tAUJanp
SNOcktRvfuAKNLcCFKgLP3xEYkBjHynlh6Q9btaEpTCP57Pm8poLWS2djHiC7JEAT8w41OtAqRqv
wW1FpDWrzbVb+4mlpVzymoLKtXN/PDfkI2Xt5Drlg6uDjjAygQmk4nbyvhoLzNrjt5ZbZcXh1XuT
FfukDheZeM0eeu96EX4m4fLFyjthf9aHs+e5Uy6FDg+5+g3ZSOHZeJuAzjbniJVbzwG5+baOwhO6
7V4x/fMDorKz4sqQ4WdUa+IhFadvuWJkgtCue1NHNDmsGU57Sc+XEdo2XCQbNzCn4ROvL7lLLKzR
CpeVY/uui8J+vrbyzqyO1naSz0gBV3hGwrxpl6b7gqblbCYIiYfrrDsYkVuj7BoYJqCialW7EM4o
PS5wK4cKJfrcphOPPEh6gzhswNWeYR34mDmfA7L1FQtFs7/wj9MbnnC452bL7WtYSKr5vbfHvmhG
Xk+utHUCEyQJfjAWKxW39UVuBOz79UzKogiVoZxn73tBwT0H5Sef2qC1jOgJAMf5GOOj5BjnEnTN
H3IaFusw4O4fQViLQd+RK+6rw6wnBCmqzu6ZSkFL7xT4yzXCRx39rS3W2njKSKB2VFL2JqRAECY0
3zLhCMRHVWsNRqLxdwkaT3EFVJt3nzTcSBMiLhZfaRg1p3LUOnyxKJbdegHxIxYaX/JTuJBy//S4
1uTVoRdk6mQdPWjoa4myQCvgrp5wXzSNaY0/UekMFXQOgGY8cSSuoG2fB8707Jl25P0l55ZZ8Es0
c0MC5Hacru7QJd1tRc96iX6knF3AP3HpALhtM7KGpoHWG1EWOAGMb9MkYDgQiB0MeA4CMdN1voth
7Rhuo56NXH6dObtqq0WP24WscxuAh7QHoI9tL5jDonteI57CpkwWQIJ/qOpjG6kcunjg9ePELZ4o
+5/Wftf/bFMlEx7ik4BabnLTz47mafxgROVcLhFnbnX87xbjUeBWIAjYWdO058t6GTlpMKrDViLp
IBdohKw6X1x2WVUnl4Kv5F2MorG6Cq2DXydxivYLBPVOm4/xIgWzKzzpuaNU9n8Dyn9wxBBYoiei
3No4qyYMptFdZxmGS1OjhFKsbkO7WzMznNXRXW7byB23A1kC8qjJ7lyr36nbJCxQoG25HVLY3lAJ
mfKBqrwRB9nSEOScjDEV3/XQA8K9usIdL3Ru8sFvV9KVCE5mQMm+DLS2lANyOZStMTg0a8OaWMFm
pU7mXmiZyHqiOD3H+UpAFJbjsmM8NADiVl0izfRu4orkJnxBvtL4tVbzfmSqYCDCUWfNUdlPn2fN
AAs9CUH/GQV2eBLIg96d4t+mBU+1mmz2w1+Jiqm3nLerVSQBXJwCwZQhsTONcKIMTCaocn2cKBhX
G2nHJAjZTKIq1yLS4QmNFxS3n8nN7EdTRcfJ84kQUccZhT3SSVwznunG5vuFFB6bEeZybJMTGLwE
QPZY3zELX0o338NAVfsA+4kYG9LtWQ7ruMd3jL/FIW4dRW2cvhZSjPNG6DWT6t2N6eLKu7rzqXIH
c6Dg9KqwaLqgXCBk/YfwPO6hQPyuOuvWTlyNYpzieIYrdi4k2FdZit+o4tXJ+LzMLq3F2rchhPM/
/pfRWlQYAr73SJ6MW5rZP+Y1W8nReEERn0eauZAQ/4Ih4ZGIjt/ZO5Hl2oj2jU2RELThjqZbHrMF
Wun2SSUnTpOcmXxKicBu9FwABe2q6Wraa7OVkRwlVBYcosCE+TrEzt/S/aWYiSWhfObrUiLGf+O3
+O3BJiCMmP721yuUaes/ylPsxwVJVhIQdmxvn+FM/7v9Qp56Kj+WY61UmpLKl2NyXwyMX+eWppmW
w9fZqnvMZZmk5cI0xq5fl9ZPxyt/9muEnOyaf3BSoZpjYo5LBpelxkwTRIXt4NGJQAJMTHMJ7+5c
lTknDAstmfqZuYHl/Aqif3gysiOAtVV8KVvZFldoe2ZKmr3K40TV9ysiw3wvCA9chnweZXf+PALF
AtPKsILVFAiwv6rb7APFMbzLzR1vytjU/0PdWF69zrCqxsmzKrkplNJxTZLm+Fn+mllVxsxaihmP
7hYZ2Hgd+CAls71vIVqQxvxHn/ScX2Yaef8bNKzFK5WILiYFHbfS6Nr2he/w3HpbQGbU6b9Djxem
00G9FrR1KrQYv91A1zivnxLMssVyeZnbuRPR99yARsg5OZfIpNFaWMoKIhpbdU/eUX6/RWz1jSIC
K4jDm2ChajL9ADLHCH80sCBsduIy1vzpfoiWK8p/OFvET0yG/aXOdRmjQOTOmPjBvNNh+bqJ5Ic5
tpHFfws1NkHRvTwWS6x+0IYcmazUkIeZ7qxe2dIqFPIBaTOdJQmBCHch2a1DNgtPZW8D4eJlk07L
3G9azhS9CN308Vin27/pw7avg0tRaDXGX/Ssnnfi6fHzp04h0Rx7gfSDJqWPtcDNO02mSgPg5viu
QPf3JYfOCmB4fknB4yoM0ZMDKz4u0dOxC2qWW5e3Xdka2H1tS+0BO4CViBNndiO+hrkttghCJZek
Jbzl9LiQr376eDYwItIB07Fp9++ERvqCO6NmHma76GpTej3fjJ5EgbUYCTZx63Zw38YA/nfU/LPu
tXYb6e030a22KJUG9ppGuQ/q38m3PeBwoLH+PPBw86O4ZtSQ0I/JjauokiuGqiWuW9ELi3dLiPTe
NoIkMY1GKZmrWH1rtjZtmOGlcPXc+XUElcO2Qlg1lgRDQCzudgfj8zq8x0pPDLxiAiSuRkuDWcaM
WyXt4mYsRcszP9hylAfDTc/7uQqon9HoeABwgBzZVsgD0B2GP7xLDucYp/2Qh4RzMPXTDnI4+NNW
sr4ww6Qbkfiufv0KnAoIR8T0PIGaf0efhVQ1hKVikcA+FSwPUs2MWn8jKtM08fBhOefvP0Aogoxm
KOPPAzLGBPE2ixvqKUE6+vy82Ym3Jz5+pjFq3rm6kwP4e+g8JQg/jSXqPTk2Ht8rktoY+iYpVw5b
v2rwvDpgb8DRB4FOAC6lHpkXtEKVXaQsVSqmiXBqS+dyYqMeFzT31vF/rB5P7jGSHw1Eb3I4FYJf
HVa/N/i5Q7zVC1OCGYcicDvptw8MjepePrkV17Xz7NQKPNrei0nLd0+F8IT8b0yKJHo4mLBXomLT
mtWTd2k4jlrF/2pYd0QTIBlGExsyMIGkEQR8HtKHEiPTQ7FDDYBoUxXOigAdXTTr1owJdKCvftmr
IF86jd8NVIMXnuwAGpSMMCm7SeDKz6uMl1hT9gZR3ZwbCrY8oZ07vFmG6y030TwXMAgzLsr1TvlO
XABjlxopjMHv7Aayje/r5BNFx/ZPNlOdBqNsUIQYZaAdCJokcVRPfIZi6zR2NOcCyYTtBGSPc7Td
FgZhBsxVEhlSQtLx57TWmULIHHwqQO58jtLp2cccTJ3wCb8z5A0045Mpp5jrBpmAdj6+aDr1J6Gx
u/zDDIQG10ayh9/BtE739eUl3k93SKdLimnsXgDSzAGDmoNAjE9rLCh8E53KWCpHKRRNNz2Mkr9Q
XKVm+XSm591p2MYtwYx7bOoBw6+SJwo57jZB1rH6PvU2blcBdOsWvJpd15nstE4hammnlT7t03g+
n4UXrZfrlmNqfcDT1QRzygoqi61FH7K9okvdUvO15UkRSupvAUmvqDYWL8KPn+mOZVjVi2WMD3At
z2dQ2VBZ7FteFVHjE8POVGiS5Zrbxl7Tnz1QoacoasSdbRfN8w4Sc2s+hVRPDQ/zkllg/NOATmQi
m0y33nPCUaSVEMCtDjI6V3OfIqmyp2WOLiaRbJWrWQrVpMjW6q3fKIGWGnSN6uUFFe3bMrFmIC4E
315+H1cGjqBfIH2n+5I4m7hwnYb1IYmeJqyvEcBCiSHjoPlGeAuFx1VPzVhY9kfOBhk7x4wt1Qfu
II9QTDktHeJGq8MEe8olqz6gRKN/a7w322b/7bNGyttjtIG/ARfm4I8Gamhs7jQtMb7ESDeLpbKs
MeKeUHnTsQNS61EbbJP6ewaiqSPw3rgGekyz82DIyPai3dJLv9gecbBUZggrcmGeQX0EutLwMUUt
lD/EG1sJRL5IYhcOWFAZMuXNw3WIVvHCsJs98dnoMYOXBZ6w8+edk748oypnJnfVMh711eAhJqgh
IQmriSsrE9IqECrtugmsiKqOqpGY/LSRadE2fGTUtgbtatayb1PqHVpBsIk8kixSHYtT0s7AJqOq
wGs3NOEPq1ty1Bm9wSq2YKQDAeERAQIjHUc36zg3VcPrFe0/shIfsGp9FdETC4KNUtGvkCHiqkwJ
CL9idWmxDYwvKiYi/8Oo3HWqlodpeJqZuprITvdAfkrFJTaPz7OvYMaDLWdSwxuy9APuGuAU2N5z
Njt+ffSne/HIvBCEJFlhJPaqpsu84j0S1oSoFhYIs35GELCZYpndriuee9MjokSPXH74pVZ5mMZU
qW+M0HYkmb6z6OUM9wQ5isT2bhbgfWZMIQpd2MiLrzWPbwGZXcJfi2wT2VAKiSUctAsZi6RUGB+e
Gf8rXwu6uNH3tNSsvCDFPmKRTcr51nkRBwFH8C46WxT6+bWbLWQ9HoyxFDKoqrvzHdp57vvzGJr7
rdBuX3aXmBN5A2oQ5KxaVlXoCGzeMrbvidJ2dGiN6S0KnwC89KCwSHWVo2ycGqba7jpDrXq3d4sA
H8K1fHDJnjw+iozag0Wf4SXpGrGMTrgLa6fXPG6ygTKAVAOng4A/FxkMP2Vp231Jr3cxE2dOF01I
yOttHhhCQWT6k9m3KgPd3peAE9rM/0PEtxcog4x/WaZGmcf4cT6lVG4MQIe3BWu/ep0B4rWfBp9h
t800lSgh+h9Sc57qW+Z/XKfl+FdkA2AbklqifldstuUKAKLX8+SMTW7pBUdGOi+y9pQGIcbqXnJg
g1G8D3segRgDMLXt1xDLfJS0YqScfhyicqGWdfMoI5d0YQiIGCsk1dj3r6d7wnu9fyNqcGUUn8fX
YuVZYnwPDMw5Ln7IebDdU0z+NMQ7OLL5kQ/pySB1TtF1M4/yklEGbwqaL852XX5LioZ+3qvDjrnB
ok3XMUZOJyY3TNdYNovASDb/VzNwSbKH+XxtMQDTVi8Z6aUexivyvlHFqrbZ2LPyvrsjbxJg2crT
SnXlU4BGhQdkj1Bfixtp9yl1uWkjpmoJepdPtQX2qFXs83TbDSKaS7Z4ZP+gVuQZP2cx6dSH15PZ
s4SZaW1tB7E0oMCkLahINN0lG40H59MmTYlT294/hjS3mPEO0XYJ99+YtadfGO6WDv+wFPWSSgUm
xV8iDWuABgzGKYJHwyi513DR+dPju3kHcADtiReZN/ReBpS7WoAEe4nrbrHsdoGp5mgaVSpH3GNa
qR3+uJzn825WaQ2KAAQJ/ZeTxE/7t7AXq0InMFv46wAIP8UpNESPvoDDw8VYUXacVuZwyHBv+vou
CIRcvILA2ZO7fvqC18/30CzytU4Czexb6lyg3omIyYO00MCYAf4jm3mXEwzb0fYr7VL7iU9aRa3b
PHKuYb81CiRFFPxXkekg7z1ioFJ2m3fgdg2SBMvFIwFYMi7paOFWcskx2DNhHw5fhcF+skf/40R2
31RF6vFqJdczVjfll3aAyP0KmMFWutkEd/0t3rQpWxywW1Uhc4L58pH/4oxImZs0Nj1WzKUG9rCl
zCjKZQUG0xH49raHaX1L+xwvvyIEdtF3DeWYgqsbBtMGjytxvDNO5FBuQFQ8JXS+Lbv/iogVo+cK
L6Zwvvwvgj7JVJpeNlAe1juG0KCrcktQ1o9mtAGI1lgRHj8BD64wqDR0H6TneT3waAzqYiRDeect
V/kPjdiimYt7X+1+GSp4s5Ngf5VGi+1Mk5ac8AyWnyK44fsnMbbVDH7ukjaL35e9Alq90OXV2sc9
jRRMWJUravQeHmoizmNDMFY313+//el+tAmhJVILkuzk3zQSMonKUL8NxMZ8K6M5ruFHNyTGzl46
W4HZaJ/jGZiBdy5ex7cw1F7wKf8en9F7JMDRGyeWg0fBrmf3ap0d5FLbBj9q30d76+ZdvJp9Di9D
cfamD65WJfEbwDM+VpwARlx6qojESLsWB60g147q11IHCpODytZcZpTY9CqGC6lavr6ZJYop5u0r
+CBijVZEo9Oga6UCz8DkzGNrJDHZb/D3HjRxw/zMCYVBG+NyBC4zEPkliR66VPpYbR8tDzKaGiw1
+2wU2IURgYjgmAdg3Hr6+CgRCl6s7LpNlqv7Q0eP/CuJ6CnDi3Hizwu1l8lr05qddYwOVzKLh3Aa
F31r9xrsvGXE+dI2WFeDZK0JKvd67MgDDA9Wo5lPUyDImREQN5M3Y893P64jHi+QWSCY8OnJZcn/
2c6Ahn1WzuI5mr9MsL5WrP4QGJHQ5MVf/6awuzmtiJdIzA0yPlivaT/w2Kk+k6fWjZomXVtUitHi
Xq+/uofwTNBZUTpbtHtGQJZ/Sb++SqCIvPqIdHbJlc6C3gJd57b+FJblEo/yUxWxHEXYC5/7cOLc
NSX2iUTmoGrQNTNYLwjpjwvHGFx7kkRdgfW3Kx6/3eQGoV55j0/XygMvEjxH0YCc0mJ5ITc2E7Xr
ooKndE/U4UDvhK/4QCK2v+gXXILVg5648lltGtjFzuasAXkwMtUKNES0SQ8jEVqkGzGMmsqyr09y
8w+OsWwjQQhgKaU2tWAtpuQmmYEwF2czkM7623FkJUU70HSXhPEw4BT3tIJMvg0xtJgB0DtbQpbX
Kgfy1To+GFOdYNqWPoKblmxJNaOFiZGU7bVK2y423Q52dPMw8shwC4ZZqvgkdoZsnCwwTRm0H2cg
fTfMKYi8UyXzLV0DADZeTEnG09WG0JhJ6QHtE92/x3GIxeNX9CgPsTNi04UL27nmSwHKYqGRWtIJ
wSIvJY+nf834sB3r6naFl84WKzERo0PuRNJ8QEajyxFmSIiQZAIGMdOeb/4TbEERQNCQsBIW25HM
eEeyy4ctZLOQZCjLjUTr5BEkqb1CYq2Lm1BpqS+D2lNnhak+SvCBZ0yY+stGq4lx6LKJQ8ncc+kV
okGmCJDbmdj8KdbUEfBnL4GK8A0et/xNtDnr2dbhTDRkKnyILjLDZ97X3DX845JRwFn318qjX7lC
gGOFTM6+eE2NcCutdQHu0JMQb+bdoro+25PKTHhkdDXJG3Rxh05xWNdO5sGFMzDbISjhbnK5UXbJ
EdSZZbMfWKDw9MT25BWUzqXRLaOx8fN3qdY7/GXnEM13/zpOrFbiMIM85H0pZe3TvfMvcjePc46I
9FzmcxI5GG3k8LuB+aNnPFsGwUlDS4yqjqE6pyhBSdP0zBZGvJ9pA/589SiTehjKvYaByExJ5et3
HJ3FOzivZq4pL0aYAsF0lH/qqk0LwtqZn0Jg/dkGS0StqLqDWKkwXs3hOrcObLB2vUR0C12KaeB7
HaROiP/BBiq/6BymOCqV6Cd5VQS8GvaJjyzvw6nlTYqfopnAaG9w6Qc9mtFoK+0GMxJx8e+F7ppz
JKGlU8UIso9p+KRNbv/eIuz8TLggNxMEUsZi9PUJNMIHWnK7wemMuu4vi4suIhzxQ0eGVGfSr2wo
c9lYk9V+638zZE0v0YMTIhiV5efd/K+9lt23jM7sypaYm9OQJ7ks03myMUY57Se/INpHzCGlZRnX
GjFQRJA4RijI+J7la11GcAKwTGvnkwCnDK8YhOhEPjOT6ao9J+EkBkHW0DI4/9gr5B69TXN7hG6i
tTEyaD2Y3UxJkOsPOUow415t7Vb6+stANXQUC8oMDZNYic05Cw5sIEcEix8bJqMG17dMpnf/cwAG
NnB+nd8V5GNmW6/jJgiG3hOd+xbzGoV1bf99tq3I6PJ072EFryglCC8wWtLOTOPTqdwEFS+eiKnV
P9TdhKPbXybUy9slO9XrAv5Ns+hDQ2VCXtrFwmxWP2wFXV0ftltZvy8Mm6Cs4LU+u4IsTtz/2jtB
T4kwUXFakX2B4Vq2MUa1J9A//R1n8ckswq+NPHyJjnVeijmRJ4B4zSaqaWd7OTtfCBtj16uIJ7Ym
KdpI+HlR/BAIJYzm60/krDg1ix3+hvEGtCAWmk5aIacJRQjsGhwLHV/iOETgNrOAOBNkZi8XW/Ov
S8LHK3ANQyZ7RM9rUBL5k7oRoqcG1RIy6AJEP/zDxlM+nxAj0jWTskNBsQmWPTD9S2BaWDdu0rRW
P/Ch8Y0fuTxn8zZLIIdnQdUKHhEUf4DczqV5yGeKjJVE8zCohk1Umvo8lO+QKKvJSfbmC4IsJk+7
cQswftJI+0qry3czpPz/3ZTUevzRjaD7wrdRLq6sztxoBGD0bqJfaONJ7Cf3cOA/dVp4b9osUpQy
hI6g8eeR9VG+1lUVv7b/+hsWV+exR7a8Es9P6vrDFbFBPHY33ucNqrTGoaG/vD/FNUZxiLCWmGR0
iP3MU4hE+YjUAtjSbGhOVgqRUoj5sdY+34jU70doDdGQ3CgXC+BdRiM6cLJz+P3Z0077raoTj9d1
aefbthCvqe0fvxgMJYlJtexrXfSFh+DwswCsDgzEztbnYJF4DZw9LjYWu82BBmeP6SxBlT1znQ7e
Ww78nGWZgVPXkkMUv1Sz0+Oip4/mQwGko+7Le6n1M423oB9Wq5Y0YSyB1+EfJbCZVLShtsHz5jj/
wTKAPsYB7f2TKqcDAms6jYPjEhT2yCoszyOSp2noum/zuBH+Ekn+JzyqfGfNlE4aPC9Ax4dPgQlW
fJhDlaZ8H/HfLP5uiMlv3+JoQudRKXwtTp06g9XtEvDVIQid3dTyitZ+nZ4rtPYQ09sQbcKBT9Ek
UoevtjiTt8DNx0IO2M60DrA1oG/X1zdYqc4MGVriXzTHqXvXBLSGuQHDu01rRhG1X2POg4/zuZ1E
aJKlpwBbK7Al71oFRzutgverVIw/M8tp7gqRseLxeJRHBUjmayJcO2lXZALCYNYwFmLazoYpvQEo
+V/lFC11uiqX8aOtzyefZxQNVsqdfA7WHUyMZFdEIASOej9QeDC0zl9rRmycPqD7VPRVFscqOrj1
OwYfVoph55tWhfdOD4e94LB/lCh1BbG5OxdGsfNhiV+goiQY2V7aqg9NSOhJNSh9VeUnNW6PysH1
pq+I/U6vV68g383u0eO2dtx62LkFxfzcqYjIv7l0uzZGutWuQVnHTULRo3bnNyzuz5ssQkw0gn/y
4ehFNGj1B/ecIxvZ6gr6n1/pVte401ScBZjlOxBbGW4yzPTxUDg9Ooeh+TZJRclqS3FaOYYymZFX
zJmVOLBCeC/7q071JH/vVD6cuzw+Cnc7oQPcevNFLd5UOmvhXt2391JhvQWm2toXGD2fXsS/O1sK
WhXCCQsA6szyxRqISXLmBCtLwPODCMoZinCtVSJZq99aT8h1UaxFKmFtiRwGe1aycluQQcC/yiy7
OV/FGCv1RnOoExGs8FlGhQ9Y7xTY1bzMWo7MoCN7dzX2kZGRkxXsU+OqfHKOF3KmaUyI9hkYsCh5
ehJPa12dvhddGnZV7iNISqdSB0Ne0sqxD6IftIvnzivEef/s5AteA+ysZ1h59TNDuqJ93EzXZ/lD
vDI8N+X3JnC5JjWcP2eFO2hju6QrkCdjBWm/oaa3eYyK+sJyE7A7PZPvo0gj21j9VrFxQwRagZwr
VsDqbrUgnbRq4qEspWcuoMxlNObm8BhCCkIfnUtEVJgVE9evzd2GFN2evhlQn0YkrrVrlSU/2eUp
y1pqFSEoNWOo089j5rX00O0Egvi9kfv/nwkBoGbfEpgd8gBgeIdZXTSJcK06QhujYXppcf/wwCnw
yuiKyzt5/FQh1/tSVxagpc1UoayhsqIrAz8zxi7XEXp3AIdNK0Ew9F105wVCDdcyYeWmOza2e9Qw
8TN0V3Gz5rPhrTeXUTBmSFb1FkjmgOWmXywpH6AFs+h/qhKIbUhnyfjLdNa1bPxt93YnAX1OahJD
1uO7t5zqbjWKgaxEa98WNhE6cexNhOrKlP1l3AFYpDdyzPZ4KXgIOECQZq3Tp5rbxMoMh6iKTbRn
0vVKdB3+CUS4qa9ItlODnf9sT7ADO6xTc4aMRh9oIV28O2oZZmGmPF48jTOL0XPf5y6jD3FhlCsh
rBLUoveTWG9nH6vz9gEuEbpWifyRbDR4nk4ljBkY70hM767KXwCaMxWI7RwokOGihklgtbNz32BI
vwqfj9+Fy/BKcV+N9SRS21kACp/8Ya8pakj2HPQXCfDpZslROBMqKT8A781LKgPu6lEWwPIXWY8D
HnTow5tDG9qW+hqhBjU/oRXV1Qnq9xumQvSQ6OWkLnnKNA5CJTwSeVh34Ue36SppnuZQFhYCJN5/
ybaajSRw8inxmGCDBOa2mrvu7JySrqqx0sHHqNS9UKcRrooeeeb0vfIrjFfouJr8xSw5xYCCGdoZ
fdDgybHalko/CgwUJFrtfnkKfdigR84Ku0qo9OBIt8+u7RU05pQHJT7RLy+EvfuffCHY0RQPNfPs
XF0Uy7XdR92nrQAWhvkd5u7tCxnC5yyvvl6BC9pNONUt8A1LXm704zusRc+358lVtpcYE1wyZ5S0
li0/OWtss+Z31pdmcW1pBfvb7MdCq13cbf6aXINDgWn7snwZp5KKt1v+/LuIxHJJGS9MJBYHDjER
fKsOspyVFVK5D2MKmev+iZl156VU/osS/pn2xpQNu5jYEzDPDaVjE0nO5iCqEJOvJXGhNVXWh/zX
o8+Cd67lqNIki4G6wX7sSaSTt3GnlKG6NiPftStz+M+7zkgtWSFIC98Pr/qxRNjGlY/34JHQ1UgS
Hqq2mdMAuGvDMjHrgvhm8uGyp0fMdtbxYVKmcOyMv+pqhThoi89YEdAzAgRAsn5vUSmRuiHoXKr1
Fl/k9Y9XQM0uMuPVTO4G6mzEt5a46BrHhuSvoax35zGtNqrhCP0duW56FAA4cCW7Bi11/37rkvAT
H1JjB6jQekwUTbbv5dS2Vyoj99JK6hB08ZbZnqoGHMEvz03Pe6gyLTA9YXfbC77BId6nMmVMaAPi
eijwJo9bxyclSw/gZg2G5p+bCFOyiKlSKbC89gptq1zW37RHVTQslvT+LRSQjzE9s7aon1OGZurR
zsmT2/e5cc6wRndWDupkzjeRrnuta6pPpUUfbNVZox5Zqka53ONEr1orslvAzEpJa1tUWWGQk+91
l882grO2rw1jgVAqbdGRMlwKlNm/Vqr/wiEyyrt81EIIFdJrK1WTas9cUwnOJfALTzBwBhKWmaTh
0hTNjcAl8tEDHzJJZRefCD5bCmL7aRbhztIy/QDlcwIfRDjBbzoqP/cWq1MqNQqnmp0yhESUteMz
8b78u9JBnJWfQ3CPDD8VMz5ml/rkzMuayvdU0/f8lJBw10kwtdNOyZR5Cyq8tpJzV/fxyW5dwE1Z
y+Ukvx0PPQpWyW6SGtBsRf+wVFFMK2uPPyjeNpkm2i/ScDGH2WskNMvDN0THknQpmgitoAkfs7tc
+A5Qpp/VTmFW0ChgivoyPzCYRE98eOuZI6oT3zBO78wTMhHoJXnRyjJjKx5aVZao8H+g7y53ckML
hnHTRpy6c0faY6FTrYqAZv/nt3LFemLOpjAV7keeKSvfl5dBId+KNpB/ftOOZSM2ZwWrszbUoahm
3Ap1Dvdwa6HscF24D28kBVMeiPRCvfGgVCxEQUigug7cNtukucC+UJAwXalFVM0xvihA6QUhS0D4
ZLgKRQ5vv3UJaxJuI0nawPX4dQcbK9vcHlxnYJIweVnZFL4o4KH4K9Dccu8u6XQiOKUT1gjGhdwl
6Ji0NFYxvVMiU3ZX8tRGPVaL7lLfie/jv0GaygKqHGD/fid+Gi5RCIMP/S7OVP8oaHhvVZCL93Qz
PM4valsWxdg4hBmIOHgbytrZn2nH/x0jbJAakBIJ3UbSDhQ7tUIkXqgulzQ0/59B7j+yHYjlz5Xd
bdzoFXzsP9tj4xAzYzvp3ruRH0xpoSn3f+gwcyy6Xj4RVyZyWOtz8RFtf+id9cnwzNYAX39tX4qi
q4C3i+kV6+s2HY/lZtPANmhIzHcRmVerXKeSKN2htgFJi6TGqZzcHnSALmsDZIiHi+ztWwDkdjLy
e9Fsv0zfeFPUl03kWjZfO+EFtr8DSTTsAeCmqT4hD7RIDsCZhkK7a1DlAg1nrCYqE2+yr1MpYYyi
hpc5px/uCY9i+RZjSKsSdsKlcwaCZSQwPhcvoAf2poRFpqaYTReELciIZIj4XFZNpfKgxB9JXj6D
TYk0LDWrWWZM01UZnstlJOeOp+B1unG43L9jFHPspzJU6c4P0XScRmtC7SuuvgyyqdLw1Yl6TGae
Ijv7X7JOMoPYaie75yl/IguAnTX4EUlJdFsfn5Azh/mp+HC0JTNp8M4bCJqi2ykgrnc2o1FrxcVf
JZJ0e+OcuiMMNW8n7HKvrBvkjRta0y4iaQq1pwiEPX1364zKXFushAoZT3nAhVH3VsN102n4FqHX
mQ04xZZBP35AN6XccFXN7ECv6iG+knaLPVnlIzS5mNFpWys7JsQPSumE62k7njyrYpz4HHgyZJ5z
8TPGM2FedP0hNQGKYBCxVw8KvU1UTTjjlJQ09jZvDt/pyfb+1qYS8zGy071U45aSAL5hegDL1FI6
anwdPbdEEWYQIdf04xt/uGNPXSvOONaWfMVUOfOpQ84LORA4+y+jWvjtyxev2gT62YIkxvFQsxxN
yhqS7Fz2fWjX2I9whmrxkGghB/9QWPosugOmI3OOThh+EzmckoovZmL5tMzi3yi873JRKm6CreGM
bEcI2M+GE1nRlCsGsHgc7gTt+KYUzAWjI7ep+7Jy8Q1Z30j9DDUTMlnoVhNVTMuI94p8EFSWJaXz
ikCB2MZI49T2FbxN+6kwb5+WVa4V6pKcTVSC/Czuq6oDRNGVAeg0zoE4XOsEFkWrS6jdc2Ny971f
c2Mk7X65I175d9UEpwn9ZwYG4MfxCAKW+GXSploZPyZAoP+wD74jDWOn0hrTNDw/wzZOpsZB6x2p
bA1ln0xnMePfc8gSOPOT3J2k/DyTv4ZILjCRXUlH2ynagglW9EvR7WVzMs//z9Dpoos7kdzxzNeo
Z+pAeCVMV2T6r+p6N0KnZIZFgY368uICxojU7UhGWsNOC9xKLG7obwOwKAD/qfJxfcMUhIKdPyl2
yck4JmUT4yYbAW6ZJrEfsn1WlcAsBh3odYP0EU8jp/e0DoG8o2gGMJY7qofWHn9IBAWTAUcDlkos
XJI27sCfKL7o/9k0+NfquSt5UoumKs5e2xWpEd1W6Klq6lBZ67OC4qMiAxed87wf0VIW6GI9r2QM
DUnFF9+3t6GzEAiS19V7fs4ZYumRN5cqJkkvHX+h5XG9/5RsPLzR0WdVsU8BMX+6fsUnBQRIQvYP
9YNor2OAS65IrdOCg/2TrokRAp0QLVEfCUwCgGN514r3nNVe8WWbLrctJGSyH7zWxWnfHRKWqwNK
9+yg3Xw6Ppsag9mUljGGCX0el0+YJI9WTx/8mxwjaFG3PkbnulGEy7aP9d1QrTPZBJZ97iB+Q4Jx
8GIxUvmc18CFpZW3gH6n9BvytEHVGNjnnP+WvRNIoi7ZkX26V6ukUeQKG5emptnPpXlealUjxNFu
hfTZ51Kf+wZIOdDtRKJYGMdtXuQ4JOZloopXhZkY+XABCCX0cZrXQLiIz8/Eja0LWPIW824FPnwa
y49jtFmz+RYq3hKqj3EICFQMTxJ6QIRAWS9+Nk5fMvkJcp+zRnMjpPbY2vpexAXZIpZySJedCXJc
DXke7CaqhXiH0NrJk3CazvnLb6SYePz0XF4aawuJ0bp2Y+ZagXLF2AjRciqxJZTmwbqhdFCXjZlL
Ow+lFokmIjg8Xl/KTvRA5wS7wPKN9fW8n3DXz7cal5ppXXBhZtN/Z8ss5H04y1aAdzS406CnVGin
A+BPEUvF3Y0aVZxN0iLCIX+OFnB+AZaLBnk6tbIJ8dnKmd63xdXHS+xmaC6h7dAN2WHvfFIWXy+r
toIPRDs4AibrfGSHm7WZOWoMTEHzlzB15xnw18AllGtlax61AQnAej2bCDvi4YPmw8Z0lvB9NFx5
kLXKjOt6oVbtyowXkdwphNwzl7Fb5N79HZWX3mEu/rFqteXWimtjVZEcTXcxezsBYq+/UzCaTfEw
ckItwAHPb6How7/xYhzqKnXX0dGAIJdMwpdxb3yFpJbaj+sqWDTkh5MxHUX2B9ueQZqpX/VI4rl0
v1iH7qy3fuN8TEQUlbyMkknsnsBZZUR5sKZWJaQASpSsxgeVlyQScUVJbWEhft6KtNyopne9Pbfx
8lV+ecSnJQiSezMmZmIgRtdGifzcFyKCYZFQi9Q1OJ8KEbwZsnc9S6kHMfu1OFL20SiNz3nOWdpX
jxNG0MUKy7glDkKIxXSCu0yQHoE2VuAlMXQUn8qW6uy/sOiwA9Y3221wLOr/StTd/npx0qXqMJuv
EXkGwOUBuwrfYVIyZxEuCs26QGle+YSZJYt5tE53fSphHmCdpglmvoyMDsFRXA7o8a1Xu/9QAp4Z
vsmripHZI3jCFJkjfzaiDR056zMc9vPHE4aUjEuBfkwYm5Yg3zpACnHMUPCknTIKAvo70xVrxcch
BL5Z3l0UGTampb9C8TFfFrMF2SburdVfdzoc8VLa2nfDiOdJIwo5eb1yo93L+OQiZ9AirJjRNCk6
0u3Auo4Ims/11oHnZ7ljgWS6z18oGScryL59vf+irCQIhw3ZY1xWr2+sDemB1FLkHJk56BhH6VES
I+wh27ERXf0uzIPuOgWaEIpKnVycY9G3kuj9/T2A/oZfyVL8oj/sjfUM21Ig/lDq5WNMDEODbjMe
/RCxk0UQC5LeeOJJwgvZq77I4lRg/IsEwO0xgC8yM9UBhQ3M3Qr2dABIeFT/DiVI2i6vO3104VoL
IaWdtpUjBLDCAElf82ycx9BwvmKwThJuqKRAX/u1FU3DrFQpX7RaL7yPc/pK9DBJx3xoQ9Vv3ppe
aR4Xtrev+yNubd26F0R58DPgum7syFlKAvN5/kqZWYhwOgljW3Hmmjcj1xYthcLpdC69ylYPqKtx
gn1mGMFJLw5IUg7+tfk6+NSBRbjkbikai28jJGapvKqSsU3wP41G3aoNs2HDzQldAHmgMY2fHWJP
7o6sfbVAZKmGaav3qeUw/kE0kTjwxKh1U+z4B7fbPym+HxpYG1VNETXX8G8vm0W7CbJgJwuSGsLD
QNaMxU2DjGMTfeUE0u4/a7BiTU64rAicRjZXf7nrn52XXDJ21GnAF3hOVp4GCrpowlLc5v7fOl37
ECr2oRQhn9hVUr7crKBZM47tnxFqpP5YVb/AucfxDolFGbaKbSXdv9iepqm6JYeNZM6ceSgGOMVT
v2T7D1GSvyOlVc8mkxHkxS1/VFeJfqP5t+mi3zfp8l1iYe2hB8c2XUL7uEFEAd2JR7WncMtZGPWu
eTyfiC59K0NhEbVDDro6HsNmoi4BCpwrSyp14lymSprDXBmITbMMc1eAKtqsVUbCqIW+J86royyo
EZHNVhBM8UneNzlcucPpTKxV29gppv5zJJVhUvJi2EhYhdj8gKYMnoip2U2/cGLbJnvGrEQb0nVe
nDikBvzOKa7IYEuldmIvg6e1dQGFd6bq2tTmUON/1bG1hXDHCN7sTb/17SEA5+K3ocxNTqRUmLP4
N1LMA/i+wzjomndHYbjw22NxeFxMr8ItzO4ILkAiKqgZBZK7QSYATJ8yXgWbx+BkWbn7GQNF6MWv
bgg/cKGWZyaIW/qXBWi8HwPnXJ1K0cZAul70Z4JZMqUEGXGd0YDaGn9KKgOXcgBCghOEFLm2mM1M
8sc3jVZPxKeCPLs2LfeGOVKQjlZcnORkbC2duDdMYlKpH7Q2vTq1znRKqgeh280wJOSBWImPJzFU
12jL4gE9EJCC68FX509Dpdid4YRb0/JZ8Q7g+Rl9T3vu0z8pE4yh5gODzKAYWdvV7SE9PWODG+Tq
VNFMgTiDyiKVCJ5uk80YWgLuImW3wcuPmpdRWJXZP5d5zRXIJ/uumG1G6yDNSmCAAfpyRCy7L9re
euIyrpOTrMh567tLRjcrjYcSg1PpNhXTpmUlPVmUbEUg3Lzcx6Y7umwGqaCckalYSdK1N4Vb5lVs
L8yY7sVoXedJjL0jFYqQPbw8v/HnsiLcI4bJpe6mEFONspMhASvatGyFWAFaTqdXypoV+pcwXij4
Xo0U0TsmTC3fxb6ZDSsKCxRaWu+2G8FruDIomtFaN2eSuI+fT+uI7crx8l8a9UxtDmGIrF4O1Ric
atDeM6QCqF/1BhEm9eCXVHwREo4Zsv71vnqjFM+7GM6v5Nq5+ODmRzjUe2ah7xExJ2MynKDhrD3m
4ul5WsBs54ADmKgcstTPBmf52mAYQXMXUG1neVPr4BsHCAsOo6KoLIDoFQip9JqvKjfInJEd2IjQ
pfQIiqefau++6A3h11lqcBC6dvY0jn49Pn//lJj2yLVTPxgrFPAhhjiVhsiQ/ISXUhd4q+lpI4bS
/YcLgQ29z804jeGjS8y10jk1mTqGLsDvH/lTmaQeADLliIXU68+gzRK5xp2Q4DgES2A+EeX56/Ck
q6hZuP3hFN4bcH96eztI4/oQ+iR5vyQHxxwC2LSFmR3snH1SCPIHdb+Hot75nGn3lNDsv3eNTkIL
EVzdyy9zqhY7DJnkMKO3dhRp21QuIq+9yHpSkbs9jwHIrAumQ/hN1tecKsvFFjLGhuHupVl5RHs8
AfZiVZuaMJEdu7sEpYqUW8FOHS5s/88nDRv3WScoEutmLJ0/Ufqj/SOUCZq5FrRINHtl3eH3jdzP
y4sd3PRGuo5hL9OisfYc8Sgck6QiXzfKmMmi5lRWp4O90/LHJDTT0B4Rek8WE4PDA+SKCKV7xpRO
ljozigQx9NxTTNZ8IjWHlYKjrxhh2wRLcH80YAIJMggpzyIK+lLCqiKdvnhpv5X62ElhrjFBDMzf
RSIHebcfPL/lkbFw6/JV4qqtYt6Zg8M1K4Nz32svIrrYrnC4fHkRIA1ykBPL2kjhydbMkzqRTjjQ
Rr2rJegmZEkuP/ABvcrTi0WFcbdNUWf73d22j6F6t+r9KKvD2ElLRcJ1nVWpBV1pL+Dxu26uWb9T
drr9v55z6IfPUSyE/EdKvXZ1zUKUHc84cJZL9bLhLwUGF9qySOPjyAIXROwCtTzQQzmoIIB9il29
qs/SZtq5UdR/8XippFAR7SdiK/cPCTYT5zvLMgm42o66MplUvjlb8Z9XxvaSI4HJJsKZLwQe+Fj5
cmpMyCFojT9GsGYb+BtRCRxbDyh9xm3WtWTaOgpEkprfbBti62ZtLxz4B/ooL7NkDq6Bg51GHthl
s94XhVM65ZgLPKFIxGmzinx/xpdu69gY3yqA4d1hrfKEbEhMCnGFETyzkJJVjVJUy4rOYLAh1s66
U47Yqm6ntqhgqW5DfwylYOmosFSpACumh1eaoxCcWsZ2cBbNhRu9SVKXz3EkrFD1F9ogUFuWloqa
OPdhxmmsyXrrwc8x+alN7FCrOmEdSI1MpGReDi9T7rjMldNkcl/TGAwVBGnlLBC6pnORRPFzJNYj
UoHSHBGE3rMGeBw3tO6NZOeVYEyD3EWjiYLS4mL5qLMBpbmEB6+Ub+pXwRGqHh8k/Ml0BnVfqjra
zDnz1gq6EoNz2EHVge9mAXfcD/SFebO12tAgA+xk5gtt6pBZtY5KMM8VxhUSYLvQu6NcGfGUB8yN
Jjvupdgjo7ItBZAHLxVIqbl8jC1CpbS91TnW1r7Vk4nq5wNAP7PtTb1/TccXCcfDtODiAykJWoj1
w8TaVkk0hxWwCyZsr74ii1z/+o86CNB+aLJISo1CSH0+jI0qjNK3d3QacJE+vY0YwcZCzbRDUU+G
pqv7HioeZEztza2O3oeaVAaEkE0Y0J7Nxhcpc5lBHrIxBt8OhEAyvUu+WPTZD7EdmtZQYvXEn1nO
pXhaS6YZmx116FDWRZmBB3qilRnDesSt8ICLsgYzZFKgr5bq5KsCsWGnyoquUWzXRt4tanHK3NAN
3eQegwTsC5WqLlnbOvOXoRGXzQElrYjHeyt3x1EDSD19IltJ7LNptX4Bgn+rt/+XfqlykZo0D/0H
qZ8bgJHv3C9idjIr1a+IU0NDp5O1y3waeDv7R3zoNaxY5XwsTv48bCjuozE4Gnwz4kpA/NzQF+zK
kwRGOSWxL+RfYQr86liRJXWg23ED+0M7ZrnW9tgsHYuJa+QSugwRw2/XHqhnLwiWsVf3X+nD90vw
3mSIfpW28UI756X800Oljh6NNhwtvlAiG38OPZOnCa7kx5HwvSDmKOsYqf7UFtlsH7HCiOYMLps9
3miI0MeXWdLy7QiYk26sxo0o0LqmkDAtw8FXBdSjxV4E6qoKGsx4C02ifpQauYFjrL5Ku2CZaeXM
juGOMWXzcuDawZCQWOpNj7N7YKX4BIWDvL16upZaGOdzzeVvVWIqJGd9dd6R2ms6P7TB5/A9RoIS
Z+Tc+xkjkWCth04gvzvUG3jgFCGAozLnokJefvIstiah+7FKWuOKMBNaDP83CCq1YxIobYQ/MkdH
T9lNuYkk85bhO3E0xKbh58/jXnxGo0fikeLoAzQf8Dj8g3FKhwm8uDnC/SsGor6MZVLDNUacBeE6
kmtf+hRXSA5knOpK9o91BgHBDAXsW5BWOmK9m7lqZroEyLMEhFfLP264Zx8nXvRDQu7tkIRDv57i
LVKIZCaMcA/rp/mCYI7NWrt7rxExQxjqKQHl3m//WmseO3no5kk9GbhZ3qKuZIfNdvfM/YWgevrM
CSTiJbJQcT5KN30sF0gGz6/3Bfok7+rL8FTdgqDETRdPO0tdUzjDHm/b4nMWlPQaRBTM8GPMH2eR
ne/T7KjDQSo5qOCyzihVAMVT+/G0ZxIJ9nnOuHN39En5ZjfM6U8c7pnfWnvuu5YTfL2M211WCV24
Zj+17XBRYG746/BOhjx6GAwd5/Hhx7+47fldIp75tm9EvpbfY+eymk6Pl4lS5rmcmJCuZOEfmde4
CFSG6MKQ/WWy1j2sjut5T4Sg6iRkLCvWxqZWaDCJD5XZ+qRCSmwcm2kH5+2LiIjmB4TKegO2eNRr
+JAwnZOedERAKV8kOHzX00292ST4nlJAMrxex3PRHCHuY/Xfz7gDQ3tnZdgZ2zyj/4gkEfXcF+Gt
tywt+Y0j7tPc5XTPV7lYy37u1cj57Jxvdkn7ta84BJq6pImwxsU7FI0ac2H6YxLrzZfL07ygEIeT
HTNJWaNAEoySLyCkmn4wzo7avffosfkGEzTpIIh5UQc5VEw2EieivFnv+5De3TXORozujvnO8L7W
XGogtB+MhwQhfn5DzoctgcahNHBXvl6PQ3RkygSlGRwNFMrzY8kRaBt3uBnYGZ+seTimeXze8RHx
YEX7MCI+rOU2374Luaq9SvM6NBfqdJYoZlFlJovRB84S4aPIZMOI/3xdICZ8r30wxZB9tdnlcNfI
w1xfQ0thPZ23vl5S/+iSolLubQinBk4O49TmbvCkoHMujdbVN5wGNcWEjU1pOIf6XgJ6MpAdAwPn
ZrvXviXVBTWETP2mq/O7tJv5MwaM4Bn4ALZX1Whlcj6lpi7CjAJa0ibZj60YPl6O3OVCJsPU9Sww
o9zM9LIesrRTGVP2qOtJAO5Zu3QjOz/mh2rwnbzZUiW/qU05TIuG/26kidV3vm/incZnBGq/EsCZ
K2exLv2v8PXtXMFpY/8byJm/RZIRs+8xVq0MBwL/DxlDYb1+jYthJ63Z06t9L6sK6cCMNXMoLE3p
QM6CJJVR4HppbKyl+a4X+U02ITUt+eEkFOneYvcKUYNzdIHnhVdpWw4HK5NfuAVQm6VEeCOq+jMo
eJR+0DfvSyGonFiSTAXGyRLFXtAZBa0shm6sJouKkGQRSaF97Mtp+s0snu9VC6st6PPsasEVqPzR
TNxHqukWUS8CCgpGXRCQl8Lyr+cZpjdaQhjzODgwFuqgeHFDTGqrPJAi2yiWRBd3+wQozqehO2Gp
37KrCwmp6qxRvx17xQx2RAVSadpYZRj9gbSgI2lm7VkpvQhjfugBIymDYT/+WWraIpkgYpazBZow
TcguOYMRgsbtbPTCtgbaKE5G2kD3e9vjRuoj1ATVtQn/sv/co/+3ZKIAGvVDPqfOmspjg1vk9htu
3jgIazvM7sr+vye2kZpGGevNhHce3hKokbvvBPAy6njBgXyvRQokGy+BEZ8uvrxRGeNKdEk6Al17
i11jBtJaPm86NydZvPb7gzFhHA8gBWxgyzD0KKFMryDPdwxdbAEx9UMQOYA4Ik2WOVgOWQFaEzbk
Es8+MvStLjV+2K31/H8rFyxftw8JVgDpEQhpUtAsu2s1qlF8OrtMVTWOJRkf22t3b13AZbQ0OKaz
du+VWvNU1OpOALWVgXYHaQYx7rgfu43plIXzFjxfArp4McTwH/dwEuFvD6+0LV+WgVAQ5AWaMOQw
zXmq4HzgiX6C3sYosL8mHPG+QcyeKMk/3ZuT0zg1UNQJmirKd95W4FePF0cerQBI+GkP7o+jwCfi
zbGrUsM4NoMDpFexcSkblcPBy/s32ehC7Yg5HnjnwLsCs3MnK7siQTn9VQEZ7KS3nwcuzQbG+EuA
he0dR9MPd0KInEFcoC84k3mTuzU3OO6iAqimJiHpU9X/jJ92f40xEwGvmWPcr3GYdHpDPOBitax/
aXtsayI4X3DZYbskA5P4XwpzmPFZswENUAh69VOgnu59Rd0UnyjV9DoTX2oNw26basbZ2pRPJ5xx
u3XycK+64JWDF/a03DqjDhcZ/l80EK0PZzlAcQfS5HYGH+KmzELRiqMevEopJdxMzI24Ocd1WCND
yMgOQ1jZw9mldEaS/D0eWdZ1jdwyaW8VbsPCSaNLFXaH7neggsIRym2G0W225TC8YNC/HBifG0Xw
PAf7i6xb5o4W4QH9OzXkmZ1OEpoVfdeRzuk8NiZVDLGtS7VSREOBTXdFUGgGTTQjQ4+iuWVnCfz0
tl1KjXoJlFFaH7oe6yNlK7EX6wZOaGCvVgEn80QFa4E7JkMOyRq9lFPWIA61lzmoiIRKQNlBZf9V
fyZWXBnEgTuazKoxfmN8+Yz6wLSMhPJKNydX/z97k1lxZpmOc1YUSFrJOkdo6lVJ/QSBlsikUlB8
9Xn6VAJTS6Xp8bwKOUhjSnkjMcZWIZvIjYuutWh3tPmzMXwn4i+qyY/RNpdgyYLU0iHwqOpdiWCw
WLaQiZIy12dRxyvk1De/Qk8TiKUC2o+S4H3UnLm20RITsXemmU9ZloOIK1dcF4ZDtvoa9+913kXE
/PXx6xCKbjYv4lhToTcqBN29KhFXo/vKk0RJjOrJp/ZrxFEcMI0CNIjvkGs0hBjfaNPX3IvsDYRx
3khBq1gsSK7DzI/K8blntmiW7nJguOtivE03k0yRNpY2fJqR4SbtBmW22Z3ftHWuEqitiXfzw7wW
Hop1/M/WFFbheBqVcnVR4hvaA31pMZFBOaQjQYD7dHcp02PBF21hH/WJAK+aLde61XtVUPFNQVQV
Pvnrb8bF32x9fPAozYTySWkYxARSdjq/gTm7JY6YeJIB7L8cItdOfzcIjJZRGXxn/Zil/Kii7iNu
FwoGK89+He+/VdFAR/G/TNbLm+aLzQ/XLrYtQI2W067iQthRiJZ0m+fou3vdryP4+IGuKVMekw9D
mNL/p2W3dnC0aiJR+89v8GolTh5M+ONRsoleyGvK8CXy1aaDNdyfS6kv/sBG11mydkoaQng0yyWE
e/JwkRrZw6irUSQU6tIhLr2pnXrSzf1fxWqMLSjs9PG82xf5XiVZ7Uf0fieiAijkDoKhg3mpeZqG
rSx97yzOBR/S5atnko5acOcQhwH0Zi5e03SExRcV4oOMLdXWREYVfhVZ2Q6CD0MRNf1V0+TH2S8J
Km2O7FD/9gcn6Qgb7n/75aRJFzbjSqL6hNnJx542p5MdUqjTAqIsBFjKtGiT8S921Nm6mKzVTR+9
+bn5cfIn34CTp93mdTwLGdwVBGxyypD723pQeGxgbAsxrzvU2xld0M36QpNylJVu3juS2RXJHtKQ
rTafQfLNsLZQ2S27P9q8GXFRqIF5uFiySatl//3xGkWmxaf3GhCY9od1G+Hd6r732LWS2NsIDwsn
njPeqvSJO+iNiGmuaHaEWrE9oL431JJQbcPT/UzP/MqEn4u+o+RcnaEeHNNNdewhZoAVag8rEEoW
X7i2rCoSvcibwesn9eq5HQ8ffvUrB90mPsCfi3pcPpyhPJakWwJbDgNe3opP+OBQhDUYBPtRVMT+
LPQUGz6Nn3LOYy/2GlYqq+1LdIGqfWvM+Le2CEizbqGKOqlcLuRNqjRs6QIRwZ0+fJYNh9Tr+HOh
iK44qQ/AYso24t2L4n0a8F8JfbPsJnheorx5jre3Mk3OKV9K8EVJ9TeeHgMvfa3yFq6tV9iTCqJf
/Ust+pHuNAhRdXBcRQioSVOFTxi3FxePEDdsbZWDmwslU1Udf8gW0kBfk0T30wK9ZcXO0Ak4HFA/
TbYEHc9XpvFH2dIz8w9kPFpwnqzptsF5PRUi7R0OXD320Icv2IH52OuXb7ml6uPd89rAH/1lWiLS
1duAxSU9WUipGtloEW51Wyg2POyVb4Ox1/q9AD+eUBz9Bn891lVarkNVGW51M7eDhVkwokk86Ig/
IKmRrxpu4o8mQVs2E/d1VFiIvlTfPYFjoiWJUKY3z5EDgSpTOBU9SYilUZHqO0B2ubJnbr2mal04
MnIbdXfvR4YkZYEnK0ZDvMCnVCgm0iHCcvvJ493TdsVQ12s5Bleop7oHZNUv7Z/K1g36L2zfaurU
Dl+ppz8TdwD5DzH0VNuGm7iD1GN54k7IH2sh10m+5SrYGewydcvSMK79/62Za35/EMgE/tfe3prq
BIXD3GclKcvgPGlsSAmkdVkT3X1EQm6h5530eFEGProrcKRUIS1aqT5iRbgo6rKJL+ODSJ8YAIPV
ewqaWoXTBQchXH12ikSR+0hZcOpl5DSYO3kmdBT3SyTdzdc972iZoFlJOZTrrBz4MwU05M3sa5+d
n7Hso16GICRdt0N6byq10jhnjqXAbmu2Lf/jgT3sasl3y+dn6PGEmNSKg6DlMRoBUQNyLlSt3Bdg
g0YfR4POdC5j0RGGz2l+Nw8ia28AwWfSbs0r1HBpAMTtwoCovsLGziaI28FSLyMZzEVLlj7hKuJv
6ZFF6jzUSqF3Eow3H6xEC/gbs0LXCXWpgv8dzB5cdB8pWbL+hI7J5PUXXx/oDVm2nNRd+bt7D8c3
GsJwzpIa4aaoTKiPsg9EW/tdOWu+T+uqcrSj1cngNVgTjMuPllCR0QeqkE5UJ6UtrY2dhdia5kCs
0+R2zW/MruNalcHaBoNthEu6EA5tK4djPMZtDVD+3as2quBKjPGP79U6DTNUcIPizDGgZ2a8D6Oi
I8VwGM6oK+BXMNaX8TMwuIiEicakqfqzkACYQ3OgtEArSoyuNeopPaSF/n2ek01cT7By2Paqpvm6
+XwM0s7Czaekxst1lE0npxXb16qogRT1FhUm2XVbhD6e6JkB2Tp8WgKQ7vPa0qPZm8sCp08q1/Or
BfE91THfnBnt8E046byJgn8lnrK2ap11hRDuL0I1YL4evuxhmtAFtl/LZlkrN+L20qKdDpjW0Yer
RXcqrHtYQDkCebjBM05HeiU6NklCQfGgvAn3YQV7jI1d3zoiK3gbsBBMZql/Tl7+wehpIPOCF7CL
l8zCwQFvGecxdoLvSRan6rJkaLSs/rgKcRF/GahWuRLU+Pc/c50fM6roLmQc5jonPDpIan+2e3dn
xPyNAQnBqBh6U3c90G0sKHWcX4kYQo3qrk7LioINBMDwC7TxqXpb/vtqCxUSa/y+sS9M1vybw9Ev
JMwEo0hkXiUsS5R4m5No5xvavhzZcH56jssOSWDTDRHaRBDkZNL5PHOWQYr0dT6eElMjtpiU/gDq
+39W20rgvn9U3bIFuMKBUsOsS7VuxSyCx5SM6FD/pUSAGQrd6HGQiHEnAtET/wpeJWMMzAXarIfF
099EbXLWe+QFvN3zUb86oD0qIlFi7nEEg3INoaoZ+ssK+qdSOA+kBaRCxQsPc6QYkiZ7+Qt6oA9u
wW8eMizO9v8GSFLuSnrU4hCBLtQq5KqE+xqBzvZLMYBSlMtdfLKNyZb7OlTM9V5AMBzDQ0Qf3yow
gc8NDCYjpMF1JrvEI3G52YBAEBlGIYMmWXy27raQ8aF+LsQKc13mT1iWo2Cx6YNb0Iym2STz4lqf
bQfINL3gxTkV3zeqvA5MwnqgNIh8iIhVxGYpVbG5yPr2Rh2xAw0XFtw8b26deabTOgtVPCjrUpcM
8HJLzD4b4HzzJt+K2VfVIO/O7WZfBpIzz+F+L+e1EPOcgfiOU3bujZaBj3CqA9iR92+ywwOb8gRt
XeiKNtMKhroH7qseNLpB7iH6XxcwA29hhXA0oBRJaaIUlHX7qVsJoRzsFr8iNP0ruhwBUGTvcvz+
D938tykADuu4+M4E90wd5J7SsU3TSSSkTcAeupJ/EJxVzLRz+RWw0251i3x5SwEyPgwvQj179TXM
svI6S3k7AAclp1wVLFoYPFuO8Qman2Cve2mz4MF0x/TAF9LAU/y/8hkfLyAzT+jwYw0NnJQz56HK
uM3k7s9M7N15i9uKsD4EycARJUvrSw2vgUmVk/XN2q6iv86tI9mnGeO0wD9vKE+c8Adz8CVtpvby
BM70WOQtRvJiPSMro1L7QeDSYB3PTCN4MFtOxPMqk0ZbzARwoqZT6RDvGqHaWYWIxNx4us0M2oBC
EmEjhautedZEhisz0Z6lmBo6XN1nO0rLb2RExPnTsR2vTu9sctbA5JJmeBUqJO1qkax2CVACn1Fk
ocGLFeYLow4bqwbz/Wd3BiC9eB6MNp8mKMWItGmZacqzNAho/KvsJWyTIGfHY/wFnCFWw79caRSF
zKlhT86Bbw13qVq14yBgzv7upxdRNSYPeI2HTYgwStXFxG/acscLJqkRxB4aTgQNEWia3VI8gsPe
Baib9qhBOmYWCFEDADLviZjZBTcMkWK6sSxgUiQNoHwY4yLX3A0lz8FbFSo10TGS65+runwUCEmz
4UDxPK/TM8BLWuVhXuMffhajnguqWlUpYFZWYMuuOGOu6IQPUr6jT1nnrHghY4/NX1EJ7P+EbfBc
VjS8gK8YKyJV4IG08UGRekgqqY5EJBAgVr0gDSs5ZwBPVxKQynsluZkOWow/gjSXDwjPW/0hgLI3
570M4dnsaoHqEtac9FDKV22Ab0QWtsf5jR8oNbVd/i4jUv24z+UAkAqGghjF5v1aIVQX6ErAvJDI
O5zrUlG0FWBs0Fx/ch9EGE9XAyogwTs142n9ezvIWvPex9DChsGpLHHRrF6f2Ql5Y1DjoQT8zKJh
TJ6duSNA/N2Em53bAOocmk64s6cazrc1ebWIk3rdTBd/BMmOG5tZv35TePXvcznTOJcUWmqWBEAc
XDt/4D+K6fbt6wnrypKfcqO7gt5lmCKZAB7g19A3euJSg+Pxz//zG+XQbNXeNAItV5B2yvJxcsIc
Vdusx4fdjzXgvkXKRBB34NZwvtaTpqhUrCptggvv6OY+l9F9Tm95hbSvV5G5tVzVkQ2eGFmezoz/
Rmbhkq7lmUWezimjBjliNrWxayScySKYl96wIBkmuOy4Ncloh7ktLmqjG0vR1A7rL2n1I7SRUNhw
ktHavQ44NRHw2cygwgJoX/GBHUtIkzC2VJoNn3nQ4RNaNfe8A0q11kqmh0LVSjJK4IS3/13HWACD
m7JTzXZtAvZJ7Q3caTlm0xFXv6R4n861m1ot1MYM7CMlQX5tdh2FzZ3vEtm0Fwci/Y+t0V31BZvy
f6ueF9GQozXnZWtHKTgyhmLGUYlk0PO5p4ePVIZADfScIAlduEQNoIMeJ64Guk2pT7QUhrmi+Smj
i/7t2TBrJAKJF+YcDvl4519XkoHtIyROoWFA+iLjqz6YRauEaLUVtiDTIsHwXGJ3JTr48CVW3U+a
04mD3yhWyyD6ioTzSqDu2ulWCNSd2tsvEiaEzucvIIvqPgPZjAL+LSbDiT7vJVlJ6yVNCQojZhop
iKiF6O/DI+MjGhGCl5kAIMgjuNwcykT2AXkXCOMvN+JH/IrNmlMA2m1fzzAAp/ANkzxqMlH31QS9
KyWbKKM0QT+tAxdT/5hU2lkYnUuntufJfKD7f0/cOHSsz8NK8PwSog4apIYHVOKrbC1Le4clpzN7
5gBEXLy94NZsbPFiYAHgbJZbgf7DZBJmgcb6+w0hg5A9nm0blac1wap+gu/vjZHgWwYQe70vjnwU
a5wE7k7m57XsuwVfOAq8TERxOGCL50fPzhDT4BP5Y9WxcbdPVcgQd9oI0JFQS3piSW8AQFYC6muS
zy3d1EqkjjA06OLJzZL+gGrEmQ4NP1lJ2T45E3FUdJP5qAKJyFjDD7EwbzJ2opIJBegIk6cx2xRg
wfifoXUeDy3JFLZPgAiK6pg3BHFBhKeOOLhJ/J01vHDYspWs46qKHBIzP2mzABgObllWsPXIRKsZ
jHNrq8WFX+CDxuFGG/W09KgoTU8GV1fGv57Ubohv1whwL8dSdfwo312eE0+7SRhUJJpjeHJ3t3En
6S3rClRf1WU0QqDC49BRzNmpKZt1t09qnyb20tkR46sS5FlRvpy5iduEba6hpMQSmnhuvR7ky8ku
0HJ2D5rgdXGiZm7jNTFSqyBLegDsIqoaArCilpyF5fsvsRJRhTTrNsFhw41yprHZYzAhyOlIuT2U
5KavGDSvhGd7l5JsEZMR7IjuDbmj6ocVUYiYNzsL7iNJgQ3I9a0V23HW/qTT/4Qglo9xpFKfSEAt
W9iib0U/aQJUrvNyY1D0+vulD1+62XP3AKCCgq5UKNVYI7q2e2oROR2UJb9d0+eFFc2gWfD3jxuI
tzAhojcX+9xDIpZxnS6TuQCS+dmMBXAmrld6tndK/olp3pxGZDsfV/OhXXfMzEyWIix5ZbSgkKGv
GN5NJBfmR0AjmGjIkQ3x9Pt8VuPcr+CfVIG1TjYXCtIMClEtCFuP0Av7cCrc24eSX4TwZoL76jkA
lV+jprD01nvJ2c0bZhdpD//niBb0HBYriZvLf/fn6WDoDGKkGEYY0VIAP/5BmnlOv9W8nuLGuJJ5
AV9onehWuLnSMheLYhu90FaDcz8nFR8Lq72nkZCDUvhvJfTNNzPH5k+ij+mB452D5ZEc082cc1Bi
FYrXTupxl+s2OR6+k6JxXFjp9OtICmU78dLQ+xS45nklxFGZYzm5wrgNbfb2dfINBNuNN2i6HTXJ
sYvsa0rpi8VFqRT8kE7NQHVYY8lowt+mUOdD14EosstyEMDEEuCRp1Zk6UtNB6e90GZALI4yJ2lI
r6LiKBAhz44kkCtrQfWb0GFjprfdEJveOV3NspklvjUSblbalwjSJnzWSfzauIlQnhZ8mgFJ7xht
Up3U/TSnVBG4qQEDDhFRZKK4pqQajYWE1Gx3+hUvIZgzvJmWQNHgPAGJmy/2Z2obbRHHTQVF+0eH
Hm9B6s3pk5xQAjHAhZWTJHqRH3HQabwvot/ZIcptOkUBTshnzmhtkBk/N1NpIrCP/vljbri+ggUT
//XLLWw66CHL+mFIP1pufphS324T+r4+7f/bhKdJuCfVGK71jfk+Wbdg4HNinmAtDFy/TO5O3KbU
8LZ2GaBg5GkBzY5kMTNK6+gzG5PrCLFMNWHVYMV7MLjwuKeXAXh3/JL5xi9uqksSuVUAEJxTQh8X
O5L8WlI+YyO52itTCZr0oCXNYsYJ9g58WdziUk6hs6gm+3joeZ8pVWJfZGnZn/rfcK0xCuCwhudn
0jc4tsXBUB+DBKgvNbxxbcySRBA9W44KsevhG6V0wlpk84QqHr5E657G2SPvWlwh29YNTjXNRUtn
crrL5Vo7bdQ9CrONW7O/1Lge+RSfkpzTs52AvcLyUkqvs+nXqQDVxBQ+9DA89Kzz5LnZP0JHpvWy
iFtSDl2Gs68xu8FtA/1oh06lPoC6ph4e6Mp/Is+VJxY4zOYPzcXPdEz1z34zncsjIavMcm9uJiec
mo/ZQq1XJxVcLKiBx+axvCm3SAC7j/6cCyclLTShQkPy+n8H6nloUaH6NYq5AVmSmAxJHncFy4Yw
66fFwOqKy5AEaSbfQC9JXK34CRwpciU6nzvB1y132WyHM5D29DfFXemXR8RfiKZBKJNGEZNvTOv7
07pEOPwwWiO6G9XPUVg5jpLFeNlhpl4Go81gt5I8TRZ3IBBBly2YOmcBhKyT/A7XSO6rvvCISGTa
+jRvTgTU1VYA4vFe3naGcreGBDpfSRhg+5HmVqNzgqZkvyICcnbrgPaYUpL8TxyLON4Zxh5gMuO1
M/1xpcXO+3eimsrhmvprMycu528eSsHPSylirkOAnR5As9ISriOvX/Sxdb8dvJi8u0O60dG2Eh+F
5iukQuDRnkDUCO6qR86/4262CyETIHipK400nR2MHGuL8mOTbpbRDdq0eSbj+9gxv1QS6h6/kKqW
qIj2T3/PhhKKtNkn67PD4yV1afdQqStvce35rGhgBmPIBLshHfbwOOG0coXmMEzZPYzUcpp3eVX2
CrGhFzXcFYYOa7UYHPd3maGB9/fgyz5aRHb8Pg1cTgovadJUGEQNjDgpK3f7jbtZlYNs1Y4urUuc
PAlyIT6GokXl1DQSMn7pUUXBGK2qbCJ0uZU66RgzDAlHWikuybxxhBWWd4hymTjcBaSyFIC7+EIQ
HLljQVP4DiBjZmdNL4KlYR0b4BWDB3ncUyDKujfAm+XhPoE02S4POICX5SuBn8qU349RlO8f7PRP
fQdkF/0c7qXZ9vfSlgrTm21euGJ4Nfw4xygnnI0eiCsBFS+dmrTCMvqQlW3WPRQF/2/nIUrXPuF0
WCJUOEUH1Q/nFnI6k88Ig61kuoWIb1fZ5FU3CYur0huuvXeMZpJ7Yd7Ff1gZDKHmGBQInLpuBEqy
F0KGjiCH/aCDviM2gFG0LrvSKlO7oNHcpDaAh0SdIoChnIfeGg/uzBn24Yg2YameZblxJneHTAmT
+U7aJpdSjaosPneAHmZ4Wp11HJNehFOyx7yCajk3MW3O4VjDV0A7jhIm0VLRe+6wgXdwW0sDDM4l
fxJGe2lEwX5tFnj5J0N/Py2S8ntTakPg5GOZG0KjeVnGd0/NR+NFHIvv//zjzfVNSCTpP0QGkjwU
qoHonYEEGEu4+rB6hw7JcazDc4b0ZNeoShRiFLa+09zyW9NZm7YzyMIRkiFLgoCwjVWTQ6QMCHVD
VIBhv4+l5a6LKgEQd7w4ye9zgpvy3sZyEP1rc/B+xbDvAMymRZYpJryl28l5ac0F5r7x+MSyjrcu
UzGWJPFm2wDnGGqjWoqIUoY1BKqK8GhgdSrWvX+YqdHhe/KyhOFk/hYOmk0DLtM/tEvAYO8ceNNt
P3x2hzUzMBCRwf6APGs3+0oKdpHZ1rU5d8NQMx34uH2xi9qJugBYvvEogArDGL4URXk/6rR5Ffxv
PP+v4BRUwrRyKCvs3tWBKsba18+2jyT2n96Mo4/begIpLC64277MSBZ8DZ5QaHomTI0AWSV1djd6
M58VzWK8m2Jp5Up1QXoCn+vIsc5BrPqE273dCqzRdocskD7mAfuiuV40OxL7cLJlzW44OTGQQjff
bmMIgwbJgUl8dQkK85363d1LA6fdF5dxbvOstq8CiqrI2pClRf/bGz2CXPWxwAMrbzJQM66sflSY
4dhcJLZvq2CwWOJSNkAaDTbd1NBXwalkueTbA6tIJj7xhqa0ftAVH+NwqBSQUUeH3P8w4PzxetGZ
8WvliriMsRRPSAhDE791a3UHO8KMd+2rkzIl2xTqrYSUfitKUhbdr16hLnrGpdRP1xkUXAb8Ksf+
au1/XhIht/wmFF96P0tlb/OpOvtLsNfV36wePqnCuFU2Z8DOSWNmsj1WO+aTXn3gPHxiWC86M6by
ilwC5itLHSSBWrC7GNblRnDZGl1nqlr/nLKeqBlxuPN66Amtg3C/anGCe1DTLRc77aVApQHZykcJ
hAe7Wt29xOX0ECH8KMj76OdOggUtf4pePOCjp2Ogg+V7lkRaCcuYVP0hTKa8cWHo9RqstlluG2kU
TAf6DSChn8eLer3Wph+sqT4I6xxR/Fi1ON194trsG93CzVMz7+MIyCevnbBVucNwNdV0668SK5vl
DgUfkmreCcmbgyl21gdeiOYbsyvlcZWVTBjLVQ87ue/8P7/xpJgC12GciA3uXKEaqgAcwT8h+xQJ
suAG0Du0LBGi3QARUYF+wUKKjZl3wbeaTMZrLPRZO2a341taBoV2C33wWk8UGVtcVy3z4nWNlnyN
jGKQ1PwGsAiPwfMX8zZu2uenF616cnwXrp8nIDIhwVinR+jlDiGb6F4Tu+jkAEkdby6nAxMSAZw8
2v8q/YujxdPpX+ueuq6Pbkh+zuphfxhcPWrF0E2zMX0sVC8cfLDWU0EapAlblfUtbe0IGOMtqxXf
/XaqLL1IBU0ou0bgMOdrV/6hbMrsWv/AHlNtHCQ4f7egiMrCKqjVlxac9CdhPWalx3NVamufJgp5
jJU+cL7vhi/8njpfVNEuiwUZtLsyjPFmfNHyEprO5nz+Dfe3W5rUJqPO89estGz69q5tyQG/UI8y
+gjSBoYvcIeQf17Ple7V2Icc9zxczh12a4R2ijMf2DFINrQi5oUJqoWjQdCsVeIk0bUmJE8LMr24
7O3E9unRK/+urP/ZE+zxlGc0fdw4ImRAs1CDHNhKKOTWTwcXqYXG0IM14sm6X30QSpYvZrwpP3dm
q+RqPc2JNqM6Ib0wRj+wO2TWABxy/tYHvnRM4Cgb2uw6bbkAW5Yy1vBoN467EvrDPqM2k3y1s2o2
yOWpFQVxa4zpLI42IhFqq7DN3aBXxPsiS/SJUQBN348EhWBnpl6rbFjniRa8PTcy8AIcbip8uWPZ
IsggnJzEW07Wk0jHHiEdXIyFW4Nv4z4vKk0g8XnZnesTjHUpPEFZmo5APuih1X2h/xT52WjZ3UDw
cv5RDlSZRVLNgRUxTOleZPRxHPqWDi4K8PhxZwR7UW2rjRE8Ca4iDJVqk4UpPAsAsBrRUw1yl3FV
wzTTi7AtJJnDH/fkLJmm74ZtcIddzygcXfdwrbCDkpCcLXYlqXtzT6SB1ZPFZtxUUtzsgKFZcnpu
9aSSEsahjW1GeStkt+2gYSgxJJ5XsS6EnkP/3TS2tXWet8vOGqHT9M4ZQquiShbCuHeHsWDRx1hq
IYcnBRHf69aGVkMQECx+ucsMqaYP6m3ahCJv50/6HWuVM6lt0cD0anw8eDfXYEcDhfeHKrUFgtoX
R3YHLXy5PJgCMBfs4K3l/M0izL2j2OyN43XlBbikpEOGqbZ5z6eHhTTw4D45XrAnuXGFfTC+J3xU
V+DluZZ8DLTkCs0Upv76ghri52jtd9amBPgcVdy+RDzwXGvsJEuAob+BjR+KqfLbyyAmu/Rh6og+
gcVWVdW8KnpJWPhXzIKEWOtOfby9cmxFnbiuzwZcsmNtKNH7BT1kx3GIP0vjlGt2nZuCyiu/lhnC
ZYRnHO3zI8tF9/fSDf5VEgpjbIbf/j16681PCK6s3+D3HrcWdp35lc/Gox8Lnwpa86lGHAtGKq18
9da4jMuoVh+WfwleCU32vuDn8NUVSZg5zZGervoU2VHtYulE80z6wtz7ZwVC3K1MmQFirye2lLvu
Fh7+YmMCSWyN9MAbNKmotzCd/KQgrMytKzeb3wIuF0zlOrNKxdQRJw2s8sfnrOQeupseBdk09I3L
kuix5sJbeEamwNTaDrpIcUDxlu/kovqvWGeO6wcl23TNQCZ6IHc64tBwFDXEEULXd/7RBDZ5Wmsd
NakmTRdbVFWzrXphmDlV6M6phJ6fZiDBXagaqI6onFubotQEkw5x5wplJMXy75EfkE6Sc3XLb7/n
gROGbQtNx+KBm7BaClQOS4W6BbzzGYK5Bk+pMX3HV/GGf8LOmaITweindPyKYgRpIbwWe8HvYndL
bfMICe1WAkNj5IT+1CC2JZ0oZCt2EwBRIlAmQZGp2B2V/FpKXkCVPMBCBYg4we4kQHecuHsD26kr
DH7my58ew0L0O6ZSjLIaEdHFkNCv1w/SVrIUj+Zr/x7LntQ1jHENMwH1qrDCvWh95LBEdtzel0oI
DYA2X3e+JWUeJODnMddXeE8id8xRMuUXCe2yEonomRYxnQ2z8FDPfaLe3z76cKtF+MyjB44hQBA7
VMSunrnQ8B0VGdmlIdQT/QDpW3yTeHVIf+vnR+Dl3cWzpsiTT/xruGER1mM5fOEcSMQuoAsVNrwU
yL48XKSWCEJjBHUB3Muml7doMRyX0QlCyiN5kxoGIVlt/lpsigTsWAj4IDvVRku3QNebhd8G+pyw
Bo8p7Ldvf6utNrVOE4oKWWb7xh2TgfLXuunStQAw8wM8G02JcdYeNf8Q4Okiy+HfHfbhdgvBtnUs
VPCOlBDM4UTQLHfzzUPe/VfNgqJourKtCzXfu4s+J6Sji+OOkpy7fYtudxafQLvpXCQ6suV5Oe9m
oKKk48G47LSI6bjsqEkAEdbAklQ+5TGos62YM72+Ac7BNqetw2oyrhwWGrALspVxi4J3iLBkpDSS
GHNHiKrmfXviD90mISB25amzgKePA+lGOxw+O5mFdCPxBw5q2Pnz5UmhjR81zkRrW5wMFtzKTK5q
KTlckG7Z5wcpHSG1VSK0jNBbkJlfB2UAhKHn+XH/Lbs4I8UhqzjdB6hlMfCy8GQ/I+y+fdcTEPYg
mheaaJmG6nzV3McKgGpv4I7TEQGWM9AItKXk2BFkH/rVwEcIGkDP525m4s72yZyCl6+0tP+aHXtz
wrBMtc0YbkJTUyw/IT6u3Q86vTAnPVER10GJaiWtG9D5NVEcb3yDJn+l5yrJg4UsY8vNoMniptmm
mldFPSr+bv55vRwVCB9190EPtRUomlimPhY4DTubgkSr8M3FDO6nKCeN6u6rv2gtgNjMtnI65CYg
ZTIFH8DDDCGt3BJ2wL+UkMuYQiVH7Bno/HY7JjoaI24+NuR2bYYZdXgkUAd7GesPOiEf6uSRQimw
K484XGz558F7W9QUzav0Gljn8wdX/mPJ27zSx4KeK4RtMUG9Og+ic4BflDxNJ/BAPTKi/C1HyDFv
ku6rlrJK3DQBxp8zTsjkIr8Q0xyS6g+lhFozCP8GXN6JC25m/kAiy2hcaeEy+ItEtuMI1TKo0ZCO
tfkGPcTQemKAqqO06+xXCx5CmYmmnOzbqsiJwIs8vD7VBA8xoEkM/QysgjXxjozdSz6LnkeXachX
d9vQkuzWOxQjXjXBgnUtAm/94zRBulG3OgeI3f4JzNCEGh7oRkf4OKA9JRKZPvagUFAJg3Kgk8Wa
uMK8/F8qZN4zFeqf86ul61WdD+4FkgMqChpuqrQ4F48RxkUdgAG5lR3sG+O1u57waHpjAwLBph+G
QoI1KfNUm+6PHBDU2qv+anfl/cDjFiRW06ol1FJS9AuzuI7EDlDn7rcnhSwvYE67kqzB4hreLnIs
HRcTyX6GVq/YeIZR5HGlDHq1eqgE66SYOjVFa1KjPAK6F5ZGH0cmTrKfwVf7SA8b6jPRIZ0N0++z
DCrHYJuFuU6kONajA4T0lxiA8IuR4mmXRx0Dgvk2AviCzKiH2FeE/KIJvBYK5wPVIHsAbDgIWeD3
qUwyQ13t3G7W29ARUByVmWAWOV5TP4avtzbq/5VHBwAQZFs1blAVyBRJDHZU38QRim7Q4cUHy5+j
y+o3cQIphuPzQcUAW+Bb96+kgWLpwbPQ+bDELyRxKuSH8SIsXgED5/6C0KwxbkINKwa5VEsR1AOL
aJOzFrj+Td3D4Zgds8S0idbjsdX2c/LsiGkbPNT4FDXATbpGrui53hPnxoWvmYgjM6wtgMP6detL
m9FCDKMgv8lyHfOMsxqN5kclVPTeLdV7928OFtVkYQ9a28bnQWiHl1O+RrZw0UgKKFuNGIfssHd+
TjkD5qRHWfgrYATHLH/9umZLrQiXL0BtlpA1Glt9pX8S3+BH1YUKqDhjuKo825lgc+AYzSDXjqs2
mhDhVj9XjPavfdzSQ13YoqrlzFXfkVwQaTh/iFmwvTWZISCC5feUEk88d6TeIHJl/wKNubUzfXn1
P9BDoR5rwr3eJ2vvNiU8rdxbB10OKl7hHIlQubq20w1SyRb5VGrFjjvJfrL2HVbEZUk6RwcOdbHJ
9Z7Q4we947NsBfUkYbxiCpJMzytzDu2b2XTmVWNc6bwN+eihjKPPicnbK5doR4Jw7OdGyd6KJeWQ
XAbFRHt7tpgVv0PRxh/a9c+oqUwt6RdsQhvO1IfgDSr46fDtvgxyiC0vALpn/X443+Y5ThX4VamJ
lq6YJpoifXFzGhJihvO36ZoIwAMx6ixFa4jQ51Nj0unYPv/eWDRqJq9k0bpwHeFQTyeurJNYST/C
1YI9Cc9pDnSqQJZiqZYYGzrpJw1mqdFXkTOOrYximkRZ9FUAd76YV79pqkXqjpjIiK+WPFBeTG8U
n4bhhIXV0KQ3Vl5JCXtuvaArIVaBQJFvD1CwgdEHCyeHCeqqoc7gYdnipX1B/FRNnD0wHoLZ0CWJ
dqpAyXPRJtj9DgLMzvbBHpbIJlPxzI/mC+GBpT6KdCSwy6kcSbsHNyteXe4CmjVOg9r2MYPM2o6O
26Sw8vVbkf4MxPUdth5YasH9164fMDe1ByG3TYzPTS6v7YcHFuzpGNHArEWBLGX+W1w70FNTW0Vw
b4k4PQjVQGSyS25oA8F/dtjxNcnoBpxDAGwgcIaMdVgKHtAmGUp5jtF/syjSQ6KFkiKzcO2Nd1uv
7JvdkQrSduhqxf18e7kBmXWLMp4DUjStD8RRnPCKNxHWDqPiEGT0Du90+NQvnYrQZpz4W7khTS9J
fVfHcp8k06ANiVNTmRf8yiYVTyb/RpXGCJzypt7yOxnH1WqfJOc3gIZ2wrePKHzWJ1xKHuAllHOJ
k2WyxvoCVCLWEV/myvICjLf5Zo6Vwc+puQL85t79RVRS16f+t/d8XwtOZ6/7GCThYus2IVeRRRSk
NqQG3Sz9Q+z4tUCfESi2tsJYtjEGMFkBuamlEskf/V4+NdDsRDEEnwlS6o1t+/Ygf/d43xcfz0Yp
BUs9b1rodlMAPVIJxSr2mqzeZR5G7n1nIptC/1U0yJW2X7xuyDfx8CfYru5Hay3acpDSlfULagLS
Z3fcvp2laxM+uXA1Ktx6wgr0s3/qY/su1fZXPLXMmdvU36SFD7BRuVjEHNnlDJ1C3dL0bwUURmqc
rCUXtLD63qj9QN9GR4OCIgs7C4H/jzvnYIbtMVi0vjFAYrsAsmlXN0JG4doCV0YySunlgFYj5RAO
Hv+giQGorLjRtcddGnw3bf8/rVFNnsT259MgLHz6buSWnya9DdHk/FUz5tmr+N/cOvag4Zclfivi
WcRl8SSbKr2SsK9X1y4a7y2pmEFyMJY7qApof02Lj3Dh4F7W/OJ76W0kqt5x3Ojxb97nZFXVyw+O
hvjqabjI2oDA2/oJ7MLLwpd4d+8x+8yzw2h4HI7h7z3mhe4l8uuQXTHXbQWmSNgCcQvF2rCIqvnc
dukvt7eVqKKmnIXMoAFaFQCEk+/JtU6u4cqmDUxn7RkCOEg+ZCbmxctNbu2BHXO3R/xVoED4expo
awqtaB5UNV89dKPZl0f1KBj4SqhFL/586oRnnc57fEAzrH1v9CA6cqvOeK4SV4lv9iTYdJz0n2Ao
FkC97tTzu0usXqrW7KLClkyuj/y6JtsJefoSFwL3weCZLkzRdMByguznJFP5vEaG7NZSDSPUgLoj
yOwFinH4j5m2B+zbrJxt5lw2ncY06Q4L8Jd1HR4h+/h8cqIuYCR40STmOWL671/B9OXGVK9xDRHE
26CeulPiw5qUpwqtWtEM4vTI5JjQmsTd01chPNqWUBeN6JQhr8z59OJeg+Rz/27LamncitzGDpgS
Gwya5Fn5TVz7KasZxj7Phr1zc2bgfmVPlf6VJuQRZtKz35CSjqwipcDGuda3PQDNlITPz8ifmLSx
uCmimxuvnnSV58Mq7do/OfZOgC8oqDO6O/it6UdMKY3pHPDQ7iMy2+rqlnkwsg/LRHgOLn8BnVSy
YOTaPbROyf3CFOE0PTVQHqu4VZxTPLuhzUiHkBEpc2QhacfZw4RJBNLZnvRUNzkohJQ7Oh2f+zrw
8dktKnvgIuXQFgGVl3YDhHoituCbFtIaFZGjraPmqCX2fYebeJ0fey8SHQDA1kHf+j4XPTjmfq4K
5eq5EZSnE0B+7SlwpCIPBSsSrtgP0JDI1oF7qv7t1hwrdkZQip9fQT8CubpEnHu18I/xiFlS4+lq
p8GdG3ip+NJE5fKTQs1VEqCATzSAHXvf+k5VznvoHpxAlOh8ZKf36OwBw801Y9XVh+zMM6BhQZq0
DIfULGHngn8huyURbL9x0BjQhUi0nD6k4FL16lgJvyBGDCmUvpEDQIBt5xVsSQoXOTU5hyH/JNLn
BfswiK+c5l8/UPDjYv0uebDNrpezidA/EqpLh+rBs+vnsODAHDBSb4+T+gylliMA6liNa2GLu3wM
ype3H4vgyuA/QRGoVnuMiDLPxkGzpLJg4UizTACdYNEv5gr28F8x0ZjbyZjZ50UHsaYnH531xUBm
erWtcuGdln8ZLrGbN50ShHQITt4knB4DXZWzMnwOg1qieEQYc3QTmS6o28WEHWxiMe8/56oToih6
j0UQLMXqXT7uWaCQ2oVYS74e0WIAlN7ViChtK8+Y3pt9k806jvvjvkDJ/WxsBQVNwYaOClpZANA2
2iXjG2ylr7quthUCaqQLPfn6ZVymCdR5lJ1X13aAKw7jRWjvYB/kLDqSPpdMPc/cmQFbtGTEahs9
n/eHsOMgWa/V5x8Ky9pCcIKrlM1foeY0K1cz6rPRuvCVhP1vGutmyCtIC4fL5YNkIirey5NFfEbc
kXOgbi4838nT6nxi6ZFqJtkOzYhi+p4xqAJdUiQp52NPXe1xdRYCWEa4J8AeUKtGJUtcdBDagPl8
pH6o28VvQOBNWx5weYygtw0VVMvj1BeBTp35Q5PBlEBfHdWZflu+nEEIHCumPWQmL0FZyi2xBcFI
1UXOGhIZI2FgribVZhSKGfiVblhaStueoLbEKn55OPzlqTiBu6ZUqmg9S5PkuQ3gRTjoeet6sJke
rxIIVRkBAwpsE0Flf6NzOJ7XYx9i49FUlZHK9BM3Z8U2/KqsZlAuR1fMmF9HVzK3doLsvRD7qGOt
7dqsGN2cy1HnrfgrW5EUq2YIOp7QoYI/M4o3LCH0NhByxMrztWhvFqoBMMB/I1r4urjHiNQryMf+
NZo3f4yWt35qv8zMfNr1qIC/pWfUkU5ZdpWdHcl25UoZuBvaJqOK4zDfgyfZKny0c8O3dUBquJ4f
5K13Kr7eNtnMTvxnbWzkAgwcmpRXKNliK3/WdAf2k0zimnOfz6Qsxh1q0YmK6UgC1m57BPCSmuo/
Qf/AyJupNjv4EckPrEMenp9Eu2GkGaynxEWRFst4+GytTym/WmkVsBRpPKRS/FTOZLpi/8dFFset
OiV2mJ/cnvXS3w2q1YhOa4DVknt7AmAiN1J3Wd6sDNYG+0wnvKM4P/Tf2l6O+TTG3CBFoDX3FjGo
wPD8XBGTE47vmSOEDQpLuE86I/4sN/bKJZjKovqD9HnZmIJOxeYIhXgNB+EijeTUd7M+d/XVExqS
k0XsrXMDRIUfgK8dO8uKR8fMhOglL7yj2jyBgGifIqAgFqpLFRtPJoEFmAkqZVe9az99hI8OT7Q6
rcMr2giib37HFon99dVXjn9EIrfzZkr8rqbb3nZYHxnTnkg4lptuIG9mB2FEc8oBf1Tw9o6w+/gB
wxeihZW+m5PbnuIUplAfZBqKcSHBWUQDl3u9xGsUO5cYxJ9A6ahd7yezMHZxW/LZrOYJxFwEj6iD
1UByDa7wrFePaX6Tl+RG8ZVMQhRIUXTB9UPx6DW8IVIi4bcBizo280UXl9gIjmmMjzwhe/PFIkJX
SVXdqVAOjb9nYLfFrXV1MtDn3O8mwzXoJZQ+8dX7XClMHjPHZsxINZJUZlY7VPJphsifjiuPZHkJ
ihM/0tLl+Ffc3DJ9qWGF8eZgb92dK+8Oo/oqjn/o4wbzMVmgIH6+y+x7v46zDxuC1Lv0ujrEm5cD
e5CCOi7v1DQCDZnSnn/Rz3Q0uVmyRolRoGUs/7fIMM5n5g+a2UaSON7HBu3N2DpnN1MKfqurt+UJ
eA4S/T13IOBxsvfpva2DaOUA4TufkNs71DDmwpnKGklh6eQ3+V8UuGSstlhY0j1Y/MZ0hr1twYBR
ywz25eGDNpgDvffMasfZlirOxb170RISwZ/3MP54Eeb6/210ktlPdq+PheRRK36/TDADZ3A+vTau
xxUfriVfyXyjwGzqFm1xrIozk+rbGSFiMKLjTrCwU5B6EXdvgHpEt5eF0NZbBnU/K4vXozhP8YVo
eWAc4XHKMuoosCCmBDOzD2C5g/en+DZfY1KABqnfuE5FuTFWph0qVBksU746e891d3YhxKsa2yLw
IsiHxfTEOQgiiEjoLgc5edVtYt3ygGozHGs7awF7Jhli9ElM/LO1rw+bQpqhi1p74dTpGJ2J8khR
WP9cG39k/FRSsWOu3rFgR3BZk4/8Q0bY7KU37nLTJKywxmPTy///YqQl2rgKGVRiB9UfdiJVOeIG
o/d5xqLQr6g2KT1hBBRgZy3WPuyZfpMB/+AGom86ZATUb2I64olPtLLbZ4Z5WiefUin/IDaf5CNh
tVQVpF3n7UP2+/TCHl2LIhGmqkW/McuvBXWctI8z34ZdSPU+1CSy9NeRBqyDcJ+ocX2KJBnYAfkq
l+k19UJD+ZJoMjug87GhVl1kAKDFuHkfZRcJ/WU/oa9/q4fQqzz9xL10AFsehX5d20iA/YSN16+w
HZuQeHQCm7QgeH4s5uXUuguIbzTzD2vYPEHNaus12BCiwu7gdsv3bxORmTQpV5jMcLKSTKNQt1MR
fQGXPxiWlwMHBnN4UdhvGLwxbar3UqqTzd5T94qCNyZRu3PzwLf+P/l7FIyT5JGbs77LWzbcsVKX
h9VNWRXIlwkSdbwTIfZH20Jl1jzOnxfVtHyz0LS9+bgk5hef8R1bfASXd0fpZ0KA4uE8Yvs9hUbu
wYZsoSOMYiB+Py2gq2j3dDodaz2ml/XNSDzeqFARCIhuYYNtTdxqou08VpxFVaA31DLe1jTWH3dG
Qur9i7Ff6haZkAgC63wWmKNRXl5oSOhhIf63Z/KRUzFdWIwajnz8Nuj5Hc+TYxSYbd1wIezd7aAG
nv3JxtpSdOyQeMxiRus5elNk6KO5ocywOnnGP0Jxex2oja2/yRW4JA0V8ZoKDeGgvFJtQyX1Anp/
mmT0lV/GDh0GIXgqfehWMELCNw8msFmcmNlFS65ecBGA+WSymPSZ65/bK0OXa8ftICAy1J+HX5+3
YXJsOW36Rwp/wfEzgVtNcMG2skLpvnSbXfkJMwUOTeaiLvh0JXNwFwhkwOfw7w1bQ9SAQydFeFCq
7pIijpTS59SKugV2Dfkrfvw6Bh57zH4jxLQpMXPO80zAQkUqRVLVAF1oNGw6lya7sR3sGjkGciGh
pov2B9I0bNUvkGE7nGqPHkPVF/ujARu0oRNnzTuT1P6+5PBlqOe6F++sboK8vp/VtPCyU3tg7s7M
l4CO09l7IpXzsS2jkfHHEvpDgo3u5mJtnUlakJ+vvKEwG4OytU+RLiV9pcqRVrS6NTZoHN+QEhBq
PPT7+a8o04Mak5A+766htuuHVdIN3yrKXeHfGsveC5AZe3rMIbXejBCRNfAjYQ9zmFMAqprZffMP
41zwRXN2q+iWz8GtJCGE6ko27USnIT931PpHQLnb4wdGeGU95qCzV/XontRk1E+jFXtj9nQGZizN
wnOg8N76y987CXXD7ThwgbQS38CVEeU2DAOeL9dqC9Rc34c4qvmqtI0xic334QArBTxVo09232Vo
UDK+VOpRmMkmtZME+iEJ6Yq5DTKRqt1m1De2d1uAJNWGSpYr+lbAjTX7C5pgLrUevGRPY/RldIRQ
4LVU4/PjDSJKatQgmpOPab4U1rq+a7WSfXwsHksJ/158XccUbNS93HEZs3mFX6DHwobtQPsFtWDm
UmQWUKshvlqpwq3he8c937J0Gecc8/CPB3rZZkT/fdoNI1PSIGv3vj5WcZlDFLDwyCcbDybrldiN
2Q/F3vkX+3MllmWhkwFZxS3HmJIFqCZYjEhXytFW8LKaUMQQk3G17jFCHVz3V1Wne0e2Mt3eifkz
vL2r6jORx0nrJs1cPOY4kt1uMNWlT2UXDRp/mocRSRDHqOYB1qup+TmiKsPnlCMx7FtmTYoGws6m
UYMx7sh+YZEyfh5SvsuCfrZ9GBMyT2mS9mhFr2CXuANyd3het6HjAbGp7F6DDgP6X4ahQWBNsivt
xduRUkyB4+ObezpoSq+uyouWvZTUCyysycx3qAjz751YtPOhbrP4nRyEqxkxLDsfNx944n/Z7ZLw
Fr0JWq0qiNo9RF5E7VON+04mgNvO4G3+P8DVVnSpXIRXEOxFyKKyY/IQUXhgo6gVsVEn3lusOdN/
nMkJ0tioHgTuwh/nvoAn7RPRqc22YjDFX5mRaghDIreNSfIACqSJK86FQVeORt0pM+aZIqvHxgK8
JRBELVvfo1cjO2wYPFCG/HjWTBG0AT7Dk3LYYv1qcYgNpmLBkujP/j2JSu45Ud0+vn6WHgcjoF6+
39rivguOxe+dtMnBPlCkSfJe1I0h4F69Hxot5Wnli/qBv4IzxxQtaqXvForQbiFryngpAuUKikTx
/vEhfpRQPvQowpP8v+TQmBZAq5w3vdV3IE7nr4VVnIOyRcP8q1XKxReOSgYdUdQLWsK3qwACZcpI
tkzxIldr9LWhjXw5AgVqmIWzmNnOaAOmVBDiBaWfbuSGSZw81UMBge7cUqeB8Az+b3D3b/dBrj6o
IUCGwj4B7rhCTlLpBl8O5U+3cF7FPeuL74PArE1Y0rOXGlOCuQiGgKtLwEvs9U4HIhO4LRqf4ADs
Z/Nep1QDUufnddRRBTCTtoM4sJuKlGjxjCv7nufxDEQtanYcF0KnSMUi6Lx4TYT9YXe0VcLyqIB9
BREBWJ5ZLjN01zeyoV1md4Ha6pgWIyK9OgETf1aWcMdj3kD04Isb8WP3o1ip+j1YP+j590OcjwDn
9Ng2AbWMWh8U5kLIVgEU1kFrmkLIBK7z4HuBsClrn4vsPVkzTFi/deQF/MqR73vgmY7oCRNKRjWE
aIM8gGjewNswhjZj6Vaysf6A1iauC3GhwcwjrgQidxHMl5xG8KO7CeQLaBbBQmAjEcX+p0aieeLX
rFR9wkASBawXLGLp7IEhUy2D5DyfReqz1rGgsXW82hFr4kkvUn7+IzMCkHxfYXJKn8jbI4JAbggH
m/6QXWVtnpcNW6PYLBBjqqLfaTdK52xgkwuU7S69qI3p7icoqEuDqMRwjMWgozhhDJ3/LbRan1ZP
iCTkL0XYR/tGZ8burXIYWhm6h9ErFHMzuuXsfLyyfRT9p4zxscIEyVX3QuOvQMS1ojJf+jeQwRvM
A0fieWezKA7DfG8rKsGPsUY38p1Enw7MfY+aGTTgzauN6/M7/VG4UVxVkSNVEQleMDdYF6hVvAYA
cvz/j4lK+/mCaJ5uY0vWUsT7o9tln7Z/bqqve3Sq4T880XDkpVqy9pagVVVmsE9ubGb+qGwVnIuD
jphhGxtRw5AKocfKSzrbFomyQyf/7QF7DL12rLOkYrFKiLZxdm3fJF87q6WGl4V/0iLwiqO+pX8d
8fUZGy0rFlv/qyqZHXcOz1I2eANAH70cNLI4/kbppTqNNuRPEey7XCTV7f1vcvXGFHCVLDCuAYjR
MSd3xvkGzXID1UkopNAB2xZTjiRAvtHFvUHwfMECZ9sjTnEEsiybFsox5aJWn92N9oVdd3NusKIh
pKa0qNovE6HwjXtKaHzXpmb/axF/CjVwUTAXyXOE3kYLbrECAM5tpRT7DvoIkye5qlL5K03adufv
lRUvGH8QrxzE4gFfqlI6V8jB6T1TD73AXKib/o0TTvj6xb4K5FV2KNwJ0jeg5OWtY9eU9yAfuqp/
ytmYdMdFjF+e2AzFeF2GbeQlxqcPGoVPpY9CkiQg3qUstyEUVtJpkvuL3GdqD8AKAP7xpWazOnpP
wjr8tBW3e/FVxLCEyRPP+YtZRDfvEopdsD4k4BEMLyc6+AYWkAL11QJJHuqfwpsk8nbzTx8aKT4t
oMG5k9muWVMq4QmS20wMJOGwL0Jn80EIvxR2c1/iAtYg6QsCXnDIz+rFokiZadiQJ/2zylNgriM2
XP5hL9m/zhCchdtBukRvPGqeGMemIFcAVNCes4AKQytSht4563QzjJV7K7Il8a6ICSUmgZ8Jo14Z
avng+7dNSOpl27VRtXIGmVxPR61x9urizGkfw1u4xzZRuiixftbpjXlxFmWuS3adMYlxkUJpwwSK
vjbYk/g6UKzgoUrRvYI2lIFrgDfWU+2IjMuj1iwSgzUjleSP5J5aKozlMVCPbtVcm0g+Xhqw+L5W
WT78z0tIkXpEhC8LqP2G1QtKwEYU5Yj2e3ptpiIaaXDgP3zj+H1HtAIj1OE2hRXS8gF2VPJtrIB3
1+u1fQ3Fw8aelCW1Hs/+1GhfUBnQz61gS9iYo+vZgk9vIUVF1pLBmOvqS8DaQp7C+Jc/W17F1Jx7
IW9Wl/eOA61WhT2+zZoheXaK+gZ5TgTyhUVTEIfNht3Kvdm2e+vb9vHDjqjTKTJoA50uMPxWvNXU
IVABRbKmN+jqutfbQfP4l9n9YN3q7KwyMe0udHl0WDRCdSs2qDFaGjwcTkRZqbAQesL7Nz4G0Njt
KC1ojKuHk0IJHZLZ2O8jruOgixLnGNWOR91xxlTTsSEYGGUwuOKgwhqqx2qZACkOYeRM8LLJJfIG
iJOetF0Vf7XQFNqQkD3lnpzvauZyZomks+t0kg7v6lbrDTJk1/Q5XV8r1nG/KUZEBm9jQ6J1ZcFU
M0elrZzhpXk8s83qCktC5r08SiwZ0EHkL9z8qe8kPCIUI6OHs3smWWMRyKGizt8FFQPk5jxcSeBr
7KKcmX2RCax32Bd6bdOvpDHWQS7A3yS24hjHCROM1pw/W9S1VQBTM+9VHeaL4QGFlIbDlhVD0nC0
2lKpgtmhUM38wPz2phUMUT48EXTplogrdBEYZghoJn/f1mqmzgTCkLac3PPbXgM+TR2lYdjoImbp
lTXVjVCtPXUGoeHj8MHUEEgK1Bl4SuGb9GqWfNsP9HqUl59j3uh9nU7wciEoAIV30QGGptVR01dQ
gX9mRDWPQ3wFusmQEczJ/unwapeRArtlzWs4KSPwKLtza7r87/dSHuH3dws5c17OyNLOacwZVFFg
CLYYRpgLkOveMKKSMQ8PUxQl9Rikm15cce8HfetPro92WeYc7CQFd2uuYQ7oZsLrVOs4iDlqx3Xv
WEbOPTM2zS28UawqkNN8YJHxtirUQTY+oDN7m1UUrma8Jjone4uB8PCo1/l57mb4Zz6wB1ggmGnu
EbyhNtbI5R019bX8y1IXOP73La1UQrTB1Awwv5YBLhsvd0PIdOzV2iedlq4TmCRyTt3157fu44tR
tlpfA7xN3KrGzv8rZiIQ3di5YtK8SbsENp1UuK0lqpzpAzt8mTDkO6rF5+6sfqBX3+NP+p2fMyHG
SMwyPH6gxNJp7Le8JDlaV2TPuv3qNkyqyLJZgnJSceK6wnETNcf1z0V3/EIrnKyF5jsYrGPZvEK8
5bmC5Q9CX0P0L3cCKguhgdDIktYvPcwpx08Smwbspog74n7PaXfLCs+mdyIm9LXmxTXdvl9MC6rz
gTmNLbuC+rtAZ97tfOsxwTSnOKgrXsJKiI+om+WibNNNr8U5xlb48ug9Wmzal7B+tMlIbKpZYQuZ
M3joaaUGVmPOWeJp7VJK/EOSZH0vCjgFEU1MuqVkH7ASSys8pQlzXvxqoA8HMzFNs2jaQOL5z0UF
8czRBS5PhzTpQo6QV0e3WOAh5tJspxVoCCrKcwVtNjhqdkrO/GQ9Phz8miKykTRsTPb91f2kcDI+
lYg+rASjvQzbko06LzJ2pe8LrrP5MqZ1Mhm/PZkHArNELsXEblBxO2m6tXJkTPKNr4pqvvTXxwSA
vIemqyklW3RMtBgsK36l6HE3+On27ukoVpycvDon6fF2nAR3UqC1UJ10pNMYmDMZNgpaZ7GJ9PzV
u2qebaw+z/qlynnsDrL13pwwAq763ovZ+Q5hBnUIGLAPG5NKaPySLg3FVkvsfqgeWU4MDcg2UiTn
Em8aIXFTXO0hJ7XaBBfHGKbvh8plWVD+FQaEEC/u3+rDcIplOLCiARKzfYyiMmLxrxqJPVvYEOHm
iN6eiZmASdFqa6AIP0REkH4TkRmAUmuvzYKR3zidwix7ltvAzBWmKxuw9htdyVcTNGqpzIX/T+eq
PTKunVuAVTmNeDZYUPQwhIEnQT7SNYt40rDPTtSeunPNWi3Dv+1v5L6APzDD4MtyW1d0RnSUnXEw
GqXW/yoYo6xx3xol0qMKXBNe8AmhkjqseIihvYCGoo36OhKaQ4YEwZBk0mnHWX0ZtNfPj5jXWXzv
W66F9uL+hSBmB3/yU7e2/t6/mzzchLG9SOSaJjJnpKovwmULY7gHS13j5AIeLnIx8mJlvCN6LxAQ
Pm8XFxuT3Hm2fQdP691hJ7tw1h15wI85jxEh9DOUeh6tv/6jswWRoQNAu7rI19UJFhzvN88JevU4
+1MgCq1CSPVef1vyoOQ/0i/PNe7JnxfstZOdAAmdA5LyUq6oZeteXV5WxMIczAcEZe6oSn7/2iPc
h6w3EyMjyNoF0+45gDgd55zTG7O+oCrwehoiz7BwpPTz+KObIZD0VCCFMY1mve32D4I6wUTeAGM/
tdZ9dcLZG4mqRYdcM76rFAgn6vl6Y/G9c+uQ5tCM9wup6hqJl5WeIZ5efy8H70CmrqFM5leWWyQV
HPmAnISlPPX748tiY/vydbNLQxDUZutaoYXCFtR9XMahtdHmY/jZyzvQLAj17vUEbZehvtfmFhp3
EDQMShEitSJ8qxBjOpl3pmIN40bMhtBC8gotmSx+s5sFJpUJJaPVqnKYYoyyWGT6cW4JbCPwvbbS
P6VC+GRcXGKFO1HUeyRfB0KWxSQ9Io4HCKa4OvmA8uW8c0KZYoJGVGnQUgAnOvzXegRBjEYJlIAJ
uKxWZkgkFQbGQon3wPrsAGRzubjHsf4MlMSk0Kbkvt0MbmH1RP+u/2HCCdgr9UNbXXJBCTdQ3xz0
cAsjwORFvTYnQ0I9zVunmYNYPEK8LVagM30cKvOOeynOGDPRwPXnoDGTFb4zbrKotF7x2+kcOUDq
hCecZ1iDj09qWqkT6kWwmbc8GweG3BXClBvMSBL+aMRzSIV21tikAWZQYbIwS1y9zKbL/00ttTPW
CcmKT3aE+otnU1riqq3AGHDLyUHTUYpx7tP0cT8ZfualLUI/ozxnzhhujaCthtmacgrimbFUGoux
cyi+taJbcepcFtZdEj2fpMnaSP9Ci+sJqq8frXoSt2GiDLv+2Q4CrZRCyZtVj1Rkl3CciNv4QOOn
QsUTzkZUVidBDP5g7WVPhJs8tJhY7OIqZWpx9U3gs6CrnbztY8Jtyr3H921dpB7uCeODiVX6Fc31
B1cdTyPyRqGNXb/5dQg9vEjhf7aCztywVORq+6wbqb5BQbaBLY6eY2aHiohRCRjUSrMtszCBLzir
WJwiuCeF4ETWXLPG3JCvqLHTwLnxTOG9K0EJ2zxFR891zgSqmzHvAoeFMnjR47S1nOTDSWzb1nfh
UQ6cUQVXHNlLZjsIbEgKYVggLf9FktaETKtJQEAErFYhiXUDRiO58HkLO8Qu9Yi+q7v/m5nJ+PjA
NOrARBlDIL9MKZahgMR/jrBlhjx6q1ryrSoiFPI9wd1oJ8OPYbDbF2rvmQNkwRsPlzUlshsE8/oh
GpjH7gUfKU4Nd93exPzcWpsp/Ja6+Rtz9MEYEO8NmfPGkrUUMugeiHxQ0DYcmzDcagVP0AMo6+v4
kIgPIiv4hIFkOn3HfdtiXdb+687q6EOtmaxcfhqvYM/+rB1ueNEmTRKKnqvSe11LewWUZ+7ZlqDM
peR02W4JCJowLA+We6Va+hl35F7Z5eGRcjlF7qRqla4Hv/dM4LqRbdJjAM4lCOxlNVI8kw1SBfiM
AZPWzunA/nuTZDfAILt7vnrfXnWGscoQFDQJRKi9S2yLYPHe4phCwJj+hXxW/WRZeAZmV1Mg/GAD
pUaCF8DXyPDTHFSw18v0wPVPBMVh60lHBG2ehAn+p3Wa5RZdgatxVGWbHOiGmgmETRerhfCX5LcT
jUL766JikykWAkc9QJF+KKVh1RHCnk2D9pRimu9inNfWoDCwjUlocKxZqI6S35FDCUrHqOGmOMU4
9+g59ApK4Eh+awvrqHRUlV4ut/Ojt54WG4+3pb6RHKAsZIPkEE9123Srse/s9KNS1j+iS1YdwtXu
0iRgUDTgo2bV+j80jHf8W6JdjJzbFpR1nTrmQheWzseyLpYZdWydHfY2obkFY/3U9Flqh6QS++Yp
ieOAKxMX4s64CLRFyqchCxLgSNL6fgctMfgH/QRIwQUuoCRb7V1dvtCuwpN00bd8mgf5MIt0yBx5
Bo5zxt2aZ4wu+LqQ9UJucztApe5QDStg3jMTCuPDBH5jWwIFxVm6QgvU9A0ZpcHbu5qf4/lWpIDD
PJuY3rBuDiuq1rLnGfU9ph03G3Tx9swgp5sKVrZzPl1X0dObFIlPuEpHQM8TCVM2XuUTiDnY5xds
OJ+O+HBqr73K9vT2MIiDeJmRabHsdjwpaYvW8PslZmj6E6OvJObXuGArOSZCXwE8MZuYB4tjaBSK
8Y6o+7prqP/OwEHQRiAnQ2R/x2Q5sJp3exFyB94t5d97haBKGfH+Y6hQO+JbaAQmPOEup/uKJWsG
+eZsl66imq4EM9LGXt+BsgoWfry4uvz0rtSTuD8887FivVsPv/io57EdC+0SaNdJIsc7k+s9Qfu7
+HN9fWo0PdZwnKZv/L3tJHsw/t3Y3cWUNX9qCryjP29iqosyhrFJI4cnVTGncqBiQ9CES9OdXlXG
a5SWqzr9uhkHGLDNOyWaEkQhXMY4aRhFBls9VT1onX+UErxQaEAG7Kla6vtI7bbPp1QGQ9HZSWI7
89Ovx3lSrujDTnncY1bMUp0Xlpq0eM7hgNaLvZYsey3q9lvXndVoWyKGdBPWN0/cjdk2BLEUCp/P
FQTLaRjUplKQhnUfPWJpZjBvrQiYpYYVLyrhkLd7oz/npMpOgjqJonitqQy6nmDd0ynxXBASQGjz
jDdJhQG9PtOyAqEXgJ5rz35EqGShNVxX28kZP4L08/dUH4IW1ljmz3DCCw2lMJOKy5o4yPRhFbMS
8kQhI81ELGBVLeaQJjRK1AWpwFVqYQZ5heqvzzbqKY20dZZzY35yBHDWBsi/4YfIcAOTQg9q8X8k
HIxWBuk2cwF7QOjGdldK4ShJ0HLpqKvaMg3UM/FSZMksFWqK+o9VKBWUAwspXsZyoX5BMlwygVrm
Zo4/YsDpfRj2DfGSvB/3bfstawj07p38GznhwERFYb5V+v9D/fxOhdmLJnh+YbDIRTwlpVj8GBL8
lWSErEzv6IOiC4sV2lpwR9YqW5KOBUgUdYlq6wiyMXYIyx2gIiRqQhVDw22FHXco7vkKzeDmkS/a
NMnOoEDQlrMUz1rBYfSSs0KNkL4Eg60K6vrySeXTDEltAfjwZDPkQ6//37keB/vXb0lzUrtrY1Bw
bVQCSZWf3EyuXEx+VDhlA0T5eG2r4v5h05fZzdDrLd+S5VjbUttx5Xdt08RcXZDipeeUMPS3BQob
dUtbnSLGUDv0PEcHaaJzN8ES+Q3ne1R7wgMHU9dhBfQFkokT/K+L+TEkzwU97s/jXlSwPYkhV4yM
jWDCS9o1GHLYJlZ6xGyEQa0h0oEkLqVW57vnOmJAnGM9tOWRPHfbYg7PiP8Mf6YhSnPCM51Ka0As
93v4iwalHFLPM1+K2gmkTiI+mcshK/uA0bHUJlznRknk2wQ948IQq485gLOQZrVbCX+t3qy64NOU
CghCiPEcmLs4K3ekq9vu4BUjjOFlVuzROKmIQJSg/5SIylBO9I1F7cRLYAjQSzwmFcY3DHmg5egR
9R6uIOEjX9puXZiY+8c5r6fXY+h+P/tUVlu81sL94vDpQBd+CGo5QzUozjVUNSQeUea1c4gSp9Q2
EomMZ3sQc1WYcPkGxqlu95Y4ZKPKhMecWAO0bJyrLQTMqN/IB3j1h2zu76U6kSb8b9g7lN/SuQCF
rT6GrVDXxn39t6KjMILnatSD4LdVnLVgJQEQHwuzpbwM0Y+AyinIJU+Fbsr6Cx3F5mUGS34H0R1+
8FWeEizBSd/557GovG3sh0lluUM0j/xW3bI+/svcvI3Vn3gs+fSEpK98icg1y0l/hFCHCIXZ9OGd
W16UdZrHiX13NjV7kREMPs3MCueHZI1b1krx5b9XsGHV73GO2IAEUYKq/xY+oppZHenpkhiPxRoP
xysCF+ItJVKHs94Jq08eLTRiAhV3vLnj+9Xtc5RgpLInyN5HjVYwX8yM8tDarkw/IG3FNrd0AjQX
VSZVNzhoi8GhKK5eSxjQr7z+rYiRA9ZJ5JHqv+nQwh4QLOcQ/cYrQ1/KRhARdnyul08D9i69QfVK
MmHQBUtGHJWDcnW06AwD0TL7sb+uDLfzGVbgErtE9xkbWkUJ21WQKxHlex/lbaWcvKV9awRuC+h+
d/evp4116vJ0SxndGYZxDMe3wVcPGmNOj2WVtI4h7TKMDloem3dBFRAVt8kBCY7J+uXP4rJ6RKL0
tWWut0vZP3oewFS0/UOW+IMh4YXIsL2tciFg9Ve0e5HrFud9jCGkIsrG+Lsg0OY9XzkvbdqMuqPx
zFaPsROXbL/O9hLiDuAu81i579gKNsSh7OzKD5LaChhuViSurBdDeDLQCRTXVlRhK8Sn0yuKs2im
vapV88HkEOcVNK0ZsYtLYGJp3qsxbt4wrewhC8iS6RPtkBw/iQvSKMFkcUUnjs43xfjo/0MDXQNS
m7YkUI3tef6HnVj77HV0JEVbAfUEk6K5YzNMJUSe8bVNGMIpMWHpfBqbsg27OWQgZ0yE/hxD/gnP
xfUVtj/jkxraoPBnAsWiOUvY+XOp5aaNh6P+3zPEmb396jnHfe++RkNyWnQzQ83ZtZreYJF7Wug+
gUE9ZwVRHGqA07+1HObSO6RhMFJWZ2FaBsk6XGCCuVzoc1nsJBGrAlHOLVWvXjnYAYLaTBQQKanT
7+eETlGxLCJ0acFLLnQOLQdqUuXjvG/0fNFDxDKupq4dIUChkOJ5pZ6M1/9iKtlvFwg/1Crs39Zp
2wOyauabtOF/jpOSYmjE30qr5JBmrhaP8vHR+gtDJ/XqQ/VPmi4L10EJljkr3PN0u4+xHd+nwIqc
0uaXeH2azl2uAwVpkEb7GDsaD0zGofceGb1kz5kKyA1JCFjpad/JjisJdq2KGAJgI+FZ8RIVi71/
gsiPgaavMJTF3xgWzcTpv6kEcJHizYjso3c26TAGhBoRpL+F0MeVsWnVYW0ApbFNr2bbKN3nn2C1
Y6CZnnj4YnUjncNySKk/8nargNFTXRCMtGddpdTqbHn/1s3HSZD/yUIpvb9gi5OEeLewGtYi7udB
bhhfuDhSlFcJeF8YwERQSE4LN6KV9J0Vl7NV3bz0qd0Yn+rhjduxxeBCNqPXCKMnEK8LD4Z+RWrS
IAKAQZ5lqMj9GqIiqkv4pgDSD9/5wVmEb3xhKVgh6ZbtgChgEcUUHG/1CIzt6ZqKh9w5PgBtcRxo
gVHf6UbrxyIJIeozmZph2NsokY+8l5DaYP2zozwF1arum3018Fd1pQZhrJ/613DQCARRoiFJQesN
iRMqaOGTOAkfhqNGM5E4Gi7m7WLsmueRju0nwVjkOeeyNjma1kY+dxMKfigGjT1GGW866B0iKoWP
mILh6rr+Qe0zJxv+72mWRs0VvLx/obGen+ahUj9Q8f/tK37KwD6jFbiR2jJr247W4Vt1s2JavXW5
Zs1PYqUAXsF79ikS7A7U4260T+Rav6SkhxO+TKkciRMrhFtdZoSFlRFsccDqhIWsaCE0lDNMR0nq
oMRYxbDRMSYd1WTk7xXcj4DB95dJzZFs+aNbsbNIp6d04IPo4GfwVgxMZ/VUchIcMD3uH+MzqjBB
lzL3bRaGS+DxcB6mopY70WuELB4MlK4k9P9MT20JqOf8/Hj8rg836pK/jSfgH0Rv7qAvVR1auLzC
CQ9V7yPbAwxNQPrLd5bBWhg8L/+7mVAMlnRtcxvY4REwkuG3USHTFtQ3u9wG2lTZ5dMTkFUgYwNE
4fhFUYFGxva3KGwZOQ9jPfrQzfnrkc6MtAzRAgxdIGOrA+P1Zbly+3VpQ2kD0WwJBEd+zks6XweR
mkD2Un0vmodOsDDpwVHKUgjIwQ4i17IjdSnBrgJotn7ORu5QAv0gc5h9GmbUUWjzcnPYXe4fHzJe
mMgYxOX5JA1snZ6m4wUuaouj96LbIrXPsjCrtwKQ079a7nEmUkPmV1REOlDxLUn88ULHpRQ22Vtc
gArIpreZZ7xsVHVLivWU3krC8EXEroUOCxLaCIFkJK3IWTtlsVCvRyknaGZock559vzFFvc7pHi7
R2xYpsS+aCKt9qtQbCUhTS0+JQH6kmqoMSrTsRgHnioCy4vm298TuVHmrjb9fLkp1wUkgkB47qII
ypqfn5jKaRP8LOSvp0tK9Z3VPIe3TvwK6YBYDpX9NHD4POFhiL19E3iTFK77oHLc6t7SugZDHgJ8
U+i1tmm03OpGGXDktvUTg2isrffYCV9QmARSfBtX1AnMN13JveZXFAjlk841RNucCREK8X9wgb8V
Rv00EcZn1/8bEwlrzjDuuuNsiX/UATzDGDZzvR6bFusGdeZ0nMfyfBqrn5eD/i2mSiSrZXoaO54C
yQW9i3YDgLwvOWjZ/k/ZiVmJ3uyZjBO9XFKp6jG6H3ITK2lhZHnMdjFll4dun5K2+lXCK/RGBzHJ
csYVOe700A1wNCwBAFw8fCZD999ABR0Ojb5e4SLJf0mOSjJgPRTJGAvHUVGwgXYedGe0/+jRD02D
aAXKE84lgAkOBi8XHDShyBEX3VodfoabtCMemcdj967F3Is5GMpaq0e3GKqW7DRcs49DWYTd+Eqn
Z1zMbigT6bMBgTAy5QpflzZHCnLlxnzVxDihr0ZsI13MloesG54eCTIw8X5+993SZEfYFd2F1joD
hacgJyZMvIB3tVJOgz4OACp+cubPFv0Zf/tGYxUoCYh1ZPd+D8ODUbOomK/i8b5ouuy/HQDHVUJN
+DYm7cpR2PnFviYfl+y2+gLl9iTb5Xdx/pfDvvCu7GNyr5586a4/zKJgbc6CPRA6+2pve3AnAwEY
OTaYYFwye8ilaOQGFnikLoEZ/+gyaM/n4lvy2coh4AcitIkdP3HYfMLnEV7NM+NIYOHXZRltBGNI
D69OrGQ6Wmwtks/RfpiVImcCYRyttKRuTmJs/62hMbZixXVVn3PH1agv3uNbivovIz+n1AsoB/E/
hHURa/2SlQSlS3mzomx+02YPKsADYoETabGweYFK2CxKUKdblAy1geQadF7+SNqleoXUO2xNmbVQ
AQ4xQJ/zkqShS1s9BKXaznbA7zZoXc2gM8jVIVhVHp9PxpRIPmnoB1TF8yYnlwkp12hLed0+Iyag
+xnJOOdLB4xDKHk/+RD5BDrGqpqP+vPfVoGKLAuR8xcRqq64IYatumLbC8cPrWcNw4k1Ac27jjy+
Y5/3GYvIFLKiFVAPqeEj/9iZgKuckHHWahHBbXUtG+4cz7VPlJAds9CmBactV/ppNw3F7JuYxIRy
BWYIO2WqxF5xXEhWUmPc1h2WLUjNhOrnqg1qCShWUXqgXOdRWK44D9FfAAAe/z4y1Ibg232srYS3
I/ztpIrZeKVnlka9A/AjHnufUhE9lhCrMe1P2aVZlDjMsnUBGEuZoj6+MEjX3/6K9tpl1bU3Qeb7
2b0CdFtAx6kUklFvNyS7adH2ZJ1Db4upTqMZC8mjdbaDcJ4/1XDLhkc2yENTyvcX6czLK0wZPVsP
okpgXivJJdWXzqESd9BJKG8NwiHW9JqaKaIEG/zC1YfnPT9e4XgYqfUzKwmT9Q6qDPf4vQRN+8kv
aOcBHV3cGesPJvJN9RQ/jSeTU6tWgis4ZS2iMl1zKQN4fv1hrFRees3vVcvlZT+Yl1F0FIC/msad
adXoL4xcp0YxsjXv2vV5nvxwXl6N962nPtfQ6FL3fp0XbIPYDCzsncOV5KyYNtNgGRpCO3doKT1d
xdYwxqpYP7THxK4u0FQHiTwsSMoiXykdHMc5aD5BdJ4VW4Ab37g0ACkpzmOrqrmmDUEgRHwehjpD
hqsnC1SA1cFfE3FKFx/eJgSeeAxHubP6AzXBOGQXJPu33UsHUytuMtvglOOEqNS0KEAzg17cegKf
/Ny+91AM4JIVIFM15G/DQvogb5trII82RlLAAi+l7YAiutlbuPiZPUlT1lwDZl7zLcEjFowRerCT
ZENFDESSsm2qot0O+4QNuOY7mxigq/ffz6NJcPuLAwuYOGlN2OtPUB+/N0VD10fjtPU5Tw13p2ja
QyJC2bOqDdQjFsX8WyqpbRIKdT6Ptk6R3n87IyVaxLynbEuYuzo/usio1t4X/Cc125DPeHtoMq0V
aMvKOYUHN0loIsqy7urZEt8e6nQKAnRg5axnWYQ2lSdpYZGe9S6OCymesi/7Qrsrk6c5WcUn1LTA
Xro0NS1GVP07ca0bID9P3H03HSJc6Xk0LgSk6lllOuRIA/jVqC4uDLdMhNlSjucJMXz1xj3xbDIj
h16kVePxJgI/6YiC5TZ/nW/g393BmboAKIphBXEUM5iWuxMPKABHkB0wnY+CML9Bzml2r94pAHhq
6H/LHHOH4/1fe+meCynpFj/sIVdLDOdU/SFH9hQRQVoQxN5jir+dXXGzfqT693z5u7ZFioOSPZMN
4GUcPEzcbJQ8GtkP8+DKOoUUJxM3Ut9Pj+ivrtce/aaDVijd+JQlMzPlgVYhxkFSqLkeWJv0zNVK
tj9aaN5eOxBEVlqwzE8fxsYkh3ajGqKp+G1Jn4h/BhVaZvy/IvNm1qXcdVYJ/E7ePpEKnELnTzgz
FfyHqE75OlrvJhOjWZqo/FYlttg/hg7XFx/TdrPaCTYuzvcyWQi1bEFevcBk2+7wmMAeOWUcXflZ
NXV52KlGvBunOycIJhb1qfl5FMY/RSTr5TiTcU8LAK8KCIzRkI59FQ8ugsnJ3KkhBcuEv/ehjeHb
gDM5qmOHkH6XHOWj6okmAM5fEMF0BLhO1VIQvU0ggARMb33vODpKXstLlfxvVbsk9glYcwxgcL4F
COdh9rGNqhGiC+/lSA9lCFS0ek4+gZxUcLXL50pMBcZ+rcCASufqHehf3l2MMse72DKVzvuKbWUz
H72rK4bjvnCqS0Z9QgxjCv7gw377yOK+/QbByJjJEyHRSo/Z+WgnFPZRQIPw/c9bdP00EmMIgCkE
5YfOyH4CuJCEztiKXU863HyyFTXy7fh/tkO68Jn4rjiWllYewMLnek7ScJdJe9xI68iZKw2KWPYP
EvrJ8kzx22lX8TZ2P82JG/Tac6ASmReFhyk5nP/AywFtsN3he4FdmhoqQFAkFkoYQciNMYQTd9m5
bFE600mk8ON4I4/mgtKhVw/sVjSy7FzjJN6+lGsU2qUhnkG4CH8mluNQTXj3p0JQyl1Xk5sK0JAg
eC7xknVaSrv0ynbXoqHy9VNdwAySbbNq71qDe9Fh34ka8YqNsiQjS0Y+zBZx8s9AO9tnPtQcs1Rz
fLXUiq3KUkbYvrDc7plpp1lLIV/DWt4IgBMBOgdkPbk7A6SLwBRNip7N8Anj+J1IDs2V263v8zIA
GVpMXazqdjgF8NCpXS+vvZsSixfo9Wd6pUaiuIVB2gsB+YAZv3o94y89YKelJ9Z9l3Q9FhXq+eHj
yGF68mvB0uIFiYd5BYyouRz/p8X53fHeGJ8PTsnZ9F0AhJ0XIYTherTYtMFv6jW2sbfMRGlP+Ym9
hDy0Mp6VHp7iMKxJOqHiPO3rW7DLHoXZIivxt/rxf4893n99p298/CM+ciTfetKsO1bzVIlys5yk
jkuurSaw13H9t8m7OM1YVGZCy7mjX/eYB5osKHHpONvaahbs1W90gmsgNB01vfkhZfStBXukEyeq
WqIZELuhUShfrD0bcxiRX4rtJEHvtOJVIzlFYeEwxvlzr9y4VDj+4bJtE7BiRR7NfvPzS+O2mV7Q
jedteh5oj9VwE35ZmUkDiF+sugwRKwYGmejjb7grdKQGsheBk0yyxGgUwDBMizeexEF3SCMM/Z8C
KF/icZTza9/iXSwgShCq+fHNAGdNmrgbD7Wp7EEa/eylKzyndx7uMWqwHFVkuE2V14DTbNJf7qnU
3TjYiQxM2tzPjfoA+afGk7RObobr/VPwNCFxcUVe1FB3p77+ltWuD/QsYOqMv915OUhEkuMJDE8i
8/qaBtB9t3xawy6tcqVPgsYKoUkbCiCDN1ORVSCafdJXMQEIJNp4qm17sKrMs3cz+DfDnE1at7SA
kW2yumjZ/iYiO2jSrx44Byk41RC82P4Aaz5H83awfteVXCVbN1oFP/prwXsxcpn1wZBvOiQiAVD9
Z6zWhPmMavkkzJyNuZfc2AAYkhPTF9eXlzuiljXF5VfT4m3mFdfd9MRbjfQVvIRAiibG9uOybtXj
NMsNMiS8f5a/n+pytmAPzLEFa+JarRUL5UUwEEL0s5OgZDpgWqiGwzV6ppUJWaR78CSBpUPspM/A
f4MxfJzu4OGeP6YPf6xlUKv+lGD+jKLyhxqfu+TMAJUBrrMTg8XeK1ZUHkp3FnWGB/ZneyIPPkMe
kLSu5Bi3xEw/ZxtUySyUogQWWRjMULF24Q0iB1un129c/TX91lB+3fFuCekSrMMPxglxLkTxnqBy
hUaINwlhwUEk/dakw2ghATrUdemEgBnwxvOstQ1iexXqseuY1z7+jmmOBu6iyY6cAJXuJq8m8hu8
w+oPEE7eW40+fadzHoBKs1gtvCabqGL/+SbSldPhUmuX+JAuiHwA6gKI1Z3U/6ydk0WcpdRQQDGB
ySNrwq1+5qM3VYD/9ETQjwV6YXVXPuscj7mv7PAoMgiEKoC5f2LEAsVNP6J3nlINpoC3YMPOI15P
dRoWAlFoD8hMz3TpWf9PeIwHhl3QGnwjtfT9Mf5UFIGNE8mH/5xWZUm1awf6d7G3M4yNmx7CykuI
M/xc0ZXcBOEo4g5+5mWg2uyqzzjPqCqHzkW8wZNa5oKn/KmVTSA7VtBM0HuqtjcfuGJWIoONSVv/
kpAwYX+m5r8ln7/RK+rHj7bIMnGgpgs9MDd+aouOKRec7byJ9OUmX3YYSsindyut5l3YlbWzkOeP
+8hs1rNN21OWn3YPOm5MWjQ4fKF0pcjP2f6wFfbAXtGhP7Hgo62n89VklOqUVdrpUx2F3z62Lpg6
DnqNY28oZuqHD1YCpXZCPACUnJMQCmcmBmTl0S7Zvsp8/lB8LRiZPqwZF5Lshys1j34UNGn4x8QB
fhCqBkZdJYVj7i1MTnwj72CeOTaIjgczzlEofQUOmzkmaS0wo2Fvmy5XBZRi+Lw6Nxx/W+f6HYcB
f6mnBKv+txRh9J7yAXh8FK/42UI7pbe7Ze7FwAT4SVY8y0k+k2UQ5gssB8uS8g/Ov1ju6pw6ZBwa
LX2/Y0Cl1pAFoKXKc5OKWtZCee9bsYpx6BJHFVtNmfLx9SKfCxtt4xJhk06ZNsOlhxtCyZrXoHb8
T40U6q9T5ovun0S70lcaPNjC0RtwfIH9l4SSqHE7fj15f/1+0Xf0SOOtPDnk7QNO8j5FfCAPEOOu
9VJAXdWWkSoDw/g4TPiDYZZCye+TKHk0M5z0juxtYG8utuC68GIe5O2M0e/00rVV5saxO1tmkWfV
ALmjDzj8REhNmuT3jRRQI4LbZtSxNOjp8q3OjEzavc0iL/Rz60ZM830aEGVDw1tyeHHsvS2DC95I
SKNmyHtjdm2uN/6QPqHpWnJIjJnnCGIbvZ00gqfVZGBUSkO5qMHUOAkdi4tGWrxcKj/Ms27jQUDZ
5eOWym5/rJQl3KIh7vRtcOUZTBaeh2z8gqlefC3ig3ztFiYfLAGk2gYUb4iOXDt8pnoCJFS3im4T
fhLEz8EG0cWlkPv8tehI0aagOxkZwt9o3YVloYuWm0SiNVcs5cETH2tLH8P87wfbCL16ce6yvyU1
yiynV/wy+r0zjVgRMJwdWyHh9g7cAbFvXKtUw2aG4PLJFaHrMepEdsXpQ5kwOIIeQ54hU0IdUGp2
dVbPcO9rVtXpix3Q6HL3FdeXOkPYb/hycU0VXKilD/dH4ODeDoIREmzuwvFpzHlpalkjd4Lqws5i
61HPlDaQsR3qRf6P5PxUCWJsW3xrki8dEKgsspVkiRcITx5daUQ5u0LFMoJNAZ36ZD5T8wo25SSq
lwRPEpUIeDMYUaSburqeDB8/aq3UkKUu/Oy+psdM1zAaqiyvWv28xUb4Ekc6S1vjrr094URII7EL
ERfCgqtwm6GrawlnBsJUHhYg6isOg0Rm8U3Wiq0gneYbc9RQRLisksmzOozdmiE+TvvwpFodu54i
f1WKWj3vTmoQVMIOmMHARosjyqv1/PNnQYOxQyblaTmK4Is7jI9PViWuFUCui6t2r9Xv073LL1K2
NdC7DzC3XaJQFQjagzHA8dKFS8plZrS7cUKbduyC42teghCqJK8hDEL20SoghDrXJWh1HXq30HCd
1OkNA53flCe5xsIGGSFeC/hD/GDP6YolpLNea5en0zKVTEtlQjrU5uAXV9tLfszKYamW5FDpLvII
NL9dNjZO9NKMxm3SszjYnti5xTzFw04+AqYEUy3/+Nlk46teEQRoqYX8EcjzMrGqOwgo1G6LKUzQ
5pUo0HeHLIg1nAnWH3blzt3IkFLCir3tC2xRsQjtG02jGGZ3rhXYLgaLyng78va2Wc5OLgql3/ro
9LUfYddNVjZo/E7+Ib4J5AHxRgKUjqH+kgMY0ta7gpwMpPAtX4UfCjpTi565shs37AFvrpxofbZV
5T1fBhdT6BfRdjSO4fh64E17eITb3BG4MgQoJYvWK0NvQD2UcQYOVLFxeXL962Xuf3NgxOIfftT6
N0eWbvvL/iiOExgUz0RcMgPnHw+833607WJMuH1UP550pJzNfrhJaqoAbhHB5CoKLe3/k6wN0FCy
YXgi2fdXNg1mLPZxOLa4vk4jtv8ktuRDvRyM+QjtohbJB0x3ZxcvTNjmiA9hFHhri+8VhkbKZ3FT
GNTY9lkncz/79bUI2BrqbzgsDnxQvHZsaeS0w5KHeq5v1Inqb3eblyPNpfZHvnadWhFKgj/sdjdA
anJCjHI3owl0ZbieFope4umzn6OJqix/EdoZeDrsqe1fHUR502XmNDUA28DZ27e0kI9Xd/X0BteT
DNpxeBEJ+xgY3m2eB0N8l+FdeAOX9xY0wXmGiuPupqFucEjqhVH/Q7Yyi/Tq8bd6++KA9giByHOu
GK5q/tZh9HNkzWXn69r7BT+2/YSsh38NrgrgJppGUCaWOis5mB6ie1eZ/5NiKo6/LFLItdRtCw/3
9mkkWZt13F0Tbqsw028nLToNaBwgTxsdXBlRBa2HDjcxpRp83ij2VXFhe2mkybNpCWUxVUqOVzmy
y9w133T0jPtOQhOjeBeirlcxALGtsFUgdnTQb5RZox7w/zXzUJwiUfPunlJL91dydbWM6j4BpJ/e
mMK1O1fMrvCQyTMj+KUNZZ7yprZmjqC4/l4HZxuuzFQCRaOJtX7zv1Gdo+hMWqBXnck7Yla5IChc
ArXCB/IxqfdEWIiI3q86pfHSW14HQyTqQtM2p7WRZiEpuhzq6DCil2HFh/M2Gi5jdCp25SPRo/1j
/Kyi2xKQlVQn9UwQ6R94xQg5h/lQivrrEwKQKDuRKQUTmGpv1tY9goNXAa2Sq2ezdNKfe5cjYTJa
EFnmHJG5vJ0vsg/j05xkmhlxSegtbe++lSPG7+18MP2Uo7QfJMer5HmqTnEZOtZSn77o4jii8db4
BgyJFvcxeqxYd8mCtcme+c8VjuBrc5++oXOhc4Ng83rK+Q+ojyRTZkbjQTjFhs4ecOtFf2TlowJN
hnuY3OKzQ881wbUsftCNBNwk+9+zFN1b+jmqX9k+OCSqNvj8CzWnUCeC+Y97GCf3I2VZrSl/l8MU
0bUjqGyon2WhyPm/ttrD08XtLe1KhoxbnJ4yxCeghBw/cU0OW1kpESke5QdbdiueinO14uG+ul+p
V7ePRfF8ZFbpz27wHrZllnBQMyBMfBtxfVz1NuwqZhV5GLtu/0QjzBnhhX+n1BazHHG70rsrVXIq
dk6orXGZdStiWT19QG36TvHIyWRjSbqFRMfTmXaXdiTgc8GvcBFJd4rFanE4WlZbeL6b4sPX7s9R
AvMxBpPZBTtBYKN60xOw2KdPVibs9ZiYbDWUZBgiOYfpnwctn7cZQU24Dsqg6MQyb7Mso9n5SP3S
W4P5jmzxOCVtfKtrfn2WC77HE/mizdsb6yv+iWnK2izMS2P3GS32mN9VobMRmQ5E6yX5YeOANNVK
VEzry0mQbLqRas7xxNTmtBtVYC7eo8x6HaTMwlXKncMxEgUAF1xkbiTXc6oew4bBPmigjTZ7ew9j
Ikv9n8D2kAXKUl8G5AaGfpMbOkGewaGgvuYBz14qaiDUBGBgiephHYalIzBatzp2VdPcufvl9l1k
spfEfBmEa0TldK7HzokuC6ASyxgfx82oF9WZj8ouK7fV4M+9DlnVX42EW+/ogcGPx7Ch4oFsXEpQ
bYrguAqoE9f6m2ocrtilF/q5/yZ0xeBsuFKAv6AiAnmV7Gy4Z5hec9x0W0AQH0RyegtZ1tXrT1zs
1y+nciOu7qOXrNd2v9WpLVtIqDqKAVtrUSJoEYJkpMSRXjctzqmjbFgUzaojNgR9g9Qwj2MKJg4p
C650lkHJVs4NMeXnQ6DmVCQhPx5M9ikvUVFokgTad3EhGgoMRCZeCeS7dnZqNEsfbY1Trl8jW7kA
6kUdy5iWlciqyS+E9CML7U7cX98uKLrrp0FaRrovLmrStbJ0l4xCf3KRhPFp7qHfvlPqv+c4YQAe
s1p4ik5Ddxe/2AO/7inNd6RtnaAZiqVKVV46yLlMVWFvNH/miljyp6Wh/DgCLLVCSoDqGNR10M3J
kWe3bd5Jz8L8oUbfgetD3CRyTRZGLJ92oxLsBtYdP8teyjV4N5/nCMIvYHVO2FGbFB+NHyGkrTZO
2QYv46Vcvvv0EkSRukPvcq+x3N7IriyeLq+3JAocukxQB6+SI70c0FAzJdcWGHuc3T2aNMaDta0x
807dKNLqByxe5u4NYp7XXx+fV+KRocKNeEicA6SCC2C6ff6Hrk1YyBrSS2vMkAeht1V5FoPgDLWP
q/r+0SYxFQZXXFy9VuJDNQ/gjHiZerFUMthKt/Q0Qb4OjDi033idKLS7DaLvX7LWKR+sLLyv8Qm/
KqSqQ2pjZ82VS80/pUydB2nvflPlaliKQ8P61Qf+fEbPYdv5+LCyc7tp0/qM23qbX0FDPtA5OSCF
4aRHEbpO98Fqp7ilA/ewSTA8d7oD9ME+W4/IOKrX0jh6/tfCoSEWuP3LBy/HsGcFScrjuqk+iInM
my1dxdg32yUDHv6i0G29OuItmxHetxupIAO1snS5MrcwPKM9d/u8Xwl+cFT1hJNS0e0Ka6xxAwcS
yNSET00qt0kSxNkskLh4vSyMXjhAxOl24IHOQRh+CJdyQZKdjzxrHNtdj7jSYljYd+oUtoCN9l18
qNcokyaO26JQaujdJ/khQP5sFE70A3NMjKxkrdw+Hpd5KI5cYa4xpiP/joctTfEk0bGVlM/hLeU7
IHEpwwOmNUZXGYUEkJBeEbSv8peyFoxezjgNMmZHWrBQvanYt/ZLA3+d+PN0j78aBhaPiVogRUJo
UrPuSyIP3+IqmUd2yjRFqhrXfk9SDitpwbp06tBOzsff+fnKdBtsRqxMUWX+jQkR2hpCfedhtXVb
Q6Lb2SGQqDuFcWDm/FytprNXjUaMewLVMYq1ZcSbd0vxGXMtx59ReuDCIWdfCadnBfHUR+1l+0LC
EZcwYam/6Z5lbmC8O6aZWmhnP4KPjJ7QTFTWL/GOkIZdjH8XoN+Zt2lHdqQ0J13moumCd5j0sJ1L
gmJQXyQAZXnYuDTZpSMnXRBKqUamYZJm+APDmcDgp/TDjW3y54+EjuK1qrOjCVw47wwEQOeGl6Oo
5xZrQ0YfryusGgdhz+sgLdcLEZWcgPpgx4IgArV4WS+rrK3t3tIycbf48E5tVP1v8nAwhhuy7S/c
wGTmlGWJZTOY+RRx8mzx1dOBJLTYPnQawUbtNlHwIgoEfLTAQ/ouX37D6RSK02hyLsPM+1b1D+JT
+NsXRp48quk7MsA0agPbI/C6kxnMosjnRrSejIDiprDXNfmWeEmPvXTaXM4k7y6MTKSWPy9Bsusl
R2ASeL3wzPfR0USPTOqZL0mAciEvM5q25DTFxDA31PIz0Q+X9iMlbT6qmnndAEKdL5Cjx4w2InXI
5DoEV8kGYVYFs5222eZb6PZ9XEl5fivvQDuxtBO8nMS3Y+t4bZ+9JIGENfPIqOyNnJuZiO+ON6Lr
y8Pj7EqQ5x9K5FNQMR0h8f4prV0sGjnwxpZ0JSjwz6kfAZhtV7VYPWTNwxw5iOseBqQOLJRabgjC
uHruwEcRO7wkaPMQTcmcBLk6Ji0Y8ZX/I3xaToPeZVictST3h4+1066fbfpMiGx3eKEbT8IG8Kt5
cfZt+TA0HKyN2FYzAeMbx/IDJ6mct46kPtedOBl7QAimyNSS3lsdxfYWTUn/cissyLeGG2akV7go
dMIY5W0fLKQKJdTIyqF0zMEO5rQcHW72bH5qHxffTKsJ6wCwJNYjVML5+K685XjbAwbMJXFCKt5s
EvZwqfUsblI2oY+HwacrzYRjFY3jyeFnzN3lHT7qpFZuGcaNw9YDRZ3N1qtshxxJpz4oEZSgCjpw
4ETVc0NNmkId76Vn3BxcGWK/xsmuwaaPSIH+7QfyKGwPkTpppAqrPiVNdDu+4fMqypHeBhL7ukC2
+TcWhjc1eM/OxLR/j/lSlNVR7tiWRzD9QNf9GFkzFCi9aa8Qqf00BVlTT7WOKakwY5DGBqxNaUae
SGHPhJMnAyWhqwKFHCHPPYty5ONkdoiiNjnntIEMKUKzS5fMwJZwpRNXuxG7deShjikzEZJK+cKZ
FP8m+/c0H0N1MY+3fOL1XXbkB6noroz9ADnT0oa50lDLYTSt6VjhRw6yQYiNag7K3khafaq0pBSO
A1nIUdR7oGETrmYFXZ+HFZEGc+xYB3/tcr4+4c7lMxkDfPMjbLFGI7LubC/9h9AvUMmsj4GNT6ws
bx3Fsw1W/g2u8CdjnnIh3/Agh72ry07B6cGtJ7hDw7F0hgsF2xGyRpAvb1Hajbk2M4zga0dvthjz
akD5imkHWwSvJ+/mzOEAMebkMa1tAG+kIGnWwWBMStOiXU5asj4gbmq8lOAZ2v30Utqj3npc4lhI
967O2eZsXte2nTpAyLFUld7/vk7f6/rIeABI89x8pazfCsmTSdesG+M9i9/Q3NhmUAahRE+eSO8c
Hb0G1Jd5lt75Us9ffMRmElIaAESgUyPEpinVugiBcTvmJqCljZc7hjeCwafkvN4pj6JLsyylnlSj
/t8Cb0ggM4ELBh52yQuWUbJaqfz9tGjxaVLUB1rHwr60O9Y474pI2mwSQVEjXZgnrV1bkrO9BMbm
OxIFcbaVI3j9Tpa/s+alzxtOTynWN+2u1BH6cryNW+F1FelBEGJtFLXVN51VL7ki5DQKTaT+i0M2
xeZHt/tGAu+THFytX6jczXH0sjJDecfSawHeKCz75rERGKGcOl1H2Zqd9cnVRny5M1j5gAo7i2y3
//wY0wx2nZ5GHxdKiXwMTV0nPw+Pyc27yNKCRaM3+298trsxO5EeQBrJyerIG7Qkedopmd8eO1DJ
wpc2g5Z+gvSkQBJLcQ86RD7ki9d1ZJdeX/nzN+5O82kGkABIsEXHO8pHs5tCv6kFRyUSBAFfzb+F
hUku/TuBBlJXlEgyo+231URnX/YTCK9HsPx5Io/Y1WsOHP9HADeG0qxvRWrp+mnHXoCAriyXjry3
KEyoQYpF2ssBltt9mOCyCsUkwwlcI3Rx2D30XXkZTg3+HDgGwtmOGYfjrm1BP1goOL9YsMZPYjsf
MU8sqDAMxI/OwKgQKlur9shkEAJMItC6pDfX+y62M4dl7adI6QgGVrkOoQa75fxGLLQ2lbaoY4mg
VBf4j9c4ohuLR4p5BAxXWj4MEnLKObeDpN3C0dkq0cTxMHULN9O5HVaCy4Ye3SWaSJZsvz1f1xlX
Mf8cdUlQTvKjpv5XXaYuZ+Q0E4Zfa3dOPBe560BGoBBCKVm/lVQWI53SjPgvSCkTnEfvOQ6+YWNz
XuNPgruBvVCeItoRhoudM1Zz4eJB2felwKB1pQY/KnTb94Sdje0EZr+f7v44E0vQZxcvc1mkfABK
o/aqkYLVDWVrOIf6gxIF5eGHMNgqcO3led53kCP5WGfAz/DzBVpaaIGJIGRzE5/c5tExYW7MkDgk
6UDvb5YjHRuHupDeDbKUyw+50OrS44hTE3gkgb+4SDOxiR1ZFmtlSPrhZhQcIPDyyU28P6QS71SQ
awo15b6AxDTbP7oXsjd45tr8jnQJHv2c9cUotichxRtabISzFLh99EyFLvAkKasN0Tkt13GFSjHv
1zQfj7Itv6Fy8aj/sqaoD0BepSPHA0Cq1fmpR5cNDq9J2CvZul0yV1dX/p1k4xfKIDB8xqzDAZIx
qY7eaPBqdAtIUQRXIyNPUWHtipFkfABVfEU60SJw1vKjWuTffJDDvgekTcoLnS1AnDP4dxXMqOdL
g6XXlYU960GRsHjVK3nHnPMvDj4TRRVhPkgEGGGq84n39aNbF/QFu2Gq+8h7O8mSy/E1eKQfQMsf
XjNkhFP7EXKZXn63PbGJF5+o5ueezVdz9tZZZfpbiqGKUL4bkwxE6j1cFTw6/SAOg373VxO2l08x
AN9fLrGcEp/m+ej6jr0amfvME4KfqR7SH7YpgfvF5shtU/BCx0bUKxw/f8reXpAuRuV5zhkNTY/E
ZZJAc0Awe4eWztMT6QSQd/vA0tR5dEmWESl+lvJRhG4InD2D19Qg0eiEUhdAq4tLlZGrwdclwl3v
6sq9d5HKubgxm/MJKmfNzcM6CavKMS9kSJg3nlqO+KNxyR+dvCy9dNQr7ZgLGt3pOuCuMRmfdQTK
klteNeKpJW+tBO+Xa45FRky3IiEcPQ5FQsuhqaPQrWgVr7906pZ6wlF9E0fvfh60w++9z8y4wpLt
MXF5zo4rtl0PsqcXsf2zjS1Xro178cN3VZ0z+Nproser3LVi2opx1wnm7fYQWLAxHGrdSj6s/rQi
sVyCATABxt9bZA9XlqOEygkoV2gKTz0lidyyZRUJ+DZHkdhSJ95oD+UpgqTYJcPFgiTIo0jGakuY
90ITOytTLhh5T1BN9uQRztKY1a6kXfpD3+YtgNLjd5hzqpznRpDRVP6kvtvF+PV6juwwMUSQf6G7
e/d9ApMOGeUByqzQBR7rTGojSJSTMcxD+oSErAJgUSfKYq9u+REgDpUAM1k8xBEa7JZ6wpkvcEMO
sl/95C/LETfaCdvflUb/gpfelhlXh/W6yPrF+EXrH3/dlaMUZjabvacNfgZffjj28PMJIjsHPYXl
lKyYxyzoo7fnX/tbSwl4DcGmKcPHCHNB/K+BktKgUZ5YMag1Hjl1rn0tTsN+ba25dg+WXk7aAfSX
ZNpdtDBj2wKtpQ+y9cGRDiBDNNno7MsKT5KABt+R8Q9LBu4lNFyys91fBaezbvxh+ZdBpMXhpL+3
R+ehRT5S42TcXDX/r7ziFyFlE9WAb9rOmlM9YDzZ/UTkrel2w4/KRagkhrHqlTW/2MKrzkV1aRj8
6fSsyvhyh8kHGVbs0OtK4GJ00Dwa8kJiBmg8xw0k5xIINgsW2bHYunrlumYpG8XliLAc+foc/ppF
h20ZSbGrRVLGPkwpJ9ojxqa/eS6z6VNeDW79WLYb1vL904FX5EIzE/nqhTEQ5+n312/R0k4DzhSp
UUfFHC+RoxMaAOZn6MiEV2NqG5JgdmmfqjXu8o3X+l+tVhBHshbdylOtUDo+vKuYNxUtbhJacj0q
D6HK5yjAsvhhHNjYZPnXK/jzHUXT9o0STIQgOtq0yPnDsqQVdJjykpv6wkY2xoKAuDwyUxjztQvK
7xA9r/lxhPReWPc8CGZuhpvas/kXmCMVEV37o+5+DQ2ut8xuNNPxAkpZr3lt/MLW6WZJkmSMaFq4
E6GZJZ7N6YrWmCfPvAmCNKOCePPo1M3/mfOuh+Fu0lwvOWUhcGduTrGQHB89e+2NSu0mQ+sVxIWT
qPvXqb1Z/tp4P/MA2qmkb92C8Go2GrXpNUCU6NkxSgnA2NwJuq7++a0op1fJ9B/sAowwABJuC4o9
jVbiyECzMqop5B9RQC16rgLVbFAdsTJwpfD05I2/0qb6K+qASqkaDyn51J2I6CmPyjXw0Gl6sC02
kBGGr7f7B3A7lmmUnXmYxQpXlPEDGbmhKHc8+lYUfvuY08CDhBBA24Ltf70l44Odp1p7wadWaxPd
a3gpWFcTMyKqPsDjkS2EzqlnxuupH1ABCy418h7x/4vnlMypGpDwBQHcV0kEiwdFgVXS9yJdcbQd
QPSvTsnEdlsLnv/PhvGQNuYyALHrcBmi3LpmPp7Hdwiit+tMbVLfoWp5MR97ebefJ8UeaZA6JqGQ
vgdGLvgsDoOLhQIhykFlg3VNuQV/6vO6ziiF7DBd/xc2qjWARRl5B/D400lw5YpwpyhOdcp9KV96
x5JyZ9GxvKJccBxH6YJbszOrkr5nWtKAv3zR3e/RkhSQowOjGEco9WPv3X1n37uTjAUYpk8omad/
GvNn4ovtBqcHhq1+BS4c0Q/0ixZIbLTR6+XFvxiwswRHTPnlTAdvqE8mZGuS40/YmWHJVLyexiw5
J/G/abYsjMEmyMWpPD+Ifnn19xsxn6Sv1sA1J1NGlAeYEyPU/FeCbW7PSWsm1RIu3dGpgqbSE2fI
yJFKhkzS6GO6uYaa5m8Lc+iTEV6PYCYhX+Z+LGaBHfnygxwE5giUjgPQQnQh9Dcc5slFDbb1p40s
qvgqx25QoY3o3k3LF3WjvEKAZV19NrU18PPQfDlvq+VU//RGvLKWOQdN7CVWiEQzPSuATM/bagUA
JGfSPUo0gI83mY71U4b8lfES5+43wD2otmWKjSX9Tg33gSKjbhF6ukgk6OepOjQSftj8be8G899y
KPHvjzyv/SCOAfML8Re1x5bf6PAFllNbfHp4CGD7u3xIyfFucAb9R+178/1eXry5Op+Y/GCDfAzw
NZoPJYA3uBGQicM5i/RRaGpTgxqGZ3+f9SiVDuYYhByzrtfr52UDD2999dNpfg9d2pygXPDOnbue
GulLkNL7FERDQQ03uk5dsm+u9l8RR5TSl/vjguU3lTqxFvlK93Lav62ne9ycmJ0FMnmTrYL+rpIc
qmOd1NGMu8tdOxtZTbJC+4rJQ4n+l+g7ct3DdQX334zeRUkmfAsQbcELcKg2gRlI+8qb+qhMwRx5
i0yZzu08XHaeYIOkVMUQBpsdNOtFrXT0+ovj1MQSE8QKKJZvuXX7HTiJD3ORb7pJwOYPradhn/EK
3tYgixv+6G7ANDbizqhvg7B2kXeoI0+TbQwjJZ7z4bV/oFf+OAP25PCFD6/Rxf4iWyym+O2yv0s8
ATqA4VGgSqDHdFFw/vQIE0AIyigAXCDfn1IlIaqAFHEck1+tKE26ZItGRXNsl/j4COqWpxtcfFIF
kUCg9HQGfF/ta7GL1N9P363XYOUv32139LxNJeJF5e2BOPiQnXVq0zp8NbKXl7lmuX41+NEevwd9
wkKVF0UP5Vet0PJPCmzKvLPwPCK+/WrsSzwu+OK0zHx0dibERajjPbq9cYIdSPMm3gjx3X/OmdB3
sO+FzH+yHgSIUGfoEKU1LhttJKaPIvt/I1LTrx5KwXXxDc0Zpo+hqp3SuyCrSM6eSEk9yH+ELDIU
6642gXrAft+s2lkbACdzYrTpITS7e3SxzqhkxOP4Wy/aTEy/9HkefvSgofywTFjqsasm3SpMNk/j
itCx/KUkGn9JrVQBhMkmr0dMDnM0063waoE7lrywOAIZ43nIyVz72Nb/XUgGbH07NTTzawSJ0Vts
IlEARurtOhk/BK2Ms+tUvViy/hHkldEtYsEXgVB3TQDBQQsMGGBEe6lt0twS06bWC6ORbaYzItfZ
W2wFZZEuh6j5tETc2Giu9pOknvXqvSJg4zdZt4E5qPCUbmu3u2jb798UROaIFgvzjDzh7sxCOyVR
FED5LPw6axZOGVp44CY/XxGxWJ3xupc4owj8GzCyMndNMyAA4y6IYqLhHv1Cz42k1TdODhb2Bat4
UTUeddW4/m2xAPYrss623Rj/uASd+r7I6FtxDyMJp0qkQ4+DofWcJDUK+PMKA3I+X9JJex+ynEah
1H/gaov380cZHQCeYzfKr6jwOC1xlQna7jYiYu/f9cYqx69wbsFHnhN+QnwTtGKRVJFQaXRQRu1c
gV1fcBgcI2V1knsIwy3WsA1fW77D7/mZt96/T1qoy8we2xuW6WA2I15CIXkqInuIF5YSJ/mj04t4
rMk5LoMIs+p5umzqeJCsj/q07fU8+YAlHEgadg6OsYpio/5wYBUgG3k8NGbQlolvdRHywh2V5Rp4
Mqc+fIkzdmjKFdooxr543kzoD246lCtF7vIIBeaxzR+7gGcfa5n7SnAYnty9RLQZGH0Ty4k3qlWK
nZov+9IaqyooPonYY/mi/1aQ4yGd4HvbTFJGG5LOe1NEVvVqcc+edNdlZG+galrHowsuGyXgCUY3
jtSOTeHFfY4C4PoCH//Dt6MD7i7clvrXHptKCZjCn4L9Ac+Kw2O3+FI+Ky/GHZoNn8TNxOPNo0cM
61MzkRa94qsbInDoxvMwSJV7HVsRmakKkoaAoF9VYDKkcPvxDLTQqQtV7Bi02oUsD5RdFi2KoyCf
/bBZ0xFZ8zKP549WVwlFRl7ByEhRSeBZGseK5/h3YxL0TvRmlogjT+kJ/DE3QFotXQapOq+WvIVb
42QBDWlMwxCechVv+FZLDYj3IvelEwXj5h8bgrR32z9XaitIbpDqZWmVpRcfQKo9vMtPYLWUW4ca
0CTG93nUZxyuX+aTAwebrmRHysrvEXZJolla2W8RfVsrcYgtPCXyDM3YdbgwCDofy0gDFnTkfnGf
iUscZQgLUOwrHN5+5ig6klWv0HqriNHvecg2UV29NvklDJjlugzq3klEi5R18qSUlEKS7xD59XdI
DevnyCTeBNXWFmVVQl3xoN8RrPm9txRVGqwoWUB8j0vmsuC9AoMh/vnDAwAN4TPM2OnPOb91hMci
p8e8/erhFbjwq9od2iLv7MbUxOdMHjDDSCR0geII+A+1g7tiJrU8OHsEaXAJy/hWBU4zVGMu89P9
f9Ux/EkEmv7LcQUNOT08YbrvwpneoZpppYHmtov6mlNFotAnLA8yuOnQDrwst0yCPCsimig4yQQR
eHCHGOVjfWps2GUXoG3ufQJ1Y4rq5jMez7BTqjG0lh89mUCiHWi55itwMENfWAtu63Keg5JIwmaX
xbGw2j7z8sa7Cy4+8g3vMfK73q06G/Qd/5jWZ6d8dCMEl+V4oql3ZFwoEiChv8TdZ7aNEY0Sh9qy
HyF6yVx8vnS3oYIcmiVfFcmQKZOqfpZKsj97X39EXtxtBkEnI8tMW4TjZFSMfd8POnsJE+B6UDc2
STlCWNwzn16grxQvc0clZq2bffCPtru3kMSeNcbISEJw/D70XlreRxAY5NQuDnfX6WOMZNuTo1XU
XaGkI9mdp4iGNjbvZo4Js/AlTN12mlldjLY0OTPFqZSsVy25AkrKwCkH5mjODG5Rzg22WninDtOX
BY3ZbHuiwkiVsN9uSmLWzMFWsdObdCt2YP04HhlPZpIKylwg3Z8KQpzr5Nv73u/oniAfMlV8ox4j
yaO0DL2qmv4b1zP7m7RvrjQUORe2VQvEMfTQkCVzfw9QNtP7p8Uvq56C0EBWLef62vL0np03fhlz
XED5UDBHicjvVrieI2DYwxiujf7e47oIbTcqmBJLlVOxiMDGV5b2aDDGVVpa+EOJbJJdmovxA4CV
WO4VRHIZ5Z42OxP2nNYUS9WEs1Lya3qdEssuO5gWYwS1L0VByZLRTZ6+SmE3tHj9+w1EWQPsCyj1
aHrbo9fBBs+FOXvQcNB/ETR46cRF9I7/fdNdB81dNF1IH/9JPE8FSdlAmdR5vZwtiyuzahs86UzC
TwKYh/k/Z3TGbjBXEdhSo9ru4GCnrD0fwEa/kRGXexBgTHe0A9TJ2xai9dTzAzYEgbh+wJdvfVS1
tgBKYuscCSpiuN1m28HtyRgW3Ctmzf8yCUXJTa1/e7p3/qAX/dOdcJd15MDEdaHlkZXFiP8AGooz
Jp6amOOQf6O00QAKzGbJ1J5/DCwSwzzXwmhR5w6HMGHuo8omzm/kx6aCml3khggZ4Oc9K3Otauk9
e0mrd1NT7pVkYMDFqRrDuMcOYRkuXS4t0GN2g7fnYF3n9/w7sPbCayhR0E24emZx5/zCfwFhEMne
DIbSOBWlqKR5R6Y180aNcC+j2GVWz3BWLhvdtEdIy1HAY1wJL9sYwcwre5Bld+AcSzohF1j/lsza
RKMdk0oX7yATV5BGWeh1vS9YOdJKKTv9c+0Z6yGLB2/0p74fNQr9cvSWPDKX9W8H27C/ZFfFTNG5
YNLL4hLoiUqeDLuJkteXp4JDScYOM8T8CbeSeRp0+YUQo0zoORze2q17Dk5TWOET8Qq3sqIoC//3
gjPwFcLBOJdFsVsIAYCpPKruRCYSlpUl4jg+J6NhP7ZF1Uga6KJEYNHa9FM2hHYrXarVBT5fbpxN
nlfM4AMTcoLe7lgNBhyO2AQkO+w7Cmu9PDD0X7gnv9sPkqGPOSx7ywWqNOq8Urqt7i6gU32EODjz
NCxqbMZnXKIv/ILi5c/oLUgZJI1KHf73vYtpaCj4CT1lXVXd/BzuIvf/NbFHXY94rgMwQLHxFmJA
wujDrNRMfL0s90wWenzxsDubGgPd4UlEvLsSiQJ+2107RENYxwcy8zt+16fJqLpGP7dXPOtpTSp0
2b8VIVqpHDbS/LQgaDYVPOtwt7BD5aibT+9UhacqiTgZoiwlWARE8WQ4aBTt4i5RrMnnzsYQ0QHQ
ejRZRj3kOw/SayisLIbkbJBw6mbsBaFJPL+rgRZb8pZ1M+KQmCgh5IOz5/fXPklKevgJjl/zwPkq
rsSif91hDnjEna22Ll/cmVdULLvutYanX/CjSASSNVVZoHfFyXgzhcFaOEb12Nwagm+oB7Pce/ZA
vvUqVDyin3Dpoiid8qLEEqIlfB1WDNpZaeBiPGIqUBobS4JSzd/8+9R1RHKeXasEoPI+0IR47Viw
uCfi7a6S2guwNKrMakx3VI3SXLAuGocB/rRH9pVzuPIBQKU8d0YsHTkJq8NzGkGRcCitJZyp2eP1
PzOnZqCATStSgw54cnWAiKxEUNBYlziS+54UZ/Mvc20rJAFFZiJfVeLgxeVmgZW1w0COMb/hcPlk
Urt81RKklsuZSQpTMNjUzf4TdfCdGI7vbVv/2dvADLKv5COXBInEX9UXvb4E3Id43QfOuHITMJ2i
1CO4SjhBFeCc6dvGgKuxO3FTnJvr+t1oPDqziW0a76CdJ4RfQy+lfTfXzV6txxLYo45UQBYgNnlO
azEPg8BveCdmah3Wh2FPxTNOYMxBBBrTFp2FtV1/BQ4d6rss5vAbl+5X97lKypb/0gOW5j5uDCbk
oAQabHPxeU1hf4wYsrYEIHN/nzpz2diqI+DWPm2zhnX6IFqaL2HmYfR9J9EIErt2Qk9cJq2cX8QC
T7Q2X4iHJdBS9RbbP7Iz64R6Dl5Z7OXi1CvZoADZR8+EdP6yCGbPCMa2lTB4NbOiQ1EcFuRhs933
xDCFmzTXXXm21qkcYLOYKisAwAvLzQVt8Y7bS+w3CXxZb6C2ewjbplnqIiRSX2jtWyjIoM8kHcq9
+BQKQfrtruYKXEpAuFEZrKuDLRAs4DKz4u+mq9V0uVOAF6Gn7ybeVVlAIdmGiz2jcfp91nPFfn23
NkK+3AwdS7UwiQIOdzPLwro1gwhivSnlFlcfuUIrQ87eIh97sI0wAZ7+J0maU9Ul8vdPZkeQQ7ps
57OlZFZ5hch2I1ATYyfZQ6JLYiEEZY5ajsRylkwYWdJB4PaFY6+snDla3VvJu2ra1wgZtakU7MDm
JyxaeaCOun+or/Nwlb/RR9781GgAiQuegY1W1IjS/Gq2uINJmHWRlfLHHO5xDboQ5J79tvh2PqV2
J8O0B4wqIgYSp0kpbER4XjFvON0jZx0LTlA2en77jtjLvW7UkCHsgpnwqkSAKhYoktU1r2vl7xTj
aklzfQTJfDr6cWOATsgi/MIPfUmmTAssnUsBCwMQXT3PPh0a9hqgDB2LFQPSwWFRo9IGFTAyRPki
96HMxi+ymGnrMWo05EJ5LpD3e8lA98RrxbizhOZm0opMKTZx2vqNgA+/EnOzxeOBW+VLduXE53Jx
ycNo20WGqgDVKInoH6jlCNBDYJEueVx7Nge1qc5+gDYrS/Khpfr4DD3mU0bMoeH8++soCv+n4IPX
6UdmSu++CMFVtK0JKcTPqKhUKGpLa5+U1/USJLFvIqEdDjxAqUih/iKKw/TPN6N8hqxwisckmfAV
pIi/bfvDniyGhUPMLUtteLejyyVaie/20fh3OYvO5yRVqDaXt/F3NupjycWkuTY5Pyu+ShIFCiJJ
tv4kB6sjioJW0ZnXs72YykPIVB2h2afT94APEfXvvB60CCd76Ess23Z7v1IldxflRw5CtvdQiYVd
gNFbt+HQF7yjNr43yzbibQqYq9wwwrcMsHxr8TpklwlYSAr7yHsGwy4PjwjUCZjlH6mgWhzhkjWK
1xP0BHnZ02oY7F8rgX7z6AOU4y1cKSHAdNp1SDLhAM+mBERKChoW4BbDRZBKZyxE+3RPsAWKKEzp
uS/HVh8W4sa2i5CjwTb97/LMXTHJj68itXnat1iUdIPho2RKvhP1HyPO4iQYh2JNniYtQ4zP6sXQ
LzULtz+QVjyFKKeUNxHF1I9DCQixC4Pm9zLFi0Dx1NQ7lCYCz/HDTX7BDQw6Td9+zWL01yrgiPDC
YfuF1ietQc3m5O+srRiabI5MRaymmUHVL0NR9T1/Vgcz8j2I6Yyy993HTacGLYvzB/F137vQv4v1
r7y3PHDPjiDNtTTIfxx3aqUlOtyXVuKeVp8xcYHpEKjiYt0InRkRtwKHxk+CcZUwtqCnp0phm9yY
vEnybp48RG5fWSp21lMTxJ150salHXCcX9pw/Hph8CQOoIhq30KkE0s7ZxajDb4eGTNSEMj2gbHk
IX/W+4oam2DqYJ6zRMo+tv5F+oIPtd6zVH49BVZOfR1TJVeBVZ3A6lfNqrNoBqaIIXnMuIBhty3V
qx85CCX3Q48aEl8SWnkmzZCJhp6hYzctyuPGyb8qhWsg5U7cFngzlMqguNgvwADSU40Xx1878OV0
YbBxEJE6iNsr6nBdt28KqofcJaihjJJCXzEXvnLyoq+8sn9FMOvK03su8rSZSCwsWgqWDYn/uwGa
01NSzoyGRvRNa62PfQEd4yKJQfGgObj6hcuzrOtb8z3GoiugUd5TsIpLA/kp4ZIowPw/l46Mz9us
AXB6RtuA2GtIdPOba5hBUvO8CIAM6pkRmVsHp5Q3eD6KidJ379icoaMJt+kpwPNteNXVl31+RAoL
cx0RVvlGnMw12FuZW8MRotEeazTMYOepB3aUfQGUV/73DiYXOa7WCJzzXkkvFjgGVodGybK6ql+R
8XCBekQSmBrqmoA8eSYngz0DIGmMm32guM6x2DmCfFethu/FeDACe+8Mvz8Y0LZpdEOiO9da5yPL
BRWMntCwbQSYw874GnY9jRcdwXzfMU+LjLEdum/0loFqzSY9pTGDaPoTZQFJKyu08e75zfg1VnDk
gdLMAqkq9tyjwdLEJOFwiyY9mIfO0D2oLwtfRseO9suT4o6kwQEKXElJ65SLDRX7buQw6sWyVjAH
SNv3Li7WuM6WgAbDQVxo2Gex9LhArKGZP7eFI+rYpZOOHdxCQuI0BZ9TCo2sNRbYXLR6NG6dvd2n
4x45GFwwLxTxxBtNadlo+vNs4kpejGkeODatpr+sBFhWR/ZTCepkco/YpvgWV/bufofxY19jfKD8
QnmX6Y39M0E8ZJ9kpWpHFT/Wx01Rb8lmHk/SHUnve4NOPBxK0R+GkC6e+me7b9HxtbUa+0fA+W4T
06zyzJ51QLZpbpwRHA3oynhzP7/Q/B2c2IuDGvtIfsIDXk4pf3fTZXzkk43blafvFBIPkkKg4raf
sB+r8L1uzxT3rXv+f2Efwzx93VJ1TiB06XU2Km+4bfJXofsMBTgcnBqvGpaY0z3dSmm0xgI76KIZ
duloVSjmR2IUEy4ZSa/LbMolySlbjfZ53NCyreOsVsPGshALZAqOqR9S3b0uM4n4snvevTEQWvE5
tG2x3EKm5da9KqLtro8bsmY4lW4BY+AMUck6iluHPMBxLzbeK8MJKm/8jryCrsZAde1IPkhxixAW
Hjqhc20GDnZgE+iWZSpfezL8UuO8sbmK5abkBLMTSGGmV74Udd2Migv7TKELkE5dPgBo6W4CEd6m
4RXsnEF5azeCc45mQadkD+7vVy7h5kD39EnnvRfPzTKg+AzVfhrAKDiH3d6rhz+XwWhTkRKvF42S
ADJ6uD5J7DgErvDBJP25n88tIk7sb7Zd7Pfn1JUaUvZRXEf8E3+za0cxgl8e/6A8fpsBsfW5zUy0
cMbzPajg79xmoA38RQX4OUX/HPgevAQoELH+BhifFTJlp2Fbw9t6mitvHQzylh2KsPTesYd3WIxr
szOID/+glf3yy6LB8/V1pBmW19+ng0iwmHDrnr2iEWL6qdO914AU8F+isoxaNY8NdiflRlopHEZc
TKqWvrmATSXbnKVuCEjyVLlXsJWmW+C68vUQ6avGnVUp/0JpavO9emSRN0CO1fKO0kCivh7zhSl+
pqGrH9lT66+xcde+RZJzj1h3sXP7SFQ2GAwMqHpstok+U3O01Y7t9lz26heFzvzOPag9260UxCk1
s8rTll8pafslNkgMup6o7Ag6NIXJhh120cz423GsFpAEGJPxHPViZAgpjWc6/nqr60EBZXbiZfU/
cr8mIZeiq9y7/E+amqpV495qK8xuEM9/N/UgmJjZPYeILgKd1RE3uoc7FeMkUsoBDmzK43Mrguq7
2p8B1c/jaICMcJzvuET4jW06M7RfjWPJ0nzVjXFFxobXfHCP8uEUnHQtdFN6P3xSr7eoKUiIfEf1
XnOaFdpjR1vEua1KpzbCyCT81T0OsMFjQgzPL4/qyA0uncfOsnqwGkegKuLORNGuxILMp6q7vQDb
T0LOad0PdWqoh3NJJesvjBP0tKaeUEuX8LzrqWtXEymPsT7bRF6649hXTbjtSxB5zA4F3o8xKSbb
sXdZRikGOlR2U0o4a+PS/Pg/uQWh3Ehsog3EiEsP1A4BrnW5kAq3lFILunm22+29ojvEHgF1eGQd
+wIyJCdUY3iqk9nkkoat6bmRIOTj38RsbwqzcQcz1eVtRkoQt0tL4QUsBTmIMmFfe0z9bZEVP3T9
I13XTQLVNgvYB39q7Xu6wSSwbkFve5VYP2xjxZfqeDvlMbz/KogXHUjVBWZS7MyCSJC+Yvxp6X3M
E74Hvwv/ZutXQWogkZ+U2+LW6+VtzEF33YVo5jYwUQxrAgT0U2aKghzJ47kpV3IS3Md9WIUbLhn0
geJD8vqW0TmGtLCs8+050EP9NoMYnUhaaK+vJxxXS/lKdTjMk1Ma6HrbEWyBTyLqY7PFV4WoEPSK
5fE+g9Yj71ZKiYmGz6J+6QXHSikete+E0WT1pu6t/b70kWxYRrqzZvEJ9X7ecqG0t4eboEh1FXrI
Wn5hFA84ToYbQZQnvWQ+Mt9M2yEjtlgI8vaTFHFyn/5xWUfSNx4zdv1T/FpT7ODBK21CGKuVACpA
bFMar+0ZiuBq+5HwV4C37PEz2fPqzoBp4XvpHsRmfPcHfKgvK3Z/i2jla79yp8dVvE9bN+1wIyAN
4DWsDC6k6ez6Kd/ly/ROiZJIeuCzJz2grE6KbGXeKtsWaHk7UnvIL5oCrpG4CTwxnnFuPlVkNIhs
1nw+s5evZMzt2NyDNe3lI7dNgFc5ON6jjOSsvEkwY+Cp1JtWHl2iu+Fr8cwmdZI9vgD97yUXKWn0
i3FfJ83s5mrlD1tS7YQiaAKGFd9rrSFQrW98e27RQa4w6s9qtg9cO7R5wmXzy9y60tmHJk9zMRjO
ZNeTaQ/GkVnwyp9Ia+1J9LF9VGPOi4WgW3TuI7cn9Me7xT0YvO6vrRrnib73qw9/NWsPlqsc0l96
532X2P2dUJPlEwnCsxPwL+nJDFETfJYO8EHniotkwmjqUZbc/b4ZA+Qt7eUdzjn+3XDDsNSZa3Yu
QfGSisFaLJpaJ2gDUKFj4yV+58t3Ced8JGmELtsar8htC+HgFP+GMwsRBtC4tQf15UM+wyrwJCw8
WrcDyhKqUsUh0rCzvezZFFSPG2N4gigmEYrtocDqiEVzVou6wtmoTaRf7TJ8IPkL/vKIf9oN4sqe
/4ozOQvWJsNngBjaZPrATgDdL0ghYrNnmtmGFQbb13j3eW6QmKUng0wnv4Xx0p537Nvz/JCaYQo+
1McFLLgFcPCC5cMrBld9h37ch/zJnR/6awf6Oed6os58YxKVHKhNyMf+iQh1hnRKAbahA0eg73h/
7HAWWU06dRn52cXMIGHpgGtrO9YD8dVZ7S5I6Zw5CPIi8Yi+PKuB6JVtYwZ/+gCrDX2ty1OrVzoz
7qEJ+J6HeD/oNiOJ/vCaFWIuNs/fceEeL/2055D6pc0TUxZhzmUDjo+MHWGJM2u979VUANqqPrTx
SApSLrZOGBoa84tbfB4l5Gluyu+CUnmX7o7Sunj7GA4HEPNE1y2ImPljp15Rh9iNnT30b4o95mRQ
bGNXpe5vVbGUIEcEn6Izu2+lsYnn3IMPqYCQICLJUtO0+X+MXzlRE0HzblgN6i6Ul9tvWf0oZl9K
zMZRHEk8Hop16tUVdu0EWNkM1reZw8AQdiJfkPo8QnMLj5aFab7MvFYkcUf+44VrNok9HZZv7HRh
wWJlG42Baup4VGWrTvZwipATOUZof5yQbiNbjqmqD8GaV+I2tWN3yqcNowJ+pMIC/5+Mh5dKy/K5
Keg385n86M6GJzk3LsfgJCj06YJgLMmBGc3BGwEZVbBqiVndlMe088Prc2a2ShfmIVuwJLavczJg
hiPtrPr1ZZ6cDQe36qdXDqHNJmCtd+loV1r7oElwxKT4QZEHveM529UYpvy9v4xoUpDzgSguovOZ
DDs/QKnXnND29t5a0xnscibRol5UQGIgd46CCNnWl1OETJN8+qhzV7rIXLs4lb7Uk4UdduDZH6BG
mN6S4VHvZn9z9J37gyv96bWL0czP1qEOu0/xeL0SpLkQTnNwTKzNsKgoM2Mj3NHFc9krr4W+VgUd
ufguaRMuxFL3GunKDovu0TZzqBUYlZzXXDBXOeoWZ6PLnrCgG8xA6Z7v52ccFaghT5FQiHg2Ybni
pnL0jVqfRYBw5XxWOhpJd1oiFdtJHKjn7/XMUB4SFLHjrfNz9EqtgQHkLoup5crHJzL9ttbbSeGh
Rxs7CyTywc58nON1cnnV8ls9quf7i63gmbC+QrKifW2j1+lpgZ1EzdL2Q413y5dYsmAQ1LZZr67W
dMsyaoJyS8g070vUSQMiw2if3hQZAMyK3aX+tSSU70kJcPN/FyaGY2RFCo+6t/cHvJGaiPrmk6ti
aSMcjDpT+fFQtnnFImB27e8ytOdYKL8pTWju4H9Z/omiiCngmo2i2RavGysMYOYbob3v6zVxSsX9
3nJ5ZTN77pxcbRqJFSY8NoApGFkRv5EpMPpXAH2PuZ2IQ4dVPGGJX5Rr0HvbhLncQcvXUMG9pKq+
hZg7zWmoZenfWYySr0Fz2pWFc8H2C7a8NTnq9cSG4k+37St0ujDgKsmjWAuiDHTFPui6pOHQY466
q/s9JOqRr25CPC7QhwBAPKdEGoQQepqhipZdR2ZrBjFi+JH1OiIZub6oFY1A/Wo6v9IYqHj0oH3K
Q4vp/Ky23qPfgDJPP7zosqk+TvaFZXsvs+n/nzRXdetEjcULHnOm/b0r4GDPwD8s5bz8tkyCi9qQ
SyiEW7MIk/bJDyEx8bF7ECcz46PoZWbwm3p/4wIPardWGdUH5ACq+xF6RCN4jkTPi8wTMeXmZs7F
2x2WF9zZxYabp1jx/YB6YvwHO5/S9qEiHp/b1Zig1kbrMxElwuU6cikXZ5q2wOO5U2fNc+HCd6v+
my/62zWEn3IaFR+o210Q6FRAO3B76CS0c5j7cwjiHfIuFb8JsmDwgn7qBIljuynGZjBTuGQWXjgg
YZKAV8pMiRNsyGQe/LtaVJsnOFZ2UgL2wNSm07p/TOCEcSBW8iUIpq6f/vaT51CqTku72WIaiCl4
mn0rPzoCFD6wr7XCuJl8mW/BGOeOm3jF+yUVI0rFEQRrSfD1yzSvuK9bIJhgIBF3YBHkzvIEDAI6
ZF+rEWkKJjdLd5TyCOfAX/4aYTPoglTlALc0YQ1X1owyypvWxntmlNueNv7TJwhlTELqtmCTA0x4
kkTNL7bPfMc0V941GYmfr9eLgpCOljb26EIdKEFPNS4HWDnYSW+Rpz7UF7IytKSL3KBrwITTsx+a
tQZxoAUOX4cACPZGZp35K6GFcfgsaMzTWc0BTY6Dq1Jqi6Sd61efGK2rrNayeuAQblMsHECN8LJO
e8cLMb/CCrigLuyjA/SSWRF8eZc++6OFoQ9oDCW1eoRMYCDKVXYfqsNHB/sezk/o9BJjktCONLTy
DaToILrhW/b+C4x758kKUv+I3dR68vnhE7Vn3K8xJ+UwZj6PahsQhaMvlVwd46/zUYg5b9tWGdyG
cYKJ2yS/aAFbH4MAQgNDs+ZyHm0ipIyMXFl8SRqKmVg5/buoQIEsrSK+a82F3jar1Lktg4/9cOoS
gH4Fsqd8VE8FOqRIH6Wb22zccE2QXAIvk4c9Xb3SwuSYcS3qEZ6qDtIAOHn/gDyQ3tu3OYAfMsEn
C4rQ+NwtHgYakR3Qafn6q7V4e2e1GpJAsoVRo69aSc2KzOcILXPH2N+E3sKf4ACmIuINUa/Ybxs/
a7lff0wG2oPbc9OZOArMskOUcD9SGcu1acpC+F2KCgpTdAFc2a0BLpt+zTr6LmkQPH1pBJP67mhC
eokLyJeYsgLEIk3FPD+kJBun22A8YUOirpI5rp+WxB4e75GVZmMgvhCeZSbU3tzu87OWeJDrwDGz
LlQHfUVUVqGRko49Rtl4Sa9Nqyj6w9t1wF4M2Os+z+QLRTFyyxFPMsozSBfpsvHlGIKbHIlNZR/n
hAQ/KsMFljpsSjiNMzLzHs8U9I7ipZuOyl++TtjrrUCObW78EsHAp7UXQecVp8tSDo8oIOk0pxG4
1SLhTfEOgvWjaftOZlrru8hoRiFNyhuuPev2g3WXyWvIyh+j/NJPSet9t2dMq2fe+xJ6Cz/EoDus
5E9bUv/rnL2zfQ6GBptKOmVO6hxxzfZbpskzAHJfkEO2M0XlWsbjdE+bPrSjAJhLaceTNethP9CI
6Xhlc3tz3FLOlMojeBvdqy58qDs7x2ngZtV3ZLrmSW61zKs/Isvsl0bG1ccsMV67P5fsNXOLQVAT
pnWpAdc7MRbzCKZg8viRoDKefe8u8zXEsdq4LThLm3ucSumpboE2HanjViel43sp5K8D3No+VAel
9hL4ZU3jivUcN/RxnnD+fA3qMGxnB+lsD6b/NBYuNebO+mhfgunIPkV4rgbTbZ9qx2vpZxfaPkeO
a6GAyv210xbKQNIJ3i/EKmR6qgF3ucovk+VXOAxtlfTLODfVcixTVmg5cS2BySJgLgXcnsSRwxlE
y+VVy0mbueUbwEIhA/pJbn0C7FzWx3POjMQxP6MGe5YrM39Frh3wWViBRNsaHU2bM3dZAE0oG9fo
34SM75RSy4MMwMWGu52KUGaPIbAP2WZDqk0igLmbmdJxUqh00yrxnRj0RX6ABZX4VQqEomdba8r3
6L8rB9GwgsuraqOtE0oyRs5McVCVbSrRFY9wcU+i+h93KlyPJ7wqRQP9jFrMzQgYVck8vGlpH8/T
E18QtWRixmF6ac2q2wMwyZsl8S75itJiY/foXo8IMIwGXQ5t7vPn3vC52J9Be4uWvo1il3Wq1Xa1
EuJQZK9/u2h4/VV82+WauE9BujOMl4/j0ENoL8k5YjJH43nt25KyeCKeqGQYnpe1PDZS/DnNF63w
YzmW07Bn1AHZtufhNVs5Z3KXS+qmaLSiCB52C+PTfvQZJOWoCj6ET96kNhV+TTFLyl8KcOcqm9IY
XVp7vhJtIf6rxwZt+XuF/J5sAxoJK58Nz1n+T+TtcDDkn6PGEFtER86hCBL89JJe17wFtYxGbzAb
VLzqoGkp7wcl51TA67fIbiD90c3oFa+XgomvjhQYUtx1VsfXC5rglgzB6PSs+Za/CUtRRn9xE6bG
1apGvD97gSIvLDgBzRYX9EX+FcOSlHIMKjRan4Uf7gFMOYxMkgWHvNR+SrT0LJuXL6RWOsM4z3XL
VCtEkFKG6uvWUcQtePFyS7hARhZEJshCbE2Pkgr65cTupMUPq5GjGEEIpo6BJWrVxVLYcQa116m2
gRTXXvKRNz6IhWeCVKPHn4WzBDc0tvwtQYW+XVrFNjtPMLHR/3EljR1nntlYsKg+JOnG+zpRvJbu
Kf9Av8qgXR1nawO1IPxwci9K/haYYerUF5UmT5p5CZMLY61IrtvfZS6hZkRWLnKIEo6bTneWhPak
3e2+MW/xx39MdyrE2mNguGO25a66XMRgnFCPiLxlJRq5VZjob3Z/rsIEd5aMV/wWTmlm4a1wlc+q
v+E9eASYVA9M+OBoL+43zD2HLPsnLVumQaCNlJZfkMY4seEml5jcMLeMXHdI8nWnSO+/6goiXEpx
6xL/IwVbkQ24ZhVjkunSRftHGuC+gWiSEYuSqD3192phS8qKiV4DBikpqNsIeX/13vetd60TD7DH
U6hfsBV9JDw7eMFcucF0G3g2s5ajy7milCr/BM56FVuKyFmIFjx0RrNiXwFXZcTvkk1s45kL9nnD
YNgUduQyLt66ZeBfT5dYS9BKjqEWM9A2FvBz4pswd7ma7q2ErTj6GDMHnmc7kqIEWPEG44bhkfqv
+hKhbgMBdAKTihnNceJPIEhdFOpencd0XFs/YTAfyXANxNf+h+rKvgWdcIFJThiGpJS84X7zQ7y6
J1IMq8rLNccYKFWeXH8RUP4E+7mPe7Iz0TVomneBDODO/lFFiIva28WIMWAMLcMn6M/EFct5kTW1
+JNqm8oOHC6or0gtpexHROJfeZzbyH8XwE6VXGM2LMqdRgKfGBICs1O8/zMct3yI+FKvFcTwFvTN
TqRL1KTw8aNsE2Y6x6QSgxUIVDXsC4RzwMNOu5XOLnV+MCjQWuTG6L93GAV6I/RJ2DJWh/OLW74d
ck8QjF1yEXLj3j8XeAsDA325pFHNIJn1TwAMfvL3/WhGFvcWZJxOs8hKv8pGmFCAo2LEsXz/04gg
jKmlp3U6LMF1IQedJwIMI7EjM5c/rWPcM9cv1U7J/DZ4AJeCfLaFK0Ichvf9Y4UanXpQDqcYlESe
bOL/iOJGpm5dwtEB6GdIIog51EZ4atDpm1GTOVgZroP2+dVwXwJVbHhvFAYzJ/IVJjhqtEiQA+Tp
aWd9c7Zwlb4yHUJ9MgEChJ6yB21MPIajnNcV7tPqihgQ18Sm3jHKv2dgixUGRIFiZlutUZhDAH/s
nTRzZDhxqC3Izpr/b5RCftYA2li+GqSXuy+ju0uY8luQura4AXrRl4tcOE6/YLQ2dmEc5QR5U0eS
0Hy3RDTd/j6W6y20Ulx/JLxY2f23y0mMG00tWfCePMDP82i6M2yxN1gBFZRNZbaQ0nytv0HG9PLB
v3tGi4WmKnfT6V9Rx51clOgYVA5e6m320Wpw3itPDDAoO0DCmPRTLzN7eB3wmg/+sW//lktVxcdJ
xTnytxI8mdu4SNBZvjsrYOhRUVxrPtE8wyMzPUN5ee9tYMgeJeIgeXR91TwhyAnHZch6BiMzr1bU
5B1F44jLDF9/xE8ro/Lf7huNiZinqr6qVFt3gAb6qsqKvzfkTaIvv7Rlo1baBhm5nTMxoXRQtmiR
Qt2/cgyK95s6C2TgNb5huQNWJvC7QtdFUz+xUmY/zdjR+XrkqYMrwl27ugtr0AcXrvYyYB4XfDZ7
Q3MyXguIT7IADbLlu7UAsqy7d1ONta6d/1mSxJEhCd41TEpHUfXd4RH+2y6n8gzOHjYHmZdC2snP
fibzzA9PM2juVsT8zz3OM9qTVJDq8z1oYR1iOa1ITlrn0vKqSzP7x55lA0gc7vJYkXPOqoluTra/
kfn2BuDnBVpQ7ka5ig6ayzP/F4Zth2o2ZeJhL7m+dkem3r9B++iKHEctqxUesVxpqhuL9Dvflyb4
39g1rWZB7oZs0mK3S3n3fwOFvoY73iyO9OUaaD1F7cBteCNDpyhJoR/ihk8I3EsWccw9LnOvdgL1
t01PUAARaaLSWBM2ILB+58oUSBN3+gMufPtBH42u8hS2IbRZ1fC8oKBdXrXlG4r/ZCUbvB1nlNgc
3RrfIkwAAlBSUO0GfSge3ADeS5sPgDen89+rfVc6BitQzpmgI8GPkkGmrP8XdHPoD9Le4PF/XVI6
rZtrkycqzGRNTdlEuH6bQfXsre8sVj00m3EoZBZwPY+FYEO51oI3IY1vpmZQj6j6nXNldAv8/k9y
UCqKYyzdmzVUwoKpMh9Tvi5lOgRjcaBG4jd9pZbZLzYq4ielvQKBVPuFujnNl7lsTuBxKEkPi7X+
s8i5pMqpos9iA0rrRBN5IDmgCfNS1gshJhsJL6LsKse+sf8GZYqD9H0FnvJe9IUT6g1br+zzkVmT
eLn2Y0fI1r9KPR2clHEuRa1ErnRIcuS1JiIUriZ04wdCZTfJZxOypr1PFQ9+YVM5PlU3t/EQSPXK
VEbAN5FvycFiJUdQZLzEGuWMN1ztZlQ+dRtoeupOF7rB7pjHsnn8jyQRh1UJzrnW2fIdOY9DFivU
uNS/kyZX38zGtNRnB1RGMHnEBbFuwGUQbfj/FMAVWiSZ/7mHsVWsNllG9yBIBPBzR7+58ckMpA2+
WIwMjkD1M0cC6aCgDRRnSrS9N4hUns7SIlrLpdZpRIGnu+jhhVKpzSv8Aad42J7J/ti+a6Xbm72O
hjN5tOI1Ha7m2xkUB9NUY66U/tF3+qoMD3OO5k+DYf5iSxb6gWdZVk7WCQEHoypBILfUzn2fCuRw
u+bg3o4bD4vx/5vRZ88GHsZ0ACIV537FKWG9NaSNo4zJX8OBUQDUlJfcESVL5dFr42bHEVc6/yvq
OMidfMPGNj78BJLMvGHWxDkmo1sPUeU6/LDPzmGcgz+J+zl+NRcBRYn2GNOVhTPHLQG1H4u24TfU
0PVfXz8ahf6ZII8C4Wn8V4pfXmF7+kjaFgQL9tDFJhUHmqeqHN3L/29ZLG8jaztX7d2RGcyCVDAE
H4illKOl5p0KEp6JPjnVgXnBUtdbuS17p4inNsjuhX5MLp+fIFd0IMhhZfilqWK4p1FXDGJeP81g
wXCyXzRrxht5A+wjLJxBVsGZOu71hySGTz7KxcH0eQuZrPOoDpqoJISuEXcxASTglcmlSY1Qs/ox
o05YY23nwXYWzX4vI8tNpLLKygQwaYMIRXgCddEUtE4SJCtaiez4SxF442LO0rogetX4Wx5BCEql
w+dkwxrwtjHFjCUM8DAhS3w3JTgvb7gZhejI0B/hNNQ0mM2EUT3o0amGheaLqiC4Zm7cF2AWfIW2
j10Hm3AsXRaiC3hm1NQN/yEN4j3sZY0kDX4VrERczOBbUqU/M8k7kuSJ19+x+MmyX9UeoQsxOVcc
SIUamdLN4tIqnmoeD1ZHSSbk3yjkU0PHrgTTvhimUJMb8mWHh8iaiI+Vac6RIC2RHkoU+KscQ9hw
2Xwwh2GwG0+4M2dLQ4HL1TrFBA60qgFl47zENkpeuP8YT/zAq4seUQNAbqWGzaO8tqFpyr4VelVJ
kK/djF/rWrrYa+XrY+SrkpLt8IyCBM91eB1svr+9+9izOEiCZHeGHCs1h+Yf42CSbVHxefvplwJ4
Q/PbaIhF8OZjAI51fD5U/DpJa8D0Hz+VA3qPkBEtsNTjVB1/Sn95v5Dihb3SuEhTnIexx+KM27z8
hkDXsLgeZpUThPy0roioCOix+YmjQ71nM0u1SISHFaqH2+B36yUfZoXOJ66Q9Ps6wTt6hl6veH5m
zV7gRPK3aSMPugfdvYh2cbe5N+Y2Eo0xkzGxSuXiDpkynaoP3EuF8qXlJQIet1Xxt36OtSeKz0Da
hggge0haPs/VeW5eBCPqZ1rhctp1seyuHkCNH/F372mqd1MD9sKjog5+vf3ONBgtv90428I7nQRq
b9bXNd7ax4/u9EMp0y0WLOqJZZS4zO/29ql2rXw7s7hHnnDEHbwDWeIHyS47xqIo5QfMjFSBu9Ug
gpdAvCv6A19C6MvHZouPEFyVOvZroqyViTz3lP9ubl3ZaW2ebmN3ASU15CyL5N8yK+D4QOTRmocj
+ZtDOCqHDsaK8HmXqpZBP+dswm6u+ZDpOOqgzxbv4akHyN9rVReI55Ny2ucNwzVIN7Zzm3HpqymI
hn73Bz8ONKdkjDLOrX2gIRbnOim3M3i/y7F3DAWcI1P2RMjm0hnrDwTpyls846YqvbJsE1rHU4/J
IpNg/633fRbdtMk/Fqwp2vQ2vbFuxA9bh81XnHwxaeOHT7enM/5HmJ396mDWtWCEplcbEI3qtjda
+7gAYUdl5dTq7+IvUWrAxb1SdNvBLbaFjQMdzAjk/lV+nFResAiPjeLSRwvsNnKllEkzuFruBaNx
eoBF8mdkiqgZavMOQ1OlVOC2LHnXzsbL4rDI2Mxa2CmZVVvu/fYq5FjZsKlntWwD2dQETB7irOei
KsM3hsdmoqQegdBMKzeO9sP7luCrYS5i+WPSGIA6ZSYdCu7tH5s1KyG0vu65LxL3Wisj8BLYa5qZ
y0YD3W7KaaMzfAOGVI/3hRT/UMAmoWq5b6PZ5Z9KdJeUFU1O4MybA0YX9C98c8yinqSlkgnWn7xR
0owMClf86xFH0Oehf6lt7l8V9AdYYYfi8vLqX41CEq6xy5HZRNzrIY47+Ha6nq/7MuVxOLSADrDJ
WPRtYaQx0rAqoYtLJ6rwea7irj47ws2dpHWbuQKTxd1N9ihDQzeLDn6Seh0RpW5Cu05dEyFGX40z
xaELDy1zZ/Je5KdMfMx+CXLvKwiyM5kwx4AfGKVc6qCbURF7vuYdgtCVpOKOIAp06RQaZ1Ovst6I
rIDhPl2dsoYxiwW+ver4PtPivV4HGAVxyxstjbuZfqL3mv9hADxnz0vlhrqD8zqMn6NAVep7Nju7
7Ccl4SIn05Wbf/qFLQPIGYGAGASCNY3uX4P1vMvm4zJ4PgqltR/8ciR/jrga5ZcYpxgcJYUsruoT
PIr9yv4kCLuDrbOste0JnTNGzF1blSFswEsJqY/TxDJe1lP7Wv44iB0YPUGqIl+D2w7TuuyVMNBM
XuU9AMy0erEVYi/5ai9KbEyBpcyrcQgvVjJlYhJU8tbS3o5VEkoRIXAMFtB85ngwVvvB/7U3MCw3
4a+hD26fB4UNUeHkEzuf3+Wivs0Vk/BgP0JfunC0QpTUVglwgKQ4eVhWhMSMibOYplzEZUrvDm3C
4I4Kfhh0JR3ccG9Za0Mw83T2UMyi+hLyM9zeBZdR+ZPK0Q+98y/Jur5y+QUJEvvPEtqdK6hfYqqq
WAGn0dYjstOWzkfE4EBk/Utgp6JenABqZaB/fhA45d0UJ/JhmnhK5pVelLcwTAwK+u6h3JCAtIc5
7FkcZNJO+OZgPMO9oXlyHqS7Xcc59AjAgUqWHBxdH/Mfxp6rCkxZjRWqv8EeczuD8owfn7EoxR/w
RFq4E6aCKPvWRtj3S0DeFD5aTanUuHwVuXpyfw+Z6yUV2eoEekgRy6PWjyDCh1xTB7qJMdrLUFca
JuXxOMBtAjv7LTEcKLGq0zkOIPsbY86BYSI0XO8PNxt6moelB95XEwTjBY7seRNtREPl1L41Whi/
ueNSTvBgOwruZG4JxP6kAwM485BLFJL5zsMv1Sb8+bOALk4R4lI0XhJnDycaWAh/jv2MeGgE/z8S
sU+nhM0xVXMuDqBcn4JJA3UUhB+KTGq4cj/svsLRYJCUsbo+C7W0KDnbmqGeNZxxYBjU9ryrZXkP
Y9oZEzD50zp0an7t2IvJABu29lrl9SONVfitZ5HsWc8cSt0AxZgZ5YnTQN5j0sNJVlb4eFIiKguI
pjToatAgMgpom3yGzvoTJIq32ko9Zav28KKRmDmT0+NWoclIZvBeJ9X6HmmOaftJabv1Wmju7uHN
YlVjd3iYvPsGO/in+xVsmgLn+6bGmgLv1TUijzZysN69GI9f2bhcRUhNwmgeiyFOBE9ekkKrYryz
Ck5Fc46oR9B7qpk9kjB0hopnnsUXRuZfMjHmLeAC7/+y6ZbuBK6DVLCt025/U+B4QSg5OnPkUyZ5
wmiXslZPP8aFGaFx2F6i8P/Hgm1Si9X6GBn9DuxsmEtREvnwZMeDpZ+/OfH196xS3owPFt8pYZBL
ofIl07TuYcRZUTE32DD3JxWikBJXzVl4qdWk9qmqjOSXbgtmScBlb+DczkB0A5e+601zzZ5/umb2
fAxZ0SgE6246Sb+pkoAQgeH/8wE9qo8EpE4MzBr7JnFhR8iVGqI7A4oceDPhxymH4U4RUo7uRCll
p7TJA1QCK/qt2Dwu/ongwXyVST1zIR0tH5PF0xvwD0zR4uZdC2bYARb0E2GtO9OOm/O8YtMZ6NNH
7n4ZEPYvjxWpbgPLi/04i0iQHnmsDf8lxi2ZGOjkrwtU8qCUURyc7Xq0XPke35j/fc/Ug/KiW7lt
lk3jc93BVPEW471OOXCmhSKyHGh0aJzgFTorPCIrvShCdkM1xuhEQaA8xHorxmYRLe7Jq2THdX5E
O1I3IUFY1Icw8AjiqrAy74K3LG7nDUcm0wLLan7o03sSj4hPtCAnwh88N/otAGLAb07gko1zGLm4
rXgM9uGsCHVwAShzQ3dsntousz2W0j8ErlW8KcFvT9HZA0pZxPa4EaZBQI7rbWfU9nckgXCy0x0d
ym8jPniWEtJhMo1WRSEJLTLlwW9Xxt8dKgGLispoY8yQlqPw6uDfk9InWsORjUCU0eYB/OvFLbjO
2dJkNjZpkd5onWh1hIqCAf8zJtXR3TVW0LtM3pK0hvVkGp1uNeUljv39PF6uri/YfSeF4Pg4p5Q+
W1PHmoeCi5EOYbkPAo3G9tAIXCL25sT+TqRdS+E+oMy/+wfdzKfWcMBehjCel3o14EfZB4OXqn9p
TuH/HFOTnEEuTSpO3LSy7/3s8SHS1j1uaoIQE9XCVGAWtr+Ttb6SmDZUY5nSGlT2IGnEcvwvYBJ7
wAf731//DmhGiJFqsBiRjs+vfC5jDFFlQej3wCl8J3ahSL+LbdQNGMS3VksjSfJnwj3BID4QHhMh
pxfq04npWAklE/ickxeTJUNlF/V30GFpGWJ9FFPty1vS45TqLXJsCtB550m3jJ6pewoHMqXyNFYD
BPbFEluxqodbIcNLdlOx51m79j7z7fLwP1hy03jteIxes0FQxZxVo+spPLdEAbdLM8DjtTjY+2g/
RT1VeNExuGI+qsz6r3EO4E4Ne8kyfe8cSGl1GqB6F7L5QYTIU6ZuAvlwMoqGT2ix11luMyoNOpoS
ragMkewZJJdcypm/OTymyY6HG3QHuJthUTMTbSShfklinTu+sfOFtxmlEbJZJLgWeUnw7RtYjbb6
b6WxAV6wc9Ukr0xKJpOEdLvLjaqTab5bUYkt2W6Q7gFnanDZY1+stMjdesbRwq97i5gU75palkCg
soHbWvP3GLcZ/cNLwvlVzjwMcjKh1UA6ev0YdaCABZNBG5lBUZ7XmitGicY/3n8w11RFhSlCOWHH
zaJJ2ot61l7cCOu6a4OJFCf8vORtpkGaLrtSt04ujVdTfb/t60Dz0zJTBSaO8wNFTSr0tA86g5N5
wYmjx0U9TimHurRFVjxaYTeGsZ2iZkLSwin8WAzxSrp7fFLYPi3fX7kvRSNwg9oLzYSepQ132EtB
mTpQicnBhPjA1mvSEVIgzAdzlN7CO1or/ZmEfj+AlnSI72qSA2DpinQuYy+F+rl5lwnHe9CBIjKw
xVsXnBCTY7jwE0RX2jCpO8fMlvKFVpX/4pHfG//sFel/CZ119xXeX64ukyFwLcgnzACSUHQIXE1z
Fpjtwdq7+wH7YJv8aUrTy8aFVGMgj9zvVEa9vEdfr0l2BFBUldw4JJfVBCgQcH2lgvi2/rstDc5i
/P2hkLr+278CKgT6WZ+5vli3iTTHoKTlbGuAn2Dg6BOk4ArO46TlYJ/axURKd4ayujpQlijZ64+T
RoqUuanOoPAS7bi/FP8RCWORZ/Cd5SF7+StY/CKcvmsCjJzaFHD1TNoirCAZuoKZxOpFPo65KF5y
mYL6KEuXPsSGBbeZDTr4a13oZ2S3tHPrV88GkzHG7YzuqwZdIE9F/7o15qbIAoHNKPRGQeI12VZP
QRBJac2PPvHWXEMBDtCUaPwOj0/pPBH7Vmzwn5dO7yDfh+NFD7qCZXENbk1Yb4uNVVZpnzGSvvmQ
E0o1gKVCYvTCybE1K4Dm3eXkNPB+O5huuMgr5R2GZ4sBgGAg9LOstyIwz6CuqAYGheH3abL0tR86
OHh5yj1S0UphQwjd/okN8uGov9vc3GsQ3/u5VdB861b6EUnV1vYaKeM8iujBLgDIOE3pn+qo2fvF
+hN5lnnnM9uWvwR1XKLw4PAG2VESYUqgdVtFapoZmSotBdWJzJFOY9urS/ej2c9/tpn9Tu1rD7T1
P2JSlwWIfah9aAxhSKOJ/tD51N+0vzvT556hxW7l6WiXvkJHDq2M/yrPznUDBmSd/Tf+95+eVffs
cTViDM+Iwby2l1fNmLWpdig8t27kFXupFAuviu70hOf6pjtgWayLkDJU1Ka+lPewDQcl26drm7Vi
lxehsCraDuUeKhfjPc4MWris8yB0cZungYphHYRa+GB2mq/Ja8ByfQhr3tyqKxi4B7rMo33CCFiS
yOdAo+Nyn30vsqSCPSkD5/Vx8qV3FFXeZuZWKdtM7i4D8p3cxKpgsLRXE+LFOZDNLyIzDkniVLYJ
XBPsYYRNn2dZGYjEbWTZP59ljbxrjLWnek0XtBl/kD6VWnw/6NfmQIlhMr9fXnD0wLyQE+RiT9/f
k+TMZkewy/qUU5Kv06UVoOFFlKq8YTc+xM5ROk/Wa7mXuefDCR1cAEnFZ8+a30BQlvqwZr9ZPOJ4
nXDA3chyM1+BokLR/vAiV7klZdZiS+Xjbpeh2bljPdxAL1KN+u2KLqFK/JuekXKLp6qRndJit8Jv
JvSx5cD/2vNsUteMGyz86eogFHi1VhWKyk/AykZ1lniB3/YiFOBT1RpEpEdmsVWqVZieTngg5qKJ
QeAI25/R4RpewbPmnJN7KDuleQAXMhcJ4NAOuaHbBS6xYX7weUuU8v94QhaSFQKsjty6TbTnQGSN
trhQ6NL8uHvEzDU8v3hvshwVqt93qlHoDgVRbSbLz9tg6FrWfA8CCXuEkE2M3eKF84o+O7jrItGf
WB/3w0SF3QkkGztTTwYsScFXlpWJYinRJhjGAAx/hZmdFyU4LqDDfh6b4TJNwQBx+yLuJDEWYxWS
T7g7qo/jvtN3t7EvOHDAwJiXOQR7SQROivADG3weMpWv+jtJcBP4KNDS/UYqr2bxnsryAnxaxtLs
ouy8XCG99rbEWgY+ucFn+1jU/HXMMR3XDrBODgeQMTCXxpvCKc8DjgXlH0+GbjDR+kr5FiAzHu8I
+DOFebjeFU1CBt62ZageUEQ8NfJTEOf38o2jxuwR/dHYpfTLYs6gEVR1TwQp9Q7KqG1EkI6rS9hA
874CqWBlhBlajFbHKotCFkVW+RrgUiB9aVJhvBtntSC38UWqe8l4CqUYVnIv6jPZcgj/YPDnuZME
WixRvwB/0WO65h0BCDOGvWYukj6XyLDyP1frevEISsQiTDcSLZh96vTrLwpZC91bmCF23CHYqWNV
U2c39XMpIhcJaFeXD/CA3KiBhjVAoCEHLIpZa1+WCZ89vUnIFlLOzgeb5cjy87Nr2PDrQ+L2STuo
epLVR+LnLknKU8YYL0APXlpS2v2kLqAY2q9GYH18jZC7iWDc3H/dhDj3MB7I+jhLPWRKLgcbjpbv
s8aSTjsMPOWRwe1tWeyCMOP3LJCbfTDQSGVYa51pVVP/kt6UpwU+Cs4XpQ9e+hNbRD1U+y6EmKH7
mhr9qXGsSoAphHUuVQmjHfpsVntBz0AnlhM7k4HEnml0tXaFJoHWJvLXco/iZrNpZ/jAc7iBqWyz
s7H6edjeT1PRzi7JYYBDTmec/8Qyiafdp+EZXKA/4/CBSE+30vc1DR87b50ATr5jPUUT+kdG4KH3
+e99v2mEHotpE/fV4Ib/D6qzoYkg72wuxeoCH37RnBecCOV/WuvEr/xEi/nzgqcT8M9fIjQxullu
ylaoTG6UhpvOvKGCq8EolAsnE7HV5J0QxaeXYfC9y9vBPVEPqHb59PAATjLgsX50UXmXirWp+4Xl
fPyOHkwIDaIBwajFpusphqVAFpayRRzqGoVSXtwN1OYk5xDiWz2mmzko2qi/UEp7YgXvDnwrXBYT
8m9wN4tjFPm4fy3ta0koWElcP8fYUfeAwPlwQYWBgDxZP3I9v+d1Robv3tC5YUKKTNMDJd7ZcWFt
SuwSArLiVJFbbn5vXtorF50JnyS5dSkIW0s04tvCUxTiTw4ZPnvG5wnF19NcRUqjSys8dDv6CxrS
2/XIu3qnId2UzARgRJboIkRv5s+YyWK1NRn3q5fNpzGs/xiHOrsXKt6jdBFHUvaTkyZHSfHmeyLt
w6ujgP3xe4z/k8EJ8uU1jFcq2j/WE8GRzGcNlrKT/SsKERGKUZsIX3cetONmkPWU8mGOVGrgA0jF
srsuADcVkjr9cnBHeF26heA2yJE6mvT9msVR5G22kZ0rSmrZchzpNrEYRrXV8TuTYQwSRUGUQpx6
J7eExl9grR5luUj6UfeocdmpDFC5UyKrgLuENLKNPsWoabOx2uN2KlXpEfgFOA+NDWrvcIZAoJyc
yfs43l9D84MstNhuX+L7Sik0sGjpkIsmp0miC+TkQqiqHlgOkoPJQQOYY4yU/jS53N8oL+GVtKWH
z1zXQCbaXJV00HEw65sVmw3ZwykyDcQqpJE9GeKLGnj9mNDeXXET/ZQSgl2K0LcTCKM31KG4NXyE
gaV3k38pqaiyxp5H4ULN00dbuxsbmHsOsqpPxOx/j3t11vzy/yxGCnIbXFZkulClz2keFsm2dOrX
447JaY3XRQVu6Lsur0/LDirdo3Ptnw2YUpZX4cEmteQqNIzPE283dqo3L+nReiLZ9sQv4Vcfmv8o
BcP9wsl/ifpHQ5Zeu8aisEWzdWM0llCxyEWzDXZzLHf3EBRPN5oJcCRZD054Yo4xuuvVlK0IwWMw
cZ5qppLOMZQbH6t/x+MXSppgEf9U/fkM7sASHPsAUicMVZ1lLl3SFM17gfLNBXz0pCE2Z0sijLcY
9FG9ZU6kzJGQUDph+FleXp10a64dmD+v7GMWKumfxeb6Vu8/GH1W6AGldirUGAT3QBZC77CtrXqf
Z1BP6tPUiLttSIda2J0LYQEqFb1Sw/R1WRMna07fDd7LfUuhoBnkDtaAYKbIFvveKAm60uCQcrZ0
l9kzSSJZsorUIM5EJSOhfIjFDF8wD3tPChFyWMFTM0zIfQa38B/0ClXVc/NMdvGaVY/zugmOjhJe
H1zrC1FEQKe5xQhdSXB8tsuwqUGqfI/GXxfMK0M2IqHMRJMUHxgUd1xtpTADO2+t8fNZ/zyD4e4h
Tkkvvn9Ytma7GCOi3oRxwwb2wR6SiSJEgzOpIgGbAOJ8fasEXlqJv3/PYIKtl0tFkAzGGAFaPipl
0hWlF+hl7mK4qrY3vYYqOBU3DC7W4jzcooG2xfJrjiDLhA93sxXHazWKKMTNQVMp86g0DfIHvEmc
BYFy36x1zY4DeG6VdmN2AYWOOvc2NCAQNPDw6yqe4BP+wCovje4Fv3b3uRKaFlJhqQGHnapQl37k
5MdWjIvPPOiSviFa5gn5+lLbEM+35+gGkx3yUtsz3NoUht7wzWpvU2G2uVScrBC1+WhZHX/L5xCs
ruNjgWq3IWqfErh7nbEsL6iRZy8IWTz6VLBZRFHH6xX4bQ7Q3jSbvkFIxk77lgZdka9sOCTE74z2
g0+ausLSqWNxtwW5cbYiqTZyr2ZtXL3muV6GeRKYC+ABAONVbX/28aX2ZgtvLvsln34A8Wz3ZBei
Zw9/qknEsuZGJ2rEzlGn8nz9GS3AQb0SreHBjfo/DtSL3Ct/f3deGBhmhsBEAPuNupAw5aX3Rcfq
gQsHgivFBshfzIGCs9kwESAmtC+GlOZD1F8wofKVZsdSwTfWSJg+NfnjJZ6o96T5UvwSHC97NUPE
80rs5LrTdsYZZaCD4Ayy8fVRdZyK+ZX+3NHhsaROFvOCojUH8OLf7es0Aslp+xeh9ceG7AaSbvZj
h3w+jxMtWwp6w9ajmqSnaG8Nrg/DHXJN5/tIuDpBGElo8JnWMZB7sXL/EgW5vas7uwACPYxaHAM6
HLODz5zlktIW7p3ekFjeLOf8mNcemiNZC3i/SUd1Y5xs5J4cMxDftoNdrqGE+lqxbQ+ElTlE1xFU
xLh7HKpcT5Cf3VZlXeKwXPld4uMQZ79Z29/7hO5nKJhNvfX662bwlQOhQn+9AsWGybeOsea5IFrA
SZ5RL01lznZ2WCfk1HucdNTGTc6ToPNh8NYseZfOR+Q/7NRfKkHmNbQhS5DMSQ342jxZaZajr7XO
NkfwIH+dLn2ZAVdd8i8lG04RGUY50AIEAQYjZHY574To32W+e8y6DdpRD+gtK22kbAuRhnkMm3iB
+lzTz6C1idC4etSc1sTvduI9kX8zD+2W3E3MupjJtLgZqIB06uJQqNQlS7V68lNxt7Wr/SMfX2Ab
8PVU44FzmZOMAjapjwMCAdGtrQfnh3a7mpsEcDzF3cA+DNQ5c0IRV4GyUiV8ktvYgvQ2o+w7Q6xG
Qy7gkrLyb/tRylFAvFs5/5sCqDlwRWmwcXCpvVxBY+JDoHFsLYAoZ6koS4IlvZ/EybsJun/we4hg
+jN0JZG1rTokaOIuYQrt8xuzy5jAq/DiGWQN+a3b9yS0VusFzjiYeZQgPNBFVJWvPS3f/+rVbH18
fMCTSyTOM7NBSDY4cXJ5lYJbjNk4dyG1sSY6WVkkh93+U2FokUXSBZdCOkjScd5Zc67UwsZSOimP
hzDUCuudmU1KAECIIBPpuY67CpzGSEF8P9aqcheOu6HtSumR2RJVvoCtqPKWs0/aBN6WpahpZ1i0
mFn3JqDWB8hDPW5NBy7Bingwq075xowxIWjQXazkCi8HLbx+RNgi7Zgf1JUgETJK4vYEz/V0mI/l
/NxFIDzqXjMlJ9GA/K0WPqNHjlk3H/gupQHQgQEXHVbXyNly06c8QeBhkQKlEyVflJuLv8/iTQDu
MrXUhLCGpkRwxtOAtUHD6sOBJRkvMtY9+jGfrmXgx1FdfsfMmvxApQWEeDR5WEkMkbrfZyikEkFW
A/G5SbeVdYbuzgd0qpHQlC9mQw2ojlrQSrVk9eeGil6JHNASya2rfhJtdde/831Zk+MLGe8HfcNW
glU9PdGA0glIsY4aZsd/xsq5IX9RLzPerD7e0ClQMv+vIN1MCNsdMH7mipqz57HkNRI3GcEw25k6
XxOnRxxtFvx9FXD47LT4zcU3zrtFioQ1lIFVgEIwMpIPVCHa0qO7EKDI8Yh0gU+BaY2rYaU9k18S
oIYFPOijJaZW3/4iVCTv4jtwMqKCoEhfvgzaip9mK9UGFCNP7IeEVbgS3q1HrUQo3BpSDlzeLIx+
WwGW5p52d5JJmRI86Zzv+HMuCkjcxB7c47KX2r/lCQUAsaErA5wmxUKdBSKN9polDc5K1RqQVzjz
LnOobregCUx9ehTcligEOhpvxw+/GsgtuQdB/lAxQbPE1UwpdTiu8F5ZX6HxTwTt37yIMVmXlDXG
eWzg9yQKPNn4xdnQk47ZlnCSNL3FG7cKtcbCblXsIk61qBjODxFpSaRlmsWBuTU2S7wegMUHdO2H
XyX8Sx+tIn9cXv+xWHeNiQS3/EiJK/l56ML4zYY67as4unl3GuFvoCYyKRLRZQ/knGOzGytHwroA
Yb8JWHn1Q5U0BErh/FvE36UcEObTsj/91z61VnE5/hsyesQCUIiKIeTf7N57ebsTsln/4fNi1arl
erx/mdaJ0TZ18wuv8OHU5mtyXFK3G62557vI2vjZIR2QyljEgaCM21wwXrayePZ265YLxypN77K8
9ky7IG6v4eXraCYWzaibk4RXkNUD0s2EDCnSkoO8tHrUUeIK7rFdvRMzuIBSC5HUgUELW5cMQJMB
BsBhc1unUkSSnDxtEJMUJTsUKmAfw+IPkCx725Y5Kk3OnKxT8pur6JfW/TKVTXHjf8Ejo1jW7XcF
RMVsSZ2jwPbDBpb75Ey5+oqIa28ebZzteqj5xTNZ0jBaYe7ohzX5+0wOikzsO7BMik0KCw1MhRNy
g7Wv/EgOSNUGuGl2J/7bqLCEFmIjmTerxyVkRjxUpPeOZXO177dOw1HKp216ziSixkB3e1Uo32jT
htTyabYfYIYjfFFdCoH5D8D/YijDMYvXDvZNDr2XClBvNvkd3wZtkvL5Tso18yhlwhLTeqmPsnvl
KilGQ1H72aVWUhNkelyjkf/77CkSjigy5HSxy1hbJWAqw1iwg1VC8S3cq/IXUqusj45zmtTj9HRU
BCRBg6DlhlqJoJWWoJ+nDybmIII+GM5VTAj2DQYp91imDX/OCOq4uYl9Nv41LhxzwKud8icVwSP5
CxpE6ezKwr/Nuvc/0QpaXlvjXX+dN1xtI3q4GAuwsQG9NnTF+JlESIi2sz+tDRmyYwhMvtRoU8aT
Wp05ZcFUdLXf+t+jKIN6kbbjx69Vxs+RI4BM/u1d1wTCi7ZOnGISjgB12Sjj15n9OknMJQlqFRZr
jfothRIEVzqV+7QIuQScRP2fn6jg3BoNQ1+UeJ3n0xVc2w4aeNj+ZNbRUEQ9qmnY+dtAMdYfF0wo
YW1ieLqDIx+yCpSv0y/tdi2JnXugeEXspn8unT0SVGRhk/738g8qnuVprjvTDKCbBGSJVIVYNoSM
xTf83FwDtp/KB7s8tDL+Sa3Wqo6ocuObE3G9XeMQTGFqcnO3Ro6Sk0SECkikCQDhKWt15WfacDlg
J3+uKtumwaF/QtyQ0TW81cPK3C2mjpFQbglhaJ9BrLtPjDEMsbEX2+of75pVtRK+Xq0pgssWYlfc
b7xD92fDLugvvRwY3o7JzWHt24cg6b7xdfyMabyu4LAb6L7oQGnXR3IBVxZtSkMaFrymrmQBX5tW
jZ/OWpzrRx9Oe8SP0RipR5IohMsPeDsJN/I5jp9yLlPXuIMMSLwSCVLOZnyTJcWmu5xZwcr9U3KR
kDeZ4U10eyygbmbum9h7uhL0toYJEZa2/CJIWO1DseoMiNq2GFS39H/33LsCcUFYoqQkilZlzZyw
jR1PsVu3TfW+ezTzFg+93POd26W9hjvKEbLEVmsw+awaAAEqD5hY5WIdJ0LhAFj/VxA3Gj2pLUR/
4Rsv8Ayz3riNwTORvtpjAhZAYyY8o3QDVMnSVn1aM2M6ZMzCygQ1pmBsZ7HzibKcmAaHrzW4uwjQ
3cJHOSw7M4ZUYdJgqnw5IfvwUZKNWxBCtGHMJehq5t7UqB+3fdksOWYcUEoqEPR8/Xo/lIV/7hPC
aKkB48AmWsJVIV97D8QfwtP0VjNECj3T9SLBY0w2x1xhGym9KobQ624xJzbD0Ma4AkYbpZ8CJL+O
7cdNm4jOZAp5y2CVcVgiRyTgdGAlgQFenk1de9cjjo5+qWAo/FDjIYTKD/TsXGxQ6byrSkZ9CVsm
QmvwV2/deQLEE8qf07bYU1dDoysxZQkFo6T5tC/COzPhWJViRLDcPdV6LFTrtdvap782nzSCss6w
ZSHQ47GgTeX7V7Cuix8xixQDant7cMQnvfZlmLw5eBxqsgLCrE3mr7x/icZ6Gh4IkrTXDTYdf4QV
DyFZDPt2dVuSrsTErFLwR0n72V/rkCV8cQEWtAivVj+gEEeFtJae3UQ782kSRu8CZnUDFkYAb+a2
k+pKUNmeCt/NP578OvR5vtOCiluo/JDcqyQRYquOPN1xhYa5dIL4xLVEnNjAvoiLUuOpFYjM65xN
JqawCzGKSh916yFbx5ZWy09JSjnw8YvWTxGIGhckqn+Tevvq1tbUKNXCIAPdx+ann5tAgBFF+9Vq
5MQ6ALuak5dWATwm2ftU0oYBJ0ZU7cAxRppX1wfiRYE4NVH/P5xTn0QGK8auO9WfjignqA/471lS
lMl9YMkIdq3JjFaD5SxTqyonrkstEp00/+UxnCus54CaVf50AD9qpnUKkKV0O4tV57kdEQi47zmd
ttpzciKsCVTpGU4E2QNkwzV54pdmqoFjhOs3X1f6fma+6YnXx4cosh2uXr/eE6jc+7/U/5x1Fkrp
K4RpzSR6Uxe9A4J/CjqfYdkkXix264Pjdngx/Q3W0NDdATwUbcdxiLymZXSaB1czdnT75Wzkq7Uf
W1z1kpxhJ2jZakxx1xGMyH+B8FeyX6e01UykZ29oGcfsK7nN/1jDmnXUZ2T4oSk0QSFVIp8V1duL
ZHXW6+s1lrx/s5B5AYp5aza1kPFT5J9b7gCo1bugaMGypXO2S99ljTqHHd//kkvw5kAhfLVSg5Jm
pcqsWiIJth4ms8XadFNkhQRuhhSBT0W074Nl34/DTYVzcNjrlE/w59ISvpjBjfL2yffpxFxfLUKz
3hjxtdMEXhtbT2TbbUYcRkdrJP/Y/zAYxHcii2uqG01NrgH7B2MucSYzPgHn/4aYJKT7ByGKX6Ah
4HmQkGA0KFWpc6nS7LLxX7lOgVkkJe6No1u2u8bjcdpJu/q03y5fQlhkSSZRcjRaaq2BQ3ZAVXPs
rqmoaKjs0gRkmTNCxR89UMZgO7XloK2BCYDtZXkW3A2rPNvBzax90fsnFhDfWYi8+1pSUOVWEasu
lIG4fG1y+Bk2srD+OewqX4EfjSJDSZ/3GkNbbZ8r1hBAVZdsr8m2yeKGDbPvIkmfUkdYrwsP4jU0
gkI5RIuIcKq05txceUXG3yIFp4NQMbmtiSpYsa9sHEe4JhoWz1elnQTRlPWggnn2mqlRF3Eo1Xsg
qdKYB+SIMu2Cd3HjZ7TLegXRFwA1qphRgbzSsSjjwsZpTciHP8yyIsRt4pfgZHnGzbV4T726yxUL
Qn2Vksf5cezXHiGnyFPWM2paE/nI3UI+wRN76+u/luvV7EM2GhauffD5NHviEUcCNdVCyJ1pgr+Z
uLKofvUNEyyi/Tu3aI3H5EwkvW6U5O5nQzFBSXAPcmu3NCa43Z71mSnGh7wkkiRJuaQFpWrLPtyP
ljAV2DioYVa2w1P3g3Xrpx4soHBXKS3fGCTwFA0qzMFsViPAwEYl+aWQ7dyGRRlNVs5ie9dNox1H
kdG5+/AceVAo8aRI8RGt4crcuKgCc4QZeBw1YJT2NYhz6VSykxQi76BWv1YpMNhO+4K+NikZhqC7
dJyDJnT9SswxPjetECA137DGtF9eT0KAOqD8e/qLreLTgjcsxztA0zfZxEABjE9cX/0yFmzCJNpo
c9m72L8zdjZA7+XTtUdK1f+mVnfa/ODYwE8XZGXM03KGgejJIa8NUjvEl4aCaajc/THYYaUmyiAM
hFdqIfh+igV76RZaxv+iImDl4pUe5VWqSBrQDWKkYnV+Q2+TmRZafuZ2EA291l0Yxu0I3QPs2uky
NSGU5AR1R86OMRrxQV4KOThAObWPZ54G2Fcc5RY2JYcwzH5vDICKdTHI+4s5Zw9oEmawCAUFv+ju
jRIRbWl7NboE/SHYh0JM8iWajrVAoExGUp6uyp1xoJ8vkEYzJ0ShKY8Y3LoxZu9F7bLsOB/HPYds
TeRBlYGXHohSHBMAlNx75kfty2W0zF8bBgOOKxz5e2m5mcNe1yY6rkLM1rHgh7FMtF7ZUM1QGJIM
T+JOoidvBx8zsuj7KwOBfLC34BPCLFNyNY4X6eEkqxCFr/R+GHbXAdIhryWC6Upad/SqKSBriT6h
ACbf63iZXNsRCxVRgT9ZqP3cHTCAIg08guQx4wdAOusMWRhcA4mGg9dwbJJJOAqL3RAEzCW8PCuJ
N/m8Sxz13J0pq4aPe16RlVb299nT8WvYD7MqprR21tL3NY9820RSbq7sUfl5bw6Ts4Ee9BSJTtwr
7W8eq9biAddXDnJDLAU89NuBbajeYXRUGMr6cSMGDzEHt22x5tGWUaTxean2OXEkOflDyMfpaAMK
KrPryDJ82wmO2a85m5lHPIYwKcfN7G4U8+GW6vd9gKjX5ZmFqrsIRZ0WVx8knxd0It5KG8d04kTt
8WUuylFX+0PlsqwEfRjq4E4ynvAP0RyJ0K51GfW2rcjbvscpNnmLKJH3oCPFrbGdFEtOoGcsO80g
HJEONXpmrw6CMv8O9Q0+QWvguQNnd3Voc8RDEDMI1kn8Q+yPsbE1LnVbN9U/5dkY5vjIEzoAHwAR
aZqkumEJQ6dyGchMQIDIIbCe8a7SOghUmIGG5/JAVnLn5QFp6ExVKq7qysst3lSJxXhiEu/MIrIB
qkTaJKHHIo+X2RjZCLmHnEumN7Oqcp4PkQBOhS0X4z5oKQULixgAlBew+ETLZTAH1O7Sqt8ztVAd
aNBpFpDbagGXLgQPjzQ0Ycl1wlwoMl2sqOJORzjWluX6gVSzzf73PwQ4CJ+WGwtjYsGagWk+BV2h
VIiAdFmQlbiz9zHKRkrXj6fYxhpuvRI6oLXBWsHaxwmX6rUG5TwoboZQMudQvYatcpfACbi9KQXu
f31UQY0K8dqek027qgIgHqKtw0fE9Ot5ovqVF/lVu/SLKLrp/LRbGtanh7c0hXF/sw2qRDT285r1
8oXl8+WKOKsDdnoziE4zHx8BlaKTbQV3l1fYyyG17tBh3t8icHcCCGMFFnykMXJ3XH/ogVn11UaO
seD9b0HsrRSZ14G2KXCCFvOQRQLjV615UNVdf1WfotvHwHRE8MQRLgqQfXKXNTLWPZFo/YG8RDTT
ys+hemjgu8rOjX6Gyvy6TUwH4iR1Ipnd+xTOd4iQIht5rT2e3sB2gmLcTA3Q2U79FQc5aAx1ReSf
ps2ZmkEyWAKfUjr+EwgfFXRYJ6+aOzT+6OZapAOacq/H+JDmVVQakOCdVtd5jdk0g0xbUy+eMo96
gaQDw1MSea3gENvLDbyUl3ogEkUfI73n9YeZ4y6dNZVSkz6Zi/Dr9KxnC3NPblu1aN5XjbyCTF+7
ajPBbWItw+5K3YTd/MKuK5NL4bfIWi4azv6IhTV7kc8O9kesS8Sv+uN4k9og3CvEVjSLegnHIW7k
gcawUz88WnWZ8Sk8RcOZBthKFGbp5Jooz8JFHiC3nUTH5Gl+pcRZklVc+817uCKRcfKaUYo0VV2j
r9UHSydj4HGPK8GKJu1xHnqfrAaiiUC9m6OWgXmP2lKVzPmvocjZ7oZW91+a6lEv3etzvTkdjpW8
PWEYlKhzzfjuVULvCcc7D7fifIrKhInpbiYOuVDEU7p3UtSfUgiPSwJNA1rXmNBfUKm4Onl/Cn0N
bVVoO57t3ua1SY0QPczUpKvDDBW/j6jXt/m8U9Gt851q9hs6Egdf90tlTwK+xV6azBSrlMf8q9G9
Lk/0cVk5S35N6IDiRA85AzNxtBcsVpIvvGvRtVHdAe/GyUGDmNfdqcYQq/LchbBT70H5KhYoEFsh
/WgWwymBUroPlbua6olhgD2achyFHdyE8TrNrf5yrNLKJOEdNpPLhBXVlBKTi3cBWmCAvshQKjsf
WIzuZYd5d3h37dVvHYAmILd/3pEqBQhUDj451gQdwnts2PIKW+xjsVRmzNi5lVWPF4p2GVMQ7XP/
Xf7VEDWDVfO9ypY8iZabNI3gySTEvceJwz7+FJF3anu7foWuBbP3lXlN7Ves/mh3e+UOjploSAEY
a95AT3H2zJIvYA5RC8glzNjJYAMJ0pRGyTFxLnjJTewJGCyv+n1BynvB9GnTYBvdaJU6F5q1YZ0R
flTN/nRZg6ZcPOMZqkI3KM3L3+qogQln9F2uPC6bDRmbArKpGkH75Zixf/lldMmWwsSJGrti9Vz4
EP2vl8/uqqlXIwVH92hi8brsFs4SMOXx9WNcNtYOI+80Z3bbDWtZfFGuorxFkHgxGseEFPcej2NR
zhYJMFHO7xi2IqjvXVFdNv6aSNtEElZbOMA2yU+iEDJEpflJrQG6nLK6AXShoNQyFe+itoTxk4ff
cQ2+fYKDhfd9VHW/zQ4Y1Rhiuwm5K/y6/MSJkdHfMrDkPJu/Alxu8GF3wXsZyqDFasioW5lsvuqh
OYsZKu4nLmeDR7RF2peS+9XsNCWcGOJUaOgJJ5n+ubViQ+DepcTGYxW/df86V0Fg559RLCQOnL3Q
uF5lVKqopXyP2n+3q1bCNIxkR0p3NysTqD9miP3DPjZrTQgpiV+bKZqHNVrZZ5znAPxteJ6sOYrr
ahYEjmr2BGRDxu3iadRCdQOJ7fg9YhLFzyie+joxVZm59HcMK80UC18tIgS0bLRiiLoGZEJ4TSg9
UyghqJ0z2S2nIxfr1Y32wVMkPvHtVpNWA/NiL5qzAQoKEEhdLVgInAAYdC6fX+TqQG7cecl2g1Hh
6DIXm/v/v6d6m/+hsJnR+3C96gg7yxjc/4k8XUtr5vgjOSt8VxpbsY4H5jANEf3cFMs5bajJdErj
bQTKx4oqARggBwwXj1WppUfuz8r3MboXz2tdjXxHVIK1GA88eCdLHBXt5EFRTSpIGgmEqfs02CQb
XncqzHbCdG6IM8OYCNTyat0UrliWnLnyWknxMB/1paNGSAymzMHhmO+izmUSGA309l0Ni9D3yMfJ
a1eSpgHPLgHeAB/+DARWsUOo3IC1WVNcUhDJDCUN/dL+8GkfHqWfyJ2R1tVsGG8Xfok85jtvYdE0
SjbdR53yvtPT3jFUHgq74WutwFJb0z0u8kZdg3FQTX0pDTVIpaIcN2jUClPPj0ssb5RcXLD0MOH0
x69Igar6iW+WJIWRBVix6/sUThpwbsFXbzJ2HChk/Sw/hhgzkAaVWfV3JF1OZDUupdBHe9pziHX+
ONlBzebHSVG2x5JieivPHo9G/CYlRgSl/PNE3gzmR/E5cYUXZg7NTT8hzZMgKydy8fPWxPPJDLha
+P0ryGmi/7ynNG3cz1xGgmvl25eig15JA3IDilIKZ+njM+7Zi0zwGDW799ENx7FXeDmCu4b1IjZE
oYBws94wm6gOTXJRSv8dQOHVGbSHnA+T6BmE//BmbFXk9L5Wdv2Sx+ovpj5Oi/ac92Igwt/Krw52
BbtJzD1Z10feHClH6+edBO5DyrW0wAFa3vZGrInwKvilcJdoyflaaUgBVua9sEk75IWDGlp0qJAK
RtmBbKN62VOXQ62Mhx6c2CKcpCyNKMXLHfAcpAgspRJ9AygvsrFxQzPMFr5UnxhbYHBr4cXNAv88
eWPaJQsr4i74i1MJHHUCrPSN4VQnAoSCwIGcNN801PNOyY6ZVGsb75uMvL9rXDQmVjLv1cZaKwAR
SrLQ9jM1rjYanCkvqG3i9hBZRqNyaRP+ygHxzh+raSLZr1E35eejkYyQj9lmhxIQtjKTX18Ds5RY
JSp0KiTkvmpSN3WNWg89U2leZM/eFZbnp/LEA6UsjU4ALb9qeM9Z5X5uKEYEYuY//dxraJ9TGj6a
QqiFeONZUunZ6a2nIp90AOc/YgoXeLMqSuKATDyt2+cqe9leIEhR9Foefg92tl7/2anfT7qa+lm+
j/o+H6QgbIKr5ZWQrDBHMUs5UEVGqt51QJecsF3HykBYLGoZwD94FJie0wnwlC4ULlMPO08dfhGw
ucM/y9hRujS601widNMLvs+RCqN3I3aL3emgxXEs5fJILpi4kpl+ZbOlfN0MyilkTgsgT7yyfO7l
QRD9IsDd6sCRER+8SOuYyHORXbVo0PQk2AFc39C38yvIV0/ybNw+hjoMXcVGtW52ZddZ1U+CbbDi
UHP4xInsRSuVreeckMSnqeCk3eu06P8jqtgoz752bzJJtQUDfkUSawByOs9LEXRX2rWDTgy0VICj
gs+l6eeNhDnEfGpMVhvC4Vl2v9pxuRVLmZOiGnuXlOOAhQK9o1u4wa7hQXTil0TB3g1AICKJ90xn
pCsOLxlWjtXqMyOpsjZypzhEPtRn+ghkS2gwVmZM7rFg7xWr224BXoL4M9DlrNaRTFy+WeRH5UhS
q+UieTFbpiy09CC2B3AfnwVglYABniZ4vPAoHkj6EAGuw+xwcF38JgJubQ3qesRgO2tWO0FZdBxj
rahC1DUe4L9whyl8kNxB51L7Q8FROf5oGIEnFWPL5O7KvLbZbvJ8pvxKvW4f2SkLL9A6t0oIVPXc
r8XJgAgly5Gvt6POVBF1xF8ITdGu+JLjjovkbh5Nx7b2CfhO7S2VtW7HRJ1lXEZyKxtQl5gi4RjU
BlB22j6cIOgApxnrOoltQPZmrWgddK2MqHVzlUs9kmjvMVE4xpUK8KJc/MZBtRzz/b2UeHv87g9x
5K2Dm4UhOPACEdoCXHYZC7zSxOQ+mTR/p59ppa3gP+2vb3s5YxP/Ve+uSN34WjnpgmMLzT1kaLTS
8o+3bzfHyaB72ZLFKmJd2cFUz7B8IFIuBiBCmjXJeyosKj3zuNtIlxKZvkAjpOM90UADjxZ7eQ7k
3VCnKPRvChxEzcFpayP9nUl8TfoeMimtShmvmkCnDwL0RVxOLUApWcofT8Qt1hQr+n5zHynIA0/2
apBl4EBPIis76oBmbThLuOi47FIUYX3DGhrwfKXsWjuKVFzN71s7CZf1T7CDki7UPJZ1IL07W83G
K/TXD/rUnaH7/EBqyaI1PFn8HfeaOn8k2reJ2DOCa5g8PjBMZL9iVonBbtZaNHf5x13GMrZ9C8c+
FRY5LJqRFsEuXPjtsjLYbWWfKB5QlDJSs/yEL8JZ3mxqez30CW2+woMVtgPXyIZIO3oa8r82X3L2
2wXo6GNwr4+ipDLjAgbyXCvGkz8zkr+R803UcQfRyrTFZ8LZZUIbaQIa7UIOqSHiirSazRotZRcO
um4d+YyjQu41grqt0ZVh5lXtSv/vhgReQNnFeIjiD7RbdGkkiJ5rG7rOmWz+p6U79tlkcAoA2RYb
FsW+JlS5d3d6V2Tk2TjubO37WyeceycGbZVt27oQ152S+4taIXMJoLXScUidWwjgw4cgD3HWPZJt
ZENX6Ca3VGxh+WuqQe8x0ZDnVJMsLcIzj9X/wRTQ8pF7ubhaH/Z0j23BG1o3h/7bvPJSVU1Z/Sdp
QqFt4LTjysG8C5NIAhHySlq6TnpvLgpMdzvGpLGdr1SFpl1p6qilpzrzT6lPemTFelAja6ZTI9Q7
z6Ifmdv4JTUJtr9kQku9p+e0BBAq6uIps7dERJJp8GaeoODCn3PEqVMw84qOOsMWuPMBNp5qyJRR
L88nTkl9ueGvCxT8ScHDFLKHShZydLU7b4u/gtqG6qh9NPxEnrxztDDR1PWwAVUh88fqiNIH6f/P
CO5s/vFlb5KhveJwEtUdzWQ/TXgk36jnbhG0ywf11RZRKaF3FGNbyNFri/pd7Cjw4Flim8kgGMxH
R+qMQcbjvn5GEENQ1HMN34lmhWc1zbZ2bACxrUqZudXksdkpyFZqTLaKyV2+iN5TANgVPwlMik0V
SMfboviUsuctNO7BcMik2b1BpF6+MA/yyUGi9vfQT6omwZ+EObPYMaBrSSm+VMRD0JkLgjDTxWMQ
MQPocL3JteFlA5AbcAFJEoKlPSR3aSHZ8hcBAs7YcQU89HEIEg163uwtJhK7T4AZXqmV0J6WrVSt
m1RswzaDU7CrqC+/WK/K/WJfqR5QzPeX4x7Y8FbM/FZPH0LMCz9Wd82jecLKO3gA+06UMYzwXD9X
CLJvA0HYboJRNAu7JxD1sjxrtPhtrnVKP21Ii9OIK+AtNoth+EvlPwm7fdTmoIyUmVEdL6sYo2om
Q+yDrySvvd7+sDvVwapUMStLtKp+T4GWSqrQ25Kn+IvqMIauX3VvM3I41r43oUOQa2lruRDjUiSi
3Ow1XthDDKNQ/+u51JsI+FmiwOYMXFRBu/bIPltMENmfqNYDX0amSh7GrvNmis7vr4e73cjAwyGa
RXhtlhjxJk6gTxpet2yKwCvrq1zwMTcbOaXBaX7La3zfwWarmxNdt+Uhjg6ORw/2Ja0OUv8LQkED
mWvkAnbJyvs2eEyO+og2P0hTKisw5shVyadxg77vrfVDu6VLNaTWLERTarwE01C9pGnKarj+UhoW
N9ZhLvPvEImQjUAhEi3ssnhw0BMsnZ/S+fDVZebvR992lFPa/0XKVJMWanqrWpIKEtmPW7ICXEAk
rAeJs0Z5MlV8nomMI5Eump5h/JwR6yjou0aQH2p95mqObpSIZ49c2ApWsBn9INq11op5v//s9qEB
zrU5MbUOxfiIpgcVsbE9k0ZV+NZ6xINhD3uQYEx7caYaghkQOwnNbwxxnURTVYIV0gTCPpZKlZfW
aDnqunvudtk9j/K1O8XcvOuNpQDwJTw0pMJY0xCelWSIwLnZM1fJ5ARDkm3J920/Ly3HG+rhMfES
fm5gNLRdXpF221BJDZg+QLyCAu2t/4qUVThvTFmQpMr9FDbVdsdAMcDSITs5jWUXaQzhCvJqPEkb
Oqrhey542QVE+tCn9SO0JiK32TEck9Nh0tDwQwloUKpBcsjsw324WnI2LXeNi1mEUe7r7GIkIHqm
1YZ8Txn59qmSRrPwumGLkFddgQHNcFTzptTT4+FXHqq0FyV2fUca28SNjjNpVZ1Dubvt6SRd4S5/
aCUfDyZBk69B780oEZ4Y6p5JdCkLIFEmLTryuvFjQpLXyIUPI+6OZOb8oeEwPT3K09QlLFpaMn3t
nWjFWKODEGxXEMUQ0yLKy8kTHhWvtSogEjFxmVB6K0u+VOhKuetGaOgpIxPV8YqNvl19wPbpJ+db
0rJyVO21bW5P1C71Qi/xtAYSuTSMTj6BaJPKuG8r+GRCWfwOGieprsrRnKLvmhzjtgiCn5Vkznfx
a0FRtTO6PmAwci1nubtktv04uEH0WsANWlICV3d5jJ3ln5rzijNwZz84rPcFZXCG1B9l6li9CKl7
13v3KdESvDC7YQDLhd9al43Ewqafdt8DdDSGgzOzUahKd2AV1M7EtXDEQI8Xz/JgqtG+yYfzdAG9
gGcYkIXWQFmQtinEgEw1klpju0sw2hviT9fPQRp+xGNkhn2OFtV9yRN3tdIB3APaxXtfHMerh62T
XSt52sagxpqCHDDS9Xdm4dGkxxFMJhhhDgHWGVXTf496E6+TuVWfpIw1BEgl07D7jgSAb0u6pUjI
V0kejQ7XVHcCZGobgXwzwylO1Rppa10pYRcwwlWw4EMKpEtifTKMfploHBzk1I9wRNSOq+TWoROE
qw0CLVRu0oT6SdC5pnQIa+WJ2VsUXifbTYdXiNUPUvAWjschW5P/SkkyYAKrvpCWvM1EwUuY6End
oBut+qwwerzk1V9wNU1QluuKohl5PJAzNVtZfz9bxWhx2KcNs1AjsxQtqo2fVY78apEc3llLq1sU
3sgw3skKOAANPSN7/ba4PEiRijotoLmaExS+cqeUFfOwmzynvKbfg/S1hyCKoH93/z0vIo1pAzMO
IfefSNrLl8wNzQImMIATmALx1ql4r84e+sIzNN4xBx5qX9lpxp9nVw92d8jAQs/Ck8rxeQa0Px8x
kHEl44QAIHKnxqVdBCIrRqVWtAfi8vDyQJ9c0vWC5znANkuRAV4+UBU9cysg9g+fRbrjzfAiTwB9
Jywz6POss0JJYtJuoaQ419xe18m0EuRwpxv0JfHhNlwbfbYZD6Tlmj9YMUXPNS1Z0TESw+mA/0IX
UspgWxcvbS8kF4X6kodDXXWFbdTNI+GgXpPKs1+2QR4djuCwgOoWFtVbDB2KtuZmU3/kEa+V/tbR
JxcNCKq2KeVB80eyBbyZL2CQpZnvdUDUkLOi5Aq5oNElLFj2AWex6+96IT13e5bat9ewtipMq5F3
lEXmz4TDRIMMN1LkOBPtHQVW+z0wvTxPnWYbi6mUl/9R4nqkA86u2+rk81fsxNp4wTjSRzv0o35D
vGJ9TXhs91yPgOeWLrjDU6y/E4S/M941cPUBNsYY1ZrTvotshOQTqMQ1B+XhrqWK2bnGPGFRr7CG
8N9ZDeRMDZeFjhvH8StkJoQ9vtFRcdCA1gsnEOql6Gj8Pkl2AFD1ZbnFSNsyVmQwk9bfQBBfRR5b
uc7esV65N4b7SOjEeXYHaTgLyzGOLH5t6xwFLykX1yMxp5JMST9HDWU47VZmbMUdCmcYVcmIxsUq
eNKWG0qmEnaNjsJYh9byoC8rHil4YxLtWfnj13Pd5hvP5lEO9LJ5BFvb6vpIdNuohzqrmCuau0uN
NNC09JS9M1q9U/o2vz6WIX8oj7+O80tyYcX6Q8MLq14VPOHzjoHzsbGcBEXzLvwDWvhIA2aq/nNk
d9QT9TzLnAYWtDrIdy1V4NtXcH2NFy+FF+evNkqhpXAI4oMHhzx772QiOz3AsKWnSOwxZNM1dyU+
CKEmrm+JrViy8xF1KLNc2HFbo5dXa09f8BlCXuM91buYSeaoQYm45C2HR+cZyrRZYBkppdH2amtJ
lJ4Y2HOLs4Cn+/RPjS/GORzyhGXlnoBZT7INIRrC8j8ZXhB10SRdwB7ZsAKioHwJdGGEKaeUYUE5
itP58Py4YjfrX702LG80mOIxihZhk0ZLOVoa2b8ZGHKlk/Seo1kThTSAdtD74N465uyLdmQYEVLn
b3BK0+VtVSeFwIIX+lwoG0S1+wEKCuOy4DPo/QzOc7PRoHDUkrerUqhaCmqB2zKBTv+JeCO7BxfI
e0jmX/0oPDUOycSOx2myo0eZKlfCvB5lItDV+KJKvhTjUuDV3fGUYzCANCnhvpmJw1xXH5tGLFqJ
749G3/525WiFWZTZRMNR0SWarVfsZlffUTS/SaRA6baEnMImsPaPPU9LbkiEchyqmiLhDuQijEQ4
TSXDC9/mxJ9kZ/sx5zsafoCSd26NtNpWsOyJJTXCGfdj2qQZxN2Z0rHjAiUibEJ937Qo4EGGUro9
zZdb6MbxNoeEt3g/DpRx3DW3TGL1N57pqQDG+XTEZsCDRE6+RTA4nxEhgwQ/VcoLtrE+kvwQKFIR
NRjab07f1pTUdkrcEpQOm8U0N8pNGoNQFvk4+SXTbsmQLFnxPAjgLTGIOabfF5bWerl6a6GuGPhe
pVHjAEhDdLGao3mRcW2ioe/DriDqN2Pw1vjnrhBm7aKHh2oqmSfqnbM4lc3c5cSaKdwGsgLO/dOn
G+qR7e64lxqFr/YpHHRu8LJtAp9071fx5ormkFU7PnLJJkAReRX0QBLKX9if2caMuIdIUEP7x0JU
MFLbNsq8YliBTNN8tufvRtji5DVRGBCKEn6W7N7mHZZEysCIQ0N1Xmrg9DeON1psQWjVmwJMDLdC
CGDh68ujU5bNqEKrMPWH/vW67HqkPWwAslWPg0YGWozmVKxwvb2eswtaZpZP+Aifbg6jdJWAlbjn
0dxjkFWNDR68Z42ymfBbSTfRKA8vhG4dyrITOO2UZ9zmb20b+2LJoM3fnvfu3UkB7Eeev7bqPh0t
EEz4uaOT8iiHrNExTK5ofLe/OFVT4dn5qaqLtwB1Ss8SuVJVmZju+KS7J9eFFGvwMu68LEOb+0zK
vdWm7+URuX/Yq+Im1jwykg3SLZhoc53VqnZvNQVzQNcTKSAOK+ppLktGZ4rGhLZL/k9lypSiRzxr
Mo6kot1RdzthxwZWNXaUykeMSUR8MtY1CFNBdYun4cAsFRDQtxVa3JJM7zMGMgtrWcABhDbPskH7
MbNXbdKF+YLgZqo+3dYKOgavTear8nICxK9QqkKh0LkJgfkDi2PK7RNwAJCRpqhejK2wDuxYlzUf
L+1Lff/qbwpUL9Yp3Fba3OmkminOi4uZ9Gf4oSy/JQvBVwSKWIXT47dH8zl29+YsAItnvaCpz31b
do5pmpuG/HQJDKWGKCSdc9jk+XtzIcr0GRMrJGhpooHs3BjygKsJi3605D6fJ5Wc8fGim0AI8X17
4OWuaL/+QdKsvESNANUU72wQjovQSLfAmvL1y43jdnLaSUM5hqdvcLFjY5CsurHaYebBXO8Xmg1P
CLFBHOeO3Yvs3hN0H1nSOA4AZF4q3+G6fU1iJRxmQU/eF3g3TeH64+iejar4X+mbFeLvsbKcMo01
RfkTb/2uqZhKZUntcuzHM3okpWNJL5NUh4h32vdXSTvumtat05sfPgqiWVcRoX0Ii2dvpxq1Fp5N
K8Fa8W4Nv6mhqxpveMPEm4ZoYC1hhVc4j8ZlX5RglBPFmg+QYLm7lGermuy5Hh+oto7e6eB1QXZ2
+DoD7yyZg87jYB1r9lErny7+H19XbKLKmKiDC1KID5rPEXFcKag42ZujWYj8vK4lrkfPzS6riPxP
BtlZbq29Awzhqg+j3+HXIWSJHT0CjB17N7vf0MrfeLxb33I/strtne0Zib9KAU4acl8voVkLAVh+
X7OTjUwuAoKZMM19mVIAljdsay7YdNqa4OqShZOmqeO1VzL1nJEcbj7VqqrAdJ/bwGXHTF9A5+v2
rjvo8xKfJiN9wnQTYUMU+I8g13uCoZld6ArO7R/R2FUWg/b7hLqHhupeT3/rtpY7eayoJK0s5jt8
wYPU743kR58NLXhhooRiopBPg6UqDQJwqyRN2+XOUX9nGrz7m9DfbSNbClAUhwasKgKyn8j5zjcw
TZr7el1tWr4t9KfB4F+l7Yx43aSKrRV9rbpcDDRxOVxV2Q3869HUjB4W7d4tu+acD9JDpW9fDJHG
Xw7byA4zub2tWH9J0lSb+agfknih9FHrEOXsVdYk7X9ayhNF4GVpErv33v5edm23NOa2blxjEJ5J
5aFfonumFloelsfDkI1VNM3eZD1hdsadF7oP2HaGNFP/krjlUgYTSzk8SWh8BsXRChNCZEK8daI1
DdkdigXFqhureurCvWO7Y9MIJ1ffaKcqGBTyBDrEbeOGQC+lTmdhCUMdStLOGk61njkfQjnj0zuJ
gUfyp9YY98mI8HX+y/mfrMDg/URBQigurhW71DNjj9FM6fASCgm/PenjpU4XQZqf1ktMQ6X/NoKV
p4HwKs1qfM4jhEjk/n+feqFSSqpepjxIC82YcIGOuu3pL+yNEHNMDYob5YvwXPtgLo5Ail6+hQfl
m0nlBB7MJAcnMHVVlkNgENLbLAFD0hEI7GAvsiFmZxA240watU6J+KDjGWwp0yfHwvAMQ+O2N9Mn
49AZ8/AyB04F26h4+E800mpU9gwxRuZena5eHH0oEax41E1M00PfTaDL0fRyPedCNTDvMO22I0LD
8U4sb80zX4+4YtPD3Rjp+InMhRd+hIUIbX7r2PwwpXvKQNqahIO6BSJUl5S+Igx0mFxawh8Q7zG3
zEe0Wd8zFfSiod0T+luFyJpuuGlwJRo6CFFRZsCkKlvfi4k71NlTZfGH2px9yvEyk+lL3UcrU3q3
sPlgCxnOMAv6OJToXPmJagwUiyL1Wxro2NSPUuIr3gLEZijUX4vXkKS4WxlusNpLCH0EEbTrVVyN
7SyqFM1BxawDpTRFwuyvaB/FX5LM9gmrX2sEclHAjKEmcE3UbDlHrMMtV/da7j5e/noa9Ol5KYsU
oPP8Ad9ff264dVwnWtO04sZlOq8cRyDDDoHJwMsZylVghZe4+GXEboHPfBfIuc5bw4BQfhlFAa3i
rxjwX8H5j3Dm/QZ2K/2980JbliNHx1gpRUNK6ILcWX9BOlRmgQc/o2k0KbhzvO9LchNIBQ/TTSZ1
1MDCN4b+ESJ9DluNvpz/rXz5LeeBFyWd30i03o10psZXlM4l68TQ/u9K5Xb8MEAkmiCyP/sca1Lw
QAXSWWOnZvwNaIzupLIrZq9ptREeOp0msJvElGGhtvoggZAJREV/AdNlV5Tf/3HcwMjwpFrkxSaB
kNN6Dm3WFDp/nxN44LQRjTEg7kYJ6TJwCjGkfbPOgEu9E0mBM1i2KWRI5gHH2KjBPuzZ4fne2Z30
bi9aDdGaK8hK9bMiqk/5A7oJy7seEcDrJzl0zISNVGkyfUtgjYc4R5bC02h9lFMlvULtEXSDaIjq
5uyfgtq7u6+0dDhdb4Vt9Ch2cMovCHgp5eTRFxv4Ekkl6VgLidxXOvLxePr1rdNzub5vKkPovPMw
GnDbVOv7gMrrw/iYV2Buu6n0Gl3420/20CQ2PnBrp/DkU7YWMwX1pjVsuHEB2kDsxukkQsWCXdgf
hJ6A4mJUbgJi2KFTqZnW9dNdyG5lF3SOHk9VmSK4p1G3L/jJpkajCfjn9wJlXoQmgMD8MuSdjfmn
Btgf5bCi9xw4TPOtJNmBJlKuLpeH1isSkdFF/XOhJfccLvAupn/XoARaw0ftVP3RhAebCg/v5X04
Gy9v8+XzVSo9pdykj9QqGvI/rUAAxEZcfugS5uP7kBiN96UC/LUeZc8TgqZrgYuKcy8ZB75F2436
gTDm+kH/zYRyQoI7kYyRbf0AcfaMNHew1C9v7IzuCsZJYt849xhOmF+5K0SowsN6TZEyq7jGzNab
lSBItJf/J+XnprChKgs9G28UOi4zyDtu2w8uqvXrmPg+FXFZzSU97mrvVpg9QvsP+ZD6U7tUayjz
rwWdSgmIh4puLujE8TpR4nAaoqPEpnIaPUudAk68PYf/N4UUJtp39JP1yknSp4zuPd9RMXfNNPmo
yAGAALRVW5vYEjWpN/QgtwyPb05K+kEt9hrOR7PvhbAwJR0A/sIRZoynUnWbxIfyEMs70XQ3t4XE
n+y9YowFjNjc7ohNricP5C19cY3pW+/v3ZcOXolZhb7SgupT9r6uP/JfHNO8EwQ03qusHdoPJ/7E
3V3fH6X8bNytc5wGZXuqK2RqHzouauePjzT/Px0RV/lqkTCqR0br+Lz+OP5ABlOx44IxHWPbIjua
PDJrLS5osMS7mJSC2iS3iVy2ClBTlnTTVwpk35egx9fsRLhaWghWkOu0Q7mZ3wQX/N9Se0Q0G0/L
sDKVcOdJWum5h67uC3kuryS6g7UvwLlh/vT1h2U83BmVzxlgKBzzshTa9suGOvLJsOrdc7yO2aGk
wz+Ytjcu6tMM7Il7O14A+3mIwNnPVO/3Jbom+56vJY4j7WQ2IrS1h3erBs+qjBMbrKRLaMg5aXle
++mQ0tyfFKF11hKBYqcHABNwdEGXHYpCJl8efsOEXnMenrGZCnDOPTIHI9Vb+A7CxVZB0DCfLRtL
6ZvS9mnW5D0k1ERdGbJ5eRVycnrRZlp4yoOMNxBEZmC1x1H35xeve5Hw5e3Bu2BIseKla1n50sv2
y9wbVXzGDKJ2sCid93+xbRplk7zkHmEuXZhEJZJnHX/JjJYi812+zlgbE6/DZJfszTbwa43Zbnys
2imiI3IJXGKgCVLjfSW8lQYxXgY7fe7hLrzVFIdAnqbG+a2q3aKpFy25cDsgdJLemsAV1qWirTue
GUrhmPLh4EXYf/uvJG1P//TbGz/9BXD1BWw+MHor13XDncaYcA6qAzs6wFIHWIsEeibbjlHXw0tg
0qzWLZKk/nZUh9bssWo8y3CXlaB/bLF9ayOT9AxCWHVGJKCcOCfz0FmoXk4ZneyenO8PwJ9tXwFG
ypn6SqDDuxpUV4KQTCDNpEzLZ9H630g5v3T2Hvl3q/Al04iPbPy9JghLMt63jd/0cSRPbbZJfNel
R7GAHku+PLqeX45HjTPVP2c7VG6yL+kmbT0k+ij6H5tl0MGXmTCavxRW6MVjOVRahs8WrNsoaZ78
nKoG7jCHd0ffpSb3xGgelHSED1/8o9/E+xIDmOMj+4uxe3rePz7UJ2NGbogok8CK14u4MI3cOfOn
G9msbRlTp9Rn2Jstf7JE4YQTVtLzDzlDJ5MSR6QFn+YtZp//hhKgXfOuXJ4f0ShPlRyII6sT2XUi
dtG67C/aJhvMIFOhlab8VOlm7ONI8gR+fT6L8XQZRg2GBiQ8v04FmuXR2Nlk4Ky7UpmZq2JOV75P
dy4tbf1nXdNFrXbQf7ZkFnfXnJs6mvx4u8mvuMy0i6VA1P4zYHZ1yeuLFGQ/q9iCXBFbs+8PGsoD
wy1haq3CrMYAorMj2VkaCy4InydqcS+5j5Ze7plATtHCTuAVOGkLZP1na7yyk7kTaf2YC5NOxCKr
QYkIhIDf/oIzcMQpkRId5Tz9WG0HYqY28RtEgFDSzW+GxXrQ94UR1EAiY9oXIfGKyHbLiz/AHdoP
27sHPAL+4BU71Oz/H2CO2dXgqymJNvNt5jiMdR6hNZUgZWDtB6Y7DA2DUSuKcLFbnw8rO5TWKa5k
CeqhEb8OgBPxHv6SQvlu3cQwCUg7zIcemFE+52XOoYGFYtwn53FUPwp0gEVHj02lqu56Ni4G7T7s
pnp2MA2E6H8XCSgxHfG22XjUkckR4zdIEXUTekGyppdRCn5qbEBkPKPxCM/L+iUovjYEUhgZ+VfW
sSpL3up73je9tLN3+D7odt06l5Pv7hCLIT0ZZ5D7Kofe9dgr+E/iHPAjn9zM7RWKKJSjE0rVmb9R
T6edeabjvWzDL8Qa44VdyhF4gGUlZDDiIoD2nrT/vOSsMdhLPm+wTIOBCILdvsycFr0WSkDmIWlW
kTGIUkeBkwE4SxElDhpeB2smAQ1Itgrx7j4RItO4k+Eo7fok9A2gp0EdbPaf5q6T2aXQ8n7/H73W
z/9i/rEkH4ePGK2iiVrIXlSo3AoE08IpoBmlttJ82rZFepLXUbTjXt1KkrfjXr34yKf55dX4H5gf
XcOdW959DuiTpzwQGm+XTf+63/nmXKNXSXXY0UN4XAjrX0nYRtoDt06gjmtYftKEuCa+034enV5n
riuZLTrsXKe2NsGF7zL64/aWmXRF8cmrBPPEr6f4JnK3f4W73RHG75PgfsCSivjAmLOfxndg6p1t
nooqzTOfnCxwo0abYOsCnLgR+Do1aForbP7Vl7D4m/JlhJqGuEm1F55Z+7iXQx2LF7U4zpIpDdBJ
SpsAyerjxzYHfeXm0ZCE7Us8GGUCWAiNiAN8GPxCBbIcYg+ZpJh30qSBDn0Vqvnp1x4JRikajqmd
yv62WWfzTmQV75YddmgvbYLIzG/XysC0aG9PDyUL8+xQEZeSrrpvqZ+3JXME4mIzUR+UdCu7T4DR
BvwTEOXF73IQSWNLqFszTqVeeUexoB4GPqayGq2JK70sh2tFPflOxyJo03kQMIC2IVzfnnwwj8Zq
4tAj9Ea6HHxpdgIeUwuB/Ed67+Y9zbKhuMaxRntkoIPhBWUptDcL316OgTRdJBTEysb24empgaEJ
cl0UUq2VSFDbPXYj9FkNMHZ1CX/Dp169pggkhaBG5eMEotuk9neGYj+9Jvp2F31/DFWLoHW98gnf
gwfh7GwBM6T6T+SQ3hoWB3TknTst2w81+x9G5TGSy7RY6NKASKO6/XVbZFTvy878yWNV630Cw9oM
oXBGizy7GKgusJXRWCrp8iaNNUjpkDGIteWnm79Mi7hKdOFLpzw3YgzGmTFEd5RILAwSQQoARnCC
1uO6jTb1rudeeVr0L+cGaVkSo5wyLdYCt7t8OtEbzOFkijM3OBmEKsz/WpwLfT+8giUQLquYGt1+
zxLjaNiwtMie4jMwvx7u8Pv3GlZQz1/yibxMI6he9UVBp6dd0I8CF8AkDvoMKH+W109I6AgV/zMs
2ibrEKxJ622RyVFkMvYPsG/XQxnAwlFXv+4sNAxH03mf2x0thNKxv3d9hbWGpt1pJZqqyRnTl6q5
a1BT1rvZzklsEj9MAtp3vtSKUlSpbAqldeo1lf8AWJd87TEoD9VjdnZf76xABf+LVzQPMwW7dV2X
9iD8XpAentk4n/GHk/g4lrlAfEjNZDvXBePJTdUxjwp/Dy2fWkCB7UJwp8L/eJ7zJvt5Yu3Fh5r6
6UrOhAfN35qHgbO77oYbr99KyoGSenoKQHpIj12RxbyZEksajvwP4riFvU/wCHtltBpVK7hGbqB1
ljspKfW0mCrphEODDWcXWzyWbAYXMm+nbd91dIDZKNeTJ6khbr9OazBu1xf+YH3P0nwREvjUi3J5
1q2/KV+GCeml9Xyj7vEsVApOuyj7Iqq+wVA5SXRBKv1ZYLy7cBEBPR+Io9RxlgBuCRR/nwHAFIYg
6qClwRK6qqYFHSo4ERIfFFKptpvkmdQWyqbfPKazF3oskZ/5o1zXAkSqDJgEZ6oogGZ2uBQ5/KON
x45+v7mg34qyG57d+h47Zo+u9BKO5aYm9ti/0eihQMoEYMBTWdptuUWPZ5w1H0gKfri25D5u3lrl
Q3ypkE1trp8mpcIzAmA6Yb0rJvsm3yI6kw/5ZaT0+995eTAnY27AdCS2EK4cRLVfffBDacttpxvd
mSUjpwUfXGRHdb7UpXjG1hAhlkRnwq4TQPv5HSc8l8TcoNjHaeVYQ2bZbHW0HZPo6nGzmDGko4YA
aVBaqiaURwEjqOzKM0nulqspcD0gy7dUEW9SefaMEJdXWN7x903suNDSiYEPWpI+48mjB0PYWc4P
ykBRrDwzJJ6/S9An9H5X47CCTBzBNIGTYQXdp0H+v3rVszv5LiOa1EG9McqtBJEYHQMNUW3gsUt9
i1FWvjZpWLW3FdUn5FIlHYkm8g/0rH1xBJiriP3LR2zIIfA5FoUJsrDMVzvpmcmH2UY7ZE0U/qqJ
Eepz4JryG1WgOZqqBZanvjDNhZFByjn8MiEtXKjYPZyH0+pEKxAiCTwjrIdQSt0hBnaVdyMOrWFy
w+459uYvmldc2+j+dL3m1VUjZEilxm4vlYGpXVviACp4v2oMZ/uoUkrdfTQlkBw7Xn2cmJ5fpFgA
MjIQ++9kxCvhrFMGHrN2zMuQ3Cxua1PpNtvPHP4WCgMaYdJmLSb5WyxaSVrjAtAe7UBZspNjspyW
ZWQ3xHLK+qaZyQIz5QwrAygxpf12GhE2PujmCJpgSvvCcwdtINuCmWDaA5yVQgH1QMMdHaGS3suT
QsuuMa69fA2BHz0Jw2RWKIclVssTx2j7dpSJZO1ZdJJXLATs9BmYBMSrA0djVqiGHr11aUZNLGRy
CrjbWsUJrb13ePWs5SLoed9ekxx48cc2jGGy6TX9W8DNfwPSxWQdQacS85yhRKe9TVdMF4zZGAnQ
SkR7Waixr3MPp3xoabCDavIslCacz9FSc5tYrZneH5OXqMiPeMs3bGYRlDXYFxNmgOjRsaMaLkq1
YTrWQZsjuLy4uSqV0K640yjEQ6m5L91moe3hI+Y5kInhYQSk1VuGKiBibJ4c0ZvOfgAXVI89Bd4A
yvB6D5DX+nbMYMwBq5039/27RjRH7MKgFhbhgqsUzihTJubUVv0PY077lO6bodWjQBSKfcZuJIvz
eWIsi9/u/PpyiBEtfqV4wf39tTWCbpqcvbPDqsTVtUwYwZ/KVNSZ00hApAJ7wNSYI2C1Ci+A3TZ/
IvUDO9eDp8VmKNlcNKUqV20dxwXkISqd61nVvjGrfnQLr/LLiNYB063XXkzCxyb+accvcLgtSYp1
vXgTZZ3J0SCi1BARQC4luCPFn2qlJ/K0BFxH6fkIwlVNVCGpTBVAa/OZC29bXPE8Ebmj4icLDJrV
WWIjR5OJSDyADNki4PFAPQ8nBIRDqZg2sxKwh505SvG6xepW/n9XMExCZ2M+1O7VLv5+HlWAwo/F
Unng/WfAt150P+wvKzko/sH7x/mj07bKp4t4afriiyio0mJpOwHqSC8J5s1DRhBTBftQPLNDW34s
qPCf5qn1VmolK1eABUX2n4ppP9Sa6E9avjAEmbVPgttyov0fVgrOToXuGLqSD2dOyVUSAQH/v4Xu
T5N8TYttwI/DRQ9ZW3nTAUhhp8YxaWqGND6mQs44TQ1RnU+x94aPd8FEg603/ty11mvr6rxxe4zX
RuKY7+wBoUdenvMknP3oCE+nkgWNJ83X2tLI7bMorO4f2nrOTfdt5HmFBu5V/gb1vE7PfzVU0H7n
M3pGjDmU+btfhvs9se3I/iOizI30SzWWkn1ejZRrN7PZOgPTwAuf1dEHVGLZecBGNPc/qGNd6o/K
D2tIBjMjJW11hd2IGHurE+PsNmbtIQQJfu4iEbcWBEDQbMhlhizTzNYkK2oSbiy73aCk68qKwcpf
jrOoOQmrEC1RHo9mUM7m6m32hFpSBfv9e7FmizbG0q08mTauw8Cw10jvUF9+IdyR+paeo3Bushsa
4tkoB/w2Y5soAJFJX+wW3fwE1cBAiApCxruaQxZuhZDxylg34zefv+ORmu5Mv1YUjfyfKmuQspTi
XLr9aCEm0JHomnC18iE+jeOfeBpNs4Q45tr/RlgP7xuRGjLNMt0XnYp5seLo2JKAKD3yPblXes7s
g510Z8yAbzzfZRCGuv3K0dJaAzBClt58zh76TYZGZenhqjKwg4ze89osTceUqc8w0+oITEYJag7m
9PifPj/DXVZ6zWOsi7WIVjupRxPpdgJPabOEP1LCIMDoMYitsGeasjUNv1iA9PDS7NpwDL+FT1zX
YpZgiRCXA+5bGSRwMMkvT1pdjFvKlyBXEOPyO6Lxg1Oa6oEojC8TWpP7kXpDHCGrIcMUYnTYzlmw
NI3rPdjFF4LToZV2Nnf0fTXizWWrVcWiMBgRGC3edXPVOfQ9/guUq3QjhWiov760zSptc8za5djv
hq5KP93cQNs1wYVND1PP8Jg3Nm8lpYqAde4wrDg7ISUEP5F79MsObkMqEqW38cWFdZmm1y97xBWI
2LDKzCjpODpDT/0M7FqkhN7gZC2q4tFC15VX5UdHxy3z9bn1yrfOAUw952J5So03d/KC9VRCcdWc
p+4vtWek770W52FvB4H3/zGBZBC8bkuCs5iDSJMnz02BFWkVJMp6K0eumxJtxH/+KEMH0FwhR4CK
zWpsfmnx6b6rufUkv2F9z6nZdiTCb/hKXWvP126KmvRqyTc5D5TxRq14sB9qpY2E9e69om21IFmH
FyFXsmp4i6dnb0Mv+lj4m4TH/w9YJRyIeWbXvO9vBiz7etJh6IEIID3k7SkICO3t32QQ1cCAS1Cr
tFUEV/l/SyilD5vkyYXwIh4gRJpVuR+PXRn2UxOZQWsSDk8ysJd5CCZlYs966ivEa24G8IMVik+l
Od/vKu2bbBzUxYv2dpLy1Cv9fS+2WFpoQ7aRC59q/RR6HlmGEGve0a6ZMkUniWdm84FXsggRiP2G
3FQRQOLQ0ZWket3ZFO+upU1YlEev6Vnu0Eh+B4iGQy3y9Q4J+WhGQZC6URwY27qXx0AfmKeiNTVx
EF6wW4dLK46NV7nuO13m9W/x9JUvNK26kWRcawuwKWidAhIrM/n7Czu3JnyOcryCdRlxe7qRxErj
LjauP5V3NK9baUNUriUglh+NVSH4gwjhPuFrmLJRA/iOLNpfKF5Do1SfWlHcCLgbyK24hI0QXsko
tlz3/XMJSS5Wpc1OYSFJUZHi4AgstA1/06eO4XV07c0/o66Gniv//65ceERZ5UqIFIfbODYAbdup
FgyrHzCbFoOX0RwzST0joi36eQbTmdwHBN5YIIvRYPBNA97AvFPT8m7oGF5TBJ7aCz8TBzQnnmnI
RoaxdqGxDY6XnEyBr7kpSHMq4j8OcODH3+x5yIsCIgETY1Ba0oOXYGPCKfP4JFQJOGvHn9MBejLr
UZkeWhGGJPthWCgUX3btMyBjyBZR+w+mli0mPosQ/ejsHeAJYZTj/rky0qQQVQm/Tjn7JFqLFx3P
xpqtb0QLE5mnIftQMvgcwQcfM2TtvEBjZPt3bc1SiDyMUNizWr23eos7lupM8qxYEGFDcqYq6jTq
8h9Kcx6HCudOHeY6ITd6LDNfKvdM6OrDEv9H4jb46yiNjyTwp2zZufJN0VvVxsnJ6uVtXTKHT74L
dOZ/cCD+FvL+E0EBB6Si+JWK577qXr/Vn1VV4kOpyEWe4s9XTopuPUjiFVvvLnSsp5nKA8abRluC
fEY7XaTVfU1yfOWqE9XuVjEQNvQuturoiW92eDXFp/08Bl+FQNrMd8vs6gZYmVB4jHs48Fg9Ri7r
ET31mhHzgF90g7ze01EQCAr89PU2+eOHPIbn0J0ye7O4FbKXv4kVAnEClXLBuVHzepqzVS2xPMk1
1nUdWqgifvH/zl/+mMGBwmMeZDFsMYIKPBIXLjMOUq/sG/5uCUyLpnhBpGDstnA8aC841sCbt9oD
gL+G/4FAiWHHA/sYa+yBa248vLehbTkFaWl4YJq/S4TOKg4SubHKgsazWx2+9MQjYCv++3xUktsF
9Iul1CjaUHJNLURNT/2zvOhDoZl2mDio0E8Bx6xlnmPhCdh4WrvzdE+PXw/MdKGinmTEwEPBNm1Q
tv92E30rjHPTFDCvAtGhcLaL541zj3dNJcio9no3bLpHVFvbx1D6PQB7pczkp4KmzGnJxvc79MP9
RU527p70anuCrO9cMUgNztsgBRsA66zWPDLhLHj2VmnO+Wgv0jDjE3miygAxGRsh+0CT+DqIwBBa
G3TCUvkvG6JTMR5jJaHPcIRqBHwDdSLBa/l2Cn2WNH0PAKC+Fq5LCvkYiqnCD37SRxutQWebW2zb
oxgyz1lYmdPiFwZoLM4AhWON+u9zqk1zcAEnsmwI7udnre+k8qdSXxgw9XTVvlNnDo6ZxrN+GIIf
N43aSw0ZxlfD/SA0nixjWOYoP4koUVRXIBLc9sVEAdJ6QKazHL4uQUNsE/jeJTZu8DhWuHTcB3AB
9vY9TpT3cle0/644bL0lY4utNrbr571/yjk+O3vzK8DdJDuIzqMD9jKidCTVbijW5gHD7DHl1pA2
A2wOgpKq9KuA3DMv3WbdILeVHWkxY/xypPcN8Eir9uJW1C4EiWalU7Q/pRyCRt/QC7GD4PhqQ9Pa
luDXcRf9+3RFMa1g8FU06vTBJmEXOql+vQqv53p14t3m1nXgWsHAre7ssdodZR5qv6/O+SciZEYO
4aQ0REtSpV8OB6Iu4Y682LgtUMubP8yMVTs7gNEHrK0rECNseBQUITglWOxEqnkj//bvz1OyX/ie
smLGhCL+RQ1vbnk8UvlSYB8a5PR3AnMYt6EvvllMjAII+p6vq4wzlqeQD90OrDxgFv3/727ZplQQ
7SKPEsAPaLd3YSgrgePYEvtj8FXXeRAP/Y1fbb1h39nwpBYEq2etsEAaLAbQU7qQotGwsDSUI1JY
rX+4khN8Zf89AtpmdVJSF3dpmFomWIW/HUfAFUZcjgBpuIyUAeX8W/OMIITmV3g7Is5s4UdCgY9g
Qf2xPkOzEQOxQYDkVl6sNbiQVvwtRz/LxjMVKO2NOzZa40z9q9l7BOByIy8UyuC+nP8lmmyCJ6RQ
kxod5bSLp4JiCccTSeMozm5Kkg+alrj1PHpV1jfrQwgNeHF/xe7qelmvGypCfzCg1E3JLZw8y89d
BbrbTlrx7cozDNEa6xzzNs5RBhDvULkoCbnsxZCcoj9WUYWFLJFdkkVvBkEoKxVBBh0iYutnJzGm
57520RvJbo7g+UDMyRFb72sVTspmBI7QFs/f9qrmZuepxJ1fkEfYaWkaZI0VxmRzH+pafH3evMhZ
Vsg9eASeWwRugm12tEfuy3VRhCmYFkwiQaezcILf8RAhhDfgySWowMj/kNJhhxNi2xnKJTU1aG4o
nFeTBBwvmw7v44A5bxK3wx136Ss3oC7AcbMJzmXJ0chlotoeatWOoMcnR2H4nrfHa5UODxBxLm3i
f4A1XXX+m8V//SBRcpPwEKQrX4bG7qRHpHFTqa2zGELuJKxMDboaB+3pp/hx3luBtp5C621i8zQf
Juno8u4l0WwfRDoK7uviCjZxLP/Pq2d70pS3MoM7eD/1jrGNefwoFj7UrOuIERvmsU8TZJmOhWCL
FLBpMLQBzjVhGClRsbLpC5an1ySQBv2Z4tRxXYjs5D4fjxKxuDCtYUl7nZsVAkLXFN+ySNwQlxpo
pUEA9D/ZNI1fA26CLnBch5qvPE2Tf/mTJJXBDVE3b6oPcV50JotxEyzTnUsEGJKTTWGZ7l8d0S8t
rNq+GvEQDfxe+h8tj7mNsWW1FliATxOSQdpF/k2LgxQR/mHGxrF+x/Ov5VrDkjQK+Fq20ArP382p
LVsYDYZLG5ztZbcU7sy2PgdChbmELTKK1zIcAKI0v/4KOb/XXwhCiExFiUkUkZrU+q5LDvJtRFMA
EpNdlOZ9R6/Tq34smFgfQ1CvuOOtNjbXJnx2fGpmk8dnf55oLj2LmK3w4OpgbxGXgzE/V3po7BMy
I/LsZehe8bJ1v+fQcWLVom/QOo109OievhJDtqM98dWObiPa6VtD9uQQghKvbs+K6TPbgcCfGy+2
5OQO19xGenRbvFKAMTnnD3eKguAmm6v1W6HEraAmxN10OZ7ZPdnFEL/T6j4GYrbeums4zSWV8Bd8
O+YzAjnakMbu5wQDdjdDikqfikfKhv+n8J0Gt+TUM5RrzMo+hFFGBM8epaPnz+De10SIPwROdPpo
5s8aO6V1is27rZQmoN5coR0jQYoye6M779aZaquPMlxBUPA38Unm4BGwprJ3//T4LWjMBilOXaDs
BEJygP/IdaeitCiT5Z9aCOPaCoA6UE2IDYZinfD19aO4O9cZKIYYU3vhEpmnGhitSIK1BzfmDgAt
wAuCPP0LXank3TPR3SjVxr0Jd0iYhKsW+pu2K3y5O9F46ExeiCMnniJ9YrhSX7WoLZQJ2E1udWXv
IJjRWsEwJREPOulAmOko5YJoeIalbUn0P3N0Td34+S9B7OzrknymGO0pTSR5g0i3N+VPqewbg1Om
cSZXWAVeqrSpHuWDRte4INIvXKbDLfI+cxH3O/ofW1DVCdHBGcvItXPN9WfTgAJfUdvoKELDWQZK
miT8UyNRzzFCh+Un3n0/+s0hTf/C13sZRffmHU5aBji8TNGFOUzB5wHABDFM6F8YBnC1OQT9HE3l
kISdTWNERrrly8cqfZKnkzPPA4N2HuBQK5C/JMvNEzJy0HyH4+TIXdIIStdC/AkgvEo7hXRSBxAr
T8HBcyMICAul55WQSzQ8PSuIVb2ET6YjyVaN7/yoaGWreXBEhkJhVdLwQ8CIniRWYMrIZlCnIZ+H
WXGsIL9rA9ofVBTug6zHt+8fJaXSqEDlxC1a+zv6unvGF/tn8t9TJs/Vc2gng1FKeSR7C2g5PrUd
mJ7K7a/bepT9psSTOw60FmR6yb+2xUxqedVYhuVr9uY6j1eydL9xLcKCmYuVEzFhjT95dPnioELZ
xJLny4jEMx7GLHfOCISl8QXSuREy+TGFqaodiyOSnmlWy13Np/5cjKIzVN80GwnRzUQmdT33bs/J
e+3TmoLd0GjX3An/E/SvlFgJZV9IMSESKuiQq7gOyUKPaY2m1uV3zvuHQGavkVMwNXtm1oUKJzjP
x+bxf+Dkz3YeUCAZ6lQaXlb/szmmbSNWbpNNhppNPpl84GW+ka3a9azME5acNBCRR4SAbhNyg2oC
EaEg5+5Yw3po7oOg7EGweOjxJNmT9NoQ41tZXx3j+LSnmVSGq0igHeWc7zW3ACEOPB5gwrDwv5R+
ThruCVtJsBm3zc6jduncMVqKfg33zhUgbyhsNoiCFYw7HmWVq/yv6Wm+2phJ5xZs2A5XBOJPhlsQ
y1KrVAFXfePd2/8kO85NV1jjvXYGmbCnWVCMRN+vYJbByKOelTkrLAc/urf0R306omxx1COA6TYM
N9YLUbNwCaSLC7KOvOeREJAcXYfLcRA4MAOWyWQFsUjIb1rb6AAI3Tty3S1DIO8P9EoHIfy7sKxI
WXohc9nBF6pJxFOOWbhKCBQV/AClmrZJf1nnFog7QUhm/tdpLMx4m5nNZf/+TeVdtcXd9L2B36Kw
CHpNelj08fJi79CbEa+bQX8aXuSANrow+9Hm3blUMMuET9ykqTFsrnXjKcgn5pA9SGwdLh1lCIun
HqjAj5wJgcPjy//a/+uLgLlEkROJNUgwfuMOcC0Hkgh2iuimaS7FALyO6L5YstoYD6mS8mBuU78V
Wd3vXRCf+W/2eO7uFEl7Y4kb4fBRor/8UYCVriliLmTFhf2wFbS5iEIp/1y8XtPvPtA3G0MGGs8q
1YUzxQopDVqVAcGmXRqfsC/La+tp4js22vU67gibxOn11HKYXC0VVkmmmns2YfXEqGAcz7V+Ul1v
XqcAQv58wua33TDwyy0mCin81XLsei00O11oGVqMJbhF5cVfKi2hbdYMEhg6gsBIYGwlZvvBBjq5
FjwaERmqd1NyXRNtI2RT02rqH9hlf0ahjeXa8TiNCYEGPob/kDuyzZ59zfdjp+LvdCcdzpcR8HPu
d6Shy+v3QWsbpmF6zKPpPidWLd+ZTnwg5XcrhUoh45jQ3FNCusCRVypLAVi+r8Mpj4IVCeFIdYlb
BY4ajGzCAL1B+4JLwezYgK/h3U7e2C/F7eFLtYgvibPRvJqyhrswe0Wj1OJMr9LQPbswDYhFFfJl
/d1h7LeN2b6uefgINrrL4FcZPRqpEqrwBGiHVlOXQNGIrskQ4XTTHkSWW6Vgddq6XwwgOxlU6pdO
MzYUC15BGg+9zUzNVPpzGBQJWcph9v4q9P7Fl6gOCil3Ch++oWMsMXH+eVrNyiBSNu4TqlnBRsh2
ZgCFTE54nV+7ndPV9vZMEZrnYZJxX6otN2lH+4RA32DvZBeSON6gr5x48o6FaHvDKnpcj1KYr6S4
5zfD6t2z5tbnSLfKZxOd7UeBXtHgzik0QEj6POheLQTxcxTcuepy/iPXTZ8sHjNY+1azPZgxSN6G
muTr7V+lyxbz2djZtrgfOicB6f/SAQZa2HOV8zyjyXU4wzJGZTF6HwUvzq4p1+rQhiQeyIfUpWZU
R2orsLmf3R1PnnctEU5vqzMs8CmtJc6FdcZZnVctqeK8lku3/1jukrh7qtCPRMJwfCJO0+Og0n5l
pXUXNTsfwJQinr3ZFTvEDnIpMBCBxgvo9QgPudD04KD3LLEfXy0GQS3XGEoMnDkRltez4F+axsEU
HZQhOrQlaF6g05uK7mqmr/3YAyJb+qropz27wXVm4S9zmQf2ugFt8Cs707os6fIK5KNs+OlABUU7
2wGSE7tIPeC4Aoz1SgvfRIey4DU2+im4ZcuZUH3rA8C+Zlch9qAlqC7gKmSJ1Dr6RWlgMcEC0sr7
+i5amu13QAaJwxUlTJKjDZlnTOrdbqTUvUWORM5LmVVyfH0mhe/Qs4qQT7HM1MYtJdL8O1stpnit
elHECMib3u/D3YHLX5DGVDyCElOpYKgf+2k2POV+WYkG8N27P2xBwzTdBRe1vrr8jBD96gMNXaSc
FGM3lqdAfC7UkCaZ61qx9YjnpkheNTxYVPbBdhz+6II4trZAmA25hCfD4jH6DILSpBL1TNaH4O5F
fgk+vK/UridbVYnVCw9ZqLfBDArw8R2DJVKwVfbfl5lq3DtmLhNlKc2M7AktsPKMXS3lO2T/Uc8f
+ORkdOzI7DZxHntDZQDK+QuraJP4vvD1Fs7hMTAi7yuB5KcXDXBGCtYFQxQvZZN9HMKPkWm0wF+7
CI0ueZijnhnOtotrUEQHCbQ6uuBKDrsa6QcLRaEjV5mvHLxcS9Bw/1RiWFu02JCD2a2u+T7Nr1Oy
OBLYoYS5jIA8SKfaECMBaFzntJohgzo2X8s3gz/iEQqdNXLUbHiUCLfImVm9HGMARFOTnFWfnET9
wXFrEL8xGzqdNIKBSdwFfd+ULCYkluaoPLai+dgvomEg6nU3ZGRFx2ixcrtUhyphRUR/3nKOwy+e
d6ctknLsAYtsPEtoKXsmEcl3rLc8K/DoFMMbfjV4ST0FmbrZKKT2k9NYiWcD5QOpwHlCoHYU1SgC
JhE7/u3rJj/hfKanvVPThhJxPfnGXeVXN/ePx20AVhTMnC8V+Npddvex4L/Zo7pVn16at775XGEP
42voqACQrgJlOGW7Wog+eSciQOeoG54fyUm5hIpfCbv29TKXy4wID9ShMEDF/Rh25g1ZxPDhkzQn
IPmm8N5Gftk6CwVWwD6KBO7PJtej7siGsnb5AjlgQ2iPgsuQYRUYrGAAh1zp8GO4U7PA7W9LYjQY
EP2pIPCHpEUv+LelB7Vjb1U5xycq0JHBZjqRFR/hlaiQXSq+Su5nbDQu5x8TCXFwrg9By+Aa4r9d
y2l6AZDgO50qw29Hng2UqygvqJJTYytNroNBFDcA8b77LNeHoh1e7aM9WSZqyYWclvWevbllf3z7
NYFv/eyMzhXEaA708kmP0Dzws1JO08TxMwQIej7m6A511YQ54AJETEIEyhLeV7bMt0BPbsDPWuJK
WPhujlz+6J3tIZ8UnPgg7bRdOtrng5hI3gYZ8nG5W+TILqU8DiS6BQujjOp1gZHYB9ho5cmtS3KV
ISjHbd+gAaoQX7C+t53HTsgjmN7ZreUpZreyFps7vkHa1cZNpf1C55A6GNffN48aV/WTCrnmuSoG
lFcwU/Xn264wo9uzKAwihUF0oaa/W7FLTM7YG2rLLQ4Z7XJQfUqCMvt7KlIqpA43DnKE2VvhfJcq
imscTvOfLTWlK//B1dzPU/wRZnLgA4wItNqwXrazyT0AR+JuZCi4RecZA6U5lCkizOrWZV3+phWG
LnxLGABzISY+HBw6YbrRI9PFM+tc5/tIJ33rNYmwFJG3EmwEZWl7D8C/jEmrF5XDwoUktd0EUz81
tmPrH1K9dBBpIpEX3odeeMyJJzXXan3OXdpPrUi5PnvVjVWK6iE8kf4OF+hWPUj0tgexz68miSIP
tLjbbJWgCBsxBOfHMPdr9MExnhRxqBI+e6lo/Rb0FbiN0JXkqYYzovH/zrKNQHMykstg09a9iFm5
Mz/fpPoVJSzmFWmO3KHzk5urGA0BtcVF9dHAF58UrfK9P0D5WkHOMJWiMF1sOdMJYjomvNgqLDkS
R2bSY6aovhCtES5qcVVTSWJ40MsH8y9bCIcqLwYRzF+7VmnIEpvOfAzFAurIBpv3pcGtPoGYsAa6
0ml46W0n9+WuWzSC0GuB1SKyYX5u1RNmQAsEhIBWbFF6f/C45fEHfoFy1GPyh1pxnR447Tk//Fxi
ADBgDNUXTw2QYgO08JPvVHK+lz7Ye8OGvnyhFOakTC+y6NiH2NuV0BK8/4gLrREc+Q6qwvJKBhh1
pvrNT/B7c4UF4QljsifvM+i5sTEaTvrzOSy4pfmUhySLbzvV0CkGYOjBgh1cafLacVGMRjGG0SyF
zqXOnxLpeLblzBsv4o8OQqHdWiG3/wHZIMbJDq8wxJbsNaZapeiwlLDazbtOYxQbpOM3FHk8+s8I
3uVUQ/4mwoFE0WPzA79C0c4D1Q5xUBJk5e57z7f3JlqLDEoSlSrHAQ0Pjj6cpcnHc4UNefu72B9d
twJWjYupVVT56kt+vsKre37nLqEM7R/JtwuxuCLjq3gVYovLj5LCuzs8ZyzDSzx0Pe/QeUNJhrWi
rEqgY5myX704SbnZgRKjGu/Z4azJCMYrSOAUh07nejQiCgZdlKEo1fdchwOl81Dv9UGq2me5cC53
N1A6ZSLH5kGpTQqkuJnfsk6KuX4cwTLtHCaqRsRBrsl0C9f7a0jOGtu5/F9cK7N4OFy6Lm7OXr5H
ooGWVNpg57zfUtuvuj8LChEZ4mw0jwZ+DalixRPDLuCs5LEwDQXEDmxieQChFzePiKqfwncX13FB
FgVO+26ZL3JEuEY8l2pMC7xGpi4wqA+Jpol13b8eBcc4XkDWM9wRb3nfXSPyu/AMbCs/di2o5fJj
h5PZFTvidFUpKvGTN2czUcTKohw2IBFF2XIO5T0HK2djdTShWCnSHYyQCRpi1tBu/jklxK/0sPCW
Cn+tBi1VO4UmLxd3SKJAVh5BeF4ZEcp6878RiU2BKPZ9xwNlmE0yafflI7e8sSClpu1qEExZICUK
1OCRoKxsLFh0x9TUs9DptLu2SWObZG+oQgiEsRQySbFZoIVnbxqvZfZGNAV3huylT+s9MLpjWouf
CmE08AtAWVOz9olfpc0geNLscuAb3/l0Q1v10abjJSm8+j8jyI+Ym/5LDYtWH7yV8H0N78mYwvtY
yaGysZKm48r7eRYZgw9OOo1zOguhylqckTxnVLQG+/S03+nwDLnu3VNSIZu9wOJ1olfWwB8qWOnZ
8JHaXxt+bpXl76KicH6o8u0KdL2MumtLjKjfCwaMzudRUOkJdU+IrKiTVU8KXm8ovbQYKBnNRT6n
CFcAdAra7DNzOsIb900qnwSgffb7d10ayjPTImqenqInqg4zPGOxB5BO+EKk0fNqpvBT8F8jm8en
+e5QGDPC+SYajsSownwSP2ElHvBoE8lWUu8MI7HCDGmrYdLjv2YJ7dtdyOcVsSgV6fC6tNVzKUkn
UqTPZcNywqZY3OUir8T7MbPMAJMHC6nWnxalMmUVLV1G7X0Kgo/1pXnwQQWuwraC3QVOntMgMZUj
3P+/PLEeXWo61Iv17lNTpppSu34X1axRlaGIFeIyfXLVgra0eHtTyVFH7D5LAv70LxvS6W+YhiqM
2Y50NTt1zH2/ZZdF7kBW43TRMIWl8yypQroDSE9fKUV7mUaWw0hqGZSwRemK9irOGDYWhPh+P9a3
DUFTmGKbNqfLTDI6N0627Imh5K10py4ggzTf459l6xZe8ccsO/aigYrKKDuJ5MJLCMCj68E64Ymj
fH0QTMrg0f6F7qgtSkBhCXSZ6r+gnn0MElVnKDhUlxtuuHUUSeGeLdhM0ByTbMpiUF6zKJCRQIaR
s6BmGxf2DY+1mObC2e4i4zFTlax3/c0Vl8/s7XgKHJe/dTs8kfM4DG/c//Mv8uDAFu5pWTbC7FW+
D+dL07M3WPZw3jLJJFvC3uzSndMG98fDeDBqs3w0sNK1ULyV3I4Hw57lIX0+F0/gzRcclgUvO2oV
sZreUFE1Uid1aXwjPZBbjnIN8lE2jW0od2rcjqhb+Jia/ZlnJKg459ieN4WDjiCkNXdHFOJ4mfFc
nohgv2cegXhJx3XBnWWyRsrtCCZORTiMhw8YZqw+3eF+WDx5vt85CtyKwA4DQ4HQ78lsBdG5G8ad
PIBnhW+WNajdtPe6KIVxqaNZqA7qsK7Hf8ifPSGw+QCwgCsBq8lQA+LSzMyeKHygzamTlREmoRKv
wlK3qy+CMiZa0VCcqn2bullDIPRsHFROF13le1OFEDpjAD7lZRo57wUC6PSqEYCmlYkdrjwc72pr
aednsJLpLKF6OWOo7/EAth1bKH1qqtkX9m7TuPuQ8JU7P58W7B7Mr4UMuqXP61twZeUrgRWjmE5T
qsIvlI6WXw3r+Nzm/oYDK1IFipybxOUpvyupCbzbHwp3PawbBeNJDHWlB1PyWDgN76QFtQuylKJf
4daGw0fp8CjHHVRe0x0LkWKw5fKu6+Nrrb8z63Ng7F+3KBu9zW/UsLGtru+CbENvnqCHy99KfdWB
zuv9/8ruSlSTENCW2e7udgbY1Lz/b3XldB7I/y7ETm4w9Y1anZRJrK2MxDzyme9otKwG3Vbg2Pzk
4fmbQYijbLwkpzEZrbu5P6WPc6/sQ28gV88dTPauWmCEHgz+g/1JsUzVBFt4LZCxDWSYZGMimRmP
w+zRryNkEy30UeQNB+6iHMOf3N8rpH9cgjSBbvHc/exLXuZbfkrBLq7f1aXwLPtOo/bd6wLvs1NE
DF/KfaIf1xhjgwzeSLmz9anBJUpYlTR61Mt7wO1Bk+Va2tl/isK2crx6eWQYO58afrQh85ARGm+2
Z/PV7YH/TSGLwFYEQ8rWbPCZYr7K6wcleILQ86BsXg4eMnELNxNdUYO9q2NcvIG52S6H3wvhLjGM
YUCiV2V62WlTlf8khsqCGujgvWX1dLMhp2j/yecK/80Tpo5yj5B5gqo1qkAfU9xpOzxwL2L+aWVM
RL8i8omPN0L8x57qop/Oj/FJYxuEaS7yoEAZsCXalWfnLfVH871PYkkpM7Ryi7zhGGm2IvCzz2Gc
Z9zTSWOvsYRemte7u5MWykXQG0oom03YcSYjyJP35Nil+HOcvOgitjQTSTQGW8UwVfSrtRWGF8ay
Kwnli2EKlD9m+Z/mYwZRJ9pLBZOtSD/udRvrtfzi/f4Mjd6QRkwIvOah6Le8B/mZgn4L9/CPVLvr
fNJXMMSBXG0ykYfpoiBkUa+xoePJYolh8wQxC0pQB14A6xWaY0FelRfQj/yBywI/VnK5aE1GXIdV
KwuP64FRcKIQBXhMf/V/L4ScEi1LCy01cMK/1D0GXNTbqm2kn/DL3VY2OZE2POZuazRWOQ5hgfut
PilO294zScY58eW/jw70oqgT0JNYF5xonjBA+jInWF6cy7aEv+DHMkgVeX/HccDLv3UsgKNo3B7Z
DJvBnpxglu3FMhK8ZF96951uGvTIv7GcCrJESTBx4zqIcWr4PY/sxz8KXLxctW+rfNosBprmcIft
bfdauFqTCVw3iB1B93stZQDn7FPNYIAlbJL3FfLsxLo7broxBcrxRz3/huXz/QbADbWQ/OcV6P+W
kl3BRBPWIGtOxb5kTtSz7lnwA+GNPulqeKjG956EuLZ+0FQgkkjUVT3Esk0pNG54Yf/d2lA6P0yp
XfEhcB591ciGbLbIeyPwM2g2mNwv21r5n2IwH3do5wh4+tVJftWhcgD8bT8VK46XY+md+IaZSBKO
8n2Xv5UXK5vqWNL8TiAUHl0T/brDh+Ad5nXNvNfccretsTAmbOatgJfXKZGGvnwtTNt+syFiOCS/
CGGMRWkD8Rfyf38q3mcHkTaV02M2NfifqqqHU0e772GDUEldn03tntiXSnzTBQqXVKmyK7CQ1Bny
ZYzTc4djJZzsnVaA0FyKd1CdGUxavMtjhiaQboSs5/ngnW/x8cmopukCEmt8eFbfCKh+uYzYuX7D
g8amQ4vmhPLPBQemfkfA4YRcTnPW4c6Q7f6Wg7LLPoudMKg2p+LpXCzo7HftVV4cO8EibavINFjh
f3a2t+od5H7/VdBGzYm4G2vHQ1twqTLWCx72tGPbxdtg3qNQDS5XXGoh9y/egSxgonaqvilQLwg3
4IoXMuTGG+AscpiK4cQn9I/WFczGRkz4G9u42HUDOec2vpUsIGSmU2HLg4Gq3F7ljtPvabQNFEhy
oPHGX/HoGg4Jc15QLAzM5XMkEBerB6YIBMcyKgl2K99Hsa0U3aE63Xlk4ATVXYy38Vmw3hwKjGnO
DKmQq45HBJ4JNjGq3kWTNFZg9ieDWmDwCe2Q9jMgwBq97Omo/tGImoxjneCZetJiAJXK/uGBzxJy
B2gybMnzt9Wp2Q7cDqoACBlhHmRwCIeLhAC4kaUBMg1QJCT2Vu+OVXXqfr/AY+ZEQy9J/9Ct9YhE
zNItB5JCZ7s0H50VN2IRPoAFJ0ja/Iq4ilNzWKDxQQCfhnIroDSI+moSiAMXxssJliDaTXKAG3Oa
vMSgdUXePMzVTkYNCEUDjC9mTBxvGomyq2x3v33ZLLSSiBhh3KZ1RTU0A0DWi8djMSjqMNIGXGG0
QHQnJ6AbDjkOH/liD68pAI0Pbcq4D/KSqpeoeFoc1BgOTqW6NnxajEr5akTANm53M8KF3FucS5JR
gR3MxV6xtda0BrcWgESFQaU9irNBkWkMe+gM+7mGvkDTbbc092fcmpluZHC1eq2pvr2UeS5VGTcp
4XGSE+slFonWVTSDp+l3bgvrhyEuBlGxs7DTaLLJ7HfRF9csPH+CPylL3qRL2sAyGlKUPKc0T+1/
8YTEKEOOZFFCPwpGB60heChC3hgPnpitUbdPnZZYPp0I5UZ/mfsnXBEDxRlwWItrB0Xj/nftO2Eh
4hhdvlN3bLOhmBgZ3wVbRRInVdTZ85Y60BhLpDHVaj3pr04XYwjz6vA0kjhVnLuuqPQEjqTWzm89
eD7CvgNK+qy+xPYBV9h717YY8FNj6wuyMP3NtsXJle3iwEYsmpJQR4VXXN4kShFy8TZk7GRYWMto
nDMYfSQr58xay4ig3M4U5xVkZERiqWE6Muj+woUPg5O0l3WumctjLG9+DdwCjswx0IBXKbyTjqT9
9i+kiWkEymRJMyRsfmaIiGIb4CmvLaELnXdd8aAzbh6S2EuqAJ5zFSK0GM2dWy7N6y8QIPejIe5A
Lk5YUDbIo0p5sNcLycsAOPLfk/rUJP1OgTnO2CR84x4fS84b2qpmCaC+/Eh15Sn3A0QQFDoQ+Sd+
jiojtT74fJ6xPkOOTh8KYbK8Ovua8vn3A9AfTLaKU3Ffa/mMAScQDWHbip4KT7+wEVpYZ//dzKC8
DgZ/toj/WVXZUopP3cVTIjB0pH+p44rWx6WtoC3wPKOY7OGqvLt9peskxb4zbco6BgAbUZgM1gI3
Bjf2fVrYW3Upb7V0ExuCUH5TK/3loqgxFCFBFQD1X2dDJIJjZ+N387xaRykaPMpPh3YG+zBMhKML
G3BmpY4ZYvSOlvmfYrmvFaTOz1K4tR6danxR48AivB61ur2+XwlIWfX3zgojPgo0y8ePLUiv61yx
AZQksdHRgSHapRMlUYvJFUxTsk/u4sm6SN2g3cgLMQ8op8blfYzzK0GP4vZFMlvfQDkzbvPl60Uj
V5HNJ6uj0u4Gwbd3BEu9LXq0w0oD9zf9HHYVItgIfsO6zkg5/hk9TGtNnBur7ILWpTiRe3Cyu8xC
xFR3NxQk32BN61Lr/b3MzfN1QxUOZs13U8aHoJxLPmpJi/tj4wwOQHdNXyFGigvT3JaCT5R+wUbS
dyYIujnFIzlW4tYXiPCKHWtmGy1+YMbBMGuDDutQEnX4t4Zy1T6VYt5cwJEIU07eckNYQP+t7c6C
6VWaj2amWrnMrUflhWF+28SZAmOJTJ3AkJcMzlA6QQvYW5SjIaX8t6Kw5B7jH6bj0TJ1DghJnrSN
sSSl+grAcrNpGDxUf/OZfSmexd3cquC5QA871HU4lNOJbimKXNNLgbJPjIs58rGhoDfPOx/bX+WB
SYU/40muukLdpXmQ7d6FgE2pO93Qe86dqHwWFopnok7Qana4JSFnYMr1etZFSyBz8ImuTTYJLmS0
5hMVjSEgiZ0J6+gT5uLDmB3SjtAqZqLoY1M+iWkJb/PS4AmhTYgsqw7/OMFVNw9TARGiddzD2kN4
hDLuvoLnwFo46Ew9eO3XkD+HmKTw1hfBvLEmIsSYmjXM8YUMGeT1Mlf7Pms99ktMvvd0g6vudgQ5
8+b+yj/j2P4PDwVP2u84S7TGH3Fr70fn8NOX0zAoWvzBYHUtLOHPcSVOHzva0L/1hbZDs5/lospl
UM9B+mPsdll+bhkUArbdQSLBHMWGPBt3sre7Hgl/9y1+54o/ov18K7uhq0/B64iy9WJjBbsApg7B
YcJsqZcV6KXK59Q6Qb1JD379G/1vpwEj+pwzY+MNeIvcq7R83YdjDfiYVytfRpveFq0WxvrK+flh
0EuFcT/Eupyw1GVlZawHOx5+Ceds8Y8VF9T0GZzrZNhHg483EnvdqC2Rouuq0ozo0cTrESN8Eskv
0zgGt1hwrKnlrGWOMNtr87FLwxexkCZYxpSQObQKKX3TrtQYEE4Pl/Z9F+62OqezK2dbf5OGKBh4
AP8kKycm+CYygbd89CB10cU1Q5qEeNMS9hmtjg1wYZpnibS2FPKySK1WftVuWFRfyWmKzF1caT5E
3V7N2/RAm84WFEUPAETyOtJJOEOyL4E0VFwrvKmk7iPGsOWKWKy4ln8QEZkB08iNdaQkuV4tueRO
TWl9e7vZFj4oc9dxmH8cXzqR81OADo8+yiGEntr7x/3BNJUkKLfhoaJESk4Qu3fhC+ENMCz730DZ
iYElm38Z3ZLz5cbHvFuHi3qvrBLxGcW4VgfMsoNrr6UhCN5qVX/SuIxGTq9ig0N1lO5cEeAeT4cz
88yeMju35hO3MnisBExl8vDkTnXdS2gb3cY1BZStotjj+sP/z3gDM7CcnwX53E9bHV7VLiSY3bBI
S4MbJFnPS8ySxq60PFtZ8ki2SXYjlforDEMPtaE+obU/+nBhsx9gd0yJte8ssA+y4D3jjZA3GPeM
i9iBlZSmUFeH05EUYtQjjE9KD89CGO9RPZf2pFp+Q5ga+ApC+fXSMVGYzKsbPLiJVk6eLPkIuP00
l+87/QqBO55/8Z0OJXERKHxNxHx1A6C5lbUK1Ga1MhFcpaaJOplWtj1iC++O6it2Bw9d1xwxBSV4
xNRyDLY+MAoB8WE3v8foBnsYureIkJEk7Ejvt2cQGAUWWA5agVMtgr7I8yPlCf1mQR7F5+37P/dP
NiZRYbvvVJ101bI8b8G4nuBlMZ4HCVOHyWR0BzGgNkPGnYoqShfEbtnBrgrleKf6YCsjpYl0tcBj
DGv6X76dSfFNmvXYhpsIyNCGEyftcktkcC+4gwOaJsaf93n9ngqEICeeBRcY3/KRUmMradWrYGyI
apGmFwWEOXVNZDTb+svqha48jBTPrp+/SjuLgtjcvI3mOmAogG6X3wLDvXaJBpgQOZnhI1IydxXo
JGeF0pIiNscfZkPkHD3Dj+Pmifg1k3ErecHh26v9d+/Owvvwow/ZnqQFzOCi7/wbd5fvURjYTWC7
z6HpAfQ51NS3y0oEieWeVWuD3o42zbtW/xyOBCWjWRKzgrBUYQYLbNMra69WgAFMIiSaRFwyH4Jx
YnIthbuNCjZvi4ohtJXyPcKJ2+agQtwaaO7ACEnfk0PZYtFIdbDi1yGDye2l9YbQCP2aTZCTg4Gz
+c+gvmRiS8mlNW5C9/tC1E8w44foqt4LyZJdt5PFxYodXhwQ6ZkBKB7uN/pqtUpOEn804MswJbzn
0Ub5s5dsPeADZXeG//RDnVgi7wSyjCq8Vs7hLwVstejMSvz/UWNgM8Z3Ys1YqLM0/Z969++zXMNz
ZJdF21N4zFVCsW2SzJ6y2Jl3+4MTFxKLRpPM0NinNzFTU6Lt+OM5ioL5/wG/PB0yWSrFPS7xO07E
KfTYO1/830Qv2zvlILS12bkyng5Udt0yuSFGnMill+HrHcEEJpMQhA1aRwRl40joryeJEjKH4NHu
wgzTAs3DDRzh6/Eaxocirq97+artwwBZJzmNDMIJwjzYVURpJ85SILwbpl2XS2XurwYsdO9mcIFp
6FfBcBDWHDILM2K7gMSh0d9qMCQBPc8UvR4F3ky5+dJF8ZRXyJumzgWp+llrAQpaUk5GfjzxTj9d
qLBkql4a9Dz4LvIkB71Ele2XjeFAK0cJBZ45D2Xy+zsIenVhHHETIJL55Xr+UwibRJxd7Fs261+h
QHKOPDWwLNyWivnBLaPWqWFpAwQRCLrm9E8Te/YPFxZq+L/q7KZ5dZpH3cKWPMjQDjdLVAG24pXl
03LLmK3Hn8kQm8rxbHEeLkZzLgJhAxwVpC0x/GQFoTy0wse3MgVd+YzwId9jxIvx+P5xO7boN17r
HmPTe5LIKBcPBSBAqu7nv2jifg+SzKGTqXEuPqsXzgLy8P4RCXkPDzTyxOiL/l1DNqL+QxNeh8+z
tbPQemLMXhQp+Z2aHzbdKX9viuTJVzLIXLYmnzik/a8elo8LAohBxux3SZ3/Oo+Ow1PAIiYQpsYC
YznNVJpWBz+X5ByaMluEhP/ohyxMFmwhPIeVazyuxevuXt5ECLpuSrqppp+gEbKNm1bh+TLI5Ywb
d3AyMdKOmURIdgfotMFpNkqpJapJCm6hqwmODeTMVEMNyzxCW74hMbPUbwD+C9RVKRgVhvqJtF7h
tJ2lX3da1f5J+kQTu8YBUEsZ6rCJkkFy+YkGnO1y9tQHlj0uWs0ma0wlXXaULItFKfnC0b9jrbgf
HNRWF6Xvmor3hspzb7GXRQJK3QzLzzmpU73J79Hc+zvZKTxbBTZdCuLS0YXkFMVYjIfdAtn5Wyc9
n3cDF+A0/bsRwBjOmEvBHJBOuouIfucfpcJZK8/bfgP/tSU1UNrf8gycmo16y62DRn9Wnry7pteL
nlOHw/rz0ztmqSkUuyQLnM5Ci8u+bmKNom0MO/6Na2nnhh80hfLH+wA8v4vTwo0HXKKesE3CxX/i
BLLDhZTOpgAxb74PsviHij8uZ1/3aHpKSWonntW9Qq+B1pKTRqiq+ok2upYvWU5U/OCvRWl/ztKP
4lS4Czazlnfd/0/TtFYeAvc8PHeUAprZY0AqeIAWUeZM14H9EAWmf+U0aPT4UF6BJJs/uYwDUwKb
RGk/+88TtFUxx1XHC8oIEeofIeZ4Zx8mIFULFvEQ+odf/MZpoh5YlxlrIlwOvPNsiNUsCuDDmaC+
ulgPlfuAuosFKGbRhmwylxMeFITenGr3xAu1WZF+vjPpg5/AjxDZkmFEBFL+uBIe05TL7oz/GUoL
mamPNWaEDv+pdhitFtL7Y1I3eq7X/TM7AL4KdN6Ez+BKs75YmZALdMOq7HmqiGyPY3g0f5SMDVq/
Cjner62PvwEPNDU7lxwFfcFk3w3UYjXvZQjaalk5Yco/d8uy6m2Cm8tCC7qIu4a9iVuRFTIQpGm3
VDfv9k+bS1UIXA88mIYWNvzXGM19Pa8qSSl6TPHEMX5UQHgYA1QZuVk9XofYKyxOcJjlyyoqCjV1
dlqHkHCKS8ScnqIHsmLrFP+P88GsTtu8OA3QoBeww4PgaJ0523HZcZvvjwjZmCGG9cekO4vZMCNO
yihxJqVQ6Bw+GYQlH/U5zPuv6MJbJXwO7OYKDTDasaO79lRYQbzahpTLKWNzQ8FaiFoiIGNNYl3W
QHIjzTOVeNe5chcV82fgtQBc1hGbYTapYw9MEjxzyF0SwiXf0MMvPWxJxrSKcTEOfhi4HNv0VmSQ
1pfnfob4PjRKSV8Culklshvd3H+G/AYNJmLgFeu7r3sam7PsZqZDMlM0Ggbzdbeo0fki5wf8NJD1
xmU4Rj0n0itodJB3UT+5u6Eab57aqGXhsJ+Psty4P1lznV2WRcsLBr/ujm5XKurr1u3Q02qRlYwm
c1elHBqFkzaRrCIZinf1nr2URm4NcjbHUTSfMd+auN62Di7dW80xcspC17oZ6fcpgoAk1/3FYjcW
qVUqHdpEBJ0n805XLFdkR5KTwQNFJk6wZxwH8oLI5dUAko3PAqYB22wK9HUv4o/ZMGpD0DTyzXUZ
clFb8qkVB0uBLswFEvNdV7Ep6dtGEG9gjSd6AWIuCSBTps3nNs8GxXTqDOkSFAqlL9WW/0dE47ec
SrEkz9XfIbZwcVpwaq/I312j3AVKHFsbQID7debVvvZ8HiSgeZx3K40OZTpzzqnQiuECxcZZ6mwO
+0A+kLWL4VPzXXGqSq3DlJ6pEbQZOmhzBGkDmQoyY7IiYD7LqlPCrdatbR6hNZNTQblfeRl2KsC0
WX04fwhhWv656LBf69NFqN9OFPe6rmhZ8Fij/thV3dSwO2MqOe9GUpM8CFMhgC3j707YpJlet0na
CbIHhojZAAdRWsgLMGVZ+eam2MESmLLubHSUO8Lz2EE53BAnjU5pHQNXdl+B+6txz3Dd7WVm1SDP
VDlkhIwu4rsNm+evdKvUW14RvkL/ujRvLFDr24wnfrzSuzAd+EgeDcc2Zd+ICact32bFIyPclXwI
QmmK2PrKiawSGEjDl4zTNZygWuzWGzVmc7LlgCtrhd9wcubnbg3pVME9V/ltSydWL/XEiHcZdmfv
vsarul4RsxEsl7u/eATYLgkxY+rBKJN5FNTj8zh7HiD/682zRDoXX5LV+D3RIxUS7Sm6o45ekQwT
sVKB6wPmgXHApG2JAVXqpPe4BK616M9J22StTlXcMkIUKvAChwP0u/Q70I5zDwi+i+RsgC+QufeM
ut8FIoj2UvnXvWlbyO/2+hYT8/nWv4bho6Q6Ixj+vwVLPp2KipxhD2HAg3LRP/h1XomU5OtVFOtZ
Mjho672azFw1eFU3WQ8hkYZgRmrpQ1sp+buScI3DGGKzgBDpKRYCAsAvzvhZ7GDt0jFgJy6nW8N0
Vcep1aLBCrDXho8zyn5XxS0NAkTYGtaImYmCIh2g17Bl6JWFktNWWGmw+AqgEjlEqu/5GukcfL8D
V+xhi0XhzflaXP0tWCwX1/sEBMbHBRXmDNx0vLjZw7RJ9bkpDQvOL5JioJbp9GdBQwHEctUWH7HS
8ncda1DqIuNqB3QUhsvLNPrZ2PizoINyFI0bMWf5HmhY/W6tlfGz+PoQTwafLJdtLzuXZDuA8bi8
B4LtlxFWcqqaxIzyfhe0sSi9MQQWfqh53lT85jXgNvtbJlEYbD2z/g5Psc9eEIJcXkBdb+Vab+ed
ZqiD58t+Zg30tW+BC8cmqYf1ODMigoGZ4FQsjB1ZiDbi2ZxShCnin3R19Imde16N1CDludVY2Pti
5+dF96RCcN3fr/yUgC2q5kwzbPUN6lPbOtRnXb63EmMpnPvf57AJC+i+PPYSYynKt6KO7VpEu617
ozhQKnvsVdiQmlKaUSBqWeXuGhdIJPJ49VFkvNretU0oCs1wHhgdq8YibHUkoLYH017xn9WkFhev
8j9/A4AXwlObrfLWo8ga1HQYC8t42aHJXnMyWsnNs4dNHfbR4O2j2DqN9yM+l4QZtOXuVSb9ebCT
bwqdkn9XuufT0RR55MusqfZCUwXYi0aOFbRLfDc06PFWLuZ5k7dWwVkKO6USlMa5iSkxzEPxoU9d
FpUvZX0l28RyiZqOl8IMqCkGSw261zRcy63TBX+Z00t2BxU1CMUiBy4xiecIotSKXk9hl1c0IwXH
UDyev0bbYx5CS9fNXQm/IhYNBSeVkI3axOceiXLRMIynM4rojraGGAZWJ4b98EgngRhvTt8EGEb+
kZVkqn0g9+fg56xyv0EurPAeWsJRqaUdk63z9ebuv3LY68H7y3b2EPtvS6zK4rq0HI2eBkgHWjnz
zsaHzfZIYqWUSpPy11901xWo/R3W+J6kfa4qNADh5uGcxUtWfAXCdlRXP/PtbckulBHnJ9ZgZ3qb
lgHJn7zuOrVPAIqd0xaAvacm6QdO+gvyiYdYbPCt7pEocyQ+WTNwYOShVnGq+g24nzRRoeVZTw5+
+8PXHWXZUkQGpl59bP0GCBz+lT4kq7MReqKDKgFnnjpz+57p0dJ513OBBIf2bUfDCmrC5MA6vzgE
ovNq5ozHeOUMmEP8JHlYtCzbEfq66obZazv7gmltimj7L9blZY6FWBrdldlebqZtZU1024uaekw9
h1JAKi6kM/WcEldC1jgheV0JADVcbgUCQAvruM0tE0pIJWR+Z0OORlmvVhrVRP5aBS5hyUaymOd2
+T+azyefHa/yKSwr3HcK1ssAs8HwBToKF2misE5GHYRiI2IUaWwrhS9CCg8hdJbsw3dQS12KmRs6
oZTCv0tYdQYaNTORHanwNUPBMzLkPPbsBlodoU+uDLcPGctZF9MNfCSKL4qpdFmyGc14N6Seuyt/
eNf1V2HCniv/uC3Nvf7luh2Zt49HJXR7dwROZBOEAkVkFypzWPwovb84WcWP8PliKqwtd4Q7JEhw
mhWJX4CoMUSmDMDZvtQKFO3W8SgJKMki9yaIUyBtKp87eSRQoJJ2XhS14LkyJ+5rm0z/ne8wqbGi
KpWOvz+RihU3fECR1cxfOT/5YGk/pr/sC3B3l5SkdpvUhkYiflvzTMJSNMW/oymrDJCui33O0Wu2
T+U1yqeu2qr2N3+JESAq/I4MtWnh6dNIa5Y/qCT749dhBW/m3dsenbvRUShY0Z8Xqq1n2K5qyAAj
nNHOq5D3RBUJe6vescR1AtE2qgbWTKk0GkCmObJswKjMLsTg2CVsUX2yWnkwG2leOXyHNGLvRkcf
mLlqP9CZQ3rTQPrpwYuNeA1j2mBn1gH/b5FwC8R9TxME0pnG1AD42nZwqXGqKfzGrzl5Tv7TUUBG
mppwRSEw53Fsx9s5mm2KSGr9OANoI/Smbi7P9685/rwQhFBXVg8YY1+rJ7Vv8jhVBuXsC4oQ0lx2
UCgCuTDX2JfZyhEOVPhKHScNCgf7WzVz3OuIVBgASsGQnx6G+xTpIGr+V5O/8AME4/Y3h7PoXq5o
5h0wiaz/8ag9vHea9k1ejQUbR40wc6AUGcNMNpR1yUMiG6ecje3en9NzPzy/wq0rCPu+Ygz03xwM
IkcKdoWb9LNuqjrputBju2yflDnXWIzgbXnoR1teeWAxXyWYdfSWZhkb6KA0iiO9bicuDwuio0+g
cL5vuhZlJ29yvttS6BQPWEGORnaSSKYHBw/7d6cs9tQAucLkKhWu9QQ7AMabuhCaEjAv2C/91Nx4
IsrNkwFHDUdGid9GHsRWHnEyS207qCe8VSHI8NGRQAC732qQMpmLYM7A5RGunDjP7cJeTHHQ8dKE
SDSumVTaUjdvZIxzviy+lWC71Ekf/Vl0GIU22XQI2C3ZsMFdpCDI2ooZaEQy9PNdEf/ts6UZsTRa
efxvKPptQyILebHdwHvnkOkrOxCalvhQy3Ls1vU2v1whqpJGBjc5CTu4xHPAKDjUXkq0/kHRkfHz
FhTxMK6m1G6HEhNMrYNW0nfYxrMuLCqqhNLIamsnE82h2HzWHk8iBY3noKKQ1DtzT9/dHGqjV5hS
Am6eTjNEfF7JsAgoFoGEfd2DKRYMBAFw7sknZLJSGZgaExkhbSiDer+j7Wf7TOWinhMtXpZRZbuT
JOBFze8aeP+FiGXcXtDcYp00HPoWDJmZzHy2SFU4vra53FHmaJLbVYBqbBFuU1Cd3mRQmC/NxJ1z
g4Z3gAuGNAezADaA6XHAFx9HPMdSIOg44VZsQfs+7bta0aIFAZE2yFuCkE7Wc5vEjBy5HnQixMPf
soN9MDG1rUYp6hSPwmf94hEt8o4L6lt1Eo9eniYZfm3vfxVvyzQjhGFyn/Wg16+p15QHqVIl/Oqn
TUMbzhVLDFV1YMPYQ+jSTCjk4PEReQC6hAE3zxh2DSWWCEyfbmu2dEiIYrj48sDm5ypYZVQJHoBC
WMBUROLg1YQLGlKXk+eqNb2dGRgFnF/pgZGP7Er/q/RporQuaAcwLTMzGvnbIaugE0wrJuij59fv
aIbvobVPGXD/omgE/u9rD6PJShCekK1pucFn4tL9yUoyH05ZfW5dbnYDu03brKltilVpzw3SQEDm
/Oz1zMiFk3H4PJKIdxVqh3hQ7KIuQ8uTc50FgPfDO//hl2OF+D3OfNI65V5Z+rj7EG/4gOt8wnB0
Mp+M+Big6XL3sqsUKkks4YP+C2spMmAG6pncXAtHNU7SjLqoqpHA/Vx2Nd/vP03qoa4wGV6WINNv
esZ8VR1qsL8qB5JpdhXOig0EsCHpAPTI+Mh0IPOPWEXutoj06thNIvNomSN6vNUses5lI5Bv2ZV/
qPV5SP2iPeO0HT5BqmcneI03UAxnUyIRW31WjIhPBcywzaupazKiGyh6CLVjBrcssB37GtFzR1af
pow9VFFoPkXWq6w9wfq+xoLcMPioLyclR+0KkYhoPyHQMGTTSmDQVAVCdwLZmjKDOqiYEZWetYrG
pmhERB/V4J5nNSwbVTPBjQsWAgKHxKR/VvSIyjXNY3gULw7UBlQVG+IeLp6trmu/jDXeYU4ZLSF+
9NRBvLbG/W8us6OEe0llEdoTrNDzVa2AZcltt5R+9tIot4pytD2oxcJWaLaWnIeJ/UffSsaTx4zd
3CeXWC69IQSVj/EJWGEaMbrS4qfHGD1tNKdw9BqInKgo90vn0UAsDrGcqI6t8qoE3b3b9b5jPl6+
+D7A/64mKjXAvHhtHgk6gC4M8U+VyNuTVC9FEVGBX6y15pnK4zOmK3uplVYAf6XitXOeK8CnDnpi
7IA2zXmcnS8FNl97Nlc/DiDrhFOpJHCqwO76GLdyyL/hcjtdGpkKWUqNQD0XGt7x3UjrWYoCyL4d
rfK9I5TNZT9k1gyoJRuCs9Rp2ZtBfyGNiljXIqMxdor11u101NUpiyuaGJPcfe+HAC+XiS6s6DuQ
B21mN5BXxFEr5rg+UpzxBqKnxOzu/pjSBxNXgKQ6Z4G9J5jPHtCytxhpTxrLZqaZSW38SEE8IXYG
iLG3ExSJV7oVCsQPB6IyrSozwquz5bYbcz+qGcxrajpwyQlU1dV32n+eU2hRKmxB2DpMdxqHXnla
r8dP9cYw/gnm1bq15T2wIdHLRuettoxARgzEOi4MGPobyKDOSiw5qsGT3JU4f6FvkpngwedL6CGS
U95YzO48GTBqyH/wE7aTp/a0GgcGi06fGmk7jLh2FSql+VSz1qRRw1GiNHSXXyatqZfHVoxO/l+T
XwS9p16Piq1Ub1+65UhLS68mKAVv7Q6mTp+GvQEXtSSWek2dYsd4stgZEtgZQzQWDtyjTenKANJz
sAUsRJYcef5N44nvFTZbp8niWvkER8A+VSHlGZXbk5RQVhmwvdhmuOyPLPkAdsP76SdSVhnJP0tN
/ry/xmZ6kczidDhS1W8asRymYS3VfA4VffUuws9sZ4bHaJnvZ+BGSmfz41E35Ssobpv1cFMjGFFQ
6uCa8FitLddHvSBJ9/853ALfROSOxNxozSmYfa/nvf0UMQVpyrA2/sYawsxq6vR8bFWDovzTZEpq
ZAWepDbkU8L/uM8L2jXXg4/XwJsQmg7K77F6g6b4p5UA0wGTgpTgLfRdIX2icy/3UAbTdv4GZVob
2fQfeO1YJeeURl4C4UM+nfx/vmjg7nQClJwlBu8bPaqAzxJhDGIiOvKF5dchCY0mIy3ESoYoqXy/
EOi6oYRL1dN4v6geSEmg90Wz/h1s2lLhN7P/Zn9Omxn32FCqppqUQbbTeNZTSyHlUwj2xxfumfBs
In7JnUYTFJ1EXymRMHSCXwlunE7aAXw0tL6cfc5LRZvSxN8aGlL1wNTQZc/tXuxt/4amPIrxcdJz
KcQV36AvEbXRI09LA8l9CTjHKO4pYwGNDKJrVrYd6Xe5B+0I6TR1LXdBEhUCJ8U4SJUcgVKQBAPG
Zt13+JaR6muE9nE0s6EoMEb0HhvL/KCyj8O11XwHhg5nTlTnz6PcYJyZHvRc+6RQJRd8rhJKPw+m
YHFTA9cWQKxKBajBLOWYbMvCBjFcABYwnL8gMVzBuK45QE1U1QmGwZUYgeoi5fcfP5atXsS0kb8s
mm69+dAEjdEY3rOWamjdahCP/iVfH9IMOv0DA648F/jm8pDCkZtK518/lUPrU4JeAbUaEJ27DXRj
+vGsb5H7jG9BJAJhIF/vj+3Idd5440qPxolUYnbO0dI7iTcxAxFqu7BstTPUmJQO4wmnFdEL5teS
/LCs/5zm/PULBhG/Y9opEOFykKaXDx+fWWfYUDgoSom1OKVkxytpJo3KE0sXk2yeOHJUNiF1uIY+
nwEN4jr7MkO/ldPeuI35qQNmiEyDxmgn21E2s1YYba6q3SlE4u8ywm00G2OLjUlnSJCYTQpEJS71
QhiKOKs9vUP947hGGu3xsJqBy34SZQEG5z9ZxS9oO7H5mu3vaAedFxfhagXneT00PfDHjfv01FvZ
j58VpHM3fJ0H9AdZkyuMdOrVuGM821iMWhaoJVri1E/Aau4t0us5B3ilTehLVbXaR2nq/Yt5S5yQ
FZtpcHHLDUt8VENchNUX1WLTNQs7YNkGaX7tpj+KEFZP/CFLbi94k3Xd+mWTGn2j1s1ILMWt/INy
4NVfcWxjJUD6tdhGO1pGun+qwi/jhVXrXHFZsl0NgMm3H9orj0rC+dqqXyq5r4ViVdiKC2LSfrre
0zY44+LCv3eZcpQud3IFSsLFLpFm0UZpsUxZ1aX28aqEmJl4HlgzpqVqGj/xJkU+NcS2Qr7ChZqX
j1PtSkycdQYZLmd1yBySpRsrTDemxrDmPkK+/zscCsKe7DRgfMBN8e/uwC6e+6mbPQr2KH0T6d8d
D0+HaC2jMqT2wF3FSlnNMe/2CrboYXa3ynqT2FpcNN2hxG3VK4R3DbUD9W0bqfEKTJODbNT/xplL
FLZPL5iQimvUkLbpj3MUpr59MTWCYEF7l5akIIESHNYRfpUHXDbQyLW7h4StN9moGvvzUE+AQpYJ
2vQmogBXlXev6yvJ2JKfwAJQl6vXvYZv6sgCHrd49GpOJAshw7dqoiq5CwvNHy+hBED7FB+PAG19
twT1Al88MxysFU2mv/HBB75eq83EdE4iNR3fhMF1v/3ODB3zc0HesAb/5+lwnagspnIPCFOIH2Y1
90qn8NpmmBujoUnNdfsd7bFJdTy+8kvfjrTgVrAyKUav40EGqfv6Y+vwDiD4jkBSg9NWQVMpYS6t
frYVnf6Agcj4RWovtv69pjPfMMRYDZEYM1jjonttzMBKK97Skh342ulnX2x+OfTyZc9vsyMDJhZ3
o3Q+r9ERQLx/K8Qt/PrInH0hyOJTkQI6/1PuhwpmW2y3ek9ZiT8GIZdiEN8EnVRR7DCuJzP64R0/
dI/CYNYYg31VlBQ+FPhh0RbArjvjLFjfkyu32bmqDfQFd0EoerZYyOiKOn8Bvfqnq594153Df04G
QKvumOw5FXZfIZ+sgx04X+OAnhEC8tHW2+UP0HlB4KVzqy9QT2Au9ghb5x3JBcd0sLyQuQU+wXl4
DiSuoWYWbEM9dFKWrvnLfc41Q1x/jn9e+084e0byGI4VjQQE+DWtdedXIYe2BwE9G+rhg/j/y9T0
MinwFY5oOvgPq9+xZ5r64nrgllyz+ZB1ZGaJvMaG5cYxRBHULA45m0/PYBTIjuUcfO5ykNo8gT4S
jekfbzRe7raTlB32kP367o1QdcvO6pYgcSCLj5p+u5/DH4OwCsvfcQhoGWxNkB2+OJTFIqo7EpRG
1xp3ZDEcSWsM6Zc2XCq3x5KJZcjNkqTDGbtNxUaET1qxV/qxKgrKyJDyGDv8apO7sYeEpUlvbgK5
MeFry8yRjr32ttKzmGeqA3UEWySjxpEYxsXunxpzr0OsTLcO+YKoEeCQguCeYfTWaVp4Kk2drWcC
rPzUOfjrFS+gaMjxqCZQ02jxTCWCkNrguEYi/M3L1TQAMdIr5fmxciSU1K1hOz4RivmIposAQkXy
dJi+9/zhOnKegr7L0WbBmQaxx/pCiMtwlDiTaVuUaQ462L6HdTagB6hMDAftb/vbTK/sf78Wr1Pu
zIEIfLYiKDq5dI/32D87Y+/qk3goOm6tJTpYfqCZcfbFPBdLnkcZxw/BDlPhMI+4F6cB9GFGL8vW
mWPBFNcGAixk5FgB+3L2OrSWjIFo8DXFKYv55EAJlMFhqUEvaf/+02Vk9EtDndntzm03LdjAF8DH
MPLIOhjZjuy/sIDf7fsAVOihgpltMGO1Kro9FvekzMGbNHACABNv0wQxOcEWNF+m85RJrT+1nZ6h
LlORjkyQ1ow0UDW0OR82SB/8FGeeWnZ9RgoYkrpQr6t8mCsg70j8XMr/5/5n/myOMCjvCMLRplUe
XXrjboXPwyExiqKREYaW+8zAc663OJirqGV9OoWSs4pLcbn8Aw/pn0vC6GeTWd+j6KkFwwmw8A6y
MnlKeOerCRrI+vqosGCriNW4Xe1MkeuneuxtMhETIPTjhaUfRm12c7oarwPB2HZOJRYIJ585cP17
nX5mvD6HVvzjkyKIAKyINRqVxKSzTKP0byrvJcQNnDuyKHy9tMziC3UgMdzqBe1P8n2q7HI9xr8e
xcJcPjCYT3f+uXFDrCohdNDBuQOaFmNvPNCkXaTJ4er3li1aOBiDly4sK+1CiWuMWnW2pmOSptZR
oD/cknREOFjUrC7us+az2D0UoeY4HwpU5NN1KnLEYZJchX+bs74IHLiq2XWmj+ElncA9BJthrruf
/jrSFcsJKYTRuhsZia7HFUzYmEOajl2FrQitYRRZEdj9kD4XeKh+Va2ntWa3eeup/oj+LrhX7Sxx
RC64Fq6t0ePfrZPAGfv/5HIRhjSEiGytn3vpwkBk8NsfqJcE/SDOs1wIKFaX2qLR4MthqQl7IyTH
5koVoDo3fZXdwoSu9o7U4Ic4A+12NsNYHjB8ntFFRO/8Sgi1BD6hf0cv+NTcEVnatEO0gavrpWa8
U/8Si/JzkRlL3nzdkyUVYtVezqrDcy5PJg/fUbLgSRgm3FEz7RIPMvVMw8ZlLd4WYhMuWZzkBiKS
Goyux7Sot8B3NqPQHv2m56FntCfZ0RYBK+wQ7l8i8Ffrfy1PouaQG/Zs/jSbxfqZZauLnrfNxcxg
wt/SEFRaIt0JvbC27m8/6dZMQx0I1yRhDCgUvRZuzLUnuQMorzb6bm3iwVJGLxyXOIabOGj6ReKU
l+rBMtjJdEVafivwj+uECyBBfKBgL/cL0tK1kzVQk3KVOp9pg6PZFPSu5/EstGHG0hF8bBNFyWps
befu2KNCb3aHnJF8Xed+jOYyuBuomHkM+QTMbMiXQd3EpYo2Exs1W4UqBn7/a3Hop4kMZZmIFJA8
HywC0mtj82Yk/jApIMDCByYJ9vfxJYTLh6vauWgu6QDQH/nOFXvjWb2pjN2mtxT2RsaqMdOanYyC
I5FiIdokuz6DOWsx+YYoEYtZFD6nZQEmzsyTDAN6/xQ4xatQtrS5vfp7Iy1ih8wVgmEs5vu/wrfs
SX9kC7oW76DjOiaDxJ20xGzqWoBy/CQDgfVbsJLiP835q2aiD4yPTuRaqWs5N5PbWVC0nHGPwOt9
26drQLQFznVLXgx6iMZ64aCF2TOTwa23trEKZwBdhxo1z8GUGptWdC9YhpNvacEpm9yd0SKdYcel
Li6G8nunLV/byg+dIrimNjgkWcu15rr2mq9n92cd+ZBjq6s8BbwpV1mPRq8hri6Qz0lAVVMcvLEb
GHwoRPqtDOHQFbnK1gY8d30/CheOVGO/Y6eGt26YMyTsOV8L78ZA8aKs9T98VlmbVX2h8ieaW1I7
+bdvxG8PsSWKFFP9YQc6sWmmuc/DaNZrJ8SQawz/ugsVvOgyDnp/a5R6PnUJMivUkuxCuykySpA3
21an68Cyd5nU0QnDKeHtqpStxsvdgnrhVASNtouxPkG5AiJ6lFRZcS8zNCfBOF+bLUxyGoEFuwSq
wLBXE6GXtYVg0pL5mLpwUAFZgqAaJOD/Nhn+Kuv4PnrQaH4bfdqcIPgEYPSlFcfzevauyMZW7oxv
GE9q1r0EEN5j29vH2LGNhVNVgVteA7Dpye77zZ4A366fAQVXb63aSM9uF+JgYqKhKGzTSicN0II1
ZeVKhLu3NICFMLxhyCqFiXOpxtQoWbLOWpf6zTHdYuaCeSTpoNY+sAyN8R2oXIyBRRCCITlzbE7U
zmeyfz2U84DOSdYA2RJ/lRxsmIgWprF97JCr9xCMd3UXf4y9OfpxG4+hIvc+w2jJinCCJu/zRrEo
7wZUsNi/d/DB9CLlb7zYLs/u5CpDcNA4tJQtdCLuWpW3mLiMNEEuyJkCsXmtHn3z1uDDvRt8xBle
VoOs+PDBcAgU1SXkP1gwhaRiTrRkUezJ4jWkApn17TXmRBVF6p8nJHeqYAMeKjrs81NDzrjBsMxf
+bGluTjcV7NZTzVcTZdP25V0+mZD/B/KbT/Q3gTKfUCXNOg9kEvIlc8WGEM1AQ7KYfPSwhxUQPOy
2QIN8KbOkHuaEmpV/Exr/OgzFZiTFQYViDWBx9PShYeQuMLoM6U+KUVyXmwQckwqKHEcUP8c+3B2
X1KdjqMeqNHuF6PRZTwaUSD/zPpYnjqpuB1QvB6KnYbgSA0qFhJjz8mJYNXuai8DOux5DVt+O9Yx
mvQ/9hr+hZCMKzO3RDTAZVAUY654+nUoPzoOE1Z5etkxj8m+ZmUkRGG5lGCS9Mdboxx0q83qJHUt
s58OOCffTySG0cFs+vnAYT6kYdPfkoB8zrWmZJQcRq2RJfGF/3jkYRXvek9bEL9xurdqssDzjXyt
v9t9JKeS2DOEtKLtSMxD2jhIuPzp6vtTDglXVMoHwAAUH+PO0DLedUCMPT3PPmWeoftl3uFnGfUf
rnTIAoHolMBNLbrsdWYqtSmQtLeyuxPxzhLu6KDTpT/z5L6sYUHMxTwyzWIfGEGf/oLaqeM0rbev
5J48H3sAEZ3YsWBUUe4OxJGZWlPymx/645VK6JNJ2RPhEE0upImEKLMtZnk9MLHGpzqee62wloW9
BTF3F8CG3qAtvvMAQiTfIm19LXIZY6JVyMNj3db/nC96JW3L6OR/fRAJEu2OVcwJ6ydK2NIE9Bu7
emJrGWMWS6AzDyskhF7uXDALhvs3oRv3mXyep+eDtES4Iao9CtwFTK+Dp1aXCnGzc4apN6WfzZM3
ZtQ6FfRu8iJVFFTyDJ9xbPRtHcTcVuLQ5mowjXvQ+lLaVTEf3T0R6XMYXX+VwQnoSxWaKMXgahWF
n+hnMrTJrhhAz0RhGrfglalnQdz7BPMnJF4O6X9tD4I+ZotrLBrqyfrF4PKhHMDQCOqhXLcKaJhc
wZVW2duSeDopPOBzIKilO6HEY1DZPp+pBOu39K3i4DwbIVxvwE1cji7qeFy9pdGTTyhIqTINKnhm
OG6SOfqio9qNVWa+o2Ljdg6tobbofL475XuFZWB6mcALy8XL/AhA6vvX89h5ju06uxELkd/SWB0V
UWhzZoY6T55FUgH23oGDz1U2I4LaQzMaYwqYp1JXCb3keI5R/PXcXU0337uDneiXuUwRx8Ora63U
KXU44Z+tUh1jSCuJpB1auJK4oFaighIKUwGhWPubGU77NtuV2GR6LbbC/8b5sNzU/+UsLRlI8NRi
09nVVnZQbLhRE/XLkgIlprkOgTFcz3iVedD6JaPPRmjRTUyop4psz6hEsXrD8fpPte2RSH7tI7vT
MVzP+s8+ZRVPrqO6Fw9Nyx7cIIjlHq9RU54dKfJOVD4PCTQspVY9W7gFwUJFNoGP/4+jCTOffq73
qBezOxHREAoNkjrX9O+fIlEvbmRqOlbADMWlaK+dthzSge3iKN93kuOdhjTfOIxzYbA38+4NCj0R
icyspT5Vxuo8yOZ7elprkKI50hX02mAjnzu22CE+21uEqtgn+05SXIANYPIOvUbukatNEDi7oCJM
iV5N9fQoHimRS9DXaN9SSUf37ghWCwo4LXKurro+SajiY/mZW57VPCEsoH/yXA5piO5UCE32tVut
u1Cpy5yOrZ4aUB97F2hAKpSJVTJ5wVeijQ03aRE9DgjPYMKP/BeILRDp2Yz00rdOePjPMyOf3uni
8FsqMPSn6TBVLM67dBpBqmbSJbVQ+0Pcn/mgqKD3mCnP3D5x7lRyFqXlHvQLk3CkdQIzUJEUeSPI
27q7y6+XUQu1rVHyiHRK0UpLLnrfU7A43zHs5Nl8f8iWLsmwVA4ava4GZxAX6PcFykGzVoj4chVW
sjffyPcq2EzFdC/6wXNgwaL9hLtZ2MYRGX326gPcRc8x376y0W7S8yssv2zNNvedgjPa34hJVNON
G4uh6ef0UjmWu/2zi6SXR14iPOfGydjNt7tjNy35rvYtLxv5UVLal3tbkCSrK/lcgFjZMjIfr2RG
L7bvX0RQmYxxyK0Pu9SplEZfIwdzXE+7u7ss8wdPIQY91CbAbNEmnoBZa2zwkxwtbelvuPeeWM59
2wxuWlkDjID1HO/BvTUDxJ4qW+vfTELmmjvCp33Wwu4+7rbS2ndMVdMe7AXpJMnZCf7AFuicDt+l
0S4dhkI5uxf26fxf8ih3T62NKc7I2+HqszIfsKWbe2RZ43cYY2FwUBo21G/9JmdoNqUz+71z9nQR
L8eDn03MgTYb7F9UHWULtZ3PoqITz4PwFwOxoUpmWDzuK315JU4mZ3knjcsRST8yi9uK6Og3IUJe
nqxE5N/qKxbOnlxY7+q/Da8ZplU1bjRe/UbbHIYqGYZu02fvIDQQLLOLx/jm0mv3Ai745PNVZnDy
EFlUSVPlm606bz+0g82w2/M4qmIMglZ8F58F7seepHihknosgnWr5l2WkrITQEJ4GoSCnRScLbUU
+Fgd7BEjKULSI4/OuVLLcbb0Y0+wLNtGpe2BvueAnZS08bpzg3fgeWyuqWWIMXQexsUUhazbm7Qg
aZ+zVzzR4qplePdhXibnXT40xV0JX+aa1gqZZeOwOeU60kAMJPFp1CWzTYCRfBqmzj+eayF6jBxY
Vtu2RDnd+3bCnIL5+Dr+5OIt6sWD6UzqSd7GjtJfrSjRzKFRhn7lhDGlCBl72+A8o4tY1hvkHdiC
80jSFcfyI3ZNLJJJwGjQENXWMZPyZp4ep89N75GoceozZL+B90xlQuIu3Ij80iHxZkKoVmLlRsZm
sYMElKBCc6BV1Xg1EFlG/wRUNkUiPzQc+ZcJqrJ4W3SskEuUtNIg69uufWqDL+vcgxE4C6VHSfAS
EaCJSZAfUzZ1qeTU5SOWk8lIqsiFGJgPdbtiwA3uaguFln7k2UgM7WYlfrs4rPBtHlDawTryECwD
YNnr0N0inF/bwMEuKJm0bpyBIKhe1RsnxxgGI9seIju6ecJ31pIi4Ry2+I4citnZKlUROduds/ES
c0KnBLaU3Drj7fLCfc61g+1fhdDVVSzUIvbHDx+OKNbLJ52je5/b6mc9LlkLXikU4B8vyvgIgwXF
Zm6mhtXXBP8X8MXNfaed8gZCT/YRJP7ius+nBGi8hC4wJTvUmnW+pqWkui74baWtLC/AcPEHL3Y/
ukVljcQnUQtvk9tLBMCRCsf5hxQV6pP+T42EmwPgV4/jbhb4L7h1kpwFNJEfgCLjnfTWA89ilTOU
mjSOvatcl4EdpdjzGROoYz2piK4jeVdWaMs28UydmJ+zLfyV5YKTi/nOs+boV3y46L1wDH1b73IO
JV0JY4012vJ/QAxCfFGCYUMdNSZBPet+wNedpfF8ZKVsVKrCwY+QZJJKkfxhZntyGcEhDq6bWdPE
GfXSnDNrgQEWIzrjKf4pzTX2YVmAgZojDG5f25dpqMQKObQOAzyc0rVnSiPnrT0/F+l7VrxY13v3
abv4VtMBJOgExNNtYbi6XbfESyPLo13jOWyPySdHICB/8fzBdITLHAs1HA7WWfGNDugoHCNnHmGV
e5AVN5rBbHZmJ91gL2iT/GPp7xoUtuH6CJxk0A1dLyQaRDt7RK+eAmCbKBfUI78tpdF50kOQlDgJ
jij4Qh1BdDhMdKk3hQBRuLKD9Qr9EebCzHEUvXSSy8eVtfnu5MO6NSqlc03fByprDtts485b39ln
BfQLwQbB8cpGxOL7yGJuquzKkl/3I7uazWcefnJM6Ti+OBb0lX/BhfPTy90jF1s5ovYzVGra7OLh
HkOO83Czt7IglOm0LwUCIARjYqXTGN5ycVKz5n82XwNaQmrQg9sTARg30E/rjfYw76EEbf8rN+B5
VKveHRvzS606FXfU2smkglDZDf0uMaFz6gjyxFQwfqqjRUoTpRxZK2pTDV5N0gmH8GBXhkr6KZxb
usuOjAyOwHPQD1Z4IOIT2Fmk9PApNmkJZ4O/BMcd5SkXOXgVdkrdgW5A845dTBk5H77YBpO+ioRz
rMtafLig+D7jYoCHqjo0qC3f0IWQa1sB5g/df4g3N9zgab6QqctoCjdPEpk1m6z4t9spHzvhcztv
8hyWjxkWmaIHWKDSXIsjuaL8SmbTWxtmUie1nBqNNgtT0/1zkT2k1UtKMw7I8t35BH9rlHZ7UwZ4
GlW0p3eqhHcl1uqPD0WB72+O6v6uUy3xrd/LiVzy18EPQSPhRLoOhNqzy7UdpEzM8zqDC+FRKxY9
Pk+/tHxx9MeM7GZc0n4OztVIpxU1mZDNnatJI8yIpVYVpNwmtaFovDRdj68PLF/PyZB+5/Att8MN
kA3bH1zdViHnBttsqA6tZEPi9vJwva4mvRhwCgJaR+90SCL0Iu4N3lywGQflZajIl77ohKrJ5vVX
/OmyN64lPt9mY8ldXsJX+WP8FTq1dozvyfymVq/m1tR93ENfTjmCwFkHtGqTJ575YjAKDU/C6FHq
wkqeMFbOE0Qzb+JLhmcqKCsFL3NLoLJCzAfPaeiouHm7nxT1/4zcjILunSBzH/qNAnRwbOpIExS7
uEoKAYz8kMTb9dSMO708S0S0z1Cep8ZWFPYb5A40qJLa1xhINEapGVZTHiUq0pGYNynOLu82V4v1
pU4uFT3CJ00qmDVHGMBYHPojMqyI3+ZpX3sESO/oJpxbjD+yaRqpztseQJf7lgy4tVuDF9S125to
SvtSONXOKfmTLR/NKl/ucDZS7oO6oE/eFLGwY1SfFJdU2HmJNhEd7rIf4PKKTp/gJ5DQ6c4D0MWd
1onSM3IdKOdNH6Ji82L5L83Iq5xltKLcjWzMoyg1NYbfjgcdtAsnGWWAU03KqkHi/n3aTLhO9PZl
44IRY4g8j6OAVpTF/KclOyKag1Wzgf/mOtzKTBDH3fWjUuXIsOl7hkOmV+JxKT2YJzRQM+GPilmh
0oKO3wzOen5PSu6JUj1TcxgDyCU2XM+sj1UZecgcs7JCh0X2LUfbRJGrCHTYmr6+4KIqL2Af2nIZ
smS7VqJspAsxnZGbZAHJA4M+fdyJnmUhsCSQ8+LbdQ6ZjZh7GY40ylac1MoU5JOiNmW2S5NFEpcJ
mo0kM+gKxbZcjIfOHzJ2o34Xnf6OSmrMFkVBKxwkCu2OdbPqVcfi3kCrXxdHgs7h5xfrciOXOfZ1
1rzfRISAvVWU54XYUs5/Ndu76Zpr9KXkFbik7lLJegAc8ZtE7DHCKx9eoVw+T5KVQfsPTBWWCWrh
JFfLoHuDOXqzXBdkF20sFOjXAw3viKC52eXN1cZIfAPWIbrxmMoee1o8VG6VqOyI1Iyl2WcWbhYE
N/u7sEtKci1o0QYXJjypfpHPJlKq7I/zM9oQO8MsXwJG3o+mWhib4TmkZMpyBT6WkJ17k5lpwzKB
+8DYi6jhrFj1JUkJTynWomevr6CUxO1CkicakXfpeCmpH3eCCtb48EEN2nhVscuw8WUNKCE3fMIL
DbwvmbGCcqXKuE+K8dbLrRcYP8+EJBf8BrVqVJbiOKcpV0V5aWbN++Ai6iNlSy9OGwHjIuOFoJlN
3UygDHsPwKZd6DGDFjtsKSsIlWRx4tz6MpGz7bbaoley8aqV8Ko75L7jmophA6rEZAHxJ0YRbe9W
6H3KuMxtTLIbvw9hdRLxWwgrlV5Mcg9sr51V6MxRS4paCy+NFmnDHjTf2A/3KO21ab6pY6QHZREv
30rHEq6EpkO1ylVuopSYRwGDLOMQsSSlUoKkSfDk/n/l7ELbztDv4s24ocibE/uPPk1rtSkcvbbv
uHEc6KtAXa6JMhdoHK9F6ftSAn5RgZjKzTFSKMCV0h60re0gPmAxDZW6oUy4J0NScPpSvhT3V+xr
leMFF0VbBp7IvFGpL2g2UEAjCUeXR6tYZ25Cx5m7J2z8q+5flyoK/ZMaK7g6hvYvZVJCo20FJurs
ydiz+ZrlV83EbS+AZRRC3nJ33awpTGGfL6BbxNUOXIgxtejcRRUMTzeUaJWbEyiaa/2kS05NgdaS
hU9st1nwysrZXnrQsyI397nqFkP3zw+owcHEZIQlBQWvu/HYExWFmGymMTJzbMEvIppY1tVnJpta
DL2K/CJFYcc5zm7eS1/KBZmCJRg9v9K8Dnm4sBxgTlA3vbTSGBje/WBm3aklSwAEGriqDsAkvSpZ
OmSjcHZrfobEvbxDbXEUZ03PR7+dBbP/CWwM05u6EVH+VZbMVx3w4SVroD1M9Xy6IyW57r/TlaBt
VEigiFepdrQnnaz98Rkmuus2beIJoatnnyGPac+CoAUTSKy0zMavAmQ880jR8INxHN4iYlP9OW2U
HY7q3EH+i5cI/Mm5ouYGnpd9sLLDlroJYaR11hSz5UOR0HrfW5ioGm7ILU2//L+FGYhoSx3oxVPb
9dmgtB4Mh9EGdSlza0rzgiBYAQ8zRABpxivxPbKIkC9LUfm3qxt5ib8Zv3Pm1MHanc+KKr7y4kWg
0KuctJV/ymR8WlSdAbIn6SCHPqua3bLVLb0R7vxyEPtL2mMuK1DKz1FC+ozgD7JI6ND/AXBqIntc
UmqpYMa9zanBwp8GdVXXMS8DkXFrt74VWfI2iOxMd7aX50ix2vjqQnkTbECGdG2V5xR/cYkVKAEB
K+b8hcWKqsTncZqqqHCSRVpEZBS3TFkbq1j/AHCEDOQnF96STBg65yL3FZXHDcbGBZa9qJjsnzo0
mhrT131GxdKor+dozJIlSW8djpbUrSx5bFg104UEbIHgPSGtd60C9CIS0K5Vc2/DfjqZDVjdt0Dz
1VC+AyRB/+CvK40ShRPyrh48vop/9rS63/hR1jGqs0wHjMWH88ic6SsbBFcHUIIJu11Pwh9MrMfQ
bN9C4WG1OHck8YrV4w5bz5yvlNAaDDdI2AIkzz0eA8TQgybj+82VQ0JLsSAy2NHaIzSW7HnYYZ+n
cYE+N7V4vzJwGGAjsdFEUO78ho4ixeZQCTA45l0EVvUdiczlTgLgD2pMqmBGBvsnfHAX28UMYvJO
cBH4y0dbchDFr4NYulJTLS9hSOGj9u9rKFvA+x5BRK0Guav/dEAbBn7PatVG0bMkd0GQcdrG27PU
HaJMiH1CHEO/6DvJUzXGhSIhgohSuA/OYirJNSJOxpr9hEZ1tB0zKOfJacEhjfXIrHudMHh/g3bQ
zoYJVeY4uJmL97RPi4Jjgj5044HIKwL73XHaRyL5a1IuWr9f27AgYFyRTRUZRstgqwih0Q3dSSQn
oFTxmh0TIs2NAHag2ywjCO1BU/Nkxg6a0ZjdWOIyMS+evvt2YK1QbSRD1ZIiw05tE67A1h4a6SDn
pj9JPj+dkUZ+p72cVgqL08KJhJ0Xo2q6Fo9924+D6SJAWIWcycQ+H16ExvPI1Pgph2d8ZXwi4tDd
QOModt7tMc0x2+7sVhysVd7xZjY3LLaFIMvfRK99rq/GBQFPEn6ryW7fnOxkG8VgNCOlz1SFaMc9
ca6G/iNG+nxl68+6zhOUcHJyRyaO12OULb5BqRUL2L8Xo0ofPIK6WzDFhSjkWPVNW4MWDLDS5Zbl
RVm/Pl6Xecq63nfwVIQI7eeLJJltvwsVguG2eS8L561WhuldNDVCP0lxDDJDh3WrPw4y0pi3tgh0
DPWw91xmy2pkbt3HqCuhCepgdqgLCk1jrGIEh+Ch2uoiTzQ98sAfCGAOWUib+VBorfLn7zYXYr8b
6hu0PI+guTKWpR6D/dM/jhJ7WA6HFOjXt6qT04kRcX571ojr4mc2u4zzO0qmwFGEv2kx+LtMixgx
ZU7owhMgSCldJFkL9q6asB11E0obpvu4rhsLOJNaMjbxNL1sqK78SJbUKa9n/IW5TtwmgzHoCacW
eA8YT5tDbB7yuynZcDOW8EGuwUcsd4rrCP6R4PyqgwAn1siMl6qiKTUDhmanRM9czUKIsdxIYsP2
HpL6+8aGTlXiqER5w5Ip0D1urSMUfFfWQMxC24dzw7MGjQoHASOnzGGh2H8EuSu7Lgy04wX0mgup
P2EDfCw0lfdy6LV0wysdwjqC0pMVOZ2ChSyT0CMcLyGlvAQeNhPnBmw8WnJmv/rBe7gXRKROmaNs
ecmQJmhMHmnHuY+V0xOU5Aujvr5OYY+Cy4c2JG+Z/Flhs2hVKKeXeOfdhgw4jdfEYtvhL0QBeJ1L
WiqW+msp1ebCIfp4b760oC6eccT6yFrbeRvJ7eay+Ada4i5dR9eJZjiAAuBZBLsTY14WdDMrOWuS
QzAGbx42MAjGU9ar9xsNfrxgbFJlJrmJAsnjhKL8Dypmd6zWsekyasSBY/Inl3kQyoFxbII/jnyL
oP/mxCn+ktTd+x+P26rYhoIg56qootWeGRriA20URbXhjpg374qr95apYxWaUaHzXNg074MhHjL5
Cm+xqmvZHuZJ0ryXGPFbeqgLVhj7UfVbfVjUewZaOC1wBv++uN4E2afTB3Ib9HHi4AJlgKz6fQN7
HIqVNCrdacV4lnRHt1tZbl+7OPDAzedALJC0MrAIDkC77FocannOo7Xg2PVnaMH/+D8uVrwpcJDL
5AyEcFnEDAXvFzmiwCKe3LLYUtqMZp3hAvcwbO+g3DY6V/l3z22BtDsBfL982hJQQfkSSVPMYPdE
oSj20pxCnaOL9j84XzOPYfiEKxpF7CK5sEJDJuQ8uOkwzLVCVDpAgtTGxKNhoL2feaSVw6farJr8
oU7p5Hj8uy03UHyqmdmbSmo3kY7E2S5N5qo3uJ1hmbX7f5F4AW/cJF9A81SS2TxanFKIjdIhinzO
X4Db13Q+ONEqRxdprMgzpY/AcagqWVzYiKbvUezTfexiwFer5XhdccnI7uCbl8dtsjQ+DPlFQE7a
OwbNcjBO3HD8Iv6L4zQM63eowI7fFne8/mTqqJv/kcY35evBj02MtjjXkGTbcgbd8quwAvrtLcwH
IJFGuI5JYFdt1aTW1F6fx/OBj1XSkHFvz//Dq2ZZKnj2gVfG62lDdHpAMAGUySevNEOVsF+CsNVI
k470JwA5AJxGJqm4s2AjUS04LTlgtT7uS1khc+jvwRFpESomnLbxXQzKZrXv2xkqKx+3ujh0feEN
pBbx+nSAsrgcnShB2/a7EQY3fiJB1z1p2KnlSbrsy3bux4CJdgSDA53hYjNvCFm06nAmfpilgyT8
3Oi8XRRXElhUwwBxlu2HssRQd0ZjJQoBtkzj9/NBRvpYjQUAnzfLe5Wt6a+h/sjNknQKMpwlF2qY
Gw1TnFndiax7UOSe+TH7vr28o+xBT7wGB2NNJ0evBWXn3kL2snZshRQCluDxW3BK6I9sjDGi6rQX
gb7jdYspAbrdNbrYR0YjaMtSwlx2PdJbq28XRJF4NVliswTh6XOE3YLf+1uPavJDn78vQvtWGv0C
IwRO08p5/5LpW/lkNYvW7Qp/X4MREl9J8vLdhKMFvq5BNRqBScFoHsBKDoOsqKR74frxFI6rSahA
JOaSEBNpb60V8p4KJb0MjPvqrTOvuRlpdAA9Blujdj68uaW8dzIoMYj8/8h/Cb0aJ8JI8VQIjD1o
7Vp3ES88MOlE9NLZb0KU0NkW66uq2PJXTBmap8ZlBnQ1VBwVsMFWUevSAGB9zkXpXeaV9xyaSTvn
DSmAKZMuTLAER5wYDVIf7tc9oY8oJT1Hv/8vMPFHupzPIrT6NKgfrzjUM5ERgXo65Ia0ErzBFrr5
2gh5Rnb42OkTnzKDTj+6c03BrJboSpC7IiUEpxJaXkkLrDkdKhueSPh2HLKMisLGil1MbNmgzddP
dvBIofGZJIYzPA8jruWh+HFlv/4sYLOaVqly6cFZ+nmoNuBW+c5pqNWMxeiqIMNe8qgzGxnG/8Wd
9w7gaWkApknwZKiFCJAKnzOK/aJr2h+e5sjrOlyI7qynzZKUn7mxuugHojBqQR3yVqnfvBhq/ZM3
h9TIOPOAIdNIcp8jtglSHQ7tjShxmHNzDwi+FyLsI3t0qHvpNSON3GlAfEeW4fVklh1qpsguRqjF
zouG7K+PVL4y36CQzEXno4WXaN2RI71MQfKFtBFR7RkpVkEtkKU9M+KuSdNVquRlxhZcfyp9Rwut
A8ahXvIDF35aro7nxvuKiyNGDoorV8okrYYWvClTYCh+GDsfddg+LaMCSvz8GpA7U4zeouFsCWhl
9m3eygpt62zlHPEHjFZWpUZPbDdo/TSyQ828EzKNnRIeH9jLRGl527ihzpd2FOOHYV5bFtMykhHq
0mW8dpK7JYKElx/a7aJPtb1Ojogcpe4GEAgkPcDY5xDA22YtmBdxBg3x70XDr3d0LGwmDPXRnsfS
nIuDQ451h66LXsGFkXN7rCRBn4x/TaG4g9vNfohgpbWvh7Tp6COY4oMLHhuChr7rQmYE+4dyoE1L
vMjjP3LKpXHv5dwbY/FRXV4epOWkB1SsYOI3ZfBLAZNyCTIF27I7vu0xjk59BZzW1KJVn2MeR3Do
v2OAvCBVI3uCQkpL9PhvcXDS87B99Nvo/dE4CAog+XRtFq2X6mVeA7ZrsbMZIrzIoWN0/Oq33p/4
lp0vQgLIgo4oE+SgduM/fuDV+UG6SNTzXDo2TG6m+Bcq2wJKImw5X5H9hiEOA5OMC4IUSHN0I/rC
c0FhbkiF43toQDCXIGq+KAHOQt3vnbSK3DBy4HZeodSRAM4SLbXV4Qk9nEXC/RfedoduINEWt1Qg
rr3/8y36hq+kSLjzmnaOPUf6Ytph+1gCw97XBaitwC/hkx35ffmH19uHms2UXENQPIlQK9BH7tDX
ydEYnTfitTQ3NYmMGVMyHx1S4lPDhufml/bY4837/jklZvG65bjuKJDhbj9eXKQIXIA10Xkol5UC
mMomGSHS5ZndDJ//BAVpr+lu86Bp05zuxKLW4O0yphBc79CNsWJe5xts4YaGzmWvl6czmg4xn46v
9+05BOVlPfD9f6B/UH0WFwAoUi2QmuD2kFnNtoWo/ehfWFIH+T4ZSHD2tApX6DHDqs/fxvESV5Xa
OKbr25CN3iORadB8M6BO3gP6206capt+tHw4A09o+Wo2qiWjpUT0pSFY6BnqZeX7YR+1PNcMwH4p
3Zr0I5SJE9kY0Kd5G82nD38A1IJw3wt5NyljvbfplPs0cJoNDyinERp7+8TVAGzhSbi1HvFZq+x9
6+qV+DHszK5bpP2q/TcBBiEiwVR4GXbLmN+fPRc4GTsWbXW1WvO+EozVgcA7iOLDZT6i3g/Jhp+S
Rv5lCzmMWCic1GvjORYkIjLJl+Uj67JB+qt+9YAol5oz1d7JXGhzoyib1NwxNoKA1YrRPPkwC1v8
DQ3zKg1IrrpMB3jEEfXuH/S0+5FIWmdn4KR8g8ABpcaI+o3TGj4RZzrPY85G7HlrdhTRWaF3yXOM
csBlTWKhaMsN9KVGwUG7tQk6CB8jTyNstQfGB+jSnIEvTwscMtb8Gddny6lhETvPnRXmKeBmS71w
IDzpDIRgrpSscG48YSRycZuWl+UVZINbu4Mepla1sQCzvWTLHyigMwrbmrQfnd0qQuxz0qFoYEmg
AAfL/A1qTJkZOmLM0VXeInUbj6xSXe89TctYjYCo4WZqH4lfPi0SbRZ9RyfdqlLQ/StIq8RE7h0X
6J1WFh7a/4fKKgdMLUrBjSGyPevj161L4KcJJwo1o14g27EeX2kEZJ93DX3gUuUhsQU/p1CKX0K0
gzUROCMXNRo/VGFTlh3Yej0c4Jay/XDaxlq9XmXKeDnmfjlViiCZo1j8UxZwtO+odP2TAXmU/lxu
I/BbQw29aN4G+Ube7liG7EWqZ7b/U3ls1Njxlx3V6tqU1UWWswcj8dwj5Xu1rGkbeGENP+GqtZm/
yoLHh9Kjy/p1geos6C87oZCnmchhpJM3i2AklDdhkFy0uus/7aHW3p8KRsmiCt+Rx76hKjZJdIp2
YJS0kMD4AF6UiTscCuQwWReubIyMHZf0yrtUliZtyyIPSHcBu3n5+X2sFKLfS3B7/sQtMMOlk1xh
NGuT7u8+UbfNmrXz+Op5Ey3vmGE3r0bhAS0LykS+aXWcBgVCwYtZym9c7mwU4nLq5G68o25zqopb
HCAjp7hZUE90uUEgmx0vY/SHbW0mChiMMl+Fw0JCXx25y7Khxas4l62ks4GavvwhFL6NCKXlVKri
joutraYZMvQY+JpGdXhWmwy1p6d+IKRs/yX6St3+cg75d5ydDdDJxGHsfDZGZJaX5WqyAY5nyd69
nbSbh39h4SUCC5xzShjKvxjESF8KkNVSHTSmojPFNgaOyYcjpCZ5hPvDSBkiTyWNh2kfONm0RaAc
nrKq+1O9Ij1FiPjdrgpOuwkxbB5OLhIrR3Oz21K9+TMdJMpOIcPreAl5gia+e82UeHhTp8xTE0Pz
B7t08f588KPnOITWv7WOcw5HsKlMea8B/RLBiCABdZU0FrECjdN2U+ez+xvL9Rr82lr78MkmWWhv
+EPZdl8Rg8dLKxF2wvEVhf+ibj5iR4Wmh8fTHFt/iYvxP9RwjdyjsheWqcJW8cJ3wH6+S0EGjQiR
28kavPSV7vbshlG6XowIb7omxRHG7a7eLupIyVfxN4+TDzjg8O2EZn+n0Ld7aTDf1QelKfx3r24z
lQbXImqwd61/KgEsXSzcbWdOO4+D9ZDeg/NiJXCu4aeA8YeyHnY/oaCpn/Gcz33Yp2rP6oegW+D9
5UImZORETleASPvksCrPtQhu+mURluWhikzRHVw4SI+mIavjespFXuwfraWBod/F948JoAv9dJPQ
aZfOYSfA3hz5B/kLHEZnQyVoyBnyhH6Qf1WlbvkUfsDmOUwIiIXy9sjRpAXbS7cqVZCvaMg5dYoX
7wpVEJKEnkaFbGtIoFklTHKiA5v5kYHFy57FQl5lJU+Wq24YAa9wdUEW8IsdibM3hfzGc28725L2
Fp92VajAHsyC6FPGBN3oSR8tVvH6uSWsiM0n8F7dxNfVlifpj2LrGjH3q35MjIVJbxJlws+iIVR+
2OOyeyXkzx43IIK4lpQxah70uYY7tzA0GynI5BYOgo6WCbT6JPq2jRXFmYlLtVFWsH0AsVba/q+g
xPL86XbLt5QkRWqCRIsu3JM/0dwNzX6PbImVGwktdkxlxA+Ay8B3g8N0hBT3yfZ3m92GxqhycusT
UUEaTOZnTBreXr/fDfidB3E7PfVaHxOZPb5Hmn/swEklDoIqh/PRAsv81gm8KIRIpR+e76OvT/lg
QL8vkY4ietbCRFK6Si/Ypjldye8UIjos8E+Zhj9BqCj94uQE73cMH/fKCnsSoWpvtLU8uD3GgUUF
QUW96xerJfoX7j74krknpRwnZfnJqUQpTihnjqe9qUGvHXhv7/RJkpxKowynAcHmZsE+OJDHlCLt
VMzXGcWONtAjzNASq6bMVyhyaEbCZYHH+tQ9rwOjkVlGConID/jEhYnyu/rVQe1taUD6RcUzdlSB
AFu9X0AmqINrnWLqJSFkeraJ3gGcWhxeFxjdxndGBLs1uESLdkt7nl5tKJL1fRPlCS/Rogc4i38N
c52KVeBENRDTByakvIMB1loknmXQFmmxS5uMxVEI366GhcNtyAolbTSpmwaCZekOpM4xM8CNnWN0
hSUeaM3GoAcERsMeSydPqNUfwPf+sGIe268Fd3f99lVwryWcalWk6qoHw3YLB17LNSQKtc793jI7
qoief4vPLrL12byXjrIo69vz7PUMQBfVFvEcOU24CGd0I9URcQRC31YjdYWIGGMPDifJhUdGAoW7
8/pfGfoavG02OdX08BsF5u+p1YU+ZIliWu0vl9yii/v9i8vdKW7AtP2WSyzHMOaoAQSCnxwzf2VY
3eLkH4FdWLnA2JcAoToxnf3nfmC0LdbANlCzVGXsSrBwarTaWYCorv4gtXmAaaBp7GQlyQwqCZEY
dwiYhCHFiVvxrYp1vr+TuTQ+saJzAHwGf2jk3yGYZDvOGnapARFusz2b/e9eHtwN8amHvI5Db0UG
SniyY9DcsLyU4muJf9Lt1HcvQZQttCqwN2RiNz5OW+eIFIBeDD80yUf9E+rpF7GcU4mTspYp/sNI
/Nwl/OfXU6puqcdLoAsgYz+pRX8p3yGn4nJvrxevouipAdzxHtut+WWd7V1IW21AVm8AMCIl0cu4
8y4OhSbTRmPobzcZYk/VGpDrYwEnYm9A5s7MssuOCFLKdHoE6VEWSNr8oeKTXoRFWH74B6cbS0/c
CbKZ/OaRIio4w9bOsfbxHnqOVumsUSFwjyq3nfhofDEwBRn3Xerf5pTvW73qCqFJYci/G+dkFw2j
isour9z3BVS4r4LWfWvBRoHO2VPVTHJX/NzNhsFWK55oDXIbGD1FifiZx6yymFXEGgUdacz5m24Z
YgmTM5Y051k+puYx6IWItVegdZtzwQkQ7n843y0OLzYlE5QfJufZJV56U4jI6VBmwA1c5mL9PXfL
E+cSajqpW0eVBTRJvTI1ZLTZz4Sk0XGPt64pwTy1prCyLqS4bRA2J3GnV7E3sl5F4leYjoCnGlGx
auKM9ZeFVdlV+vEevBFxCx8m6GK3hfQFmmGDxzHNOwxw5x0QbF1ozxf6KmoceUW2nhjGzUBVJq77
+OL2Vw3BNR9sccWZo2ycL9a2esbwbJh08ISowy9jh6fYdQR+NaYhGJQTOdlX58o+EKQrVQt7vNSy
58GDGoz+HcfDnkeFaXTIPI9l3sUUluhQN7Fy92YPllHDrUdOrSs707lTWU1ftsOOCqpLHKzHaniS
JrluBOZxgaxKxYXozZT0ujKunlF74hGRdqHCoQXzg40XLygsKv2t8DdZHoj0K04Vx4UuylLbSArQ
5p2091f5uAQoaMto7bhwOzQgy4+3wtA2ocgzAOhp8XlwRgVBmgoiyPvlcsYFf2xBAOyMSlw2lgVi
U4e7vK9bqlAhDivHcdZyTYW6i8WPVx2sw0nlItUOyWp6TtVv9WZR4U25pHb5yLBjDuVCnM06FsIf
S5+Gd8DBIjo13SGY1CqiHEpxXwzkzhDr3Sx2locQPt8nT40yq11NtjdUh8R6M0VqchBVFHd6MFL1
CxhdgEkuaYkp7dXF9L0VKzPiikjOCM57wj6PNh0kujbZ7q0+y+haJTyyJYULafzAYguEqCX8vtQu
UcuP7QAnALfsvCG9/aHI9GSQyubLH+MFJi61hn9XthgzUJNn1wSjAiYL9i3R06ah6oN/lA6wPRnH
77fxxT9oGj1ER0D3ijWiCLPGUVHRyddiFJot5hY41uemQq7CNyOCORWdUBtUb4Yn2T7gja6RTOXS
Yzjmvdd/ggV6qL94++DrpaTFWEtzZWKoI71Nkmzdib1WGTgEt2ZCCYe8Y1Abc9Nto4nwPAq2cx1i
k2AUi79gjvvSiJdRs5K1y0Z5RWHNHHI9NqCjZEvU1iPYYvNZUjojOMG2zurM+fcqA7h5D4BGRuGR
8XptD1icWzwVYoWKE0zN/qmxdjhuEZ3NNg8KahBQlUianR/a6WnL+r0T1m5x4zJv3+kOajckXsAw
3D2X4qrGpD7QTBQYzGKRkf8oMFiCsOH7XsNunUQ83KEtDL+6TQ49IopW4dShh631WoI/JnWF4L3E
PmmjDqc8MAD2o93bOyp7f+1ZS2tWYl+uAzet09VraDMCuSD62InqNgGD1g4G95mW7xdt5sMUJlT9
QteR6tgII9i9M+hgxhhOJ+lsLjcy4KWTw+HBwHzQoCvhSU/GHu6XO8NQdUAC9z02vsFpGLBn8Kpl
D/lye7/vSqdtiMiMQK25qdZodip3lHpKqJFJjUH4diJ0krqV/X4agOn4D6ecz21sAZ6vsqlx9c7d
sFCHUtkA3Bc3g3ijP1tRl9FLNSFfRMwu3dRkJIkmml8DPaW8iICPctVlS0Oe0KggjbCAM8mkV0Ni
6cNac2/uAoLMRpU7e/ZLC0e2yCVc5nzwTGk4Ziu3Ryta4HhGW69lngNCpepSPB9wOzXI9gu9ZkXt
rQaPCVlUeWKjTujTQ4t8U40L0ZbXkUd1QQtDdN8bMeoQWSrV7X4UX2o66gVu8WRBqWoWjDfSqYH/
/aBb3Q5yO19ZLeeZatMqLfeKmZ+crJJYwGApglFOcH/BzKXntiXni4VotzT1m2OqNsLl8MyRAROE
uocX6YywOdXaKMsbjVd/UR4qinoaVFEhaydvdwmENqaTQ44pMUppQQ/VSxAwBIwqvwVoZbNiIqp6
SEwJYTxykngpaRpDcvJ4EkexcMxOU6o5HbkZDHuDJr9i8stNQjBTJ0ju3Rv8MrLfJc2MBrgH8SDc
9UpQ/k3F+1jA+bgRHcWiW0yM+SDR0+vQZIluVhujCw3kH8CA5RRvkI305I46WxCLFTazlF9mngGa
+CduYWHB8ROXVBu7ZvoQhMzkww9OokliNMat3gngQxKU32NuvIicsMDy/Yo02qJcBPiq7uo9NTtt
axbLae70czONDkGzY2Q5KnTtTNNvdoqDlqwhM18WQCKBzhpnFsg7NkoWkl3fXFZB6RqGyOWSDDIn
8upyw+5GKhv5KR9OAqiVO7P5ZuucamkCl1L76gDJKsrsJJsAFHTof5QhkhmC12qFwJvNTBYOfdn6
R7zpAFCbykchpULqzQ59Vxoj4lqGv4w55xlqmbTNzZ8rNEgBgHlrJSXKLqRQkrg1T3LRjDNekxak
I9LFoEMK9bGg86ZOO6N8bvBOIiG5nRTBOtTUpbVHXps04vDP0e4ddYwYBuzhJhkyAbjHmsJoP8Bi
nyx9T5Xi2U4qcxTL+Oe+/6XRa4umSN4MwZ5E1UZXVC2FolTjn23E4KaqnuyhW18X0why3HfvBiiB
SC9tukCWtPuggnYr7IuVqbDIVW8xImFVtK/UlyeC+t3+o6dxRbCW/FHBgufdlPWXWllYtpGcLxiY
OIggqXn8k7vnagT7Cd4DzvEj1i8pxotO4VbAQ6J2LRP3mUPu0Kqzyg0ZrBNNRsM78XlsZfdc1yJX
quvmrpgQfeO99OkFHIZt2Lou9vD02giWy1zszIrNrgVwKi6aElVVs76hXyTJ7OKtOhQkw9TNuHPt
uAbWzSwP6GAKokJbvD6A37TlFlApZJuwhm/OToVtTMQhPi0XIer+1bVZg9DLY1zfnLg9+lKFXQ5F
UANvORQQ0FUGDaMaOpfgEIDeSg/1bSGpWuj+DoRIVkjtc7O6AC1TF3nSgXVs7sAx98GO4PdrlOY6
7r5FOGc9/gaPjJiD0IKHyTchHBbWoKEpdAkUcBYDlDNpe5C5IBiVeOXPCHx/NeoqHX88/Li54j6k
P80PnB4hbLRTZRf61nP38vv66GsYItIZf6+834r5eCkSmuiE/ONRWPif5uMycNqX0rmeIrrBl7j6
WY1Xp39aa+UAji5SuJXMc0DvRlqgvX2Rf3kPGKKwxhBzY1mqt5YUBEQO59tlUwGlo9dTdNpgP5K9
TfunQjnOSD8vAXt7ZRCtaZEOH6UWvPmcWYBSR6eIo7SqWiFQ91kgjG+uLQ3qUeMK2iU+4xBPK4ez
exY/LtoEO3/6O0zWsaP7tvmwplDz430mBzh56CngopDSZuH3yxCqnqrWxBViCy8geHtm/XTCHC+8
sh3FTiZQomNAp2YKvVcM+DMyNLXj+EYZArpDOGX+3ZU3IOZuV/xHsuMtE0sgEVQ2FWXD7PPiNPa1
x5G7xU3dz/ZgJ1wd4tyDvX1IXe6Vvj5WPK7R1G/fnbbYhpR8Y5MG6294RMO9l61PR1YgjE6O4dS0
AO7dtpglwk50KrlwxNwtzQ86dYTKY48jfidWrchrb1V1fvpWVeKmOiQGsq8WuZEwAXP9Mm/ghYf6
m3tkPnmnPA3ODtfI4gzht2bYkip+sbZ8e5JrHu7u+vIrhTZ6RA689Gae+Uns5I7SN/CXFm3/HXLx
YaGubaZ7akYGTzWIL+cpbqq/Vkkl7oW6U1JyBtpJz8N5oG3MUN0aKd+W3UE+vGWI4ux3V2arGw1W
6f58AnB6yK7XcZprWXlLNO/6iIU1glqslyIyhrFmzxcm/dwQj8VtIOR97heFxeHIh1d/92q3vbEG
7EHhyaGEyjq3IGqr1gQK6CeqAONMh+cHjBGTKjo6BLBFXFYi/geCLGaxoJddEtMMHsz85P4clm/J
jUsoBngBCJrSPul8BaaC0WNe+pwZzkHqn/Fbk+5G5UcVcq0XacbQjtcCKoqfSmDbuFDhJZsAncA5
19vLxQ8vIDCfZNCpqBuAbncZV3JdEhT+NYv7Vw9IGAV3MOB7mlEFPpQVddu1/KWxbkOS2+faLAlb
cI5ThzIpUXkJG5TYWxoj7E9NgiynuD6tBV2Ho3eQNRQIrvjKmm5DA8gQZq0/6LA5OKBMT/I+tipY
uWhWJyBy5erRWb7eiLKKQhKpCUXeb9BHJgRq235Jn5OXlHIlgWomnB1DMspEby7ieOw8chkG/TUM
WFXnMW2qi29WJB4r7MigN4LFQTECuTdxR+U/G2GNo5HWWnsymGjDrd2Peg+FJDH8dnjaJUDXmKqJ
VV56t3P9kOyIJqXL8nlKBOyT8Gmfrgqp0f48cpdl1s96lVCFFH0CYRM/jZP2hA0c/R4QFTOdwd7j
Ij20LonJHGCyXpA0+wbNLS7V7TIsf9C+jBpbfne4sM1cCAptENn5mYBOJYHpiWTO07S/JgLVrseT
R8nxmgQra3bkS7yCVjWv/HNjDFJPJHDyJGSJWSncE2fbMgY4oacm0fy/ZEplZtdjaxkZwz80USmE
K+Z/0YD/0PicNjO5YVGXQZTWBnGeuKr38m+yXDNFA0hkkz8/52gu5ocytCOD9aW463T3NPpmb785
QSTR1mCX6nL4/VYyMbFNK0SysEhwpJLSajaN8ikJ8f179DzRvswHJUR8JMiKn7KX3Q58nHLFLl/m
9FjKHJ9iWjVu8xJhpU8o0AIAiGNt8x6nw4XyWZ6Cee1EgElU7tuFCHNzSwt3MGWAwtfFqweQwbRS
sv51PMkFDZXghcKq+irplHSPbJa55EAAL5WgVkhYmXvHQafiqYKfZhTDiNW7DugtUJKqw8r/9Iru
NakEjYdN4IRzpYkkbZ4yfN7/iRZ6YesoyZkiqDqKBDTpfFvwXi7l5Z4EW8y5t6roqnqZ09xgsfDd
wPSmRxM9gctEYiTkgVBAZUq3CdNYlxtWxBdMr1hVtBmo5588qJpn4yYQn7CR9MJqnoCxXkZ8I7nK
n7lMRNxF2TVHnjnoKHfc6Y8lICh59NyBjdP6VXw+hGRgqZL1KUWEja7X0/joRzQlh210cQO9Pe2e
di5B64RPr1nmbDDV+t3XNwV/iLUXZvF2yPkeaqu9C5551O0g2m4IjFW4RrANuluQEvy6meARTKCb
j+TSAP/pFLgbhPNF7EW0iamNvEvjfGErec6A6tdrG6yudbC7G1D/8QnB17Gk0N9w0T+gdd5Lmkf6
E3EHgs45icVk6+IvM3mat+AB8RYb3TbnY1fn7taDaabKqiaHdkd2GxTKybXvQQI5MoXM2cSoVM+U
7EHBWGZqHCRAnBqsBlUppMWHEgPbqDuPcOpNr/oR93JldslfqIdlza2d9KRgvO2PtnPJTRTzsKpI
EuXzC51q4woz8/Re2TTeq+9mYZV6OqihmUMKWFwCmwHRhJ2nFrT0qz9qYP8gX19sN58cgcLBovXn
0mW8NMZk+6q6wV9RNyaigHrvLXdKjuxAwHoZTy2zmWYtpZwD5mTI+mgMke/yGs2z/Z1k+FE9iedA
y568Doz3oW4ZqR9J93RmDS7nbMhM0OzZcqAH9QQLg2xjSyGzKvmZWvwpB5cSfnW8K7pdD2L+WIYb
vapENA148X7k5p4Kb8D/TYrxh5ZX1BRIx+5+ZK4ZBF6ycAoK8iq43rDaA0Ye7QkB8pxt35s/T37b
w+jNgrboYMrvEMbe/EzlCfaWNER0tPPFbskOaNWW7cborxv/+jfzpIPPjEUDACbyeiWB5umFpJy/
FqJkXN3HMibwuM6eB57oEsZ1HNujdi05suLsISLSBhKGOcxu8+PSJhhOilJGgWV5RbQL84ty4U1v
BJI63OVGwqzSMMVrv286xgNjbVJLILQacgJI+6ZAgcuoxDSIYA3KkxUiGRu6ChmXnKWUrExzTdHz
G42+VabrJfqBB50AnkAKqp1+v65pn65fnx0lBKQjOmjMDp1KryIx5BeWb+oirj8Hq3tCPJvrwW8K
9MNnbe7NYz/IhFTSmv/ceRktKxb6A/Tll56voxIRtkasNcUKFTh63XWFXyiCtQdR9cNlz6WCdAgz
HKxyhmLUIO9jUQxt2ttkL+ObaFP1urgfS64cNekVtlNthTndBSKRujKVzEFuVxXISNHIZkWO823Y
uJv2lKnXGbBiqHVr1QnX9t3b/xqOP5TSfpBV54VvxODSaOav8+Qk5CpcTPhdsW2O2GgDtB+sJsnW
TXTUTt+EeO1/VI4+XM1JW0p2QI+lpHPUUj7EcLyMNovFaT87v1olu8ekGk6HCqBC5sjb3l0TOb5V
la+B1FPxT1klLa4qFNt1wfMKJCfyI3m7vdz0Jlyyr16uuZib+gZ4ejyIrMonj9fYHRgx7NYewZqr
W3/GewfU9Z6MRHcU9c0RuiuBWtgtwlAjQ/gOaWjtfuyBtpIER6zhCqINaO3y3eAI0fH8TYpr2AEa
I7cLy5Gz+zkgVZl4UYqCaodBKZOxkESjhZm00AbR+erjKm6AZ4+cWuOPezEM4O/CWjFZgoMSI12v
hALwR+uI3fO5NZB2Xi/EO6QZbuHAsOn1nZKCj+cOcHT7M5gAcgdmrO2rIEc21hUgEDWgskCeF+OJ
G7nHp8ZVLZiO4kAT50a2ftNHet+e1W15dyMgTbiNkH8u8c7k/e7y65bF1+vxyv5/T0/dy+/m9Qr2
Ma5aw4vCcW3fMx0QLB3WE2WoAIUmz0OpCIH2fWfwVeXxCHFA63QuMB76/zWVF0ZTE52oyOV1Kl0T
7L/6X80uXwC7tnwABuco4l943IQqm/YlnjWXXgfALuIq7CBY60uZr7DCiS/B06LWh9LTx68r5aH6
JRzyYOFtWDoj5HyJzQ2YN0pt5FzkMYrkp9vJxiOcuS+t7qT+vGRudHFBN/Zz0OzUJFVojcDipIXT
fDM6eGW901qq09LVroWrKkyFia6zD+794n7w7qirmuE+GsRLAA1gWUg3pS3WMrOpv3pRcseHkyO9
cwRGABWtt/iV8LPeZ7IHJ1tl/O7Tt5V93GtfqWaNnMxgLWtq/dphSKmyyX+oTmHgHTG/LD2s985s
k3Nq/r7VlN+/yQnu+xZK0UH1wNBaqQmf7COSbQoAHvtC5htihro2L+4m3c8z3daLeoRX7OTaJ0Zu
G4z3V6mtF+zphzts8Ejm4EdMD+i5/1ISK18j1GIslbgzPFaHueE50ZVIPfLfy2jzvzrfmjFn7pz4
om2naYhkJQ2gVponqvpcywuKv9aRbKwC1oGAozBQVlsv+XH9ggAcqhSA4rJ32KKzNOLjyPf6QJ8O
cLCqBOvMNeDVC9D09X5JdgUSszW1BdBvaSajZPsF7j9ClfLD7RzMo0MCfcfaMSgtkQn/Qv7wyyzV
K+BMUEXr9qnDNqBvd9ysBGrOxs4s1IaFnxVCRMCJIo1c2ZdI0dERX0zboNr0/A21pKqxqPhlVuD6
2uubyMmgP5EiKUvX+uM84gL3YDCATpaaIz25XM1KIUARb9SnZvv0mdiEkxX0UJA3lequcci4EFq/
B8TpgKVm65Hht8QJJUI1zkRV1e8i7K9FmjoWhHyZwU5oo6K7BPArjJtGC2TqRVyUxYH+0CMgqRJY
UG2iL3PI5WQXMQwAJclpN2fOq8JalqnjML30YNIK39lSLz+WDpNdMa4vRpkv1sCkoAphor9jeQbv
gQAofby0K/mBefoCB29nao5ZN8+aq0sSb7rLtiWE33QpTmsOQXN7V0AMyAU+qQK6/ofq6uDPMYFh
6f4AwHO4F4RJgEFoxSPIblhjUAIYkGscpwk2lC3YQRxW+b1M3RAtIrmA3+YvwCwgAX68snWuQTtL
uqQ+5L5rV0MDjLi/kyRjEEZDW+NjXWhfdAvBoOlR3+yEyEVVONMIk5HXjbN1Yeni1MKWYjhdqeQh
FFELbOt/PJb1Y0asveh8spHN/5EnwFKhfOCCuJCZn0Zt8jCQCPTNExPUq1W/ELCzO/PxssF4bQIk
pF/MiPoqFlJ6Ql2v41z2JznIzeUJEAqH5r/uNwgmDYhbQ6TwpXD/7qxe5wzGdExXW3qwS+xQGm3O
aV+CGc9s7kxt5WlDsRhXeSoCezbWkkfj9e8wZVC1nkZEsAm/4xSvtCp0w89AgPo8xdpuGRWwGTno
eH2wC+5koq+Dt7KjO++jlFzAR10ejcyXMYdHYQGP/toDliSbJpyLW4xWgb699Xbwt3l4QwkvawoA
7wV4d77vLjXDhunkJy0QkOIfl6SYe0M39FfwqS91LZwiY1Qj2y9Fhvum+VnDlUop7HPsmYs+UXuD
dZpeXlpOgWZ13CaayGtDA0NkJxXK1y3BJBc6xpSGATrelaFirg4JaMa15cKIRczOb1X37uhEZA8s
5p+NBRBooNc9RkyLjQNTYN3Zmg6X3ATLl0knqZyelLWfhrkTpYFaac5V6cMqzNBgxdZXW1rlyk+F
/XAL3RJHrhQenSShtX4Q6+WWZgth1BWcSJmxgdzqUI/kysfEfeZIO74nJhfSAwszqD4IDK7NAbTi
UTZF0eApv12ERjOa2uWsjefU0VVACxFy+02oRk9s2EU3svK9AUZ3VvxGOFrqM9vcJRByytyuqa4S
bS+zP8bInLkQAwd5yLkPiFmNB8muu/9KQm+b/GItFdxeZy6Ei96jDVjdf1cuclBLP6Sm++rY0Wyq
Avbd88f0Ddh32I36JVRKJaHY5q/72t6Yq1XCZch6iKH/+F8c3yasMoXMiHrhNw4qGXHXktmoyhyk
50RawcOEj9yLWHS6Qy1KQw2/ap143jbuPvlAK0C9K6/L2Xj6lgnrngpTTcLpGIev/U/EzaHrHJgC
nU/9i07qM8q30dpPfJ2JWzA+OxNVZxkVNtSt/puPVkqI1ISCKbpYPUttGvhO3MOUdG061o67X48o
JGRomqbZ1HXj9h7Y+QoN16pCPg/Gv//tZIXaWtn8cHJEJr3NBIhybG/pmRfC/X+xFkErkSAxfMhu
C3nVIGL997AmgWuJasHDF/HdKRqecAYnxVgO1ek2AlvW2l8sHNdcqIf+go8UpUA+N0FTXCLf01SQ
CRYR6yMKGI+WjVgwT4auGzHoP4KSgJ3VuRx+YABkblEmt52o6y04jCaoDGS86mPKz2L2VjL9+sWR
MhsesI9VZqzy+1ffcIsJL1yNJxUz6clsP9bgm4UHMk9DB0zRGTLjmmEiCUdkLQNOWmSsFMeK7RBl
h/F8cgZLUXHWFmtqWEaCfDwhT6O4oCboqi8kmhHCeoUc38wxSbszhWj5W55XD5tWvyAxRsq9Gml1
JEwep6BmtDTT+bDGYQFGgmV0vNwz6ii08TQZquffnJbiLHy92ueYMqtJU/QJV92qxVIhk8rpQKh6
AaasGwryLRoBtX4W7OKntaZa5CL5tShz7n4apObWjyLCq30SLjaSI5fCa1QJ/uPxa+5zJro9zyDe
BytBhoTkyQPmcBSqHZCFTD1e1yCf63oEfar+5/efsmfV5/MHf7jjNeYY57MXS/mxigie+NrE/kdg
dTl7RmKEBkhSMXszI8Z+9A6JIpzEjDoNr60A08KEmClZz0C3jhG4+ANYyml+XIOoGvv5u33e6xJU
eXrRJiSf/T9k/LlCK2m9nngQOWUCHN9yeT4wnhhx9TVi1GwM9zMqDZ2gsrIrqxW82ojiFVf9cGHk
+oGoNWAQn1taWqspGNk8y8kel5PRt0vUyr5WQG2tPAlJ/fARqYb5bDVkLoYU+dTLQXv+vzQBoP6S
YMh9d87uvswxCvN0dDfpoIk9tUiEnJ2yvu79oGeRSNNlkfFqbzfARuJHg00w3s17PznbiMvE77r0
9/ACPhcfX19UoR32TZBtvMER3PcpAkjovXVvbnLgyoapoik+nRbHmJOEY491XbtPvBhr9SmgnVLj
sbjds1atk719DVAgSj6XRKapzeV8aW521xNRsTxmSYm0YYa+pFFYiFAckYV5K/9gRBSp1GPAcpRF
AIKB+gO0mhFQCHXGGmHI/1ubnPBYOrK8b61HmYwXDD79BO/i1u1ib+5/lvnq7WxNq7aDqfYe3uqG
Q6lPMNBhdfWbBJOgzkoE4moU7nFbC9nG8f+cFXJxpzLPWpbr/3c/0zk45NEZbIz5NNQlolXC33PJ
xUYi65theQbkinPHoD8CGwiId4HZKqrmJYqPGTTo85/9JLzZmRFBqXDjp2V6FRmoDd55mHJygcez
ouTmsUtTTtiyJ3BOYe3OGk49f4B9GHWlPQnQsXP4K/5gnKga8JlTvCRasF2qc0qFO20tJuSNKOaN
vUQva2M1lBEHzc1HzFGK4LeM+KwifMr4ERhhJmgWpo3nFFGVIPntEiFsAF6OZEw7dIAMo9Vg1Nf8
eCDQkIQBCXXt9yjflWqEjec5nZmsohO1yFx/7UmSeKwElv4dN3mRbagaYjNq9dukilaRXv+oU5Ba
Sl6fqEp1CuhIwiNeHh7fa/K/lxk5u7saGPL8Nl8z6g/QcYiygn/HV9Rb+raz3w5hAhS0qqsG21/P
ZiIcLGdTT7Rdh0NYi3Q7UtZ7ROcWeTk6rKGRSz9uK8NEY1pDy8s9BzLSiegG6/OunwLMp0B2su/W
RCLJ+8wr6nJ0SV+h5ihxdf5qsY6XZ3trA5XKb19DTsAlNzfBqlDMYZ/WRz96JzLT8StoROvwVC35
a5J6NhoN/bEY+8DIqoagxtK664TVYT3O/N1TstKjd/uQSwPo4oR2ORh6F+B6CdkXKV9JAmjBKL2v
p8OFQkYMFppbVEdrJ5pd75XXyOu/+tTLORUxHqZSwHARDBPMVMjHKibVyf/vZ9JtHiSf7VwqOgzN
FHFPEb3zKwGgAiH5DsTH5stfayktAqcNBoJA6JMfhQfXVqJRnwCV4VKRJN82cwYoMSNaQCWy2MS3
W5uj3CveWGzaI7L7n86Hu/ti4C2M4JnpyCV5NIZSSmVRfV6O+3xYP0vGvBkudJHIQjuWGZUWdISS
MukyuEum2YZKtlhhW9gA7rlFG59fBKKyZj7MRQyyGTp0kNAKnq+duZWDvT09I5QkiSvyWbu6FOi6
TDKqOAIVWptdSOD8T7Sj7NnwLhFu+Vg4e/H7Heh6XHMfR2pRsn2tvz976OloGczH2aKUDvnbMCFP
BdAHLcGl+fniUwnRBr51U9M5MVETd1CogmvbjQ8EAdyH9lFle0ONPzgWXQTFu2EVUOPoCBG4TuhG
1A/Zygsef646M3QYZVZoK2tIW1kBUJmpNoY2BAe2PuvlKpULXqnOfW3JNk8Ee7mfbqYSOr0RfZ5K
dhf3RCitPAUyTZ5tZEXi22+oZrt/inAjoOB+hq7UoCwktJpVnBpaPoZoUUZwmmEyzAp9ZhCIh6+5
g9tTgR/ke3dglUXxR/9O3w5DpVQrSB3jukTEmPmsYmelUnT+QvIKeRCuzR1LxV2+QRvLkbeGzPT9
ryJZUpCife2tF8u/dYzycatkw5oLcIbKKFQh5URepfhP/DX+iFn1Qd2fV21oGyPce1xhnRNohDCN
QxGEp0VaROjbhCBFEgsT8YvANOKlw6K6oHgX/nVsz96Ejp70+2t8On1nBehsjh9F2If5VGe9eIH5
DO23NG6H0m0KmfT2RI7xvD+30rlts+wMBZdeCuGS+NME1ita7X7UEPqbZ43axEHxfxuSueOkk/tS
1ipHviWl/yOgdX7/kfUl2wyynFitcUrc+4TL/lxJTNSkr8+JNrp+OzcAnwip5OLVj+3HcabOShX9
X2L4DHFOk6VtZgH9s30mQtJXkhAG3FD+/+5XpF7CQhO2Q0YcWY5r3f/1WgoSliZ3VJTX7vCTMwrh
HgcsBEuJWlzxOAJ9A4jT5MEogFDK9srVD+Dpu23BrEsSHhxAK+d5Sp4jniy3InxDPvlNpVYRPuzA
YDdyl5eG1hxUwL6XmtGZCnBy/RUry9th+SsKZxOLLCL+wzEKBdIWv3zE0hvbp3M/FGIydkAxw1gE
U24fcYNV8sdGbLd8BgyyGbr21gjxJ+u22FDxQ6JPKEX81JqEJOLgem57XjRIQlqwZUbjUKncxkst
yLYhFzHTLOOcbXH82+EFRAJWCeT+RgGqeCW87x99O1L4q+Ei0sogGipyo0bcI2BIhC6417CclZQN
CH2bNauS8s2GXs/0HDV2R1ckaPJTebW+M3YyS8/S2S5KSQnbvCY+yJ1SFKse3jhM2cr18FD8PJgx
V/t0fSv5/Fq2OVvhIOVPY6ZgBy34i31OfSDJXj4ChYmv6QsKChCL0WxkqDaS2d9TyhvPxdNZVTvx
m9avPYVdFU7quRzp+ZJPJWHEc93kuLDOdozVgKuD2xh5NXI8YQlLC49yvwvu8rxi+Jds6K0m1KIp
7/qGltN65nTSiGidfj/ZJkVYtNBSSYgZpyHOnEFknziORB1ta5+cn6uVYeVSpNl+wF6QwfFLHSjm
fQkcIIIYxZvYkeQonc15wfLPGSGoINVHMUJmPU+tXpjci+ldOkPZH6qUxhrQzdvOf/0zfyV2i2IL
rsEUiZ/JibFbxlXfpgTnEu4e9BIRqs9qrncEIuxlAvCYgoTigcfAHA/DWjSzVdlwAj9LTu2lxyx/
eCf+hvSJ7xSQtzjQc4lLHZ4lj90J4emwSqB7DkEGdrjINNqoRZd2JzN8PY+w0GandoQKbN5RaQiO
hqdx/NDL0CCijM+GwvkPwHsWqMptRlJIQiiTEt0OFa6KfqnqCHfDno3X0sWm35g+mvizPq3ZODi3
oRuXHe1hCmnnQVEwprH48R5I6yPziUWlbYplPXUiKL5hm6rBHAyiM6IRa8OubhP621DhWkrCACL8
6Kq29dFzN9PW8Z4NNfyZG/w0/4MyKeaftRcAb2RQe4qIIRrfEJ0Q6ODgOdvvYyr9+juxxqVN8NPb
FB86EDP3AstWTY5kNzL3ZhYrsOphM7TCiujYnrluYHF5maFPmIWdnxrC6TryYmIyPHW6EgmXr0R1
FYftbTPA6q1it6xKG2A6FEPrfj5cTuY12rH3+GXVio07meo6ER2EXs5yRhgovrRflkpSHkPInJVW
nSvnw5hc5kEUH5IJfekYfzR3NJv4OumhnuYrAKLyndq7ZFL90ckofX1RAQ9B7Gm2u6s/E3hfXVY2
I9g+7mLoXvd+b3sROf3zrOXaYod+o8vygUi0xqG8loY5FGjQKvPCIAZ4H8lriLTzZbjmMJet46Uw
F7Uiv0Hef2TD+xc6FjAmYSxv5b0crX1YjCPZnLBLE4o2fYmcAX8G4Ml3Sl5I3jLf/vXvbF1YrMgY
3mEzatEiXwIO/iiwbW9UQLk2kJzYrHgB/eHou3yr3DU6aDWjIr/H4eMYrFTKfZGzz+8bP0Sx46Dz
akT3PmOFDn4YL1Bk+7HbD84XgTGMlYdBlTm4KFECRKq/pUBR2gKbq/z1MCGzibonJaDt9zCZ/Hyc
1itsUXkwBr5TI+vtIawJpOrxXjo1SM8sk0JKu77xy+TarOmFi4yMYcEY8A/wW2iKn51SWEBUTmkZ
t+YUAVttSnz50OZWyA2ZlUqsCR5VB2ue+3Tl0CFSQtpyAahI8NpNPxbrwZAcswlB02rsbOwmnyW5
pIhuDXAZUROVxLX+n7Zd/ulEm2WAx9qX0nP7Nmizl9JJsJuX3jmoERGdYnSwc8R7bk0IhrcB7pZ9
EztOZ1LYz+C993XYQX/lUmaob3+jH0Qg55CQ34dcBv13p2H8HBpGMg4VWff4vjJFHB4l+nNUnyHs
pH2qF7yKeg6Jb8Ng0I8M8lpR9Ahti5IE0+UKKVK6VAxCya/2bj6mHkA5zbJzKOFBljcMqP06nF6C
RAHJ246geeWGsqFvXBX52fwEJMmrdeO9lLc5AhAqssOp8rf/P3lZsQTrj6rEqqQPnx1hR62/eCuO
RjwrjbYW9gwzTEBAdSIs2ZolxVq2fFPT5uFXtdXjfScRmWR/pUpe0R5Yy6/fJmDoORFmP/7nvSYM
MfG/KIkNxnFnmoYBuwjGSCCkSrTiVQkun0sabw3jjve0s27gdsACIfOuZcq3GxUQLmJBNmDSfnf9
qPKv4BUK8zzFHVVH6qQ2EBaoQ6Z/7286KVzFN4d+Q9t5ryd+e2RJE2IGI2vnFTunTDzhdOkiK7Gh
ABuhcYP5LSp/W8FqchggrZPGvC0ROoblTdhDJ/zpndY1997YAt2rqbVciEmfhDmiIU/HgM9kN6zF
U93zo9c81t6UdHEsSqKWr2VAda/vYpWNjWnESyKwnQ6SO/sFSkM81u9s0BhQYK4D5qsdtrGcSrp9
UhJ52nyT+PvSxGsMfgdR8S2dgI1lx+4OLXkaiY+bMiHxmYd8UsGSmXAt2f69EB5AdM6zulVK4VLa
zXPlVweo22zRTXEeDAyKgWbWsUWsPeb3V3yZxo1LgycBLGXrBsxS7bUmiqhLwfsVNPaLUZqpy7un
B2Biaj8Rseb1U0TzAmaWkZA++GlEhA/ZOcTu2mln2l9u2o7WmiTYh2rFJ4fogfND+l5m4JG5KpdE
zhaFEWQGGcMhKsRjwQ0efBmykW2hEAqGP92Wn8Tuhm19slZ2wYBIZauikbcDU4nRuGDvUtzu7rUT
k/MDRWO89X1xDNY4Kd7EYmAJ/OTTGYq4hZlmz6TGLe/lI9tmG2UIkEwkCKzsWooRPfzPWVWyC5Zd
7mQDDZHTugTeDSyaScU6iCwZhpZ3ydYYbWAQRIE1wLj8vhympezC0Qqj/ARaSqjHjE8UqeFpvoti
rlXIOJqls0Kg081Sdu6BOBA8g9ZBHpV5GjEyVigQORd46dVXPKat2G/ZRvn1SzTkXzqUwNcY3yDb
ZJEln2t9br4GbjRSwC0UGU30nzR0X9YAA4UqAfrya4Ge9tA/uNpPPzrZL9h/tCswpTWBepC46Z0G
p/E9XhYGRVTx7r8p95Pr1OenUw4ndRR6upaATJCw2d5NFTgEReBWnOR0d4AU6aDFV1MdBO330Kqz
RqL/wqB71uTCBFDkKPZt/OfPyMl89DVxYR6RotZ6HReb3DptE8A9GyvuMzkcInyN+xEkgPdWexRd
V3SlmBgp78ZYRYJb3dR8LPxGDqz4qtz859LP8eyLZ78BsQ1T6cs3yVCeIer6xivmh/yrZ6d/HPF2
wU4Qit7doZvppgKllTGrB48CaHF2f/ecY0FTAH7mHwyMzzLkMIVzf7Ifddo39PUikF/2g05V+sRP
i/cIWIgoSojmFENcMriP1wI1sRHzYFVq0xdd84ukQhXTZdkJ85jN7tnXsh90VTDcguUyDzy3byQp
C2aVy7PT3LXeDZZwDBCJ4BF0CzHCSCGXGmCJjxuxSzL9NTahfS115zYxS0e3UG0gWqKpIO1yjji/
gAbK5SYVlGHIiRNnmOT4SnMeQnbZPooa4ZxY01vynRBk5btporeKMN62pPV4agbnC5E892+RDdib
RAa/xhQXNHrwK3BWk4V4S9rk4liVunzQ1VEXcasZXIbbLANu1+Xj0WHlQCyc7gslV4sWG4OTIzzh
w4RacIcK/+wZGVMyc9KkPFaJ6Qb3B/zNoqir88xWRmHzpq1OFHqMhwc8/NS8SQgEknN7cElFZiUZ
oklqVSBwgwnTbAt7bLLi5tvQ/itR6+Vgwqkbr97ETzwJ9znXs7QixMXyGh0DUY24TBkWRrxziB9q
+5JHiyxQlrkzJ8AeovKfFlceVRHACkYLZbNK2FVCkgVDId3MIYYoZj/r9pK5HQ5lFJ30gv8/6HPB
E9igsL37tquZtLbfmHkXMPCAhni+a9NtGzgMsdP01ZLlZZttNlfYT3wRaF6nQ3iMypQQg5p53pWB
comYq2Ltoe1j6xF3DqZMzIm8tIcOz7Lm4jRLC2PutQoOIya0w554FZkfO1e2dsRD7HP2Mtn1fkGL
/W79JHjHrYP+Qlji2trYWEprZ42CWh/YKGmQiEUo7ex7MFLaM/LtdhzVfnxUyQXdKC1S5f4X6D4c
+luQ1uwBjMnXSueGzohdxHk95zi0mCF+L1kfiX6HO7e12on01fXgvelWujbXT5edzCuOY2iZ2Kui
1DsGzpyN/MttEj20XoumqRK4dqssICyMNBUF3CDan49+Fxp6MItfEgsmk19kK0ssIc11nnKk9Opd
AgHm7PBvRslTl3dtqPh0VVtm/5bW4XtkZg1ro5pNqTznju8vXna8VF6kWOG+fjlU/YtWPNATPYfU
fWYLkVOFspL/2u2ddkK6GXDzjyUpwqf/jMSvXcyyPdb/wTFdstMOWBEF4fL482ZO//PvDxhdDnVm
gL2MyUSEUHpCCcLtuOo2S3CEh9deJB9kFy9/1dxunaBy82zU5m2e/aFX6lWQuF4Ud42Ltw17OTJ9
KbLDznQxc4HAYOEcMB7uRcSBc2YX/sYyEpYizwJ6fmsxx0B6jATL241+2LJ86/cfpzQ9bpy58RmW
jfl1ljUvcSQg6yy9ty2Y+FJ60gjOeTUvBgtl5+O7T4lnHT/2LwkQfXkBf1d76v/vDTC5y6jXQFjr
PCdBml9H5tM2hN8yohWcUZLT+fKkL3MTPOFWurQUEGLqtztYtKbmEPME2DABO7eAvm4MmqUgRhwW
QZ0xsL5g8IqoQuv6lUX9vgoDvVOc6DV1LS2X4xraPIMRw/g+W8x8mfDPAVCO6q+bYnpGtXtVoIiU
hcrTiTDHpA1mC25RI00hGy2xqboKE2BiFJpTsI+iWEfxQqg/GWLug5egcGj2ekKrBS09/SKgVh/J
RDgYSEr2W5QZiG7rse6ifuWdzfc6BjXcId0/L4TGAeHWgpsxFP8mwtnWwNUyP8qRs+F0057MSSvW
/QjaJ4yu6XAyObvKbUEJ6Yp4WIwKdfpkQNQTYMqU9bN2GA36sznws7nKgx+5aUaE7LzkbqeDgftO
hfRZEdajwNQoEWtn+IC7wAenehuzaYgD5x/LWtMH9yfn3YuZvGZEclpnt3dDvmg3wDRX/YnAK6ma
3M9QFxf9n1Ch7/54lTiaTpX46sQ+USEQ1C5r3S9cZ+kOHu3WFxeLSh7clfgHzys808sHE0ks8bh9
6PGzwo3ARyzDgQYspW/V+9MpwS6vRinFWnx6/u3N7bK9fy+dxe0KHeyEszQ/KMANVx7zoDz5vb7J
ziWAEjmBtfuZg2MeV+xeYPCTeSXzr3H6rDH69yLXyIuusdtX8e2pZIAtEw5JXOkBjMb6RCwLNuSi
2aPusQ6U6CYQnXA0gzWFIFts8x2o4siSqaFon46niDz7k/Kz2bu6zgPLzdcXlmuq9ES6ouIfL5Qy
CjVXw7SGs9FaRo2rrkp4KdUlnN38csLbS4ktx4gsLO3o5KslwB1bW1WRPKWt5le4RF3APc7ElIwv
lwH8TjHHwecqqHRaycmmyvhgrOaYSmuIuaruwPWHKldqWjJ4UYiJxA0LZCkSMEJsAe3FvHeysVXa
RiTb4rK1TIUpubjPPfJRmutu316Hq074NtSQpfBpkr8Muqw3JXTLTii7AKXTDRVg7WE/LQXksvc6
URu586FiXUpBNQabMWgckmpXHre5gfQUo4TrXopTi7soKMj7gAbxYOWclR7Llv+UGyZMTpMvHrFG
AtUcWGBrXsJrooI+XGFQQyPwfoQEG/nOLNRGTZulzx5wYKVZnMPU7U3f66U6P3dYXiai5vTuUpOm
QtY0KCSSfkYH4oBAPKxfB4Rui7DYHsEL2yeCoXG3U0WFTSCqXi8LCA6JTxSz3YcGO5GpEmCcsSbL
vY1feVZQrzeNC+CqREA7L5gHo2NxRSOzhrHpsk+SbU5M/Lu5+SoPumfTGUheOlAeo7puLzgqx227
42mO2nrKRuR31k6kKTDSNkPXvleN1faK5t/X/oTcV8z9WrhvAn6ZuMUCk6wSkD2jSWKy4EPVTWbe
hjVxzmFPDX7GCxyiEGut+cfKCmUVZXYQz7QNVoNmrUzcRjkEjQLAdS1RTMBtaFiaYmqDTPLAXuKr
iZfM5KvmzGDNFtAi5g4CrNhAw5uA8XFY3tTjUtLlp27C+N/D2VVDNB700bm0lc2swl7mL3ji/tBC
eV8wGodyi8UDU/t+e4deghW8VLXzJPsylyWicdqqyopFOpPrpljBMBhpslKoQdlNlMvCtb15zwRl
fNLhd3KA/PYHpu/95PdAoHAUA+iGqUHpJngiGwSyEa/uTwo3kedoEj68gz2XcxDrFr1OIhNgNjOV
m3XiPS1I4dP3qMI8vD6rx7qnlcTEv/J85qyqM/5fn+VNiGdTxJnp9sccG50n6DiDkejN47xIhjmP
v3lIeBe6DBzPSu4LwijLJ/3AZUt2T3+rdroi/YLy1eQMJ2SgfsIDz4IDLJJ3V5Qjs69SjGL0U17G
7rZojC6dypWyySjUmvvXvMZ+kAQpbyxzQaxwYRXJNTXW9AVEsErR88c6kmmTuLzi2nO0bNi6G/73
DNbxYht4J1BMKaRE96upzKCILOvcGI6lqm1liyShRHtE4Lp5PYTeDWVpeePjftqP9txI/1tGU/lx
0wCMCOeHh2F7ibsLEXAajldazW5qtDQKgmxdkrhcGORM8B1PUJyT5RuCdZZct4aCAHI29OyNY6CY
PHR/lNPgoOYy6R3kyWPtsmOfPGX7uSMCCgfjfj4wVePYRI5aETsWdOmEXwzM1cTlbROxnbyKWC2a
7TWqQXJ6pe7hd9GWcapjf6l5skco5fQepJ+WzR+ZH6vYKE3wIrc3qB+tZ7C379BuVFPNw9f1O6Bp
Xgan+IgyZbJsq+hI+xhAT+M+aYJ8IoTw2weopGK9dI+QDp2LxiWn99iuL5PR+xBFzsTl5+hlhYS7
n7BF02xkScSqWtYxU2w+Oy0RGu4iQiA6zKdO8L5SXA5w9lQr2GFZz7yk1bwyOaVBhjOyXLgBCkg2
EhSSursmQffP9sTvCyEX0vAZoMtF2x7qZhkutahoxTlCd6xjkA/XXMeQpe13vot68C5njIL6KsGN
wTxuWiDz2MzvHS+A/RVZMF+e6QidcuxZ5ADCJX2kjVv4rw75KYXG/DIIdbQVZP8j9B0WTsHIcZI6
+Ytr9ot+iBom4akxpkHi7ijiXkLUYZ21xkAcrgcrzYA4mWNHHq9n3OR0RCG5WrE8qZdKu6OJq5hb
3cKEVLBcMSZp6g4Cjihp4obiHE6rxfUT1z6WMuvt4q8lfGEO1YzoYRFV3kURzM1AH0+5QEQUgNK1
zZ3HIzPL3O2T0uFimDPm3G6nKF5K2ULcYeh0qux5XRuqp9Eg8vNi/NSDU7uR9Zm9Y9vX5g5HGZRT
pmGpZPkd2Phy9OBUFYaFWdMYeRDyHYpzx+fLjS1SuPX4YI2QUtFQJYrb74rBk6FVFBpb3yj/Kv1l
+ayG5Wl8Fqa1qg3IwiLh5YGEWpWApfaibe1q0hijozabnvoPJvA5hGBpFHJfaIGA760ACwd7CgnO
dp62/5SVeTONZA1BWDW+nZkSis5GLFniB55NXeZw0m60828s1oYk/3TdPvhb6XuWfaYFDMENdBiV
g92SUqTm3xNtitd1T2ym8QBv7+n68YpdKIL/Di4td28HP3OufB8/+ASIcB7joVWvH56JXnp0gd4g
VnJGsB13bJRHEWdk7NlBR7e2glfNJqJBRZgO3IdlF3pT4aX2PRA9Vot1j6vY7YaBNeF5XBgUmdMA
qjDJc4qHX4IsCciBRNzk9ukWs7+aO/Jj2msD7Igv05fhUNama6f3Yq6tbj9D9pRhYjN/2JgXQJfG
GpfaFhCQ4JVvBTq7pVSykDo5ePVJDC+AS5uYHJMxtzKYQ/DPeeBvt2ARqHWAvUViuqhIQLxx2wHh
Xju/bkR/r/B/Fd9thxsy+Bc0vqiVPJo/tLNXiiE04gBVZqvw/NXgRv6acCHgL0gsodHKpMAwMUWx
YI960GJlpwL2Kb1+/slhS7J2WErW4Y4VhfUshWw1rW2hP8YUZffzOu1FZJPctZ7XGlVw8dK6mIdw
McKnKgduBgCQKR+owcV4KNDIzfC4ZVmRXZrSLQ8G3zkNHLxH6xNPPHpgWwgUO/JLK/2I54m6xIQi
DKbpNuiOd6bqrucjDlk4pzl/+1S3bBUA6WskPVGfT7sw/vFId7YNk6lNhQbCC330sANP+tMVoeqw
67t4XJBPRSpg4nK5aDQnGPQwvIQiO30L3Irs2keh0lpf5FKgl+khxmroV55aoqPYefHoqnzl+zIl
wOWN8nO9fMrlAOcHEHeGMK628W0DevlrEslJS4aYQ+1twtNjIriqDFC5eznuDfaCOofH0ja5KPON
mhSEnXPQqXmta19Q2WBo3CBlHzK8Na7Adm86alOGI9acBesnZCmMCavpmsgWIN4ZGrt+Cw9nHeDq
nhTTbhc5L1EAH1aRBX77xc6vfznooE3cWUQD2kmooBjR8qXPx/Slk/RwQLDNaXTiWXDS5RDz5jf0
VRgtE7S6YGrOtojZtHqkiMRuTpT17IWX0yRYT0uHhHnZmBrWnGroGisnv246QT/cC1sLrSnTg5v3
gUNvLd/QeFcru5kz55TihQhIt18qKEJBQOS1Xv5mE+z1CXqN2P22ZTOxjM5GHQb0fkGjkF0uSYUi
FYuIksf7mDmMuA5y3o9aPBdZBDRCk6dqaG9ssfZY4Grlt8OdFmbPvbciJyIhmppleXFxWHShMpix
7pbt0tzC0AKgE3sDQKvGixCB9yqKBZnNpF8yYL+hEE5mcCtferePyehs3uwU30GLJZOhBHWUWDof
dCCerolMkxlfdbLpDsUi6kh/i6eYSxmZmtNykeOQDz+Ee6REGiNhrY7a8B28/PVYW7QFnekSWt3E
nKJ2klH1+c3q44o3OxfaSmqock3QYNRJ0iWQO8QOB6IkqtKYkjIxOeTADJs/Gi4EaVqZU8EfTFVK
LYFX40Y0YJcynqKwP5laoCXMBjtl7SvON1xIe7ylby8uChm98i9npenYk3ZzrRMypcimDU62lDXI
HlCy5Z5n79YbX8ufim6F7FUgLhqRygUDhiUVlpl/NHGQLbGigz7F3N19E6+aIVQ/ybxj4icPJC8V
VBs24dNFs8LAyww4NASdFajifw5EDis8jQRk8bG2ShGMA4JZ97VKP2CFmT178kZYIsXjqLg96QQk
e5KLiQkHuvcvjJTiZFzCwWHyD6GQ8U57cP2QT8dv0WRSoIRXH+pdae74FuyHsUmO4DYrirBpM68f
jgWbwTGAFQHHQhlgTimAzz62AlZeaEbyb1wk5ec0HNi8Vr62w5jCRZFo7+1iwpKkAJFZvt5TB/qT
tZ07dpQewdfur0CBsZJQEkNJTDQy+zLC5bR2HnIcBcZZR8Keqp+tJxffzQdZr1JmCxzl5tX8bFxs
6u0CqVWL2/GQrp8hFvjNQcSEOEcX80AomQn0R4sUo/LrT0uo2d5663ZsfPJyQ17FGflSTHewiiED
BHeWi9bXNBdUDJwL6c9POAPwvGpTjcqHqMX13Cf2imIoNFO5+MkUCtgPliVWCZ+d2EG/rtnb5Aim
oQxECGyGpp4T+HieeHhKILStZ4tnaBAngv3beWQ3RjFNtFixLuTJVwMsuahnZUeGLes0Me67fcPy
TXZ3XkoEiVpMcRMtjJi6BqKQoTH3LROQPe6f4erWslGXHEy1rhPuoa0wqO/T1IoITn3tdZxNnCtU
dyplPYlTCXnFmXeI1kyrQvmtJGK5aFlcagjnwKeo/HvOD6dMvkN84NPg3D114saTLJiPiYxUCL3W
hdM/29XDKFM4GHqSzgCogp6iqhiKrhhPd16gj775w55SBqkv7SSGCh98Ze8Jqx24cPEpfYGz2KWU
aZgcn/jKIPTmjUPWTvvOxCklSD/mR7xHW5z0krRABcN3QKJ+tJXLXgbiVMrTw9zjAZwXVtNKIh+p
uUxZces6SLXDlfDWlLoVIvMHPIW0+xo9L1KMWakIuBoys6X/JEAp/72lJ9tMrHpZCG2WLNX1OlFb
TydY8CBYEBVyMjJuiGwrgCRH7BUuX7wq4L273xsUqH4dbVAisBxRI9DjZA3tZFmAU8nHle0IA+Ah
vkQG1zbiRlAz2BRHFMt/VxqIp5t/heKxcgAzCo1pR7bETqDTyhOjnW3LD3X+L6MIsvVD4P83e/QD
kdLjnvUaPz4dZm0zmUNbbuwLAP9zEvpzIhUXtkbxWY5AGXCTWuOkNpZ9il6n5tsVZq4du+BGATO1
c092lwBQ9JsYcqi1bvuSV2uZaZp5/UxvXO7tUZLMOvweD1edQNRbJc4sBs+nlhWGbpdmK6AamEbb
VGrtFg8eVAVEHDZYdwnKw4dFuTmPnJwgz9tzXKnL9Z7YC2e9moof8WjGvjHpbUzYfsZtq6Y6fTEa
yWI++1C3yko4K7kOuzmCP6RNXK8aGB97x30r9CZkpIS92oqQWY//0FsiZeVCqZmlETvLrb0y0jxr
NOMqeYGVuD9VD6qLftNmVJixgrwSK1HthdgNG0LBEQP7cBz8ieOlZ5rxFpTjdtKzpMRw+e/07vMT
wi35seFyUERSxpT7qWdrQr+0qseuBjWBkDOjqz2omA6yfKIVjdaglSSA825dK2h93qBJ3vgCEdOc
RnaniwVQSh6yDQg6V6APkS3vJl9PvPw6QC/fwfGGsQLMy4nZU4UtC8zp5dSQgWejT2wuFQCP6V3b
gZG+NhJyfBWql/hLYSvkFGGXn/9Is2u2RmOtLrMU1PThBtMk7mifcEfkrdJ3ytgsvlz9TArlv6gj
2Bd3V0bUYgjtO/MPKeaZ7je2Y5hs7t8zRe1vXKNrjFL8dBxNhu2ja8SGg78lb2k3lGcDiwmFrh01
Bs9YJ9FSuesdnvL01smufONrHw/IMWdzNUlbEEIVWNTF0TWGGWhp6bFCBo9VSJTywA9cYFlEyLWa
MBTlpQl77hEbROlM6CCz8pF+IA+lXCrjbey96TNfL8kk5AVROYTqGizPs/GV5ZmojOWwcJZ5+nTb
Qg0Ae/j53g7AmoTvK71KV8lALtc/QwNHzfE1EreAvVSdbI1JlRiECYee5JypdzY74+X3vZC/MuXT
TZThMqk3WYqsKPpDkYwVeTgCrMq/uKUB9yGQ0gMR9RHZmD21Ed3ACoR3S1w9LxuKYJoMvFDe8/do
12b3ziKSvWMjItFKmTlTZ5gESDzcKYQPOrV6Mysad6BBpSQIsAWl5JPOoCXyv4Dyjf4rdkDACQTR
hazmVWEdfL5BMEzp5dLkIll/a9gdhtELzDD7iKtkOJcfDiWzVbEEWWtIu8mZ1Fxq0haJOwDGZsR0
dNeQSVUe33lEeMme22JgWGvk79Z8foI7f+SI6xcnp1tNRxt6KPBzPTiVyQbQxDuXma3skm8/kiZm
TWsh/KB9D2X82BV7UECYR/pVkmy5TBHhUY6e7GxnaI6dnn32UoH8FtCcHgyqmMZemV8CbQEH7icJ
w3XZMKGz1mH1fkgkzVSdj3aIMIl/hwaYFZ/7PIV5W1A+2wiv6fpk/bpIVb8AUDeKS/TD32R/FDVV
j2H+TJphprZ1xXf6h00NxKG/FWgHm4b4YCvO0E2gjncK9DmKCTJBk27YTBJ7lVqn/B7unofu2Adl
SjCrwh+hIffVWo2u6MehtJzJodtgnax1I57szQJGZIrdB5NnBcE+Mva55azT2mTtQyQZ9U1Oeezm
paiWTgaEtfSnDDRHwfzvueT2T+ltMW1pDSgCbQW7SZMkZVSvhfzXmY16zmGAh/jORm7kulFkPFLe
T93Oe1Dt84cpXddnuFO3TaVeQRtnG2vhZbsPMOTPbH+DcQcfAATDx9dEt70fivkLWgQDdLKSL938
TMUSeRsuncFdskE1eki/yE+VsmtyG9VFLsRloJByo8cfWZb6/EapxeyZ3Q8MvmVR/vsFUDAOGMAJ
9yJxdisf5w/dWVDAr1ZDRJ2x7ynqRgPYU4U7g19Z/erO+VfZUIs7pLtYsb+l3Csj72SFrEi75Rzr
YlVxnWdF/mMHWSdQg6MjwLpXx2hiyZkQngqQekrkGuNF1GryJoMt8LdYApwe3+EQBPS1/RdcE1Ti
qSDiBnY9O5SCGRJy/SWwWFoGVaxF/sA0qE3iL2xhjbredp9fmP0iGPqab/YK0/AM1xM6ogVlHM3U
pzn8VuQrQ91xoIHbpf9YgT8QmdN2mcrbfSirFS41+iShE4FxpWrqzeh2nXGpGFqmvbySnZljdL/J
6nNyEgzOYZoXl5ygMSqLxQhkKvr7zV3W4fCR4Gl5s12ql4VOESEX74HSr7DVJFt2tTFg6awX6pZe
IytFD4VbxF6oMUcBdFn9pEGeBOVxPYthrd0XhZPwSoZ6Zp1TkM9LN1fRkbsfpeo9nBYxJdkKbv6P
j9Es3sx89ho+l/JdTczmQ6lTZjuyr07xQD0Gisy0P3HCCE6FBtL0E3YZjyWkTBKBBBiKujTbvvoj
oNmW2mOQPOjkx+OCvypawQppL+zXoexGMkUqpaF8HVhgLZcqgwxknBptUVKqe4jwYC1RuhWyGmEB
eptbW2uv6kYBZX1OJ7afoSPtG+0vfNIAEZL1lrno/7BDE8r/I00izwv0skKDuA+c5jP/03dz2teU
FLIJVu9t3WvFK1X4H9XxfmsC8NNlRXXIyLyjMek5ruFHUYGnW61KL57cDk4XJwqkqkc5pODb50Oh
EXvbFN7T1LddrkilgjkoPPb3XQbLWfirW3efGq2ImLJhb7oG/kthra76Dan3NV8uGZNMGcXUQfUi
dOEPETHtb3t/069SEaiyg68z5vr3K1bGKCQTL/+6IDrilbZRRqDyhdwjXd4Y2IaABx5t9PX2fFCA
CXjVRJIeHDyqnSThJTDTb8ARiPpaFf4f/63J4iAeugYKHzZ9LNlJvv/GQfYgZK6XCr4qVV4s+Jl8
ktstJl3zxRjdm0X+UqJUC+ZqKdn7+hq3MmZaKPhTjLFJDIkMOLI8GEucdTbttXMMBUcWcFQDW6Uj
K5ix8/rZKg1TfwzxvOqnt7G9grteupRHRn+Lr4oOOe7uo/U9fk3nUjvbNVV0ZiW+RPCxj8MJtD34
lxUAW1Zu1cfkt0/UULKJ6CvVRgjGvHPT+PGBdY/cFGX66fmnxCtFu9eKIiP6ZikOAqg6drcmOIjr
etpEBqGcOjXv/pBTpyuxMj4KByaFonOu0j11zycfXieLsNWZ++v7ux54t1esNlJ21GU01s98qNy9
IpQyh7fRAVLp9JUGN6HeIz1bA1L8tT5aNwJ6cgxNVVEJzVIkk3QN8rhegp9/gyj0O6sOCyZFYr54
7y1wDbTAnN3JVUEqzov9rK8HWIHVpRqWd9xAjGKnAgPmO5LoxdGaMd1GkfWkldt9QKfJDTGS97X5
baVwZkF99r5kZRzYPaVrSbA2xk1ztD54XKC/7uVO1sJHJFmP6OLZTpz/OIKK3ikT3xm5qfwWUcrK
Je7+VViC/FSfbaRK14mcCHIWsG8/Z427d0IG4k1E91zZbDrCqzq2djO2hZhTb3TKOQXvXsIhv4ji
ozSepbp60R93AIDzrJ9KKqZXp8+7EWRefi2buTNwrreBmld76sXABa+kmJZ53I0owF6uyOpMuIvt
aSf3QhyYdu70g+zKDMs5+lXnVhz7JIGUVptzS6ArE8anvcIKr8DWYnSH8yv5NK/4uL/opAbxhMCb
lE1hiG0lVQjCCs35j0FINexuD8qFeEEOkf08HfR/NYMmboVcIqvAd3qB0cmbc5mezKZJNgNUUfqF
6KSOvIQngnb5iUN1yWEvvgOOVLRUg5qN9lotufOUXHNmnkccL1ODKdzgR0bzlMtptMqnhhkxlBrg
MbUiwGlVffZdp10RA6NpwOhXKIVZhjYrBB835gxedWvGdh3zu3YHc9Y2JZpmCzQwk6aRRjZ1VvZZ
laDjJqLkWc+mFFP1IPZ/w27xKxed3tnLLaToHPOtzGbafh2FB3aPRYICLpkK6nBLb6i+uOLuwGuk
jp/56RcuZbY+AL6WYRqLRLuvsGi5E8elWtJDwe71ZXixIpt3p1ZeZ/ssJ+gMCdGZbMGbvBcZp2kJ
CqhIjD5ptBvn8IHbOOaNXPA+beP/lkIGyDvfbhNjsv0B6B5jH+a+IwOiLnDRBu1O3IW12cp4zBaq
WuezRnAl4PUI+HUbBMWsH8xtMqcJzOozL3AUpCR801T9/gX9A1XjqMrTUHFJnnfc1zr1JkVP7TxL
r1Rzzjy1FSZnTKyCNLdZ4ET1ScSkERfelBITbLut9QdixEqZL+8phnqL3lCTuBHA5hmy2NzvRTQm
Xj3GOmD2k7zfVJQvfNfY+aoPBvFBtDi4HIq/SDwO7CafZlmDZDQ6pftgjgiBYpdF5Gz3ZLF+hiHd
WkmuNlamBN9QtfKV7p7uumcO0JY28/HKzBb1GXUZRZpJztnrvcJWTDfT8JhxuJuswPW2DnptHZHu
1gmPfrP8FVfyqK+0ys6uFSKivbFAgXU96RgAu3v+165+fmJFXrRXP38VGfIGOywdsDMPu46hLxLZ
668ycOEzMxArMfSSqpBee02pylFZNjuGJxj5JnbXf/TwDeCNk/XCGvg23bRsbHxiDoHgsTl9RCxg
8oaPAM11H5OGPamAvrS4VpJdqtKcesUM7qMXSetu0Y/PwOnKzTxKBY01LF6gpMKzi89LmWFxuh+m
2zSIdY8fV+NaWEPHRUa4WSh79M3ZUYSN/XbdDIoD64HwJIQ4yFe4GyjD9MmG7u1yXrtN3VDS4XhW
zJYj4YXB4l/D+SWUy5WzWX7+T4GnbTp8LksjAF02mQ/Kb2InyIU5ePlYj6NtkPMNr2p3S6kX6nmu
tLfSBeVUksKJVfJvVgCpH+ocJYKC2rk0kg+Zwba3s+zXM6LOWIF9ENeYIPoVXuTQmPBiIs3LFd1s
JabyS+TCK97QgbvxSKX8iLRvT6+bPODL8rUVT0SgayzmwMUPSHi3bxJYsbE1EqhX2xrgM2R5NSUi
5/R9TG0aqKS2Nz2hJ6wa+XqvqgrJD69Pj8yymFtMjc2VkhM1+e1pHL5CzVa+xw9vXfF2iOZLpf1b
tsb3HDx6LyKY6k5vldpCHBnc5okNBBr7160wMZUKGr9Mx64T36M+GghSkavFpnF+Pj4lL4zd/VXT
HCZi0qm0L3NJsakfgdWqegfjy85zeXSu1SHkTyqazvVztiQMnK1Ylts1snMVo6Xb0AFg8YDsbwp/
mcZtO+Trx+dI6xRZrMs1Pd9qsrQctx39JZcww+c1kt3JjoIqTxniEuux9a+BCJ6QVxhSJXDh9b/M
5g5iOPEJ+8YDlDlvZSCKMamAu0k12XEy6f+UemER+V+7V8BLxPFw1TKEC8mg14S+qYA/GQ8fDonO
DtunyIiEUH3abBatpQIHcz9eVF+RKdEWpX4VgL3DgAxGLmu2/0LzeX+qwFOh14X74ur54naoJAwi
K2EBJgmi3e02Dy148BNrAzK1FAXs7Rhl5BUI31OYAdcOwJ0Qo3qNxqzLH5HxOQU9sLlRzy69LxHz
Kuw/Qyzon6rPNyNIoJJ3jYnP+d2+MdoZm5csYMiJ/wH9sNo+JcnN46wViVe/04Dg9oHY7uBQv6XA
IJHVa1fK7mF0FDkxYybZA+i3B5kEZ6QWkutx2qXojjZBHi2vuLdH9mJh4pK4O6zyPpWbG1OnfOYr
7bry6kQbTh+NJfq3vciXvolsK4cUIV6kHRtNmyZE7WEpmJnfyzM5K++UWmp9FMF2B5bodl4BHiVG
qqN0iaaZbiiWF2aAyPPqVhj7tDKyIMHCNCQfLGokm74zx62P3/D07n726y/6rfj9nyGNBLO1Zcjy
cDOoLkWllJNdrOLHuCUDd350JqTmCd7b80mUIxi2Ofek9pTjrZXMoCmu6n9G+Jij6elaqihQnb7z
+izXvA6Rl0Fgg/wmtsykYXYmDNym+AYJJiXbkR1ANkOsL4e+jnZlvkP/zncjyQ0FF1+J5k71zJYW
SIorK/esrgghEN7wKN+oQaSMs25+enAhWAMlr5xZBCVhGQFIVQsiByaRNEGlvi/QzjQrRyRLs3/h
O5DKDNbwSSXWxR8NO+g1odFk7O9BIkpGLP5CrPCWXcj5VXnrbfSF09gCFAG7aM08tdUY0rspS/+y
sQJXyU1UT0W2p2n4e/dWkuI8K/hhHsSbc1uq1CpzorlxXnZRzJOC24y3zMoUgs2oS30uch+DpNhT
b9dZZQMDDk2Thbqc2e3Soa+txMLGwTOiaFtfK28f/QLEEKEMEJm4FDODHiOmySsAqnmLE2PZAmzG
PVfeOS/90cy3F65K8Kffyh/fMLCUNQfDSgKcEHQNyKmPu2I84sDfKTuf24YLgK0XHlNWY5eiZtQ0
GIKXO6Uah6SjAAsyagCXUVcmj1BCV/a2ZkOPdVdwEeMZMkQJE2k39a4J1+qD9Il+/kOAcKKPt2RO
XhWlYzy8JnGPql/4/ammN3EYWwIbZ21ZGsgEonApXy6mZbTK9dh4PoSLe6+HeAb+56/Ng1nDJG5K
RQJ2sIlwZcGq2jeQ5BIF8Yz2p5qPsSIh7aSQb92nwtxxNj2q/KtvcHaXdNsXk2rOfDC6K71Fe1mc
0wPfHOQya4Vz1Evn+j2ayIDkR5qtmTjlO7V0T/Jxq+rbWzsazDYAYMsmZx2acQIFVS6SaqBGclAB
Okqi3EiBt/pxEMiDjDQFGQpctELxSsujaJ5M6tpEb3aAhcG6CboShcA920vlcAayqrHOwLU8p6cH
G3oxplbQKD4GZu9YRFEaY3h9m5bAjGF1A8WtBS5p/pWxiWPQauQuobinStqMR2X/GqMbO0iAyBA5
Z/cZJ3Hvy4W78W8wKWKZT9LhNe6krTihPSALv1o5NhhOlWJoRxUecj4lTi/JGt+Nc36HvYusPC3o
DVhkBgX4RmNsTLkPhieeGLafhAAzM8iygcCshl4fbWMvm0r5ABQKQlaqvP8mtUH5EbXUL2F8gFTn
zcW+KL4g5dBF9Z5VdaeOhNBcG4ejMzC7ZN6NtprObH97Q/lXPjAnUwnEB1awrj5VMn32KrNuy8CY
kDudl/p5V2MIkO+h9cEMT92I85ynvE+Wdac/+prmDJpXt1zYPH7SrL93lDuBtUPs01AnTQU8rHCO
Gx9hkIG8yb8FwWxOqACOOh2S5Cj0AFnXbb9x/2DwRF2c4nj0Qm6bIVpUIaTFIVJ12MQAdTCHhyuA
h3B20Eraf874QslnkwG9o4t57olfX3z/buiL6J2UPtN3KiltLoIAZU0Y1UJZLpCBbAwz53IyJoyX
DK5Kle1LtDCn9lMDmsosYcrtVFCJhn6S4FMw4y4x88QKtF9nKY2nkkYM1XYj2p3O1q+9ISoj/cur
k1sWdUbEpc4/SDMFVPOg6pu4tj5tEI7+t1cI00Z4quZT/Mam5h4X0VjzvRM068+uVaT8e2CdoqnU
7uLpN74ADrcpFR01eUakBhDEw4j0wwv50gxcSbe+C6f3M4eSyPWMkwUzEkodiyUqIaTQg6qdRs3V
oP1BLfuK/yYyiV7iBuPLQRGUql0A6JDSIBE4jE1/DK2oVHdAeRWlELQwvT1Y1pCnfgdgTB7JHnJ4
GKYRd+PEj5+MK396j0yZ4qCj3JyLOQi+0+XQS0b49K5LJbqYDH1vAgb4zan3pyOdGOfNPXU021nG
0y4qlPvzEMBhHFLq/LvvrNSX1dr73oTEP5sF4+K+Ih9rKlFgHJr6FsBTswXg7mR80cujU5AuBUfA
APEUeoNtOGTOmOZ01n8+tCC8FUOhjElxZtsoNOfBf+5g6AHLEO6g6Bwx9xKEr6nXauLjjqVIx7e3
WDN3Y1o66voCoZMNbtLABrKj4Ups552/v4BRhhm4iJS96lq0VClLzkkvaWT3PLjUv6VPmK+Grr/c
U08GIHgos9fpK2Z1g/abiAr7hPkqR4SsoidzGe1QLJKv6s0Z3WHsNmDUSS3Q5mZ3D02lB6vxXVdx
wRmdCf8t2MqQRu39nfaVuYtQORR+5i98WwKJGDbnVL2my/18mozqtjIY+4QPv9iN+YjCHmXqpDXP
RY6iD+ozXn5E41axyQl/qbPRMek5PZ2PsF0htOb2z+YrJawO6Wwa51HaOB6XQ4ABSyP/2TQTxnKI
6GSB1yAZMWcuIw9lBQ364KgTwqk7JVe4fcTuzt6izjiKCh4QN+OgpOCKAZIx/ya/hMQmECGyRCaK
UST5QA/Fs7i619RsQ0Nv8fdqXpi2GgJTUNPDjz5zoTjxWNTwqF5wZKvi5kNPsBTL9fTIOru1OMZc
R4J0k4Y1xPhQLI7/a/kc6E7eSYRpqQmkkAzFNtwmDd+4jT0alP/O7f7CnjSYYCCzR1z0qQEBVVpR
8y0CYlJgGUjuYDWT4t3GgfWqxLkpQRSP0On0xenJOci8Dvs7QcX5q/IwCcnpiCo04SyEothapH6f
UziEdAwYSciCVckd+rCnHHQA0lkCtgcGmj1rNeHaBuiGAxdapiGoH1ybRhfUawl3Pe9C7juRS00G
LttO1bVAIzQnv07jMJ43IKZwbJQfaQ28BvCRYrTSfcjZBM6aVE89EGRcBJNH94HVTXVbe5ZteI0l
rV/EYnaX67qg7mBEjysSTTJt98/apPxTCvZlz2lUmIa494tDSO6s66CMw2UYSonTuIRBXy9SN8sE
GMNPueN90HY/ao5WOpii6nXhDrvyO70DPzCg5Pg4KCbm0m4wvFf3p4Slm/PXg/EHjB7w/8o6qItC
gaXiGTwatZ+pyAvPlR2YyUzplONNFA0L4Dyycw+CAN6gUYqCyhIY577Gs26DTKH5xn872XLzKEnm
m4Om3mSN+SLpm1ayJgd71DMcwUZJC0mqBrn+6ydYH6Dl4u6mdtC5rgfedHWaNiHili1dJWA/ApJ3
7Y2XHD+vTkpFIy9kX1WbSxyHwF0Gh5mSNclY04mIqJm8A/6OPFs72tRTjjOzLIVL55EMyQ53CD/2
2fFXl4hI2ZXGpdAQKiYMPkngDd3O6XSwxG8Rd4m+GVTgV9wBjQPMjAiu6zB8pZjFE/A+ioU2jSGH
nfJ82xEpPwL+Wc3+7OWXJHLbS3ezhX090ZqDxFV/a8WgW0aY0Bl8oz7aj4UFL2rF9Ozx8XtDxZwO
SDw5B8OC1+JYotaGqPtGzECVnxqPIOccxe3G22yVsYFT326z22ro/PYg6/BOQbV4ETrBWdmjRNVr
M3TMm1SHtWYVEkUru/up4WnmfN1n8cP+2qOzyXsIhr+TXIDCkjhtNOGn+/VuVZNoCqzIZFmVgqRm
hM28FAgVvzhu4Uz7YfQgj0GO1HlSGtqEsDXdqcSw3cFQio3+up+k1nABL3udRGqthg0tO4zgr+0H
QfNHmVo4SgTVPVuRHZqLMujgXOJVd/ECtwwQdG75lFih9ye3ouyi5vB60w9mf2ej7es+buPepzg/
OycFhoJKNQ2WxaPSZsHuxFSnEmeCoMPZX6uuVLWSuUOy9Og7CPCcCQO7JJfk8nQt9px9T+a3VKVD
5ANcxnd2MZ6ag9W8/3SOnLZJGcTNyznWeCRuiKKWmWRM+vibIDZGGgGH4BGnEG+Objr98+K7VkZW
HtkozXuqJDSzBIusWCICzkwgCgIh6C9RldX+mUK40yXeLJK09jhLfvhqeQHcBJjYw4tXaAKbN9e5
WCsPczqf3dDk+3h0Bztm1wqCqENo/WnMmBuo74qIej5Bootj+KI6xk5AsppB9dNDD8eiuPQYfZyz
0uk59DFWHGNaULhztbTDtZ94t4+sjIhHX9o7Jdjbz752wq4uE+/gkmM9i0LsFq1B6KSHHi0nwsNM
fr2WLP4poOmKEmIJ/d6e/CPQoA3JkF6Vz48qQRXUPo7dR+Yy3onnYRPYUIwJ4xkvL5zz3O6hGqp4
rawUF4rAG0PlJilZpcLiSnL27q41nU8YhoNLW5Z2eqPrhkBk2YbZZMp49IfaL1pACMrJHQ7HfGG6
W+iTkejuqD7cfYNpyJ0GnlPnNZrcSgTMDyFnx7DA2XMnNJMSxXtNrHhL30U3iffdPK4+oKhvLgtq
pQjf+Sj9cCE8GxQpiE1wfPNc9JuCz4KpLEdnp2Hp80f2sMINOTwa8t3NI5DIZTZ4qmGKxmuF217v
gtfFOUkBwMFVhcVcTME8QSDzPqB6xdTYUhD8LxsbTrD/zF7ouyuxclrp5S5t01eEoq1x0B/9iDbA
lhP9WTst6Pkck8QJ/9eSlaevtWNjgXHlI9ob480YYlGQ7wfNEmE22f97/vO7eOzrBTu3zkZJ7N7/
7KTc8QBLlNKCKw4WDvkqBP6KR5PgEnSK4WxfqS0WC2OrZdOOGunn5DySuBgIX7e9Juq9NJfOLdgb
D4go9PaQvsDy/8JuCm8vVd6NH6AfZap/8gT2llXHbX/FD8PRqFSlPIqfmCb4EKG+qOGSWdHH0b19
K/rFMVcITYASmLg297wjy/DA50bEgvKL/iQE+n2zGXOx85BiYDbK+KYApCyX3/FAIyZl9Oz6zos9
HN5jOJDerQJhPmWeUSfIEGHK5Uey7tNM92Ol3uR+ZXZ8TAIDz5z6CxMlsI70Yv9GdcAXAYtXTJxL
jL5B9X5Uyi2A2fQQIDAMnzoDQcTYw6AscyaoO6QDOWeUMYyJ0AtoFbaFTtOeIOAXvwZYeuPROG77
Jpu9OxhrhOQJEoll24mzHOoBDRmh2cNXgrTGrBJidbwXAniaqlcwFUE5vWSxRXTq3eHrbCgFRtz6
yrRcPbxTzORbWeETp5snAjsXeHOy2Ky5cSYDR3w2I8fjR7/NTlzQOuPfg283lWvGW4wknulFW3Ei
io097gL+baOqZ9DuzMcEPPhTy79hjKTw/WTDxVG2KqU5P95usub1Cdhu9lFm2AePFZE7CxhpfLZG
mmqrpHr1LsQPTtbT5KvIoHRSniJ/5QCxuCkrAViCgCErvSkJ+r+J5ozZOLL302nac0IEzlYQBWvw
bwftXNzLFZ3oFkB/iRRORUYrPVeltF5f+7TjGk0wOBGeGjs0BmOpvDSUMBUh1Jq3DKpDFuhbdVDy
2aapHg83SImRrwd/CXedeT14H46Spqc5oJ+a7c24QhXVzs0Eedgse6FBDpivPljHZWKkIVNmakp7
CoLcRAZZQYVQ4EBSSUmTbivVFZQiqBSzxFFNScxUKaZ3ZAGCTUjczMdUhqHM2Aij+H7rEq3J8uZu
kMBVs5SmQ3+SZe4Q0NqyNsin/P8DfrmnJJLek5nFF+/KIVbBSvAcU8CiCxY8G3TUI3Rf0rE5AMsu
t3ScSVs4nGgti8Z955LbPUQk2C1QkmFMPzKOMifHi9IHR+NF6vlw5Lh1t44UvVax6Qo1wkjWaghJ
LDR5wf0E0u5w58liQ1DMrHoJouRD4V5dp7Ss/tofpoBHAhdC0BIy9t43l4r4g8g9zgu6mgmFdunF
ZwI59xdBLysLDhBk9SfCUGXodR7CRZZk1ggcuoOCgtvilNSJe928KaKEc3XkOpyN8JULJRKZsPSW
SntAP4Le8dxbrPfOfJHx/hPpXdF2BoRtKzoTRPBOIAdJHt9EPmAf8xZo7FwMo3qg9GdZNf38q8Dy
itQ46mKuV5hnJVWGY6flEPClLSt5euSLv449Tbv0YtR3CT9u16oeByx2Qi02FB5XBrQelf1t9CMU
2tAht6hRBCoA+dFrBptKfhmcfKZD+zUbJKirZgdEh1aNUwF/rU4kprV1A6cMzrO0EvvXoBMGNd16
c8QnrBIa9BUymTecOnJvFxDqIdAlX/JHnpX7Slu9H764LAVDA6o9yPRFUXzJ+3+LPrX9pzBi1Nne
ObqStuxaes3pwSbxSH31WxSjw92gBqfXg3Msh8drHxTA0iouoevA9iOq3F6IKJ6Iu/43DqbGybDn
9V+dB4JJNJGjk+pcoPOZ0Bgt/8aIzCwrApYzg/QAOkB6B2UO+hOwtEIMrqm1Kz+qhnx/VREsWpOf
4qSYDVnmsUebncUNFzy/ObR9t+BAxKLzIsvaqRp9XJugTRtpmub+DhGEF9c9hA0Aw+phdXrR2JpB
DEw2Po5Z0+3d7zWdM8ZwsTMBnbFqqtY3wQcJjGKRBhAbRUd0/TEyGGbnxIFT+PRS9KGcGgYZBqBp
oYhLU/UMZXDj2yElteHdv623W9cLDgooN0L6Ly4GF9pAf+t0SSyWcWSCNhZw/YOWd2fTj0G0DZj5
9JwJgBG48JkFpdH5YmHMoK4XVEMTJfHvX07ULGr3gwfxSZZjOHuC7uirmHAA47S/k2asWxgZfmtK
Z9MbfiwRiM3K3SjAHX0jZlfeN5hofxQrwc/U8Mqxk0jjk3YDpobGdn8oQninvTzWmhszS1beoFNF
URxF68hQN/KQVXeEisgQLA8quA7jGa9IKwx/UuJQaYzwRNFsQcuO/bnAgTd/AqxQGiU4HT4nQUh5
4m3HpCpJTBT3bAWRqqccxQsxTCZyVk9JuUeaRkM3vfcmFpVzbokr/VBNPjaJ+MLJJ5rM6ZB55SFV
0IlmiFwOJBFL8xXeoBUXHRCFown+G9wDMoQEOTs0aS3dXpl3emFVHfdD+vbVjOsAKEyvSd3/lXbq
HnndeuzqPHjKTCHR9KADX6jeIgx2wvbNWOIOlpXi2Err7wywf3IQ4DnjzIEFYGJTKi04Ke6QZ4eX
Kx+6U6Mghb2/F9RTnWeJY+bFEA1GwmedWmqYcW0e23dL/9m/vBugVr277G9m3Wgqum4D63tskugj
7x53Hqz8g3Y+ZXt/bWYFdqMh3zGNOua3j+l0cabBBeyCZn4w3/hAIungo+2jBka3CqGeWLfs4p9w
W3R+ia89yRYghN3dBjN0HLMKTEEdLpESGg62ZmC49/4sqdWSn0Xksp5d0FHSJLZCMx/eRfejS+Sz
IMbTHZe57/O6+R6O9v5sguYuMQITfOeyZ6c8eo5/ZqGUmJObfXOITCl4jaNC0NOaIAe0WhfsrVr/
d73g25oc/KE+j4lElCfzUd7CGj+JsG6G2nfg5lGlFOvpmaVZhR7HP3w2DPemLcnOvVyg5og6oxzx
B8wJZDeFsb6tI40JDxq2BucwmqIBRH1y6hv7N9p6cnL6TiixyKEAlOKH3BhAFcQ+EeWqq1F2zdn0
VrfdpVbSupAE9ZuIeMw1o/BLDdxyyPnQUNxLvC1TlueIkZTpHtMkIpVayJL1t//R3WHIm20XyHm4
k3IMxWF0jgCJwOVcoiekl49E1EWU4K014kOMWQJcF/Jkju1hCPTDfBUBEuf+pvIQRBGh4PCsHW6T
jQ9CaCChYXkqUSZz3QDl/mjOitAO5y7LR4T+FaoVBonyRfqbwCgAgASYAli7aneDprUyYLcr6c7S
jWUxAyr2j17UCRMHu7I9mXmd6tyNTHgUvGqZ2kegB9E8qEnpdQU0/L8U36fJ8H44GO0ctAsxJ0uA
AW9dM+OpUtM37YRTlfDo7gIFp0znz048iQlQ7Sd8v9bxblNq6AQhsOcFn7wMjEtAXPgBKqmVHYw5
YEYJF/5NdwNkbdegTEklGUWA7FmmAzfAQZNE9ewfMkamnzNW+30PDutVJOj5xly3thqpzn20flF2
DTVG00X5LMK4ugT3oZ1wAuTYkYKq7e0/a3lTg6ZM49m387ZH/gChMEKSYwjkopDwhoJjt/eUHGWr
SXEU81cZ2BFlv3F4dvpHJeBMJ9QuSlItSJQ6fO+aOKIv1RTtwMVexhLdCGeRSvdu4MZPYP9tDCVR
AzRL3eswzb0tjmFvPVBdhbi6sAR/5Ow0NnX0xJzcdGkeLULXP4ChOFcrA7LyvLeX3cYZcSLno/pH
YnYdlZyZ+odUa0/8TnyNFN6v0Vq1P6rq75f3aKfu4LbWDwldrKke2ZcUCZ1ER3Y2TNIf2bUzdWPt
m13fIWs7iTR7U69JG8zHS1i36hYDRGXiXh/R1vtu90hzUK74DPl8d7VKUG/8BAJ5UCdU0DkPsxge
wBK6XAoJCT8kRB4w+S7Xe2JazWgidMQNw6F5ZKHabitqz37UHlGhiKKem3IAR3Q51XOI9Z/BeQCJ
Go5Uy2awzSXvQ/Y36WCbBksd6kSuaPv/k0gYzQNm6EJvw76NeLzFV/jacwrbg0ESeQslO96PwsfN
1zdPaGX1h1qZqEm6zqPfa6gUjyjGl/dOpuOu22EDoWuRI4foOkOvUGYwU86dwsG24qnT1ROnru1p
gXER51QbxJBltCVh5vq5eByjGHbNXF/Yi/4QUsyjFNhUDk2lp9Sf7jH6OHkHDStU8KPyw8kkemih
+Ofls1wXS+K6pWGD/VohmWnnPprXLeSIHlKvj3eV6CKbY9g4TNN+8G/HOzTVf66R4mOpqGxmHtz1
QjQYNwHDnamvhhVda/94VxhPUFPdRZg+eN6YEzh2MtOdtWIYRUW8VExFpq2Hwn3AqRQSgZIZ0xMa
+ruvmjEcdASSMGqdqt/l855PVkBcLtNFAQrHIT5l4deeK42sBmyjW5ASQ01dSOWtz2LavEJs+cGA
H531hM7sBxQv6KXH69I3MuRCXHJ2WsDaWRIKoAaEVKGRsGvvISeHBD+CGzyhaYhWwZyXB/BTb8yq
h9W83AoXyNheDbZF/bv9372yL0PL+UUOwMB+xU/HXGIfRqRFl4eippfsYD3OHz5rL0J3VTu7fkax
K3k7fPhIdtT+quZnxBazJ6EG0fN+GCR29hApLKd2lH1LC+9WSAGECUZPgQnMcVrhtL1ghGp8hUe6
L1bkUQPO4yMS3i6ZuYIzNjPHDellFLKnpgmgeTENP6O7GXiKM9hhNmU6iB8ZajFG3ovSBVTCE1CR
XsB8N2o+sgc2ZSUDzFr0/IomHbyVCv7+/2i5szExmJ+Y4N43MybUb2pvsItotu6i8LTAPcbAIfu+
IqnTrsr+8fMiiIqBvAx1NShYGk788Ui1AL1pOBEmRcPNIvbqTGFEmLVJ/VK25J8ZXNlAsSTUslxx
9QWan9mEYVr/qI8Y+mS6kmqTGIIkv/reYKjjjfUfmVFsYVc9p5RbwhAVcmav10HBOUb+U2AnCj0H
VH/oAajtaJn67nPb7VFGZMt4HopIJbEGN8w5EeHEYA/Sz8vg6Grqpo5Jcxy3hX+nwa9QI6DeEQFs
dxV+JIsUq0S8eogRzNcC9WOXlA2D/+m3Cq5pB/FJxhpGaGxI9WanS4ShNxhNW0wq7ePJ6SjSDEKM
jEAs6f4UhOJWoTF5ldhR+ehwnIjxGW3EBo2P6MY3x+eXO5g7XuKst7VnQP2eR0Y3Pi1EhpfXJXWB
Z7z/9puw/gVKVyUes7Hfuh+m3myRW/ue9769f6BKQDTGaaAxoYpokUqIMMjXeXBXxeT5WYxiNIiE
paIB1TK9Eb01+sNxGLgfQIDMbmJY/YAG9UmZ1cBsZ/TkoHUJvqr6h65y1yVk7r+8XzjvY+E+SP6H
dnhUfWtqLa/20qWBwb3TBdLSYgyqkkxJ8FTnkrUMuxDGKQd4qGZiwcR0s/NE1Y+64zTkERBB37o4
W/eGqEA1yotyJTM7l/Yco7YuDDEw8bg0m2Efl3shWIayx2skyn6XNSOVSlpO5j38KQD1PUcLMmJE
xeAzk9av02BUPyBAMIJZ3Qfku6fZkzf/A/V48KT5fA5BT02fwbDcpuijy2snZo1ZgdQ5MhUeLmp8
QL9T6ITep8+lVmllcD6mhcGF/GZ0z0rSV+EcZUuiOPqrUtrgCOs15XRzI6Z2S3PRnpMKAQFCOysi
cwaWtP8jgFeS/8fuYY7MTwAjArqDJEtAMyjYZqfMNmD11wGr6jr83Ll4w55HZ2xulZ/332rZSy7Z
2z5+IPLtFw06Yv87qJqbtLtGwc2EBTSHA/NhOX3vEdzKLLoaFIqkOLEplzjpzECcDwI9eSxFO71P
CMCjGyn9xjeX0/xBzInsvbzzF/95txskPK1UCCPlKYjdwT/459rfRYIc+jAiF4715NQ8LWkrUUun
OymtW/E9xauFW7+nBXWw1Z+TYA8XWCyPxfcEdynXbfidb+ZuF+9mRQpJ+Fedy6w/RMvvzLLH1SAF
tSTmFtFpSpoL+fFAqzJO+FihdDJalr+Uubbs+Abqk6LXbKdN8orN2QurO6+qq/hClZKX1UDE8PAn
qx7G1PxFv6JhJFeSchK4ObyiSBaLsdMXjJCxvpSG6E9dRvgT6VEjwPwBtUiDZozAnkMihfT232xx
TFuOrRLd4oUBBsQ4SGhrBgmy0g77S7BflNkQ6kPCu47s6E7Fv0c0Debx5bAkutF6SjxWfcUa0Fez
eOFsVyr514yW9yowXjEK2fuc+4p3Jb3anNTldZFw1BeFTgUyYxMYuH+W6DDSDMOXDT1E5QLpdVnb
i46Urbe+5dMbZuUnBA+myOMvxCNiaGE3CG8+vycukv3AVBJhx8TmyBq66x1sMnXRbMnx00tp+c8Q
aZhCTqz+Wl/nhYfmm4l5NzkewIhOCvJv2XeTj/ueCr3kk+ZCd4uRwXZ/UIwCze9c00BJb0LtX82S
d+aTzwiXrVd9ww9gHlCHV1OGTaBuO0RPQPhD5gmMRrEqH4415/Hf2JmkUNAqtj5/iZUZXoP3smZu
S0+PJVhasjOmRZ51DVP91//clUDHSl20kVcXqALDJVmnYUjv7OT+YaNs/Ri52TOGobktK+ia1EdW
yr5PkENI2e+kPgdePh64ypviV59PGNQ3V+BCtIj0BaqRB825i576iqGpDr9KeXyj2AMmeg5OKLtq
Oik6elUNI+ngb7i++KwfGQCmu9t8g8t56K8F8uMwiBwe2WdJG9tbEv8hOh1E5ze3/bpCKRPbi1gL
zkyBb9+zmuJHWEZgcN1u0X7yIqeTBzmQl80hIRhBiZMlZsnRZT5kN0UD0/UuLuUhML6mLCperesR
x7O73p3u48/0zfvQGbAm3NkCVM5W0NfdJL2oiNctyPTdyJBn9SW3HOMFLpBw5T0VmuCCLYy5cfVk
MqfXdB6hFQzeiK7awmv0F42HshmE4pb7zUDOt7KXUkUAQIFl/aVM8fnTNm/A1ThIl+nmqdyMlVJv
i8KAyP5U7+UcU1rsNCMLeKbtAYVCOgsBn5HanOAo2WuCG6l66rqZi43sccXe78as1FPTicgYAwOI
I6LOtT5UVL4m3UynjR5vNBmGABfOWi+iS0/jwgHgCIOm6j91pLNyOhLfTK0peXNc9wbFIihhENXU
GnqJVwqwMtb4QK8bnGPBTADaQaqFymUpCPydzvp5ZApMzkXZbLPevqpgyOrgtvAKSs15pm+s0RnA
5xTD7Gem/Gm/29uOxE0q7cy3zJYFuacBfYDGd/1JDowWsc0r5oqNTWcCJMBc5ziZqPZkh8bjx2JC
IV7Dgx+/DbxmqYXC6iOIHQcyRby6l5DfzwtyWtBdVt9DcZQPk6zLGuFAOiPMSiwRaJbPUCjoJJU/
8Oojpv7ZyJFj2ufdXCUbhFgdwhWNsoG8tj0/9kPGclLEhGCHLOdhnx/qsoqlb76nQQXOU7QaD7wZ
4SpcjOaR4QcStjvTDgH84+NN9pMYDZWedizTDlrmSxpBYgEog9P0ADgqCyRXG7k3basUWL1rzODy
N8X+jN6pzjSxoskw4exuJ3WUu4DbYwiiPvO2GEcP0U0ILvwyt4LQ/Sh/JA4bzC5kc0C9wZZgOG1p
TG0gtqn+j+Yo0Uo3GQ8pUAnI8lF95tEnxqnWb3nAdJlfqKR93yT4u7hWwugmxz1WoxM/3k+J0g77
CFkngpKImZdjr15J7v0Zo/FoVBKQY4PW11N9SYz5gF37bO8OVImtQZCbuaRzBx+is1uyRCqGxgyr
qmALTEi2OpyDxPy3VL/oJxzILndfl5p/n5DnLMn5IujUbInIMA+J82Q6nuAkjfwUaSBLMISdbHzj
n8NmbEwEgPL4HlCJMgBc4Pb+ryTTqwwDTmhdJWZML6UFXZGYxEsCkVnnuxyvpZn+sSln8Qj54WB4
4iusuPXRKx6lBlqQAD40GMSBct0lRxHhiXpojEDVH2R/qPeojZY66xpSiwLIneDo/8knVZ/P5vaO
2nGYUvTHqIwPuQ8+k5xrBilecm68osyZcD6W4eyM9gVeVKs3sF3KtNvPa2QEc40c/j37+yCgN3mG
jZF7C3/LIMwl3a51DAPDYvvi2T2f+iB4IJWeM70lmx+xrlkXxCwY4b6mRtvTV3eDnhKW0lTmlKwD
pi41sVOtat34MJZvlGTUQY0mza0oARToDNivUrpq1N43SW7d29LVwjeqKF5I1qZYSQX3jAhi21Tj
vhkCpLeWkXXrn5qYqTj9mWm4dwclDSA+2wNyYjGEUOvRAMbVTnxIiZyYFen4IiBAICCizfdpVaSy
VEJFTRI8WlGrrer2L0mCiGvu34Em7dZfCyCfVIoAX0VxdVU++dB91Z7syc0Q+PE5M7gtpw1J9zai
w87BjxDKH41KS6OJNsUEa8TfRHVu/wG5z5dtQ6nr9nUqM5VkjT3qRGsXiuJAwrg3IyXn0bYUQtzx
Ig2KqGoqrqbApOsoFUn7SDE4u2cBk1AAOKU5AJ2uf9ifRUwGFtTSh8OtQxZFdyTvvtknD1KiKHte
e+J+v6sc040MGl971rExFuHSbyB2DUG+IcRmCLN/mZzTlkKOcphLi/yK4XqNwjg41TUjwMHdIRRW
FGIoMvvUQTMwSrzwZ/J4AlrILlg54LlDLVtnuz3N1hQPmT4twxS45lj9QQyUWIyN2NVIaKzn3Y05
xav5u7h5MDwn+iQPk1wFR5GsffPGvXaj1zcZJG7+2YNohchQjZkXywo9eFTfjHGwg1/GAhtdVB5l
zySPynlsRSjNDK3Adj7cIIVSsbp1HfIZX/C3QHIiHSB3OE5Tp+/PZ6UPQea25fridiAX8PbNPKHN
JaAQlmCynsoiZ2hPmlkDtsUlanF7JAOrjzZn0nxqJ0zpP/McjkOtyAN0nIEEUVQmFzK/bvcHL2xY
d3jnTLAT8l5FKIFQzTsxAwoqVuFQect67/vdg35yQsILXRxKNCrkUSW5cha//KTvnr8zlUAp5Kxw
b3oxOCBuVEQPovixteVaQLjGvPP05QSSvkTnuiMnUZhYPyKH4JexJh3SRhPNn+8tQZrxJTo6b1aF
6ZxPObLpOlmt+RiUH+T9EnboLWjKxgz+SP8A52MiKNQdRYbL7paXFfSYdbGpx8U9RXqM0MqgSMKR
qMgF5oOleVhmf4xQe7XPDMBDmh7azUjNFYcL1aMf5t8whR6B0QJIoiFxmeWxNqhT/XZ45OtS6FS7
WkGBUNKahNJA8dkkUUBZhLxybzmkiUMZjs2m+mSoLhU0br7QfBYjxp0EtMPZLDXRv4S49PBv3XB7
PpdQvS3O6paGk5gX2Hd4HrAGW8ZobXi/C9anMl4OXdOCuBnwqB/rVXyW31jvVHXZGjavf79rd4um
Ha9QUJzD4O5st72Xun4wIQotGxqVmnUD3dGuf3OUkA8nw0oBab2YmV4BinMcjvljJZCHFwCR5rAc
KZQikNbYxouJ/5nhnC2lzN2d/eDZYXy49l+q86CRap9+NbJJH5ACJ+2KnB2XpAw58P0hY3wPSxeV
V3bciR+0rOfHTWue37KBpDvTxPzl4y/JU4gErt6coN0bZYPHOaf9Q+J7iPYht4I2tOkcBE7ZQoOQ
nEdk44QP4XXQU+3NxbooAErzwtFtxqALdpcTjKFPw+c231JtqEuPwKUZfvDjh9IVQVBBd8MJ3j2L
PUtKsegL3ZPfyav2hkDhVYSI/Ah0zeULigQ6sgwlXiZQ1SzjefOw8QcfuPS/K4UjvN7Pm393alNl
KCkMjJh7QFN7MkMWBOpltoYCUFSjI1VGAMqYDokzhOGhBf2gVyg7SEG3ZgWXcG64O7vlvjoEVo/l
GjS+qahJuZ/qFnOW86jctEeMjmyxVmmWFzXQI8tE6HSTrs7ceaP0fnGhuaMqq7pI1x/GwGmd22m5
BtOrOniiDMLtQlJMnYm8vKYz7Qe2edvzVilfMWy5dHpzHAs2y4o5SU8oQCdWTjJadAsTNtGLVW6g
1rIZC8uE869V4ln4dORCl5nV9RdPdxO/kVMUtWa9jKrwGt1ldBTVY0XZXR7GKBrrMDdXFUC0Kwc/
SvI6c6cL22VSVy5IWFm8d+HUdJz/RWFeIp9Dp5k10qnH1wH3RxY298urEJwqcQ3N4ov0kXMPWjZj
IkrxfeSRNmjy70caZxBoRQ/aLbPTzFjbp7Jgzb6HnLk5Qwh3sc76czOSYunkWQncqyI8Wwwx27Im
bBJQrPOr59w652iuuQNaHqBHEJjKct1VKzw3OA9sWJ5Ubi5UM36sawE22k1nVyCWzk7Q09cObttx
lkeBnQ1XLtPpJC36YbRxacbPVAAcrqEcbXTnc3ENttPJzzRo9Ilt+eczWYTdCSEv0D+fsknVyQ2X
Os+P8113IeuwwzR0yc7RMFbgdjbBJoTgdAz59OGkp4aN7C/g1dAVIJj2Y0NDm28+XScEXzFo6/Xn
e1bWgv9h+w1jvWihmyneap+f7dtHQud32s9f55e6Erq2sJmtIX1jo2hMAs0n0oIskrfmGUh+eBj3
AMhfOKtwjOCfsfLKnKN6h0iUkoTOR6HEOfVE8sQqhOgj0SStaG4z586q4uFr2pQ+GmkrC1dt9rxv
ssZntp2sl+7BNa5hNIhG58YB3faOBwVHaHAHQI1nuhqAAXmJPcUyP6dRc5oIVhJ0+GmEQS5VYwJ9
li2xhBYR2mnEdx9AQTnKzXojZJTeISh6QLyxzvtcK0PwuYFkOTq2XrrAiEOJ0AxLD9sBZdqCh7rQ
mKELdLzt8E5Yjl9HOTG6+LsWvL83hoj9hcqzdHBt1oQrPDGk59ZiPsGlY9LD91j1HR4pGdwi8yMu
GqydGUBJH8uTJf98PXM/oUsEO6oVg8ED/1OF0g9bxWBcRA96Isb11O5ImAvjGC3a4goGzp5eBNcb
uimZ5GqdbfP43AaqrisaH9qk5+pY/ptIYmA0Tv9UrBbnkYiUVOk6AfXfzmxn08FE6DMSJMF/gRfV
dw1wXiZhh2NWk8/ra43+omWAn5XifRctUoY5u1+QjmV6A48288FYMmKnRFaUewjMz3z/+KkAMZIh
jm5V/05c9wx0aAUyKy2fpWDYB69iQ4lJt29pmn8yxhCQJfPJlC36BvXc7dEvSbv1qCRUmu71hm6A
2MW4V4T309fwVz4TGhIQtIf3mo+D1YCbLqgCPQXP9Loj3f/oeV8UXkF6bQxuf+SoUcAm1e6FHEu/
X8R2hWNaVXVps40PMOGvo0Zmzgt2C1T8SjVTplniVPGISjid/tGCgrUAEWhMspNS+JBF0tT03/M8
a+LlbjWSGoQB57irdc7dZTWR9xBzJHVdEdFJpYeebqNSGhMZ2z7OKBoh/y/0kFNo2bNkqUPLSSEP
y5f6h6UtxYuyS6uAUqFOxkr9w4vD7CyhenmBsDknuyS0NnE3xDX1xdDaQVGPYMQl8oDbWmz51qTo
YZmLtdb08W+FPSbcx+dvUEOfbYMKve46jdmlal1wlgCxP99RHbFfcrgGMimjqXMElKDtan/SC8lj
d1lxjV36+msHjf2kqQQttHQ60PzYWnuWoBljfP94O9X9cshfLxoECqoydxZgr0GfQyl3ufP58YwI
fi7xM7CetqmluR9sRBrOUhJqrKY0VpAiJD3nEvK5LiF64VLHrPip7qJ11/r42TnIdBKBuo3KEHSr
dW+bPBP3KAo2HYjpfMim2Io3y6vscleI9RZqakwTtkdzPSBUp0NEX9pBSJJDKlSwYQWRz4s9l4jX
/8w9nFj07mkVMzzaHMXZHIzjAN8nygmNZtcqVKVIEsyRiQSK1p54uLjdcGTNhSbjIy05C8wIbKM8
4IHGPgw4hKn9WhqZiE7YkqPxWNQPTz2iIEMeUb24bYingbPBIboMEPwq5svjQan+vwsWECMUblXq
LxEKYaODp6+4RbEbbF2eC3/wWG+RJhFWWaz3tZhmjwaS4frOUkzdgGUxP0dZ6mprFbhVrep3C4oD
rZXrg7seS8emSgRWBD0knlzh1paDFwa1wxjS5Kfhi3BzdH6f3KU11MYEsWOvu45zmJBU7w4BFKya
MxvM9fY5hDR2spq1Uzay5/xJXvF2gmwe8gjqYEgdlGjV+cTzXGzKOXrzUoxBs5nlHIfuXqvuJwCG
ic9GHbYU1zSOYqRbAIvA1F9oOrHnafV2IxasOYuZ+iI45aYJcCHjqUEBfFttJcx6ykRttWCDOpJG
Afeg67tvrqpAY3I5zdVv5+t/x45OH+DDojeRS1QAw1vzeMk0AnJxrG4wr5t7kdjls+oZwf0EaRI1
K69d2KStImjeLJr4CmuDZzGvQvQAKsIbYiz9uJJbKTMKu3SWRqvQRhvt2UXbgI3OTexqVh8MR09n
QQgTFzPkv+Yt2Sm5KkUYiJvMoaiAoYMuFmQkJtwp+T+NW6AbR8MDJbejdDgMJqEONCK928whSjuG
ESUOWSpDwh0qy5lARVRRWIXwGPaB+EOvPUC6n51MI1Buciy/kYVrCpa04izOOnMB52SzED4XQF6i
7GUoOmMUGcC/aQvF+zJBwhszKr8Poc4MmnEnf7ymTRdpfVoI1ftqgpriGEsDfit6e0yMkl+z0+si
nnaPAyUb4uaqm83NemksxSrO4yGRE3qKgqksWB5EV5uHc97V1/IVtnw9a45Af8a901BgUN5VY3G9
vweLmBmKEbPb5dcG1V2Af/1GKzTh+7Xugxqg8EhFLY51Grpj9eOgJ5Y9RQCFyR+hAwQqDHtKGNHQ
D+LLrgUbryQcJBa01RboUm6UFROfmVFwDtpPIuTHsB60y9nVgvY0M2zJICsf7USvLE+A4b2llVL4
MvlTIackRNmrvEtpe8yVx1yGAgf/9qQcO3BnXNtq9u/Nl8fvopItiZhT9o4WoK2RbyOT7YrZRzU9
RnGyqBzqGwvY1pWRCT71U+bSJlXDCKAfEA43gBCmfrFg7CkWHWfGI3iD5pkmCS4fHPaWe9lF+CzV
/mvoR6xJSJXsmx04PZgh4kk6AKKw3XOjyKotrJ2l8zuokA/PD8hzY1NMqmOyrOuVA/hFnT4tblkI
RKS35veZprJVHyLRTh9lqTY79nR0xg2ckUHbcz4QYCL2uDYkxZLH/yF5jHfuX63EYOJVCk3ANTSG
lLsgZOmA72tRXeSxhlgZTs4AvkqMzBYpsvvZpdDFi2Av1KHvUfCYl6XNt0FtgaEOlKUUrWnzd7ue
EblytZZAmswx6hxdTXxjbpPcJfiNa/MU34mR0SB6de9TurdDC7vHBMJjunZ0090q6GowHSVx4Sef
0mPBXpEhCXuOiMOH06viuvCCz7LKI1dP8cy3ThTf/zcsHoBliBQBjpoTk/2PZYbW1NbXzbZ764YT
foqqEXeEsMAKm3lx64Lfcs3j3i82tlRsKor88xKD/tBDXlDD96vM1m+dYrACepJwMIbzz1RSvASV
DHv/wSaWOcmENTy4PN4qwHax28tV7ZYcADVvrYiHyBVbmtuliRj2rTGPRVE7SeyCTT+aNubnOqy6
16KaMdBYnfjW9cLAsjg3j4Fq1NhL50pUnjXx9RLnPLFyIm4TLVaS4uwJ98teS2/fXsIuMsyid+ju
B2pLya3EuxLayAhCoNiVBwOBNuNjeffk2F3HR8eJKDbQsOfUvQQkTr19EC7XCnwSNK3ZMuvIVH1i
H3nTTs9ujIkmmZbU9+V1KP8bNUcutq6pF9juIC1ekUaDjcFa558jX4t/IcW3lHLCokADpavw99W/
CsNdvnOeKjAd9UOngMl3bxpKuE3uEZq3p2OD2DqzLdg0IfC8lnO8W/pTarKooQinFY7XlqKUqMsw
OSJHirAxlhXRolflFJcomxWLjJCPsGxPvL5oDInIW2QxdEZTrduNJTidL8hlYJnjpss+jXA4eHrp
AlOwXFWn/8tg7FiZSQUWq/eB+q6eE492JMvM9Dabc7w35YQL2SUQZ0sTQ6D+cZY2LniZjNs4A0UE
4QK4UnIgiJP6Kp+OrJw0B/+7gnEtN2TxOr/JGRl6fAVjx4n5xcNc/U1rceEUjb3leW8CQg7idos4
fXDEvPO+iSQseLFqu9CF7An5hUhC2gP5Kijnh25Z99TfAclnsG90O/CoSmU2klofDzmZK9IMVn9w
aHUq7iXlq8go5deJ+DzBfqLaggf+UC6mtZqFbE0WcI0m8Q4at7RcxJU5jrFHU4KQOeNqQjUU+ue7
tpJAT4mFyp/9U41OC9JZ9vqBDUoTolVJXLly10GjGP5IO0+J0C71rHi4wF/sOO8QMNXF8wnASHtm
otDDP5m7HZ4Yxa9FnEIUkHL3X6J0B99fKT8jpJ/qqceNQ8sXsuerU5W77hCBqn2rHdfxOkQmcmm5
TJkA0QZmZPhDsU/NEekWCLGxl2sH88RmjCL5rb8o73+jO/m6cYdYoPmKfUJbBIMkBvj0BL6TU4BJ
GTOFsPPTsv8xzeBRvLSRqs4itRLpsk0HRrFVi3wEdmvVKZzXgN/K3NHCSdNymX1Z8//RWGVc0UX+
jof5KIAUkSs9XoiQwvzWtlks3CZJvkUdm5zMToq+O9hPr3Q29Ry3rlcQRx4R2bi8YoabNMWSGGzU
64eY7QJURhCTirbHTioDv8NUjhtT82yeGT0Tnmnd7MZexMXRb9/C9lL8stInz0E1y5i/JsGgLbrB
atIBU5QvT9eMOcWbCyUL7lAFPf4nQnGYIleqC7Y5aNkWV09BheKbtEicOZeekzP+QsT4kXEV920C
wvxxGDuAdUMrDmynIeeemgwku1DUUgFMpQ+3DjG/bL9fjRmemiqYSa1OvUI7Z8IxC0aEG8zYXNbz
xA3gnK7nMJ9/vpgR1gQJhveG70tEkOwcWRmpd64hCJWgaVF46yKIVsS2N4KiDadCqQfjNFZweug8
I5Y95lQbFtYjsWt7EoT3UQ+E+l2EQ4ZFo11u4NXe2bwCJBdKroqIXreiais7avh8jG991JnmOQdV
YssKhfl0xg+LVJ6Nv3/xxgvUL1oJTxk2mQI+hkXdXXUDSM3AKKrC1qAq2AK9IPNJUDYAVg2FBket
LRuh2QSmGZZy+iYSbuHhMGdUeCI1WhBo4UiXuvHpFCVN0rDsihAhdrNlT5s0VWWxW8lT2ivoM1zz
Klecyp9/1AEk/UUbyM09Z0LQaN/bFxgeNxSWtp5P8Hx+9Q2xF0RnwMrGinHt4abnyHPb/ZVLCGRV
qniFICdGGBuM5IocMpRSO1Fqlg9F1JaoIv4XBY57K8HheWYYtquUlB5xVK0ZC1bsiuJmw9apcoud
cQ6wFJxHIdYlP7cjgm/MMOPGOVpZJDrAL4VKZz3M1PjyUNEPL/rBTAXhZvxft3ABQDB5iDLJKqIY
abHxE1NpjnYrCPUghJrVpZs8lK2COnnXmF31onxg9pEH9qJHQJU1hKTvOiJ0CiyVWcgTf6S+HMEg
48049DOSKisEDUJpVewRpIPpyOcxKLl9v+z3ATFbqIjbat/uP3YUbNPbkhIi8lswYQlWRE2mVxf/
BHWft1o+vJ0XumHBq3rdmGa0SciU/OJPZKYr6XFz/hx01y3kONoA8HySJLW/GKspml1TPg0IxNnm
wvdcsxhru3INahWlrZ2XMmm5Me9rNWCdiTAAA03IN40/vjkHqfk5EockGjr+9pBMPC01tNr0UpYG
nYaF9BDkKxgTvPXC+9nyjPnbkJnO2Dwiq7uAbgk6yQp9Z2eoAMZYm7YNXgqV2pDknwGn/BV3YmgH
q+mcZoLyV77IAFRuRqBt4TrbDWhdCy4Q8kN3xfB88uso9WzVY1nlRyS8sjoOj3cG4aTBSL3FtUv3
OgqtVmVKt05zqpBZqL4eNebX2PVo5onmrFmluRoTTkVXLNMS2UxEAfDePQfjHK3lhGXafPOrVNQ1
EFMu7E7uGod3jaLA8D4NgzLV48u9N0blmBqE/OyUEfNr8LR0hZvVigX8tSMhOvc4N0JZeroBxQDc
AJ0DM8wWP2jqXGavCCi3FOo5qeVYp5PHie3KRFk85HYD5a+1Jk1J9CHoxlmToYgPNdWfCiUek4Vw
79uTVtf9LKRcT+1mp/De04EkTItaOcKqepR9E88sXuNZ+oFOcrL8M7si/oVPkbVSH1fh6QG8yTVA
7JPXVlKRGIgg+u80EsqsJgnoYDr3ikyS0QeMdz+KGIZI07EFp9WJKXqOTkbvQUogpLylc2CVXRTc
979KVa9JC79Zg83aFNvFn5tUYPQKoDm1G1l1O7pWBoQADpE9wPULWKE+iRT5MyVDa99rIbRbYwTu
pQc+NlQQ4+Z+sevuDvsrQUectEFudlH12p1vxI/RI2SHBeBBTqw848ave1og2/bnmFisJPnfWjmy
9XcU+Kha2y6yxzsN+JpWBXZe8dndFEzGf0AbfmyPXjVp4b4rD61NCQ9c9+QP0lWSYOCqZCrBf6mp
3byNY5VoC81n1XgPGcOOwZwk7g/aQ/ZQ0VxEXxscdK7bg9ejZNAgl0adJVndd87iAB7zhEzm25NI
k29SylDqZvLSps1nPiFaNcsJ/SwwX3A3a4w/nEb3KmIm+pyX3/hYIBgGluekCGZc6S/8TuJD6FpS
wrZdJnznL1ufjyJTEwe3e+Idgc0J1r70CRBzqHxjI3feUOr401TRBuYeJkHZYguNBASSzP5Al+mp
SRrjhBKvzjKCRoW3D6i7Frthvu3YgN3bjEWN5k76nTaWnM3cqSdSMTegreKua5bPSOYZ0UQTRHnI
o2TFAp4TgNy71Fm4voxO2kg2BLnn1wi21UP7XmNnkuTNKeBZUNsLlWMnM7n8WqA2CYAxCtK2rxJQ
/W9sFwaBsSr5/vUKHcGJZyTr+pzfIu06OYz0vRxlJhux7MoBzIJtAX8t++8/ffjWnj+E49ATBsa9
vzIXTr6dpoNRya1A0yhH3J2/pOzdg+eyJndFmZbCDs7aTjGK8wKI8FgBgKZqOrXz4I/koDocE7ec
+bv+lxfL3F4XBa7mBWcw6eDKWe0B3AH4dgmglHFE3mDr+KJJ4o4zw8PyuUFhnBO2QghAvEhhkNXU
1hsIw/CubE7o/sDqWkRtMOmElnZeKNBf6qorg8FP+WhAiSr5JRXAn9S3myqs3y562Fvwzkfwm1FH
RUOPTguZTPY4rbP7Te5zHplNm5lfIpdNO+i3l8LtueOZwIQvA7Le482ZaGZ0/THHcmEjNEqFNLS0
rF9JSi8KV2XrrDlzFt2kLZTYeJP4UKMk7jRp8Mm5i+DsZhQ0Jzq/n91La+f9bORsNP8MZvkNn52q
kos94gixR4jaCwJaGs665oJtFOcqjjuU/CsLRko9fE4mu+r+CxORNjSvjGnFhtHjgB30i1m4erjy
/YICHc5JKFqXXe0dDVmLmyQjUuqTybY7U3fFIJqIrw3lnJsenJEdYo4lpKw6whXI1VHLNShYmWde
KQgy/gEmOM0zXEPwUe7kD+kBVyZrC/4XQlXePXtS74L7PK1gJWdEIbaltqPU8QTrk0IrIB5134N/
5jqE0ua/RODsV+iQDRNfP7zP6TPZZaa+LtyUpEfJsERhjpbojmbB/QXpZV3p3SGUKrYcPVhnrrwb
s0M6qOOGCIlzPYFeIfar+fmAbJ3eXoKwQx4fwIqKL/4yiNcCrs2DFRVBGZADv6VmHEu+NGx/gxyC
9qZ/qmWLP4/33s68sj/8b2qN+zbHbrccVqgkrAWkmXxRgzABdtpnEqEWxdIkUfV67FHpmsO3vfRQ
EkYUFL+jZ7YNRqfX5oyZuyIoX+Z2hNOMtx0lh9hMF4ZncJtJwu+v7zEMCX8BXL/3YqRffQG96nKq
uC2RO9VFSTXDpVbkEiDvBWiPa9AIj8KZmFdIy2t7fm87R5hg8yjDqPjSo2etarl9d5ez35JnEtBK
yBaxU8lSjil0QvqaysL2+copcEFznHZ0A6GczFysr7OSDRhKY1z1EWPZ7GGEFVbhEs4VMFs+9lka
RG/WYi2iDU/RfmMVjC1GF5Ee9PYTOR5CwxewTi1NFVbzWtnGDIhrmyg57f9HB1xqW5JxmD/Rk1il
tquG2xUKCMUIvzY6uXvLpYSyamHvh5P/BTi9dVZPkum4dexZI34q79mgbSlZAmCvc2WAk7Zfkw6w
yluYroDaMg0mf9Rq1Z9aH8eWpbA5KcePGm/duH02S2Ps6zok4uKE340T+81xs5OioCPClwYvXKYT
BEg1jez86uNNKNnH9nPYgzNBdctUeMKL8unU3CJ064THcWgoeMV2BNXa1ZgjinMOFlx/S3o27WuS
kyjhoKJnwqPqTrfSvp4bgA26OYZx4zFJ0YCD6gzkWVl6fEi2SnP2i2OfbFMwRBTiiGGKr8h3licv
v2WIa1t8WcnXOoN4WoITlT4Eexum1KIwEPwszUkGj/JfpPL0T53YQIv+bkPzRz2iBLStOo3JpWrt
4mDaHugGLU6NFS0efF1IDWuJmHJ9ToePoSmNcJtS54HdnK+5BuBb9nanmuTxHHtp27pKBcdGd34j
pGr7E9PrjYXSWeXu/Ry++h9ldISlqhDmr7Ii1kbyCO9jWp6OlGd6DJJi403/MMrTtmYFdClfYXTy
q8z18dKYKDLE3CHBRmxDVsy6+fWKNatabFALeIkh/X/YpdSbj3afQ0wukUHg4kjNyraBNg1Eayjd
ZANBizlSaJGEZ8ApyruN2H8dBCUridOsJfST40xt9xcTZKiq1Wgkd3pkKr1NEVS5olcQkI5PEbo+
wBYcrbHkcUmCGYTLXTzXVUKnvQUxK02NAf9Bb51OcG2g2ko/WZMUwyoq9+J/2FYdBK/Gp/k6Juo/
urzkh/jDCYHwiWzP2rmq1qVd74/6bRzuQc3GwAZpDh8xof9zh3nW2c8rVLdzDay1nBHzKJ7kpMbL
kTwru2DNqVU3WpkL2Bv6iUP38UT+xXKUZlOmx2vz7IeJsRObd/AhaoO/XewvJ7DPIJN9EKpyN5dq
uuNryzNkxmwkvdyUZ1+2yQCg0iGng8Q5DpZ9uUafZDDo/sXqE87PMJKCiDu8heYJsgl8cobvyq8o
bofltxW1ardO0THcOmIarUoG+cORBejSDDcnTOIAhQ4nq7ilfzTeVRcxuxQ7fy5RBDbFrl64RT9I
O+pe/eLxKMrbFSj+vTz7QP2TzidIVfpZM71wwGNpgWqUyEuCO0Ke1bbjhtIz2AO0KtabijHfyChR
vfYO0TMHNdVeI1hILBX8H7Zh01plxY8AdV1QISNG5YZT1Y41zg9I3ecADggpDJIw4Bf4cMqitESN
PvYYdfMSTvCfgojlkrUIw15ut5bNpnq58KYnq7glIQVgHLt8Un+OpcgU30ZDIBYBJW3KdDjQSo5d
m1zPBBIeiRQN6CIbQsBW2folL+81f5MPxTTzxsbvNahLV++JOBIPBlXoA+gEHZf+gOBKsE0A7JQR
I1LBl98jYObFhv9ddfgranzfQ8IkO9LVbg2zTG5T/2k+/S3pkZy7j2GZcADN2lkEAEljLW0lm88j
UIHizAMcKIMrmXcmrRQ9H4eU1cIY5uueCFN4hAGDkm0D3IN+41MJ8Y9NYgfvmp62MrWW+UlsM8ee
SXsnMoUV2C19Tat8bA+nBJPMZTP6beznVfFEUYgginsmNlaMG4rmMBEDezaCklNMcvuh0nyKVlT8
tUJMqA+t2QegTu2hQ9CW/TERO6fmMFG4P5NZaZeRfpx+RnTLzB/2vosHeoLHvacR39HWZFSIi81I
IrvxxEH7G2Rvu5s+ldICWEtKvHgRvBeiR3Oe/KAllqwLnW8IDknzCdEcKHLrd+TFH9g7bFEasr0t
u1kH125zTBshVO6CoNKQyzO4TMT0C10JF0LU+yqrXHq+fKs3PETxwEDEsI79GJxprk/okH4AWVmH
ElE1IJkGiKctYSDwMpRh/XR5rMIpJgcHL//EIDuORKSMTjnSzoXBsQ1aehFBE6z7pGn58Q+NxEXy
2YShHOjvjN40h+B/HYD4JHpZUrLLiXrR6Np1ZUrGl6959CSARdcFloSTvre0JRDg2UWuKCJF1RdZ
z9FrYUJgo9sthqPht2KQ487TVNQHH2FrsKpWO/moif6gxzqhx9/o6Wuhy00t6twY7RnC+8w16T/K
0gRqtO1aJJkbqcxsKjJOQV8TM6mNqmhUXnr9JHxeBuFrOt09Z8jywjvbAs56xQBlnu/lMPE4aTEZ
MAEBDCHiQYtmIPFNluZPxs6YQmVVUX/p/hgV0R8IYb/XLfNilBlFRyUHPzmioWeyuGA2bXdj6iR8
sRix99od4s26Zvs5QuipCwIVQdd41q2dsL4JK4OTWCTzO+Pqiq0FS9bQ/sBla+XALKPWSs8OQX/k
4RnqRmR74qritx1UH/azevMWXRriAojYecxWYicLAsvy7eTR2kV4HL147y9rV+zwj9OqunN3a+8c
x/T1BWXgzxygMRpwnBs5a8rtxiUHJCm3yw036zDKES6Ca1LP2Gf2fSIqBiyU8Yv9M6NGcfLiQMFv
gfD/r0DPX0xgdrCi4hItJEc3RVllmw3dz277lJF22UYxLe478a0D4tHqOHCdGA5ff1FZjxFSN81A
w0rZ+Tlf0c0CaloGbo/YRPzh2IX3N/qQS9YUWtW+Pi82fIu7aIXcdyqauTZw+yVdXDSxgPGzJH1T
EWXYcs3Dt/V1C+1xfHE8IAc2TR9wZwVviCDcuc394PP1y5wqKyQ0KYE00KbNUY+4FIUaePs+uwr6
xeZvkUkNgV2RE/c2DP/pteuKz3unqQ0safWbsUojPZHATqzDZvJVjx/OuixqwpwCKqXZt2TnUC+h
XqxuG1cLCjHFY1g1y0m48edc4mM5v6ImkecINOP/clkf0MKHiLg3l3W8/TVOEMxxPrj5h3eEs5Vf
rOuKyFdHE9GTBkBcbzJnrM4FdF+jUv7mRlg+4rPSLpzeV4nWvL3UFtBgu1r8xjtoPcotey0Qz1jU
ockSxmHLWIJRUqf+v9w4TF1VouehPnXA8J5Ppqs+QTm/cZG89xlZeWExVZ4jakx/IocGw13TDsIS
qNzVU4QQsAQF6RVZYzOJEuhCEaZFiJkLdWArScLQNcrVaQNFG3PWwNF+u1LIFiU21puf3g+PspTS
Uy6PP63mWoYd0rgkOHPRXwYAJ50FGEKZAY7GcICpKIshN+CBFqMwwN5ftKLNjXgIB2eHMpIGg4z0
uoOFJ+VxPR1sq26xCHqCKKYBADtsNukAgIpCOS9MV406WNyY2vGnRglev6+ppQT521NlpeI1R6El
LwJizFqRhI7Y82C2n0s4uSBCsJxXZtv4TzvulxvmJDqOzJCXVSoOlbUwmKdiV/M8nIE7F/PV4lPq
NwaLwFb+ZiZzbLoJnQR308NOyvix1In9nkeeMaLRKEYNGLs9Elhb2W7UCWWrfs5iQ2aAd/eVcK0Q
C1tLEvzy8FZQu2orUsNVLoegdYUgfAnxSC89Kvt5TVz/tNKPA0P4LiJht8IcUmRdpxaDFfb0UOH3
pSSuXj/f1QNC/rmcfWJtWQpLSVk01yRe6qO3yi3erPgLt1koQ6ufcrl8qiXZKaYXyIEeeRGPxwJi
2PIEHzSoCXxuLYBvv2HS8m7Wg7xiftN6Zg9rkSb7/mqifG7hm7cada2soyhMp/rnUFFw7QDBpqEr
vvwXZsrfFX4k+6G9qsgMKw8+jTt9RnEmz9+/QT/3sBeQELlr7MQrbPZpZrLgxqCbafqLHBUA/L5G
PXZpcq7vfO8SlTvOjEmYL73bdU3/U+pDzWpOItb9VQ6VktQg4sWbDMtlNGH7HoiLbyD35QL58qpH
DNQECZ/FuWpcm6KuO9RFS+V/kP1s1n/wlyEMS1c6w5fARIoivrJa6t/zdgtlNu8cLv/Fx96V9FrT
S0ijQtsrBm8/zuk2Zb4LlXyq6XY/byfMN5B1lOFx75TvMrpYe+miON7anSrcjGia50+9SfiV/5tZ
of/INhAWACDe7da0Fyj2HC1lNLJUcUrSZ9Scys22R8E71g/944+ZuzIOL3o6DC4T7YFIO6hP2nVN
0OQUn2hh+7BVxR8zyf1AP0vtUsRN4tKdxEaVgY/CWpXB/mbLtU0VeIa7oTCHCl78lsorE0AVGQuh
Sn/i5wwqYzkE6jQ8K3+i0LRGiFjO9KpQQghJGHKXMmYm2NJqod4B8RWirBQ3DheOPp3hGFOvrIfr
5smw9EvbfzR6K6WvXHruMBL94Jg4RzwiHJncPfg6R1uAuSwfaOCkU1AtNZtFoqA67Nkd0icZiP8O
ksjsS7wWLKlbHCM/ZdPV8hiRFBQHeT9GKDKyx870JCITfhuwfSKYBSlis9kkGMmw/WzvvkFoTpPg
y3tiKPraORRhT2Qv5xfdv13kUVsaGxEyRQQFCFbhN8k8KV4TyY9P14x1WZE/ebLd0xbeKLfWUCn9
5UbJFOIz7nXR4YRxl1wR+2JlFNmTijsKx/LPvR3DB2D3tiVz6Dalut4G+ZOT/9u/ywjltzVieMWp
d7FPyP3e6srVhF4eHbUsA/3Jh/lgdVxjbYh+jTuqEU481n83Oh7u982A4TQzJWvCgS4LNIdjsEEV
PBSY/wGUrwVLec9jEKGIHfez+34BXaRYD7fh+VR1SO441K6p/XbDh49Kgx4gdP1Id1Gw/PjnYv/1
TKYfaqLGoiORJdjDqqTAswzwpPguk6gXAAIvrDWpRFh1Ip0IHzgIe/JJgo5M6C7cIWsMs8U8aLrP
g6PqT4vNybRrbDQHOvhworROJEeiUS7ugpB0qM64HYpv/YrVVLGjRk4cNV9Jn3onnjommBTlrF69
elEIKygT0NeHp6Z2v1VdDK45aAn24SKiMdxqV9DWCS0C6cv+btmrjRei015z1g7hpBbQcoXqJbY7
RIu56ChfSnzAQQgmhRWZ1YYEyzxweoi+NHRcbBKwCaxI5hsd+RUFg++8llOG/5cR+Bu9Ame+7ECI
kL+8X0OpJOZ8j8grQ5IbpzLjJAYp0hkZlTOPycfn1iPFZWxwmgOH8lb0HN7OLUOFdd5K/cPmtv+4
ij8FZTVm1Jr4TIhWXx99QYtJyTQ+SWR2GL+8mLGyh6v5FbTUejLMhPO1AxNks9+WQ6vhpjwLaj4h
TLrtV8gd9ZIBPtS66+6TICyuAPqzS0vrAFvDzOHCE8HKSGtvpJL6k0yrvqiLIqNmbFfbKCyQLAOv
D3WBguhQ6ENxhQWIWPSAd0sOIg2S1luoWjymC0ylSSDNlaKSiAKcza+wO6gMLnfudOXGcPSpACoa
i1U08rbW43kO2diL0A8qbx1mm9H0KgyTdkbYNF7r03usyrR6FYAs0ZrbJnnL46RKhDQhxbnZD9dg
LR+XVjWEMimgLj/gvdV4G9jbD6WVq3W57hjSmYjlgWZTw3nuHMxmv7YfmbsF89qkhDJOmqRcKKxj
TH5l9Hjkv5QzQc23dMi5kkgNLD4RiGz5JdprXwbGCAWZV1nBcAnVHwWVVRD3E3otYk/CMpiQqI9n
iWZjpoiTaefSvwN+ZvVQJ2M1AnA8VW9cAHyThodLzewvIf9p1JvIK7azpVTB+FxgDhYxRlbb97+k
re0p9+nvnrtFPp4O8CvTa/5vHfJWOhUMHcaaFQ8Vike14o6OhGqCY8YgxNFKqMHLb2F7o00kUfC3
/U2Jv49dMde3epWJhXAPGfttJrbzqsrE73T12EEsESpDSXXpEs5UcbFc9FB9dud9IuUmartEWTQJ
fkvh/KTPMFWR8p9Trat9ufIQYsClJrbH7HLD/SFeJWZC8SbxvLTUUqCsOM7ztWc/8dMLGaTDSuDu
iGvbx0QtsG76osgRFJJSfCfy88PIUgpdwNlyAcmpNiWZg3bFsltDPT4Dlr3YMUtWpbGp0hWkA8u6
mdauoONGyfG2Vtbdbq3ZIP4W1igUb1tuCVir9msjwmH7nRZMgDUs7BuKDHsYCR67Zx/bwRI7+CBE
qhh+9GmZD1XsDZ+gsCedtGNFPp+rsUpxOOnnGp2KRy4GsifIoyjn3QGXwV729r6H1u2oPHlwsCOw
GjErFqxOcAYIQ+KKjrpK/oTF8AymLckc3THINIhSfmwj1s3KD7WvkwZGJ0L2v87yEca/08MQRfg/
OZj+R8Pmey7l/mOdt8D+uLEMq9dXNtM33Hywr2UY1aiM/9tQvW0JEnQDIu5bPZ6ps3mPpiAMo4oS
Agw/ulelVMqXHUGNayA1JGvwsY5HcL1glIpqgt1ozrTAiuJJHxrC1H0dZIqNWaH1od0YbX+fndI2
XlhwtH6XAtySNp4zKpQdN9Kpci0+GYHvnjQeqhlZCZHshqkwlVG4URkH+Zqd+UMflzB3wYfME5S/
y0uVyHZLrgE6VK5m63YWgkAZZzHCw1QA6xty4uiUBNUAh0FYyO+HdkgiahJVFJNDXNH2KIw44dS0
Xn4R3FRxkIOFqNvm0tkVTqR8yAoJLQLedLh7qOB6Lj3F6XuhJSFvtxB7/2t1ea7+cVEBM+MrA7AA
L/Np9+61XRPqv5jeuwmLWTzsdYa2SXfeSlxzZRihVE2iESswbFZXHmAlFput9kRBuIloz8W0PH/I
MSkLFjw05/KpOgtugUCzo8bX4IOwc51NPa+BGwGIB/ok8aVNqQKM7oBZuXrVnqueS1fUJzcjVbFi
avy32mJxjsaAwd1L5IF3KvVHrGDA7z1iLZCn+mUiHiFxwNmMN5Gu/VddPZEHpgPfx4YWnMJimRK2
ld7sOM2ddCgWrIdgCtQBkk/+fMKzlOMju7MZpToRe6C+IeMa9gSSSaY5AG7tF+benCS7BKLxtVGt
T9wtbtReoNNbaEsvF1FN+11ZQUOv02QPgJ6cd/75d+8bRbKhRwRzqa1Z9cLw0b/TQ+V1GSslpGTZ
etJV9TgFZRiVdUq4lmDYKNcI3/JAb82PwGO8Mo4KJkoE+r2nZnzZKIYC7gbgYSTVmYpxm/riSZ9a
onq+1b9j7sMOr0NiSvxiYufnqSNdWYSb9bVC+Xe+ACf9FHJOLTzVP+9LXYhzKlRWHPJT8s7zm6iB
aHte7Ow6p69/w9RWyI7gjj/XjtzF4BEmRFT6sIwaxb0w+aS+Xlnu4nnyy7OBp9nAzGYFN72jt5Zw
RRdYrqY2SZ/WTOfRqqyf3FjcEdD9JytrBwZ79YIB5+/7xujSG8Rm8wtAHtwcqRvXIMFM+jOP3Zcf
lyGgiuOdUgUzh7ZvPG+PstAD94C+cyon34SCQSV6eHAWnfntFgWyzLdMqMlW7eOtFaZ4NeYG4cOm
NvGU/FbTNmHtXNjQG9oDVuy2rIrMib0GhghGvDdFkoige2isYzT52tdSDOvTN7Hxb5XZJKeuOaD9
n646R1pkeCRG+lsz5EMBoHElO6Gar/UcM+0Ua/6MZCKo1yEpCcDYgoFdgnRUnTGGeShf3qw0+yM8
+HEB+nDRAiOgjcXbDK/eifHha32BD/udCe/W+VK7BqvR9Jx91YdXq/te3eq5MulTQtSCiwGvq+R4
sa+fnRLVyVEV73fB9oMwPvBkovwhsLkQGQG0oblNKjxstZwPdaBkBF3dYX2AA5p7WnsFL6iTNB0j
Cz2L70mPPG0uH0Hd07OZR/VvM5vbmq0cxejvFb81w79Gq6FxAdLNzCj1sPEf+eD+zNtIHL1KZLrg
F2FFqyrrHDps42m1/bE2M0pPblElxzL5Q57d0R8cvxbFrxaBEAdQwxlutbpIWxdPJE1sFm9Fx/j2
kE51LLK/P/pGW8gjdGUantBAvgh4V6eesdtNxFyYjJ1/XxUdUF03DEDNd0PhKqqrV5ff6f/lFsIO
NelYUKzqOll6vCo6oS/94/w8IJS1yoHWvAwizmqr61yoR30v3DUent3kITEwxRZrzOBP0wmLszSR
jD3alPurDsti8hre/ftgOnuuLVQVaIDzpsCRrNSGLCvQjheXx5HFoJxXCXzO3XBhSEh/NMu1fy3v
W22wvek7FAHGfI3HktihJrwT5wUA58Pg6tjb5c4newBys9Uljq0+2dijBtugKs8OSZolFtD2bEPg
iwiImqoPh6EWPJB1UGvSg2pkRHgva7AvMLZE0ik5Mrp2h2xKf6+/LMqWJzP4Wk9QchU0JmLmKpw9
MgF7NRf4NSlm1Ft7pXjcfLnSVN9BVgd9ohhsZ2JBsIFEaCyB7A8agvsL44ZASIHxaRkADErlR+a4
JqJTwunIL/8kdWVbmhjc6bhWpFB5LpaEv+cDJDPgMG0sBCtcXatvOAxpF0fU5ou9f6+h04+e2N3+
Jvw+n5zOafGsB1CsVT7Bp1Vif3rZh6HDifIaFLkztEeTDU/tt4zyvmCP4B4BH97lPxmLxvHu/6Zt
9ULIyDdACb+OurWMn4wQ0q7xzqBNii7TvysM/j3+2B4UmYx1HjOhwi+HYmlgwm5tlzNF7zkorGCX
8/+n4saqpqPEMKvxymFTTHNmlus6zaYs+OcJtzxlCZ8HjdMHKBWAOr2b5xUMPOFuz9KJysg9L/wN
+MjbLVktL4fZhAd2PJfytuggg6KWbhYOlnsPECXVLaAfZQqBq1UKf5gi6JJTDxg6IjTQdY6orJKA
OT4RRwkJ7+PXKJ1LVcaETXGmAfNeDNrnmXV06GL2bolCCMidNKsYwf2JB0Ba+yHDX86Eg+rYISvI
1vpEV/JcFnGU/q/HXAxLEBkOn7eZMKyKCYJOpJrqpYdBl1VKZiA01n2eCoZTxosrfiCz2JM0woxd
JlN41Utlt0i++KiGOnEnpppvKEBRsg3KhV/AqUCnlhn2X2iTbW9NOPcO9UOd9LdiKuG47/0mzGhN
HkA88GfYCko4/sChyW1fk0h1kY2nZBRcSkFdgdvGVVzFU8RoxZ1aGizTSYtTXI61agbT8JQh77OS
bJBLu5xCGI0cjJtc1UjU0JYI/OOyUztddmOz7inE3AHE7DQ65+QljyFu0SfoFpxYgL3JM8VGeG0+
dI9tPRtpXl169PGXDX1sS5z7rDLmko8iN27B3+5bYCRyMYc5uTmx13WqkdGZT4jSAdT+5gwg5Bkt
LB3o+Vrhca9vMjZxuNXr3SYHIfbMSIEm4nWmhiww4mvUNG4EMSuIConCZgk42NjCLzCV/4MtjuLh
rW+ZEw/yJnMU1VWQUL7k2TpQO1btsvOhnRP/QFU04eLdzV0RMBfYAm9JRRmrPKBJfM3rsfV3zrYh
9FnD5Q/sL76pEvNBhAJ0waBDCs2Qs6qKMvGfuNkM0yKFyCi5ksrECW3MqPGUJueqhrSESHolnT8g
45If/7bncypFqoJgmCE//xGlNas2qmxTMpaNoGFFq7HC3Ig1yeBGPs8nTOO0u2fE2JV89femTQZl
NqL2a8nonKJkIdfT/ndsdepe47cJcx01VCPyoSjJPyCEXDz+Vha7UeIS2TvCiBgQq/3Y7niXxgqi
/Nd0yse0Cb+aek/47ClVJIGADZNNSCVlfnxkc14LuHZ8XNDY2dSSliw/NkYfdnaAEYfUz9+MiYng
FQmHoc311eZnwiaehGwKRygXrqwsXdzblfQ7FLAUaq7twhRA7IH4aGQXHCdjCp4gx+cWH8HEyNZW
8Dwxy3R06gNUjssTLX0dQ8vJaCU1SiwLEAXlcjhcxZ6GC0I3R15ktkKn3Hs2RlfTR3tTx69cuqHI
MHO4xjMo7S4ghciEoo0Cd3f8H8ejN7mca5QkyOgYvPPnmAgaZVtmpT4Pn+II2wxqDGgDJj3I2aNg
/r0c+wQxNbYdmruZeb2GYTaaVJwU17/9VIsQYJmFJfdcX1HiJ8VZCd43LzdIegAYi3S9YP8n+ywU
FuOjIMfSMF0ybcTsYVBlto0o9xIotHQR8GS1rOehCSt8NthVk1B087s5tJTMEaPhcpr7QS6AsHGy
TJr13Lu5SxLap4Rs1JMsSB9PlkPKmg6bmuHyxlPDB1TvcE4DPoEnyuLMue7ztp0IfvJVXvwkmNIo
Jy+pfWIGpOONLjeA/pmsOdrGQ5Q1yUcWvOnS9qNt8k1js8OIWWpCjZcg8/xmnoRQ2YBoBMWBNbuC
cQKm4qgzGhWjfahwATjD+a3FjjgKtQGdFbPIqYO2P4qukBkoiNmGDTGqbyQot0pV1CFrk8YuuRBL
3OjMvPWgsCi0MnQgAaLooY1LV7AXBRpdEPdkEMinwqy6Sfv1yxeEOyiqzFTVV72dkk5/UilYbyoA
O7rgstVLjj+NaWJKUo/elEKfr9sFFmw3JmHEzHlmLNo2pnagAvkZRZH8dPOOOlizD6SnA9Y+uRHv
jaCoKDbY78F7FGjZr85oCsv4XnZt0aZfPa6pRRQiamAusyRPWGxxt5YtdbSThCXI6Epzq+0IOWin
NNyGAT6ZvL6sr5JGrQCipWf/LdDOM4b+wGyss0ZU5Se+MXw4DAD97RwMolNv7FYzgVow6hNpBOPj
YVvs1rnEAjLBrM8jbXnuCTqjXI2ZmHXlOeKEywhdMK52h6UL+xaZMJkYhGXuoacpMb43dTjgKXoQ
prc2dT8wFLPCyCRxpGQNBX0w66ABeEhxDut84poSp4UAORCjJ26bmVmvd4wJoJycrLhPnID6mEgA
WyMbkXaigPd2vzwO/IsW/c7zz2GvCna1RGsycEN9cxBRFE6HN5TaKsKmcH/hLKkWqMNOsHKHTZNE
sC1d80FdqPZJh47A8AB6CkhHQFTSBpJyY+3UGwZrfyUXaXkee17nFBuA2RBabAGiK/iWFD/cfBb5
EGo9NeraOXBaPOyeh+23cjkZmjtueR5n5pbRfvFSsLao9XsUpY/ui3GRDC4BF5e9aq4KqEXLEfvr
McixRy28KMfdLekLpoTKXsjXezOcrpDYD4CorW2vofMn47cbY90rSLAHRZRHPaUjlq9JpSOBcIED
ZTr42AMQ+tF9OmDGR747E7m8WuZ0c9MCi4hQwV3Qz00OAl7gPXVEivL8zK53cQ0ojONmsDziDkiP
Lg7z9IoCCScJ07jylo8pcn5T7UtggI80Pm0ohkuGE9iZLSpM1FN4XXiyENpK9Niciy82FipxudFF
vHjXN5VRejy/GybgQgN9Bg7gwi+xnYsYuNcXqso66ENAZOe1erXEr3wu64YhsOZLu9ZS8QteqE9l
rP25IVebJrLrp1+ZY4+NvcXRXfBaLdTElaANiHarS9EJz6yFgGqSRG3b37zFqhdbw9CpnI7nOkcm
Ktmv3KjCpTzBfblazyJQI5n2IwX7CoQgBTvxIpwEHPXy7fDLQwIR5RVHXdfkN0XSaCmFdq3pu2qn
/4dAbiRLPJml453pHD8rbPkdI6M4XTXiUDF/AKwM4VUGHbHtXG9BMKO2cxqFMkbM2pFepLHc7tRA
25ACYbyWH6m4d714nnce4GNb6cgNzjF1T0oM32F5G6CrOxoAdqLfBLGpMzoGBaMMGO93HwfXhQGW
6XHikIH9JcSP9sRM1hK4TSvvsrSZWSh/DNlL3gWehQTnvDDsqJCEXTkb/BvciAuLTve4RMjBruDu
i7OBQv5m2Sqysx0qr22B8RyWNmOk4ivvQkfF2t/9OsoBQrZ7XAUvXxlfuFBrGFMlka1Dnbh+qiKD
fFBllArlP4uuwoLQPu8u1T4NE0HSvIp85xooLOm+Nohcmd5rOZkiashmh4PDWLTPiKY5Rrxp5L7S
Wdqmj5ULf+ViwXi359ACfK7P9jVVNEI2QwoDvqBKUF0v3XvH4ewYSB6+yYljuF0PlwtrtnkwtUA7
GubiwTA6UnuivL7dg0koEuLJazUMZy9Z279Sc81IjEtr4+SgG/oNdRGQcZlp3haxzGbxlGqkJy6/
/1/lfo8k3VRk0Ewy6ABv58AImH+FxyCGH7NJ2tHnqQY4ntPFyaiA3zbIpxiUTlFcLJag5MWXeGjb
Gf+BQzLoYt1d+bkcYS3MYFgyIS9UT5FtCUc8E4r9H1XNyXaIk25aNO3xSY6A2gfaHaL4aCicGr9E
pLvF6gjlodLYoONFwZK6f6+fqWjIy413elIXw7IU0eP7Z/ZjhzjoMugAT8OHxOHOk+jRkhkl6jDy
neN5fyEOUZb4u70BudvR2J3ruLMP68rC/ZGtKP1aY3n8wtxSqlNku5vkI6+CE6iewwx4zecLkIz7
1nwgGwg9X2HeZfKB/LN87PK2V8ZQSxj14lsnPxZo6IyWZvWBue/DiVDmyaFDG7NOgMF8XMm/C+7B
/1XIWYkBH6bgmEafmI1S3PrxUHZdiuMnSCt++emmfVcUgDSi5ImthrBPnUuMzqJ+NHSKnnxrNwcQ
/7YLvlH/ar1L+mjHBVEEm5cjK44VdBDnYr1Es+npgX61F///W+pKuOsHS9bm7xCHI5mdX7C6OwYv
uy3RvlxlOTGqjtXKPGhzvlFfTbcbljrIo+byxGyXVz5sotPUIoawNSF1MZ0LOsSJeJIl1RwL5SIX
6UNfQefF0yAHxbaElPUkLMah99VScYfksDfv1TxpTvpENLCKzYTXPMig/iBqHfiYkmKkjxiW3tVu
UJ57bdmPlWf8FZDZQD76lH7PDnI5dQgZx/W7HnQvvxPqi3nyfqYYiQtBjBPAsNG9ITfuXtRMaLet
zzP7UEYgGwzRu2z1javy8MCMncKcGWyCIVubMDlkpa1qPAgyydT6iN1mbSSEADqDGRZ89ef7USmr
a2du7ct+I0kQ4AGce4gWc5g0K/ccY0SLy+Hiet+Pd+h/1WVf+kdgx7MXtTG5u5DLXadYPHLXnxwV
8N1Nb4sKMAa3rf4byR451u9s7kuspPZSpN9NhpLDfvNOLwSunyQaX3xvBBxCdghhjlEvWXum87ih
D8586hVtUwKuIbj9UWOXTWl4vrZb7mlwFiJ3+BSzGyn5kPE6P9VjvvplvZmImBy0Rifisl9iQA/g
jETKmVj/rCcGwAeKeVNXmCkXCP5QaDMQfmwfvqEbVnBWQQ0IFVhQ5wTrmLDHuMrr1Z3hF/8DKcu3
hYzzyTkNnTLEidY5aknh7e71ypZ95TdY3pTj5XeKqmeX39RTG8KxPd8QDVHHNABO9KVR1lUm3Ga6
3c4FqH7O5B+/OeGKONnGqtd94GS0sSS38nXaioxXEjPEA5ti8wJoeGxnWDpA75qNhjCY9zgneWD1
6Vs1KEqFAFbX0KyCMvPZxvZnwYSV78+AusrpxH4l7ruLxZwb5u6peaLb9c3N3a/XsAUH01UZccKP
21rRuTdMksyWCBW1IyGKmiYLS7xEamOIGfE9w22r7X09pEsJWVGIy1ps0Zh9BOqVZnMt41/yfwFm
ssDXgZTHyX/y67xTAeolcyHDawcm0ZCkxsVUhHg1HtYe7Wl9TWxXy0tOMvEkakL0Cs9ceZDJrAQc
PSMcu+Q7ReYC/sH3uNor/CZ0YEDMvDMj8HDuVIbviTbtdy+q3S8qLkKD7XJiupTeyRNJXvlzpBvk
D2YxSFb55mTHzhjczx5nk9LtaDxskpYec1u2qaqyZFayYGc64KhIWMJ9Lz3t3SmuAe3FZyX3nmE2
07VkhSqIpYnAvpxKJgwymdDIrUVt/SdPI2SWrw9TJadj5mq+jVDKaAqlnregIOb/wGIm57CUkwc7
0T0agQzR7KjJ/BVWFaTkDjJ/CP6p5uOY/DeX6NGmExgBru+5kqjK8sFncB3q26zJj1L5xyvnhVTw
7QH+jWEMxjNcTjCVnB/DcgZg5qSjXtiCmR4sypAV2mLKeVUUiMWu1hT5FMslCXvaZk9YJNI6HDeH
xG6IiTo7gHfrZ+w5rJIYc+/Uy47vMCCPd09rPEga7VvqAeYXgJlNRTfdNDvIy7//kRnJKXIHZnqz
Dz0KhCeZ5HdlK5M8VOLcm02iFe3JWlnGvzLQ5BFJBVPDDzbqLqy6Yjm4au+v2KGv2XMjYKGaO8qX
eFFhoQb6j//8/5et862vTOWkgB0YxqfvOALp1Fdbf4eJ0aYfYgGUGXAdRBnwliJNN+5tXmHQUFsX
BO1rwqjU3D/RXDXgn33vMPKfvTsVGuWLPkLZ+31OYqn3egiV2b3pK5ZfT+iadJfi/h6IiWoWYgfI
hoRiPcoq4lajCtlE5I42xFwbpPjHw01e51Q/67Xo0udra18wWZLC7Dv0lA4U+/4mc0vx1h7KdNpH
WKYNnv/XZSCs2wsMfUw3eD/m0KL85Fp+cUCMZz3hC5fxEkk/1vZ4iiIbnZ/aoWq1OY0tbGYVRYaA
y8cw4yXHZrm7VtZCFBQ7nO4ukj24iXm5TInk3xSkN17XCn6SRoJmlFg8Enjww+BXjj80q1ntWyjC
xB5wQwNwT3pLfkx67pNAVy/WNGLkftA7e5Mfn+82LamQ4brq841qNn7PwSUDXe0dYJSNlDC8rzs/
8breSabE0oS9Tk8HAVLp+HiO9Sv5tlc5OpIfcXg38T9egDQFlA0DuOEwV5b9/F2VDymuz/+mQ3AJ
UznLtnBuvprWft3cAdngosuOHbcI+57GdpIutxT3I7SLKf/Vq4lJeSmbYyTPR80pO07u6ebH6s1Q
7z9uJkElYOitOm+IS9iFpxt8bP+5GxVdtjxg8AWsUUq46wrf4OQBV3JWkw/+JLhLRA7NtyFlkQde
LHG2Xto/dB3zZ0oEWSNyXVEUXmqGpkx3wOM4k+aC+kiIKLkhS1JY3n1bdQfXtTdv7MsJeCEUR3f7
VSxA0CuH82LtM3WYOusJVD4yj4LZA14dJ+41tV8dTHJGxJEUQLB/ffs2hEQTYHs/3pMY2Mh8wxS7
AnuwJIJ2IhnrEN7/FV6KJVxTNyqNcoFVcY6vn/psZcRNYNMKrZcIxl+2wSc9sYPmaOszuht0o/Qn
y2V4YHBRxpbJpSN6SuOqecF1ZxushGtwS6fELmB1tidlJ54aE6SEZciL9hQ1BhTHaKpC4JewV84x
Dn+AtFmFrpwhk1VmBGp3b9Bu7d1hRBiyaz8GV3QK4zi2w72N7UbM2TTh4a2LznEh3k94I4BveRVR
hjN9vCrsv9eSZJqgWg75KlCuJkTDcc/PbfnUJn1ulTQRpnFtji+1KZbTUe0+iuMSkSBkPGZ0H3Uk
p9XAIEKpzOZbf5DxQWO6cqNlsvgF0VZXM6hsMGm2Mdnq3byxrEmB2wkE7DPw4d+oCRn27g9NwF3a
D2xur3s9aIduwJp7PNXVs0SEDJRfIEK/VfUW+BiYo7PFrcWjilXPJc7JPO7CmKZhR4tMPDcM8ic9
6hGtVqX0USB47mgJVbIpNUkdV4CjbXDRLCpwSPcpugryAHT7Y5dqe4WGvJyKbYTPOlWNRpz2QGzi
7qhcF8C7Ng50ilN4WR0XADiDPRf4w4AoYYfwNKVTU3TO6ZEzdpSDnFVw3z0kXjlrqpwbrXnRc6Ok
C094gHRsu9QcqrKiJ+Ejdq1Ku7DwrfOH952rhMwd6C6kuygc+dyVO2OWBh4rCpaykCHnRIKCiawx
dWa+GR150dNtu2aHFMIFeNJuecwSoa3dUHUyG8tI/Td8MDPCG6CI1+SWLv73BV0JaykQr54aaQnd
ghPe9TjFPar+z304GFAxaG8xHZzIUuqSyvIhrKIYR5W75q10sdx7LZRX5I0t72a0eTlfYF1tOvB0
aoFuGKIt4rcOAOjj8c26/Zn7rsJBQicUdQru2/Zch1AnXv53WsSS3qQEl9JOU1hzxDa9qerFmu8z
pF7wvaLhrA+K3RIxcL92LI87XepMXgxsbDxjzP2Z8xnOqe+VN1uPsnmsLO8FmjDyAwTGm4fOW8xC
M0KbJqsV4ZP88ZiqtK5YFpL/E6dlo9tO++RQ/KfV/OdwjSua1yh43X9npYz5+1ndispIRdbltdoB
E6Pfg6fxnRBTa9Iz4VRJb7ghgmzNgTKp3Tuar2ToFX+lKuS2G37NJlzafHts/i5BWoVwg2ZMu5Lm
AoGh0689Lf9RRflrsDOz9/4Uinrt5S3uhw3dq7Ec9BFOCee5OsKfTAaz6EtddVTBPCvvyAHW2YkA
ilJ1O7FA6qviWI6S3pR4UbaBNLUuoi0/c/4xWlOBOwkPvkiBj+x8h2nosMc8ITqrrqBE0EVe2AQ1
L5W1kANHSeI4TCueI1jqa4UwIUZO68Dwk+VH7bHn0OOtq8CW0AXEEk3m5ZGjnoNi/1MeSQrsKVRC
zPFtkzlpVMRVK8i5jUESWxk55vOzZOUf3jZxAyMQW1pLpIJ4Sw2CEBuSXm6TUfQbOADg2BDANjyZ
lNCjb1nJCkpKWs7IVh1/wNV7ZuKfSXC1S9c2sW0wMDdtVulYXmkRfynZjP2gzb8OXFNv5ZgjP7a4
6kp+3NqorAt7ApslXDTJ9fyTps7O53DD8g6wTHBhGlUgjuHJCNITaipGXdh1Tjw/2QusNUk3CdSt
XjbVn+0+ang57C+pLLS0DSWSATd1G/70q1p3UxF9OTvc0aQwprj9pszWnIYPeAR0Ei0YIY+dLxlj
MVjUx3O3FOQvA2gYhKNHOw/Xl8SXA2prwR1TM8Rsv3o1BTSZlr7XUJrBHwBA6BaQCuqZhttHxFtz
CkDy2YOfM+OAlbngW8kpaynKs6CgFK9+abFftqYlRDb7H56TC28RbTApAgqFvkgq2T1+6cjrikLP
Ef+rCcv6mHJJ7zRAlqbkl0hKLw5KFRkSGQe/6OoB31yoMhRqobwa+M917jBjcCw5JXHwbMsUBFuE
8E9aCLsd2+kYwZNsOCDx/CjnJqtoZVRSaLjB7/P0XI3jAEHY4koMoD70dkjB2zDo/4TliB9wAwGn
DyhZXwCOxSJy4dfvgMgY67Vg9MWmnZG750P+g0IJCxzLWQyzsOMfLSR5b2sJLD0a5Q//Y3ZlkPW2
FxYn3BT/lGHJEaVBXnDjWPPdWH7jO3ccGfq7ni+8D3qryPXAGJ7H+JqnhEfZVJmKr7+JafA94VTV
BKdHg++c5Uulh5zlGFDqeMptTTfkrIHGuf4oUfLWPS83rN+cH+Gyw0jN7OAWj1YWLpNDYhBlJzrq
KKKioJbQxXEQHANh2hjj7/VPNdEsiWy0kD/40Yt7nOKuio7Dk3hfGBmWp9tHi0X8+3xpJ3fTdGzL
FnPIH/11BsrO7Xv55GzU+D3DY/4Zj967qS5gIPaloKxYaBaJWx7PldoTfNbYcG1gu0kEH+n1cr7c
+Ymne/T4uTuvY07/IZ3AoV4rQWoptatvQRAXJCTjFVgh+AeSQ7tqflFQGNF1hK9fZCq3o/0kdLty
aJlATILj0EWJ4pQ7GEj8OfX3+mJzlDWeTUQmbNxvm+Oozu5b2eScE7GTqvnCaqv44DP6+31d0NCv
iUgCCVaoGmPf0JuML8PyZfFxmsNWFHgFNyOIzB2ZHsduWJKftI9IciDmZfiD7ZPwuPhgXMFqgeXm
2wA0/+EYoN0hdthpdEziZGaVtbTGpW9q+G0vy4CnOqGCoieA9TcyrZ+l94NcItXRNklM/fXyOdxP
wUjzRd2/VyRgFFJ9c54Kd8GBm38H1aNaxKaZTKS3ya6vZD3K77BL0vO6N8XQULWQAeO+tfV6snra
hE8RQ6qgM765FasPhpu608yiMDs0sc9PVFjP1HEvmr5DyN1TivG/Vw6BLQ8y6ExirvPSqdMSpTXx
w642IcCtzyP3Sa/aBF0fHt8WzG99rcTrC54ESozUdlCG994XikX7/0gMC3BP3I8DlFOcJCHCmMh+
RNIwSRYk+uod887NitghUCUWPMR0/uVaSzUBNVPWteR7cSF9HS0U67mGVj1Ua1Hgpxa0PytsKMdP
j23eHePr5QbLaLXJh+9vd6pzLEb5y7EnKGp/Pj3cyZLX7w7bE+j230Kd4pBXYfxEkR71Thf5P4uA
0GMmzLAC19EUT0JsVgFEd673g/RTs1wp1xboyveAw4DJCeKEIUcrJDSHnWy4n8Weuv4Gu9fz5Mo4
s/5W6/sFq1VlKhfXDPUStKjCdJKpjUnmaGi6AsbM+1mGBNB0l3MWIZ0esDDLjTniqcMLrQMeJ00U
XK0KVmyDYhwlWcB1IYZ2LP5wt1I1leD5Hi8av5zswvIdFG0Pi9qJT1x3nmO9FsHqdyke7OBn7qiY
JZNl9cGoXP5R9rKCo008iBLlpNadaml1bR5Nf1WA8Nu94pFO/LHmhjxIFevqwKasSNF1VSxjsLmg
qGRFHe6AK+HCw/aCzqRR8lg8ko/+Lb7RQqZ7YKYQmtWg7JB7eI7X2zqnzMJoQ63US3V9ya7PnycY
ENW9xRWrufxy4K+4t/8keCoRwaUVpg94eFUMaphhkhUX0A8UrSZqZ/5Dw2lPY+YDKzdt4hO0OYLu
SW6dKlj9Q14udBqNqbKCR4afqwhc12xEzTDxdjXkqAGgzHKblhiaZ58JDqkRxnqrInJb0pNUFbJn
03iQq3gQOx091vndOB2pypDIWeAqQcZA6xAvNzV1ClMHtJQnhDkkbPlxktXbEkpgEopElID9Zfkn
MWF0sE6q8tPXv35ji97I1egQ6FY/zKIPn9LD6CaJEL0P/Aqdf83Am+U7BHN+GWNM8jKgqcOxg86B
zRfBeOk7S8t8mwSBCMuM77h6yeNn3cwjVjnu8aXAjP6/By0Zx0RwCr9r+jKyTaFa4zYlwnNAXd06
z5AUFGtncsbour3u05ajKRqRIKJNc86N7o4XBSewmw/zyHGXWKse4tvC+ur9Lx4/CDD204JmzqCq
CM1JXKLPxWqdfm2z2qEGT3LMl/tL8r+vUn74+FevRObik4y7e7wKsX8xoF3ePPveTQEbEkRiI1AP
acpIbGYRCyhnQUxeWcuzVMhDUg3OpS4ukWsC4KWQxXce0cFBeIukTfat1oLAXKQJmuzpWL+u1T/v
e4sPGKlR/NCC0REORDVRIqq9Afl98IGSDglhw+9edogTXCL6bee3mgumzkiS1xyQEyTBgJfejtmr
7VYxzwHyZ5fPP+nl5AH6NhskEoWjP6wnXhDZDf3NjwxME8w5o6O7kM0cqREIcPE54hUOtM+wd7ZS
8X0d4R3snQGRODGK5+zDIxcyoDXTSlOpeAfQAxunlX/bLlWY9AReClMCODaqC4BsW3Ef2pnKBD+O
83EbKEkkaQaP6B3ZfAsZK7/nyH0RZpBZzaiA11SGSnEv3TJRn2q1BNhZFhDGEnd3lB9REqXjpOU4
TnWg8kgley1ATmQcREloSjeNuXio55Bn11ol1xbZ0ccdZVZZxSbt4gHMhBsxwpmPSWXHPayf+Q03
rAgWXJ+X+iY0KwK+wfdPub0e0chZBaufpJpkSmotIDJX/c5Y9cFhG2Mj5Sa+KaFuo2mKsvgsr3xb
MN51Gh74sJK1JA4GWYWpHbhWQhrEbkpQSR5WUvcmHDOPoPYaC1yvB+VECx8hmFsW/Gz3PHoArNc6
K3ZlY3aEBSG1kkVCwVvY1KGAdnuMPj2eLTnBkKRqBZA8Q55jVaiDgXEo3cZf9MzP17GcKhaJdLaD
xRASNnggIuX2XgGZ5z0J3f0BSY+NusBgVC7fcJIYdrFuyhL/1GpcE98tVcZOEk9v3/PdwcU0J/ws
0VqZRpC6HC9v8U215TFUwiHE83mBCE/VieWAGDwAg+B/pm6VijF0HwJl0B1LnnD5na9QnLpTbs2K
/xRpL1a8QyDtAeoZ1DlmeSUeaSzZdtOoFmkUbaIXqwuZLUdGMeY6Y5uJ46eaZhijHFJhm29ldBGy
9BCAsHCUQjstwe7sZUXBbmOamSaB6Z/Nz8mTUDShvMEed9mx0jdN5ONrOo4oX2L14U7dENt+lbcg
2j+t0GC3PWeyOwOM38y29YttuHAN9lOlgeWW5t4FSV1v97Vv8D7uMtoLnm9/ua1m0y4Znq4ZjUa4
rR5/lu+ThtAixSBKJ2T3ile91JBNR6IzXjA3HE09OZh9MvuIGfAJEKrwqM2MW1t5tWENRdhQA0j2
IusfYZrqs4TbHsHix6uYagHA32jJV1nqMFyhkhExNPfNQFBNEoxx556BTMe4iiz9X0LxR1/1ahv5
TMUBETPlSRvTeemKMrpv/AAdKSXRfZmgnsK5OROSdpyO5l1/9uyhrfJGeVMcV4P05UVS0M7jwrPl
DFqQWsDjzgMjrxiPzWt7q61Mp0iBC34Qu32aNFDXLsbFFqYQBpMUisUE/QB7Eu3f4mt1osbCwj63
IEhhgRtdBfa4yskm9fjslu1Ow85WSTXfv8REZ9TpEiU0evCPzWgKpIaaJUxOAALGlRJbW17c6TpN
6c3dx8FoCgU00wHWq44yXCVZzdC6IQ+5Fjv9MhOGcW38fiRFZ9BF8cjCIxpZm4sg3ce1lituwAJ5
pStcxceCYRpH+D2xl0pljMRdwlUxExXY5eZNdlsPQob/VedgEKOmYjGnJld53qkX/ZhEMcJGwyc6
hnYxlVLoou53xVhxDbzkWYjRK9cIs7oCDWmAZUdleixsHYokvRE6I9Y0HhUZqACcQ3BfBw7oeyj2
DxLKUpGHZBD6PbdxJdQsSW9ILect02W06YaaBdg29Kmr8jjx+3B5MYCJ++Baxsbrs4gznBfuA3Nq
a+Dzn+j8OaFf9VnYfVApZG/1bNKse+NybsuNwvN9h3UVHfpXWWIK1i2Ruyj1As3BAKgboHTlY/8S
jq2wMDDdXQi6jcdIyEltXl/3Jqek+Dj+9ypO/Ne410VVZIHViC+enzUl4+KnD8Mtuhcvuc6b+1/+
QGRSk5HrfGhtHYfWaXxfAW7JSgEVZdeCuRZh81o3P/Ho8OtzYWNzmy7C3IGdPVIaBe69VOkhqXEO
GRi6LuLs8MTIXI5ZtC2WsZwnSjXn5OjJ/2OSz/T8crXYqdavFyYm0F8VC8ceYysdZY1TfxGVW6EU
sROdn2G7/ZnE7wtisJgA6+2/lUJIMuAw2QAXMGnBlMIfNGF8ENjIl6X5+/NilgnYyKIUOsoud0Lc
KPQxQn4z2bL8N65ZlfJDukrP5O3R6GHHS6FC7nLXQJuMAszMOYLas+LzO/yHsZkxcqLqWmpPUEFZ
BKq4wtzC8zwqP5+wMlHKNAkA4zszWvgLXjjj5QsTSahhsp0aK0YrBZWLn1kmj8MyImEHYyGbAa6l
LXxdeSyeb9JIGtrG3rc7HaWC5JDy3XY1UdaG/+k7X49OtFjIvQGK8k8Nx0gA/s5+XKmPCCQRfZhJ
M1CtN/Shy74pHq4P7sr4emdVxUS1CmfGdn/ktuJrA3KelqgNv6kk41fbGioEOBsO8SfgwCfRYnTv
IBYR4PUcyjLwMlX5Sf+v5McTC8d49MU1GjCAJVXO98Vsc93943TudKWE3CJdmMSiKBHi5TT0MbQ0
E+HstmvBiy8CAKFxz/JIErDAQZNgxadbKjleC46T85BqhA7GIYti11q2lGA7GTR/WqsAo4NHCZme
M8BNuw9Lapkxf55hVE5ZztuA4L5232Wm9+9s5NhNgXcEc/IKK1ZpkxXKVobXVf63fvfy7jFHWax+
3H6xYu4oKMUlxahQvhO5rLKsOeKRf3DEcMg/xngm6RIga6AzrvbLoezp9k69xSdRXrPcGahKArOI
IddfdB6vbO+rnCtWrrRxVVViW0s6pGsDDjNIz2JfswfzG85ezsyuvQCrfpUy4Nt0kuk5y0zyQbit
bMOqM9EQ2Y2nuSuMSO0NoUqYybsY/qAOASWQE2TDorLtrj5fQORgd6yZi2GsX+uVTN7n68qO/K3t
VxJ6ooSVixPiTY3XFnZOhwVcd6dY5hLeRPuiZ00nKXORcGp8xnUUv4bGziRrdfPX0KGFK9t/qz5P
KWvxaVex7JKOjl8snB+Wdhl7kXV1kVlN9Tb8yeSSaJpcUwjXFK8E3x2WN9czG2vEjUpalttBkaVr
+xPepJFGi318g2C3ZU1OlntIwMXN4krxD7fLaTmk/qq19JyEzPW0ipXbABg8jELKZWu2KrIkr9n5
fghW955DS37tCPFM6QyVHF1OeF5cL7kwwIRHgeGVaRiAHuoWYKaimTLCmSXZO/FTwfB7UMurpJaD
7q8bGG8r21LbtP+FAcuDBUKACds52gAegUdVWF/Bo9NHN24zNsknQU6x73gcfG3IsY7VrKG6EByb
BeZSc1SDCvlRzuBHmF5zAHV2btpzSCvOyM4QImx9zjf3LGxGEea9zYuMvjfs05AfqRnhdtqm3aXQ
4o9IzikDyGAEA4cSnonGoy07IPk6UX+5BQ2pFINIgmpDXsfxvwi5psUjKLDP5F1Waf7Om8/V1CSG
/CDUzrm7918tiFqgreZZoMDGAYGLYVK9UJP3n7vVyyHw9k/2TlcRTBjvmWauU6ttu5VLIDxARiDR
Z9RV2YNuEFzUkAvLvvsJv/sTsvF/Q8jDBtzLRT0X9wriI94PTc5vkpDX2rwo1XJnX4DX3SwMDfHW
ZVdYOFJiUJMGTjDtd0yP14cdLSPcn9TbOTzYM7eT5Q06hijojAqWNU00lrl17TSuK3ukV2LeX3HQ
5WpeGZUV1NNY673CJb6ONOWckuApeQBe9fb5QhROA9A8IhwVyI9TLSYaekU8LfN7nXrmHH6rDZKw
9+T8sUN40k9jTo26BRpt692N00M3bkXDzZQzj/EpKZ3aNsw65MUP1hLUPn4QwL9EdRq6xZta2weF
Sm3Efkl0ojujnz8SOYYYf3tlB0l5xw9feiyWAlG7f8tfkGuauCRipp7SO3qw5wDTsfSzWYvXM172
CgIypFGCdVsft+Vd/NMR9434uWeWkdd5NXG4vq3cVSxpquHb7r9kcwnr6S3Gykqur7LQQXVPqrkt
SFsvX89SOoIMbDNqtlZcawxR7eB1wHS/k14xOZim7dlTsQGIqXuuyBaw2CUnBy2OV0bAbHpG8BZM
Ui6loFqA810Xz93MEiAPKi4YmpQMNiTywieuQDqS5cp9Zr8ZUSu0v7dV7NHTan/cOL9/BwhsNaGU
0Bj7dK36kkc176wneXw+o8qQOfSonutQZU9AEf1pOZOvWljKAJfy+g1QsPY5+j90wQbIr8bv8UpT
d919pU4cuqheagb2UKz7AMqmK6ACfp/4P1uSiq+hn73re0uOQMdQt389TCRRxjOPU0tFd1/NJ2Cl
eVopFYu/O1IgzfNY0Kl5LrZRCH9MKt6esafh6Qxxtp+wHVBZA56Ctplt9JFm/Ewip/bol6n0ps8y
ijL6hyVpPBWDsHiFK3mdWzujgnRTytHl8CUdkaGIl8R/D5FVPIlRiY2fJehCR0F584ZEiC6zaU/+
bFzhGRWxvuuNjeRESolgEG2RrnLBA022fw56PqdDUTOVO6Rl73wteME7La1GbSlcrGDVHdS6y2xT
7TzAzPnGvDU8cwOJ6y9m4CF35GpBh8an1Q1vHH8x53R/PPlFGsAPI7w29MIhbIVVQw00yeOAybe/
TJFgCR1qUlygRwNhQspB4FmQCag+PmTn4O4PY0tdZOe0bKzAUlLqJtyoZiQKewVSzjskCWKLnBT8
nJkCpgU02f8TOFC3v9wgJzdAhXUlRtWTnwttrJATmyOG0O67mynfZOwtwYb8QJu7IPMdIGY3TY93
hMxmikc0knaCywgEVgz8VOxHE6JZHcrzV/u6Bv+d2wHZIa/0MF89tjixXGXDKgoAk6dk0W6ejnlo
IrkzCMzGYVWEcVrsxwQ9j7AiQlU60ee62uFbYgmlzKIQ0S3AybytjLATgD4OXCFwz6JIVyJhAesh
wlgZ6FaIE2pJCgvN7yjUPTcHBBuAlrncjVPN8mv5GHqhyn6RgK/MMkEP3yYBYnPY6CAIS40RmDEX
EjZA+lfkY4cPJPgjAloPGBJWf4L+4ZxYg4HPiSYjnxFw59I1MAReaCgz43C24s61d72kbhyFCjHt
qEzJigupBJIOW91VymmLgHEVwM8NuktQP92oZkudgzWD9iLN8H8UDRPWv2IIFnnxfET6hpfCOI+w
NDXc6iJe+Frh9lui82Ed7SFat7sBZrF6yRtfAl2Lxm7G0dZngX2jTYljIgtu5VQpXBNp9lbLNuwK
j9K08JFa7si6nozuwVrG0g1hrAXHGOL795VUoNSHx+985aMCcI/OH4mCWhdISfYqdGAzpD9pxPs3
kDXbjt+gzNb67HG+7vl9YjavJwjCZ6qS/rrUUfi06gqzwSWLn4IwzNJI1p4iV1tXkDcVLdnvuULF
z6N+rUhd4qUuFeV1YtzddflQLA8W8QFXd8EgVbg7moCwiWjyQle6brUH6277fEIB5SuD8YFQRqBi
MNObAwylHC52TpWS1r6h9/U+CNaz6MIjq29ma4CKODNYyPajnoL1sNvoMuf16LQugC95I30Kfknp
/bgRwvtQmb/X5UvaJOnV5VjnmWG3MTFzZ4pZmxT/Y1TynQIJyixR05EAxRKU2NO8CmSuXEqkMwoF
yPoZrozCg+iA8j/Yltf+I2n5bjIFscCSCJre0rANuo4wAaVNeLxfZ7zVbQQsqn3sfX7bSNameNly
Yu+hC53Ljt2m7yz6qxc4G1jW1J8aVC7VYWlqYLnq1XPXvItv77iaX071XC9wPWAH7mkQNN+g0CqU
MgI8OPX1RVwDPEnZpWfW5Vun33zd8uH8xl3RwbrCaVein/0+gdicDSwhr+K8yndx0UQcg0K1wEXE
VVCzaOtU9spmSkfTYd/kNu0XczMYAu6B5lHJRk0cvsRgDs9Lf318Hb//t9LWcvkrFFqEhVCqfdbU
XRsdJlHlBLvRC5N6WniCt05TP6IlYU2vzEmEToM0i+vVgS4elIPbfkZj1+gmqMyyUh4cjGT9HpWb
nufA/nazlnmGHiOVwIYw1YMYFB5LhBs93N4C5NhVpaYJPXD4XlS1salEPPZi5CBcK6IfNeQL4Hm5
o+MAS1G3O8RWLj63OoP/iRkZEj4Iqrhr39ySxWymwRx1UCub2eyVvNZWqXeiEO071cWp5eWQcP8F
CaVZhWJn8KcRp61PDJew7ngiVf4OhFzh63Ewq52KG8s2ApJG8bE6qABMAwffSNXWmsqga83zf4pE
rsP1xGdZ/VfDhJeRWPJ4WeeLiL5xr32iwlJvKKp8svhsi121tvFz/liV+u4+0mDiyceOY1cCwNH5
I+if6ytSEzzUoHmJEE7RduAKZR6sb5p6HCGMDNaNzj3FqFA2z5WcefGvqcCTNfZnKGglZI8BZ6tf
5FNkmtwGkm2F95gBTz8OU2uGMb6wKgP/VgNkM26ES9n7HwtiUF1MecmnZ/aonpv8Qv58vTnew/NU
CeeoTtfBl1agOOSiMlI29LOpt19AZ0xEwk0XeOd7sQlIdhuaS9RRws6jm9vjA4iiu4oP81eICsyT
0KxxbSaNIyS7tXXsEkBSva6VjvoA6iQpQmlDDb1yRfGvtcD/Ktw/SyGZO7tdlT7U4lLls7rkR9CR
mu4LKDLOKYLM5RpxRQETWbC4260birVxeXw/wEMSzLw/yk9x+uR9/6MfgpDs2p86rlAjNA9QnYPM
H1bBKIudCOQIEqtlj8d+SI2SRHA/1n3ILxj4A4KH5RuKiB1IIh0RTfKDqqf/jllMC7zc0Cu+EhCx
gev4ldnACviHIFPMVBcxs9Z3ZW0AtX0MCafjrYVuN0KpsJCA3aZUtMMobnwWDIpNZWk21UKT8Esk
tS+ckPoFcaJ8KTAC6UtVuBr5dAUwE26vzL1UU/CafDq0kK9Aheh3nBYDWjP5ECZ6RiAmC1yR7aIf
xzI5hBbBcq3+IfjnAez88dqhgSkBQIk5q/pgiYHkYxiJiYiAs06fogNAOfRpH3KuI8d+93Cn9ajQ
SkD9t9yidr9rB0QrbVYJpnCBqh6IMcM7I6JVbCFBFLInwalPaxbbohacuKYKwR64BKm/aetD/TWY
TdYHenYmthZHO21Koucbqw2PXeXVrAkMBLqoxEz200ClzdBiVa5EbR7mqiYrhyAHNHsdYpVuNiHc
y8HQgjgdX/zfe8SDWCTsszSGQ0ARursQS1J5Z2NR0WUtaGZvEzRhjDtN+tbtZ3bfko9psrl7LGd7
vYlq1LORF+bDJkrz+15ZcnQ1zptg5oYokuvuw9TYRWZABAGQ8ICVYJMuhXiii5JBnpdOhPGD5Kyc
m9o+0bNCbJVis1HPJxe25ZvWmezgK4oxVeM0whebLYKWMz2sToUcIOYwwOxoAoIxC+Hh7nyDqAy8
HC5psjhkE5haOX0yZfsYpHlzP0HDOYeSDsFNUwNWtA4JAf3CClc5ao/aFKugcF+4WYTBT1H8QDR2
Vrzp6iE4CXTeIcT/FsEqjOuQYdDXOIv82g7cXV+mIJvS3fzWoExY2CZdTn1iWJdCX5gmolK4IxzI
zlZJFTOG64WZFIsasVZxDznsNo6IzH2z1vFzJtCW3rU6aIRW4al23IX2AgStz+iXyi8ojejzX5+E
sGJHZVlGzymvu0DQ71Zu7mazxOJxFRkchOaP27XQWmo9zbjnXIKKpxgGYar/nRkMiqzidlrPXJep
alxQsSFnAlcxZeE5VvPZ2AzlrxhXVy0UyX06xr7JZYYt/yt8W+zcWCzMn/soMKu3RkcrdXErxym6
DJL8iKTpI7L1RqALvVLtanR047nuZ6tlKP4Z1ZnciucoKhnnJ3BjDLCOWG0OXBMPMvcpug9cEoUN
1d2Z0wpLjKENPyk5CcjVfIxpWTT64JkufnATPaHZLBrL2NVlHssupas2G0dsT12t/Mn0KIAh1PyO
ZBXFMIMqLqkzzHyK/ll0lH0mGIDx3Le3K4RK3hZbIMJbK9W8K9/00hdXjn0r4WbpG9CzTz+DYp7J
Y7iJal3PtAkllZvxBZJVv4xjS6v4gM60MqXKGYyWP3w6j650M83x9G/0BnIWlH4XfLByWxo4hlp9
VwGnINPBEFaI86jOZtbmBtSnvrpfWvviBdcUIOLGSZb5YnwE8s8u1GPyEidWXiOifRhL7nXjYFJr
S3pzuNHKmnwiOAY6IpYStM4MoLuUF5UkKedj+IbbByApiip81ouULa9+3on5QaZ5fVcVEoZpK6gP
e3XNrDrS7k9wYTXGANilvfa7FmnrkHXI+YkavL9Eb8224Ja+syp6CizmvqpQDL3cWubhjk5+zWyl
9uOHbLXxvNltIuEri/tiRzseTOr2QVUbbuwtSQMgeBfqrbuOR0adKePsEYV226E3/w80QRP2NO/8
DdrrLn1rF1Uek3CtL406hYuSziHlmSs+asn34chSdfES6a2A3k36IPh5bTs6JLm2piTuqD54zMgo
V0LX02Om7cRVvKVYU7wG8Qjc6b9WbKBPuw6OFbNkBxC4m6HZUG7Gagd5PJCHItyZTdG5SNvkc3eA
2zwdtahFQWnm0OK8kim1xrb7bEqfg3lwhgmCGeAsQ+Lr97TnOG3Eixia1iB/xkiH5161rCFYUHZC
9AjhF2sFf7jsyHBK7cBkVhfE5eEhz6XoMOZe6wxaQW21om/7fq97Tuw90995ozA35fTOsaH3DE88
n/pJnURjnnMf3IaQxUjHexRVLEAEABUlRG7Y8Y77865HuLiHffgLxTKPtaVCxNdUsWjaEEmtgsAv
gavSuj2rSrKUZANMYNOXItPVUYcHhIh/YKUhXnndFDtyk9i8IaOGFHizlAqpumOcUW/z9wPb4ZOR
VatY5uHvxuHIlLMOSChBFlvYvoyJPBBNNyZunpceCUFVpDSD3cMIOCsZth1MXunKnkZMTO8A5FjY
vGlnbxUrNIUDCucI15azORYMtGVwBeHRCitvJZBO6gwxrxkVS7Uno/fGg9nDAYH5l3/4Q2ZCAKNe
Hwxb78gJ0op1ETkHu2r3y3oPMOtoFl8cceRAP7C87QOZg1NlYlFdhuslcBl/Vbt//5R8lisSZxmh
8iPxwLE0WGsUjo8+jg/NKRKzZ0uWg5jcOXoJ3QAOGhr5eAe+o2Jfbim93dh9V0umhxPPnwJGWM7O
BPG6gTwpg8ikHV9xjRsEcRiJfY2Yesl/SbHljXx/tOM1rI+Gwurieu5vY1Ejht0E9c+lDRks2/nD
Oen/fF1lGpjthAl7a8cs05aL5n8iTwDuhdlmf7/tFLf0QbXKuCmeyDBO9JqaxH/5GRSuPDdBYzU4
sww7AWShOczIhzjKz6M3owT3nZdll+WlqxjWSAoqJAeUtqktoPzB0StQPNEW9gnBN3fD3wAvMMPE
W71NI7IFszyskWtskWrw399AH0cKl1qdQas27vtilb7W37YJLaVdkWcLWaUs6O6W/yNwD2xMo4xy
jcHS1pDfwT1ntsL0grrIxUiAAtkmurnUu7VkeNsW5L8FLDAycEa/jjMYevmOyYB2bYae2xyV1BdG
DME7bPEvjdzkluhpwexdErMUDQ95/ilRxS3t6Q0HcUxf6+XRqrYU5ocUSfB64PzcNiiwqDa544Tc
Aao2ygd5B9EgqSTF/DEpHqsVkkTw199tVyZpkrOMjuxksaEcs+pRi6UndA6xBUOLXodawnUXuaWk
mxoJd89/0pyg/vwe3HdS4Cf3ygMQX2lMMqcnTHIBULOmM7usH3H3Rdx7kT1BJoOp6yCGmuuzVeoO
UbmybTEKaSCnELPYuhngclcePTpKZfV5QqHf9s82CY2+xvtNSjht8o1QnPCEZZAQvkzgUkbc9UHn
7bdZWvl1IrhJTqwl59AIZVwVqFmQEUII2i8FIyDoNqxU2dzplq5QnpwfNP1HW3D43Yu7Eg8iGzhX
zpcTNkpVoAba0jTXFxasQj9SISfPteIbLuRIh0deu2pVJUZx1OvB7YxZp8XesMVp51W86Smua1Bt
OJMqZmidai1Yjd3AS9KpoId7xMn/fdKNtJDd/xgnftKVR4R0fA2GYooK4kS+ZPL40VcF6PaQi8m4
GrGUvce6Hnbx28ujugIy7u5/3YY6o6UvsiH3O1r95zuOq/k3MVC097scO5XV39v6NTyc8J87DWRD
/EMg39GyGQmiXvPrOgiPqED3pILAyLN97POy2oAPLnUm7AbsBJNmJxSLmmt9j/+FNPJcL2Zsb2si
WtRpe/+GYUmTfia6v084IaZJxyZ7KKCFiKwGqXNPO/9DuomLFMuY80KxChSZ79mZFCfsZOHPmxxv
yE0MG4m0CIsw3DgaPjr/TnXeEcvrU9GWehrIdiLh24O23K7P69w+2FBshAZuvDjc/H1VdtHOC49d
QALmr9q8cASiI0X2Ql+N0/oYEGJJwNd24XNVSLGu55b9TVpigmGY97TMpJdZgXBdOC8ZczH3v4wA
ciY1u5Ib1HP0fO4R8OPtuHsH9PVMjRNAtEfNMpL1iLKvXpH95XzzUVeC839305FE1xK7uda6QNEI
5zzyKUERZp0T3BsidoXcpjH1rcctZb+w2VCy/ExhUPaeYA7a2f+txbe092y736mU6PdnciwRiori
WMxX5NuoxkzhAE5Zgp8K08JyjN/2ULE3j/CcyZ3DDduFygZ6pVtaTcmjgdLAg8SJciwz2NiV2B3v
IaejkjLW8KHxy8KMud2vsvgM7o3CRc4jjotHrIBN6i+z0PW/+SH8FYm1yE6p/ABQ+Hc5exmuyGc+
pAgenJuhs+5gVABFu3LntpFKhjwz+fz10Sxf4MCstX9VTuMxibD0oXm5HCpH214DyIFngzuxEiS7
UQHfMsQCc7LSKAFAlY2FKodxlorresngZs7oz0jsObD9yK7IK0f7npe4Tir5l/485e8KhvLQgeVD
svRIssmHtR1snRKWrO0dzjveSBDMWwqnCYKNmcGRN9DOG8v2TXEIkLQeqCc3hBD/k/EMCgHOIZNw
dICkQweb3+BR46OrVd5rVbFMK8OM7LpkWAoNZvA9ef35+BayGAq3pfNcp51/gCtjVJAuN+5orVyg
ZOosfoUlwmtVJezRw55bksWjX7+Rw6vcqVWNKIxp63A/4JyRevdrFIrLo1j+d2+bY48OWOy5y+XK
+b5CeuH+gJo2rG1FT6LuQGhCC5JFJIWD4UNtMF5TuBV4unxxYKURJwEuWhJqWcjrcN/aZexepVwe
na2ZsBZb8789Gs1kodB7mLJePjDFPHR9AHT8C8jnainrb0H0MPwISMx4SPL+WkKpZZufc6vjw5zr
kRl2EdMiBELrTBYCfLuAn9A3eMAGec2wA0QiObFvE4+FLfOy4/Az6bL/v01AF2gbqmh8apWY103l
wa+P8bgws6NwYcoIArFU7T0n6vwvKcBean35ANKLdO3z+Xa8PVUdNKJjG6MdnP2DqO75Oja/jArW
Pa8UCoEgd7SZI0vfHu9Lde/EuM4gYs7sWJWqxKWRYzKgwyo3Q7s+hHpDznUIMiUbbQjoSZhfXtFk
a0enMiTyIDGoGpuncmwb869VSkbRsPlclOA9wGnObpBnW8B5Rw0Z8JmYec702Mj+/DSKNfDBAGMY
iQoF5HiXcCau65qAVwhCpcb0U68/lWzAFKq2XFDluAVexnPmIjz1QthS734OyYJICbQCHOYei41e
IP5Y7fF5FNfbKCKf7qPnXKiEGakLj2q/YT8gmAxZf2AH3N+YGVTTCR+tzBSwCJeBORZ4fGoQNkRM
CLx6RLSE+ve3BpsgePzr3D/uAXtdgSm7gGSCXeGbmf2ybmQ/cgqVUB3Ipsq3U3AcYJ9tBHj26SqK
yp5/4qbKlik4zAN9XOE9UJJ4ZYo/lSNq32Cmpv8Eu+zL0NPWnCxiOQ2RTGEEqKbLpOZzCWfaPOlV
c1YZ3TATbkcFGckzwqD4z53h8OSRgjzqaQZzYYb+8RgWStPGM8Cq7uItSZ1YG0XJdHD94jpDl+A7
JwjJEKkkM/btLG/Pn2x0tLtvhzQi2s7IHx5Qe8GXOvMA/3giWMUTr4DZxm1yRTd44aEIjGk0Wil6
m/ntHo+tmlr4jbYDlS1Fe1hDnKRPgMfAQAMRtOU6LJrDpZnhJ4DO8GgjTuY3ripWIZsKPDIeVMs5
SG9Slb8FJT/fZULaYTiOqAZIek9EJK6ROZj8U9yvzwBNFMqlTHweD876I07FRbjMWlzms5op7ZIt
0ZI72xom1iqoKIJ8JItl+Qxui2mF1zrL9riCIpQZx4qV9dmupuBzGZtDE4jAuoz04BVzKGPagRB3
Gfnuy9tfnwVUl1FjoFtk3++4J34EYboEbtN9BJagVxj9hwawN3MLRk4Ayz/4TCpttUG16kCVBNfE
EmuAq6eT5jCJ1Mp0SWtpQOlMsrdcFUYUkrlI+OqkdimEXWiveJNWzVXyofI0ZXk7y5D0BDjlm58R
zfqx3gYVV0LY46amJgK/cyq4Q9I717q7lmFS1xI4Wv9fsx+aqpR93tHZ6kX57kVUEA+yUCCIVFu/
TfzIyZunUysKdmBMRIHv9nQd92B74fm2vV1OB/hilt+XwpMKEPZtsQNzUmppquaT8Xmz+glpjxzI
bWPyVIGfYHNkFSQ4B3vu9yWMbMjceRRtAfyiamyKrNssdoap+F3sYHeIa0KTMezlxT7vfUMkW09y
ajFyyik43XwFF+9q2oo+vXqMJat0CFztqb2Yzw5NWXSXshq7b20OWLrBk0vWmdMOGEO3CiHRnf0F
dZky36TE+RpPL5COaJ0Wbbuy6iwy5XOPagdmN4nkMNQSyk+asW2nyObLADqDOBuSGWCl/Lp9+ipZ
dNEy21pdWjD7Ne6E0OdYjM+aAtWfC+nrn2Ib14BQ9PteVt5QJg4eNMFPFZZbT04yBeo0iwViqc9q
yVK5xYhsrsLkNfU5IgnxN9r/zpHGQiA/kC/JmY37RhRRjl//zJpRAg5iDReiX5lDiemIRiKQ9SWB
OYvPvaEJF47v8JZSWONJpeWK+D5CPl2OXLbA9x1EL649sKJhyKqjTtd93VwKDmW1iyJ4xxJniZBS
ZVisy/haEiwbLkxSnt0r/cqDYxiYifa/+OHW6+0kh/1A6O+8de/29nCcz3xPKWlIDAVay50uDRD7
AsVSEmTxj9gLk6lAGl2pTKeCc6KG4nP3N+v053KhMToa6ha5C65lwVfBBatPovHQdESP9AbamBom
/Zzk6U4WEha+Lh39lODLQxTf/8QUdD7JitML4GUcvMbtYQES/dK6VpK40rAEgrxT2rnkqTUHartU
r+cyNhvYiPGZaNhDG7eB8udWBApc2nMZgveOclF4Hit/SGmh3ZaMaYY7p/DNBDHkVNUX5wl67Jxn
vacAOeKaZKqhYR48UrZlOQFLK2icjMvLqJlcxKlGuwlEvtW7bB5HJdbEnNa2JoE5qfNrGaW94Axw
+DLHepNc5A2rTaXyHQC4wMpeWuP1Dnuq1U43Djs3BuchQd+vrlboPfyFAsxxVo7Bk80xcmwfkjAC
AIn7tzhodcUGuXIGOCUNsvy3LH6xgVAnAsgVJYzW2h8LKCLezLFFUk2fwIGFVAq/BbtTr8jEs6+R
5UyF1DvMOt0i0/mTRuOpoNY0U05EUZxJ267OpDHm6rcSfSOg2Q9JenD2JV4e6fGaPh9uoiLGsadI
JKHQ5OgSP0MvZ8/nVzKAPdfZyVkua44SS4yBkaeIvKtC+AwDqiw2lKpf5Sna5gxQaAJOBqGKoYnP
4q75cG7YRUO0zDTtcOlUZs6SfLhMx5Ao6qU3gh419jNYlyDZrqrZQ47hS5fg/DIQMSXrjzDgxCKH
th9zeutD/sZqKE4WOEM3+Qgx8Z663QbRJgkLeiaflfj3m8HyFtlf4Lto+si+rj+o3x8wSKo+ggbY
ZBaQxkzO3ui0X8CCjS7iFbA7RcoqrQPEEw8c7DYacsrbqVnUNRHhyYoiCG+xD4HYLN3juLmOU2EW
OfIq56sY4YO2dT9LBZ50tgknJwumXVKL+f9MByCfX0KzeNSv2zJxrmwy64jWjp9mEw43kiT+fkO3
h4qHoes2ZJPTXnm7YKORPqmT4/cH+51N4UXqc7wLLbIOOvDloGZYr/4kTO+Lhe3F9tZIQLpmK4GV
nq4rx3NjlupgITqI5G2ughRKtiyPPl6zamsqlkyqUljahbOcPhZV/dntMTcSLEhZn9SwlNE1XWIt
ndoiPGYXYWCRaoKenXYIlIbsckKdP/p6JaBphJjq7SXVFfDD7egtbNf4TKOtR5EYMKM0ORj8wPMR
z7/h8Vl7zz3L6Hj+bN27cka0Ds91vvkHkZbmBRRlZhldwCuadGIi3KBny9adHDF2a4jeQ65reTCs
WQ/H0QkbzQ4C3wKiGd7vGb+ooHf0rpB5I+iIufkrQHhZB4LYh2vzVVlpIZfKo3jgUu6luee3SQV7
CxHRn6QkT7RHK+Bsx9+FoPhVaiYXLqaSblalCFz/XoTZ7L1XwPOypjWr120iIfhtDVnDsg9htCjR
/VvpcLmCxjK9j75W/DQSimfaG7jAUjBReddvWuJsKncYoJS7NzLv8NlELKZnlubnf4ZsPgsj3S1q
QkQ+p9TxKkJfnrYCS2YWhCQLwoA7tuC8m7i2lMtyoPC8XDe3Sua9g0DMsQvrT4rpxPO1ty59Gvv0
uT0XgDtzgnB5mxRbWNk97cLdOWFhm3n/+EHuS/ieEuq5NN+f+H23F3KmYSTcIjhjEqDpz1v/bDxB
sSwoEpcD1Ec6kDYy+rP7EGWN83Fg99ewgbOTS2KKYrHQl6PxRI62RPsjGszEPHGzSM/7yRGkPu3t
KolZhjpXYX5uo0IjmADcV/wPnQGRqO8TsTr1auf7FIT4DhyKBV04tm5K0HhWumMdR3qwyyYp7Mio
+ybDBvJ46l2CA8HjwJwrhNi1laB/WbvvDsFQPmaHjQN6OZMO8R83LnpHqlDH3nlM94fcEnj/iUg7
C1N0wn/Rf3th1sx2Z0Cp3RJPnEpLtY6VO/RW+IsgLW2obaCAlnSM000COVNiDERFg2AvsH66CBk4
SvKigIQfwGtQQKDsNQjhRI/44WxxQwkIKrtQscnOEcI8NAGwsPfonfD7+Gre1A/+RWCdxNVVFPQ4
H5tTshT9fXs7Arr/E2iKLtRXcXkkgZpoqi77tozY+N5C3U2Wm6wUcWU67bjJxOduSHgaFDZCHBxi
PZwz1Slq2TqbkbY/BFLfk9qWpxVaIZF9s/415s2hb6+8Xd59Ysn7SPtlCKE87U44wxz6mNtpibBV
kDA80ck1ZAQtZNu3/UbwAO25XYw1coTbKIKnYs0uivAvRBlbiFomj6pglzxCjBx+co+1FUqOmDuY
T75q88ekyeceNzaR3QJq3dTjpE6vahqaLrzY9eTpSPrvgluOnrF5eSE1xmfbumdcA9RsvEhbzKRO
KI+AH0bc9lEsBvW3gRMEmQ1cyE1iSVhv72lxCmDPCm531wMR53sOsrqxHLS6KkTnvJPempR7I0PH
xIQ6y1nL5I3UCE8HVuuPL7ayF297K+qMeWMQdLgeofqujqlBs/eGnn0R5ckZIfcXEIA1Y3bNLlm+
hrLHak3n9UsQkjBh1/acv9UmhqdYLIzNHi5ci2/YnVsZjK0xpIqbhWtYG2rNPU1jX8p4cIW4yaie
DaZaelzA3jTTS8UWgNTvEEdQkji/3zBunMYd8nn7Z3KVFRzq/jnaGNvU8VEvzRSga+GKk+c5Vqv+
bOP6saZ+LJ3qTxiU4svoolbiAc9wIZrOmN1695n6kpOiaV0eB9iDMmaaVnbYZYJNtC2QPgFbjfIG
AGQdz4fYygcxCmob/NW3LNVSKIf+GErRJW+Rnd1Kdq61f1QRblKh01fjG3w91/0hRVZmVF41s7AX
7zRoTuTlITT0Rzc+Z/wQ6KBjJXHAOLMmWzWkOczZx+9Yd5T3Xf39kwehma9b3vC11vEfoC1s6C6E
ydCPwNnpEoHYwvxFKtCwH1ghrqyXFneTqNYCdHiNNjiTWFUQFqD3wrLsye2GYbEkeiZ+k7OZSV5+
Rpn+kt2fa1o0NKZTjlOQ9vuZnXBO+cD3QiUFBWW2FGvrIqVkwYsZoxDnvPjbFCu3b/BpLMnpxoW0
fpHRbnMROI7cpVEIGfZYQx8icPDkeFaZo8rAvuychDzRZ+pi+BncWWy49D1Fepi6Jd+xSTTgxUPv
K9WMDv0pURLagqa/DnNeyPNd+f6iB2qwF/XAEF0TbofVaFps+u7i1/XuZkyizjNPwoyUpEPU19FE
ThmhKGvU9VW5LDDntFmmbOZWqLc7sn+M36X3ApASJx49pgB53VxPUYRFjp9R+/nP3q+F+BTTtT43
jGXRq1MQV6Rr6UiJi1yk1heM/mkWOYEQeV0Hdh8z76tdX5IfvIQ8ONLlxkRB+SBOXbVaKBIxWd0S
bKj7ArAlD37ATvBj7mEgkR0ri/zx7Za3bD77rbgPiYCXm8Wgy2KkYuD0Aq2IqwrrBYescb3y6deI
uCOO4cgwJ5lWKhw6UknfgsykML7m8Q0KC1C9i9Z+vDNDE8EE1RsD44j7OHh4lkxXR4BRon5Cw4L1
uGJF/X8F2NJdifllGdJqKaXUpe3mPPM4CfAeOmqB2akwOLf/O3gRrYDFzO+8lTYHzNpqb2UfpaCq
8mN2JTGxzaTO3gqlKsY17c8TouEtKRvjJcJNYzmsK1fktBEr75zecBzqax7uhK6rv4Jhz3eIOszu
bhkYT1XrT71iGcnSaami6R/tfUP10PAFWY2EmH3y2sx/TZgbnf8ekUj4z1aNJdZVfePNoOzNL3Iz
em7aAigFCctpK3UeX85fBDXCNp/sCfhGu0qzVHV6jbSOvDwKIgaL9wqsI3u04HKK5xzTs6twUktz
SBQyLohpEimkDD7VnMusJtpxfXs0bV2hcAbOYbKK2gIiulzs0SooMlt0LW1W1B/v8HYBWVe6/cFi
avz93a6HKF91QwapBqW8dnS1C5eo/O3uPlyHgVPqSsBgTzYDIXKVobptAA8DC5oBIPW2Od5S06Xf
KFHgVhqwclc4d9SDeDiOncl1HcimuXA8rUVhEIivx8CsPuZ+jecx13+VOkbSdqkjPnhptKYm83lz
Z9eyxCMY2zVIplMQtkNt6Mi9SSYPiMkNd6KmOD8rnehxGhrd/4LKXdCmp332CWqGsH9YJtYRW4r9
f5LjCej08uMtwwShPswcphNv9bLb2LpEW0iD2iYDyBW+32/NBvNmJnBnn+c1hKg9xQac5pxCaF1e
FumP4UJIupMHXe2Vgo5LRXwDLdHITXHbhqSvCGn9FFnWxTczhgnm9qpS2Lon3Joq8P/V6WTMC02I
aVPM0TTo82g82ufa8IUWjI3S2CdHsuF4etBOEuZFMPATlVTftycMyMfIPqdOHjLkgPyL2V0fPyjP
ZgTR6BkX6eG6C3Fq0ig7cPGdYWUfFpnx9FVIsAWIgjhsmwp234/c+rI6ft2DNiV1Bz+rj6zv3rqX
+/YuoOYlthnyJc/twssRhxdR5agDggZR3m3A8IFjl+a0ddFYUwjjwKGgVdUWXE9YKQ+A/GvStv03
y4Wj3ylXfwV8MrzLmKhmeLTArjGswbBcek3QpkWeXnOqgSEgoB7TcXc5a3kR5aZ8s2eW3b0AsJ5U
twSy++yEKhLWxbFtvyalemYzVyCG4Hd6VYQHc+a1u19w+cw6ooDWPKmUOtYHKux18nJN079E9Y/S
Zk7C6P5chFUQ/TuIvZM5v+Pg2ff8ZrVVdyUeLbZgpG7KuxxGpjyVG95KYUShoZnoJWFDGSU/A0ZF
fd7acorNs2f30YyjE12QRf70HwHKmPKBbgOgtgKJRfDFjB6eGg7L81yFKYKmazpELDmkbY7A3+Iz
4PI2EPCVHNw8O4fskVuAOpGmoEPFvY/GnktI+7y3sz9qTlf/aUtujqNzJHcDylsSTJIuzfovW6et
dEhZyjw3zV7zGPL6JFgxpQ2QPYO7D2ETFDb6QEWMJMpyTx5UuuFFkzrBbODeBK4UlI11b35OgVds
c5ScNtuWSGPYsknkRkrAfiK9wx0vUZz+gFSLOmq5F0c2aN5x69kHc5pcnZ5bDQ2t8f7v7Xe/YLg1
Rz6u5eiwsV6IdYuctjqbUcg5QJdmIl+8nwvgvS2ir3UBbCa3EDTtD9vaIrqTeS0lkKtnuRmvfH8V
jAXY87SOKMQy6Yl4Rit6tM4HFNfKXvrPaduFYnl3YdqewmWWkPNBLkRI/+Kae/Xhf8i8Pw9K0ss7
g7tplXjBDv0whXSzRQwWXg9dANvvT0dMKPR4AzP4cTcrYcsUjyBahO07IIAlwBSbJAUSf3bX6ntn
6XGpCzalSO6TCN5SptwzBw8ustJKq0eTXNBccm3C3wK5vqmzBKWqZ2mKpqykRSovoX+RBMT9HBh5
Q7wPFwZapmsEfRF7roEzgiAS5oC2xjZbTxR0NY6JqqC5Qh0AHAf7N0egUnAij1dUnXrsdDO8NaFz
u4tVjaTsQv4xLSYGz5PXG/WNn+bwcIzreIwJirHl8EPvnQMoaCJUu6QASjctv4eecpu5DZAYwJHB
3zkojR254x0DoQC25Iu3eRjwZjctYMWRy13LRqtmRyFKt1a3kTcb9xwp69PKY9wdBH7dE+EMIy5v
SXLnnteppV7pP/6sYgi1Hponrwmw5qM39IWQ97vE0dmLBgNyRWhzS6W2tRntmPWDeuVRZYS1oHFH
NbIncx9pKa8Cir3bwlo1wKu9C9bYQrpIq/QGgA+Hvz7Yw2PhajrQ1lTyWVi2I7ikoLUhScOgy0CQ
cbTFa+TCeOd/0H0hIZJ2reU1YzbQN8QS+hkJFKQPrSx0ZUE7Sc+NFZqT5NLYH5KDXjgC92p1QxMl
f7FKnSUDMx5wA4M81+HuKa30yer35Oxx3wJul2MrwNoNxoBakqIyCf/i5rDddHH66rDW0PGP1MNX
LlzFgwXcmVtd89t0PuPlc3iSF07kineWy6yTzubyYoczcpHkmuatOKG0ZzVR/b+QRWvSqrMBKwhP
gduDxXsLy2pvSPqOQE7g7/mQXi0XmcuOu9KWJiERYFMkiaz3DNrgd5mZDfuI8pdu9f1I0yM6bbqX
bNYq1GeRsUFW7MJIoMD+Eca3kx4T5vJmkRc8QEaMA2h81fwens/NR9lNztLZem2gik5Cae54v2Zk
Pjd+TNB0iRQJpOcjuaFvmxrTOULQ7AqGqrXQPcjszhjnuDroaJNf0jK/GEDr1F23Y8mPcFuzpxx7
CEKVDU3pyx1jYBtucWUUq1DY/s1LsnAQSB8CFsjyi2WvFTJEuf49m8fkBn3MtRbF5U6SOI5p+38j
u1jwVnHO37HHuoh2u58R6fxM5yln/pPN1618a4LBqdfwsDw0zzlRJRMNHvfg1x+Ybr6f1RVNV/ar
Lf6QOiRYqOYRhQ244FlrmqMUJDGIVyezAlpZd9A6fwn5KFWofcQB91DXbQLRmismJELs8Rteykzn
MQ0hAm7nI8za6REvC3rmgEjhYerxrj1PFQYraZAmIxOiFpKX/qWQ55Y6sv02UPLT6qZBrV/LIbAG
YLlusbOcbXYqTx9G33i/trqKQtzKggg6jx8DnRp4IHFq2ocoUMyB0bEA2WGb5lDYA6xoE7p7fDF9
J2LC9P2vffXu5XMovpKalN0VkQ+Z4TaHXhurF1lbE74sAiWQtJvg2WutL+TCRzLYeaSxXPnFUDdP
NLQOhc4/GwRxFVrohJdKvhLHx4ql5/4gWe4ZoUSeJkAuC9tCVtEtqFgrPgKljale2hzO+8dOBNZL
A6qXCZa3T/ncxa45V/N/cDeawYZpaIsq3r5DZF0VeD+RfDghyjQV498saeoXc5F2p3IucAqVLA+P
oXwBIMjiCezqCAv1vYENBGQCuqxBW1EZGvtTMdMAyqLpyLUkmjnwcw9mydapf2dv2tFdnd6ISJ2Q
GvC/IvDBdIOSZ9PW1JUDBPo5V2H7ZmebphtjHg5VCOdQ05yJUm3b7PtHt4ueEmi2c/ivrhvAQ9ai
NSJF8XB+JGU8zPKbJ7JW7TF+Ga1bGyQNQBu996EDtnj1RQkKK/pOJAyoI+RfR+5Es6oAsP3Il6p1
M5CasQWININIX2ZDl4u70PdNIFYCG9/meLK2kxhedHJRJJKdhXbU84WNT+PodJ6nQ4do5ruzu2et
IZCHc+BvssG14DvgG7xABywL/WhBZSfhD8LlHg7TfwlIMGoN29YH757R/Uig9TgV84o0mr/q4+15
KA58o6EEt6KeAF4NqHZVCOx7kqL9wlBp6C5+gjOX7nEvbWktk/mXdsDq3NQB9RepWFkUPM7O4N7B
9hlQab00lzzWw9r3jJbg7kj7LUR1o3NNg2lXH0z/HBzCogPk6jmHTvJ0jZw9z+c+TVu3NUgaiRT0
p409qtyLKWmj+IaQdOsdwTTB7xMvTeMhCy0eNc0wAnHoAhal+X9aPUzjyqaxkenK8WghBHCeAs7Y
y9V4RxlkSuCyvI0Kv9ze3zydki/rbzTgGfkTinn3i3beGAKETrkm5kmISGRCRVCz9P2E5cymS/mc
J9ICQRkpoVrxA6uIkxGrM8Y9lzpcUUDrCFX+dErDOw7YSbUmToT9UDrTh/QI62zWt7qbwHdJDs6U
gIZiqphPMDmjE3b2Gaz/9TBrWcrBldoy65CE2/wKc0M4DoU/MwEJQSwBBVJmaf/XVT8SbuGtwHwc
oEP6pM4t5kPkcP1z2P8/5pPyaJz5q3FkrNHFegxsPmWWyEdgZfo3sL0c/gLowhXJbvvIANSjkJ0x
n4LH8CXKkDnDIRVePpkmnTK+4a2xVhBvbnXB3s+vmrUJNJcG4i4pTPUOcZ4txtJZWVzP+mVwNnYN
3++X2gn3KPRZIqEZpf1Z5i4yKUJLF8CfaTGFKOBmGx3J4hJvTdvm1pUsSU8S6qIN2kK7VO8vkjlB
VPysK2Hjc4osmre0ovQkyP9codOqbqHxSuZ1mdSUnz2BTiA1lb10FfBXVSW1dYbZMWJjy9npTOpN
HP0JaCH0u71Buosuu8NRfgdWhzShHO1BuSH7sV6pa2jwC5T025uBu41jywfnNadpX24aajg0uh5B
wzozzkxVcGhanOCPaoI3D8R+cs77RryJc46V+uAQBg0fLQ35rCXR+HtyTHLIA8GFIFNjHJdYsXKk
KfkmmPZIFLTrBRVRZvyvdi1ZKTEggGKxQb4LVZwz9M/TAT2tSeEbVlD3H9WOo5SFGnqOiBbhlk7e
IGqY+jJFzV9iB7KrPlhrf1ONA5dQN07HSPivrPpXnHdiFTkh0aMy1DOc6rm6iywOI4mbb+JFE7dZ
v2QFTuvu2KOFCWFI0tShWUSq1fgjeT+Lbrg6bM2mOI2Xv2K9Wc3DjlwfvdVhh6DuSjQjQONPIdA5
nGbQnDay0OwXxFO3fBrjngRh1pH0HDBWWEWsYlioHY2SqcC5fHI6tWv+/X/i13cIJKZK6Kt9sdpK
t89+Szxwh7Myaeqf/RFzcAb7tcnm4DidbsiOgFaevlJMF0qXO6cCUPQI+SGskcvYQjLOxRKcbCMz
ho44qkpfRF5PKpTgM6MgHNnjncvYd3hgIN2MxohT6BrwYrBMZZLAqL5bD/gMqdlW5KDs34CETJmc
1K0DQC8PHD6CnWeaYt9CVzmv17d1reelvfI/nNDJbiAttGMPnRkKJ7vD/38V/sfXbEitjxJEZuwy
ICTNjyNlvQkXehuAQUDGXERqM7DD6GCFKbii4qKwOt09Buw5Acbg0ENeAyZrCi5laCTb01Q8I1+r
w9qh8ttgjmHkLieYWLJvn0Ss/3bta+z5bGINKiEbTTV6COo3tSNwsBXYosJAX8G9lxNk97TabuRg
r0Ervwy3ryM0kFWEWThzP+b1sd5oJ+sx4cDXYZZhlJf64h2sHHFgASI9Kz5GM05SbluRQ4IJn8BG
uGlMlPwE/Oh2WAJdttBAh1iQQM94RgF0RTcDIVektXM0QPOy0nCksJ/EvXSwWGc9+DSSOsRqE6hd
i/0H1Lv3QLQRBxybOSRjclsFfHpMrxxVURg5lKkOe60Kg61wCoS+b6CLjUPX1vX99QmigR/L0/ty
eVsvJrI/W95dIjU4jy8fthgCf5FT187MnPqoAQog7n4n/1KOzdEP/86rEcemNbauXCHjhMztwgA2
XSNrRV0iD7ACEnYCYlAHmiDJRtETVkIzcs70jTDMV3hC/GrwFvV2DCFF9j4OSa0BVslb+RyS9/42
Hz/luOI8z5Ws+zaSDJJYU9XjF4SIidGa+PHKn4Jxlb/sr0ELDH3qT56uChc9FSsotIcwkpZC8S3L
UMWb5+6fABvBwlois2w7+iaOOQSMMoOENedR/D3ELD/jsAvSGySUZhBScMlz1VQm6831qREsx7sQ
bDBGmVdxsDunA/57RAB9CW9GEEm45QrQu/kw5gE8CYXxryilHk4RL0K7XrbVCz4DhFmP+w5vyjyz
KkApvwTF3nQ6tZoWrq1+OeZbMFStFpDtZlA1SvUMuxREEAyczPCsaXDdpLzhM/PUb/emkIKoAwkf
BPzm1PN4jc+oC23rdie8fVpDJ2a5QSiJpsQvWXHmJZG26kTaoippwgYB7v3XNMz/Gu6dpIqHBqkZ
LJ95zvX12cXVoMXO5lyQ64B8OcLWnsd7vcYNj9dRFNQPUPiXWYUMBkIr9acxIaU6tN6QRYBDUzxP
2H+4/YzejlQxuYTuNMKI8ApiErYaevU4Sco2YfzFDIrtAqExPCHu9I6YD55aDHxHZEvjInGFVPWs
GyF3eNBIkuMdBUDwT6C4wlXu5dTDjAWIScQsQc8uHPin/xpg3iaMnm9zMu0PW1COl90xW707F/0N
nbwkucgv9b+DPi5zx/TMAOFGq3eLVfhoEdd/0M+2s6biz5Lepq9Fq3w404WEuEcC4D319Vqn3ltz
Ib5sk8lZU3VjalZz178ssWQGU3koPUq3p8mbvx4axAt1dV3V06UuPb7lr/pAueBRxMIc6gx+teOZ
JbFA01QiwOVpMPQa3HSGoshGuA6dZcNRE71XVVozlUlUMah7OocsIBpEbpCgUCGiX2bXwgruBHGC
U/0L6i8ABPMsvykWfx3r6WuVEFmflR/nartbLZoUQ3mDAYyokWTD4Si5DLNn9dTWU85+E46poSjn
m8NEiwuDfXNNtFSuoa0RTdrGdO8DIkhPLuD2tmr3TkyMYZb73y9nd+g+TooTg+nLkzW72Q/FSfK9
vehHzIZr2QOHEVxqTqjVLL9U5uQS4iJKkABO75uFmpz1cfP6rav8XMp/XUuBEPGQ46WHuj9TQTjV
Xn2pSLz+BnswhIeSI3iQrB01h78qom/p0Uqvn8YSnc1FIne+ykGo69fxEG0kTb/yCN1yXAVysPh1
Z3r172wdCYAPD2jHobWuDF2jd1jeSEkfiD6C3+/zzkLVVvac1zNtH2fRXn1+npnYiKLGvxqRw/rD
MzeU3UZ9eHtw7iDr/hKdlgg28YHX91248+HRWFoN+jJux123F6v/uGuiSN/AUS6BR/ravhT+GrFB
lpHfnMrD8iznV6nRlQ6BJ1es0a6SYGAlnB9i9urfrJr8LTntMl9HkenG3bFzFPE94NQhFMFJebA2
DIjn4dp0Y1McThrWmS2/UupqN5HB4DddZagHcOHwUonwJ9gljBxp6jLjKmluzAICpRF3rFOA/9as
SLwQVfpwcpjorJqW/mKeAqf3x8gNg298pvH5DvEoohJ6LxH5ppS9QB40m0yW4qsJuFuT43lLxOvL
LRdfm2CZTXfeaCTVD+36+h4Gdh4VUStfS4/BN09pN7mkF5S5DuhqqpIOWfUbBPYz9PxP0aB1h4RO
VOoPCEAAgb0MkgClARY9eePc9WLvXPyBjpQxwmELiSOJgrLS06VWh6r8VzFNGg8lF0Nbh/BvkUgc
H8rot18pDdLVfQqBIAYlUVmNz793f8kt3ApQ4cirkCMaidA+0wA3ZrxnIBCDBUCjBxLUDPey1G1f
ftwXcI93NaYeihtkI1Qc41G4mEO+xhxKRaVZnJm7DI4SsQiVtjiSuV0p89nntzht2mlc7FLRtQhn
lXxe23hiK3BP9UKsqGJvJo5AEHGFE6j30SwSrKSNbEGVo674J2sZ+Ac2PfZmPDiqoa/tdoMR/1Ep
qyn34QDejzE/JcWd1+LB/mbH6ZUnmKDwW8RRiucf1W3AFOA5Wfv0UUTQraXfK96nHKG79aGiHKPJ
jxfzS4fxWPUOaWvzkfGIB93jpfGQzbMKkRRG7gwWXAVEpTpEgtwhhOv4LvweK7BCb4+a+YpSPqS5
SgIh3efZU5TMI7moUrH5CA0p8iNOEWkeiAC/kuXjbYPZkeSqAdYPSHCQLFW4SqZsL3ZodPizqfxa
7IWvDkJjh3IVGrrozBzOyvDx/6AA/epz/Ypa+hrDnr5t/ujgYPu4sVtdJDGj1IthbI5y9uS37hUo
ELJQ4rrCMOH5Gu0F3kn+qgctZbw+vcu1i9kLJ1CXR+MI4xgpS03F9NT8xQ5KFQ1BwXibQxlL38oH
eeDDNUC82hZDaFQyLccgNOfqwL0uOdIlne/MsO0MTik21ySd36CFWfDDEHXcVuNOTvY8YXelNEBH
kH2Dwt5TSfABicv9ISnNO9VTGTN0jnyIZXkODIRiytB3CReAI+ihb7ISnaWl/WJFFBWqBK4LdjzE
H/vxf5xXp9f7QgvDece6T8R842wSX8+BnYSGp9vMxSQQuP4IJcYYD6WArzGi/R+99MZvbBhF7mkH
+4c/cVnTkR2osbwzZZhFNJ2Pp00iYh+Wn4o1mW9Nw0+cGkp/KychEJA16LuEA+dIUZAkvtnvWsxS
VWxTnzWvJTVKTNkl2tNyQd6MZj9/FUSCmvaXGk2phWDG87pWYJJwgP88hc4Yh58hQhRZ+yH61Y5I
53Md2xCp448SR/xmvTnFSfaGxpB/f0FO7wfofW8VEDC7R9Kok+DwNGKd1iTRTjh/YS9Vx+J7YJnZ
DULxWbuolIjzeElshwcar5txQUhOkIH051LL/AwZtkH6C6QuROsB579jgwSsr/nS5OrKrAyAJuag
zoIjKirAG8h/O8i4NY0SjzkQ9sd2aYkK2kCJXTLkmdFrZl8G2D8ocpP1XzDxtYsdOd8hsqhv9lkC
8SMM21FNxIrvQt8Or63AXN4wjPTMLux4AiJqpF9c2BDQQGJGShjnoYAGB0eOQF0f1vohREU5uSGX
zLmIun+T/UfBLkJ4IHJVeZtroDJfDhdLSwfduSKNIdlb+v0Y8XyUVlLBCZ06tH81li3omFfNxNRI
B+FVs5AfxM9shTawz/+pz1eVuupyb9wF5UWQxNVynpX3PvYJGTff0BdQ8lEhtp74s6ftmIzISDWq
VsnyONPqgaIOM/6EzlTB5DWo0kom6JPI3EVC8BY+iC2CiOc7f67yTrjY/282wmiXybwNPP73Ug2O
YtWipsfoAm/ygBh7iSlEg7qYNI+q88s7GnXWZ79JSuRGxHrwu08hdblPZV4UiPj1rcOVysGQYP6w
WN6C8zkMQ0c1eyp59MqypK4w84QupDxpkoI+J8cpfzuZiIymxkWfJS0/KwBpH+BdauaObfC1HgB4
lMFe50xviSZZSZcHYW2XjPJl7nvJ2gbbfDpxLrgPPN2lL5r+WIn0E6zHMcf4s/CuP7sENpLVsXaW
h/ANPtXTmw92UyFXGXXoG+q8vC5jBbKlk4XSWFa6rC9z25fDisRstDFOR1e1B9mxn4KVBXHB91m2
lKnYhm65vXDnqU2vpaNrwjatK1ul0deRnjBUiAZwcJb8zZn2rKfU+qVlWBuWCKTV3a4pPbZWErvH
x6IiKKLaKtdgrBnCEx/lWbzTdvZsrziev1aPx97VBDBBOQGQWGUHcnQ3a02vo+5aJ8svmaV8B4LD
m3d4kjMbIgQ0IRYwh/I7+GG1oZnmqTXSqzPm4b4+ot4hkwpUNcGWpLG0TQasffQK49JJ9EArYziH
3dxCJYCEs/wfAg7eKCmDF01w1fk9Gaxq/bOgZB7o44B21A0q7l67DVQS/tONh4KyhtM4V5vpFUId
Ii7FqH99r1UeOgEy0vpzZx58IL2qV8abXAmcG1zq0qlBVneQ4uQDRerJyC63Bawv8fJLT+WS7Sdj
F3xeka8vXIHcDpK9Yn2CA/6S5xXbyZpq/xtttCAVXhqU+/p//dl4bAqE7U3LjKP4WyuEcLBwy4gF
cyoFCUUX/QXG73OEx6lKPrCunrDOWUWW/YHhGq8FXwqhM65pt43P7dLrTA3HGZsJD/3GS0IVPA4+
gwka7uiu+QfIEq4csszvhus5Hou0lRkuLYlTK+4gyZKKcN3s03yt+9hDm+zJQznYJD0798P5SDnb
YVa36PBQyr50smc/0VGGbGML/B8aSsb1mKlxmYvl7hNXJqlYNursuJtk180FaHCQNka3Ey7suN+a
GANfel4W70+gSoFfzu79YyZpIfrSwiCnUjuhQaFov2NXUi7Lfs2g/iZbNyGHYLUqkoXVln8LL2XL
Ct7qrhFs3NtN+bJD7z2KY4qgEMQIwONB3gtkhBx3NUOOSTiXnw2BxQF7rtSZl0x5E+pCAOthbazx
UQv+QOFIqOLzl603gwZ3lxGVezmCucvDfiKLtR0awzbt+RXMO8AFwuqvX5YQp++ywRlnGokAVXiv
HxAZq4Gt+suhdg7NMvnxiIxxJkt+ZdBZwzVZXdUAe7wJIc2A+dbYdZp7X71B+xRNxMnNcq/Uu1GD
Z1vmHLQyx/zGLwj+HFDLeTo4AHl6mjcQYKtJx0ah0Q6eA4qGXEa5Z/pPbaffNusMGrqYfGSrBNiJ
CNZB84euwuLRI3jGN5IMbKS/UxTBU6Fqyc99tOyyCmg5/y5F9X2wvZslN3bgUNHZo9+uwOGgOxWf
oP65o10gA5n1/XCAJlMg6PXlNNNn+Cj6+EivYE87KLn8dEUfjE0CYR8y2vw5U3rpci3IfAYJ9uqm
NscIHIBfBtJuZ314vggVIVxQnfgvYOpJ8JvuYoPYl3Vb4Au+25dG6U0MQu5lAN7K72mwFn0fCP19
enhyu6TD1mo0WBHCNCPPjSsTBj3QHy8Z+I3m2de2qfM/kvUlvn03cNRpUcvPRZxcHYprvWKKq0GQ
dnoAoT/vH3sh0Fz9cSuttJmCtAhF0nIB+FKD6K475i9ELVtVlb9SsNJDi4cM8TBeFwAwDP3xYt41
qwXrdOjYGoIz3z5WBLI15RCZWaXEByPVbJu3gkDPcVaHlAyonqxuW1OMHotT4S694XQicmk0Ady2
QxP4gjp1nfRpAFjUKsECYOVlcaIXqiTwupexgYozRDfB22w2dcqz0qNOP60MoZxdhn2a58Vd7AeX
XehyFsg3q9wcoM09MaJrIPHNnx050p9u/pLNVcZiAnbWcatUd+3aeqT59xVn/lJOM2Pr/UABCDd4
USYuSt2dqXQtix3I4BcIVOmTRE/mIAIdo/ecVRuUNKqjaVP/PFnHayEOk75gT7ohFzg3VvoeXN4W
rhyEdM0vgqaeBVyYP6DvDoxfi3iSoUa0YQBRpjGf9tfp2saMQmb39VXmoikkD9QcLNNdnN1kzf4P
Fv4ESA0/XrniklluA4zEI5pi7cGjFN/VMYzF4+p+/irikeGM672zzshl8kdjk5d04WesOeKg8LM2
DZPup1tCYgkoF+8WTs+02EZbtfJRSMJqXBJeDqqbcGThfeeNDY5l8FbsFajZTiXBHFVTPgC2UM2t
oqlyqVmmGPmNhGogtZ0pOAHKijgRsYVOuZpnIc7165bPjDZ3olgeNsrrAwn4UyEF6G0llY9vyNYE
c1ayvJBEtyYxJxVzaeyyZbL7MIIoaVwwnk6fB3qc+sYmE1vb9pJ6GIdLlPeYbwY42jnW4ZCQhzMM
d61xwjQ33Q3kCSXrcS9zikXVGSPgA3uNvaA4VeDpXxfjKQ0Jw01G1dgh78qOWS5nsfV1WTY8M3wT
KWkyVs03XG8baijGO29N8lEXEG3qrK0CUF7wZi9SXW3hHzsW819qdjQ2vVek1I/N5iM8kWhDqNur
Qn49ELKq08AFCjUhUwD9FbDvbbJVNY/eBMSldA2ZlbLFTOgVvs8II7L67Zh7OrKH+LpN+ss0APzf
PbWAd4idN3Jnfg3rjzTF7b5HPQLM9q2RyfKWIfUJ3fRaIUiTGU9CgiXCssIKN+Es5MdU+fx8G8re
6OLRKNYPsVWMW+Yyc1j+OTCPK8b1GP0tP0XwcaVx8jZvaVjslT8BPgGi+3W9rTCKWWXbLAAc7JJ1
+I0zAnOlc+lsVSR7nPrZhHTZsHp4bmKlvRBDbZCRhi/O+pVUCv3UAK67ClqYUjP6Kk9IKYwyJwgO
RhVuMc/vDRKQF0ITR2EGas/E/rDLqEY/crm1k3+UeCvtZZsWJ4Gacvfg4QlaCdqzN+9ZHah51bTN
iMSC2vxqi+AaFsnmynx344PMNmL8z354L5JPi1QCg3nu3OXdgwlKJ7w4CNjTaVJCe0iObBX8Do2J
nfhAVuIQ66NTYQ76e5icrT18JsskdW2FRPTEgNqxN/vjcQpHp4loca3W5TOPD0w9upKeXJjl7jeY
O0DqJ+dDg507WuLMYDbLJdwRgP2CUZWN4LHpHwGJSa0mYiprT5M1QV3Lc4lFULMdwjfkLCflsk+B
vKSKnkAj2263QjhyxAv4gZWs1A2DsG0M0xvF9bIU+GYEjrcRoEOb1W8fbQo72c+Ji53AzCaIYc62
GZTNiAtGgIxv7wgWwbN1XPLLK7E+RCeTfXZSZi2qb0QUTXptVOLYKFlPdlRIZdfOTnyaapAZT5+y
u/fzNE67RGz4TwszSvrcfbz9lR7oaEnltrn0hah8/N3rWwUXeO5U0O3FYsjARb4rwHsHdq9gRO1T
yMsL+vdY6UYQT9ACaqxrf0TlWjHjmBl++LkMyhwp1NBjQ62xZT1NG2zDZRgfceiWfsNrKqj9tI9c
AwGSjmee1Hge5ehtL5OYx6BktV7T/tfCcCrbqFmF9StTSTwgDxDAmOuVo8/s+XG/nEoZ76UQYLa6
8t7HYEOjVxDoYIDtZjG1+1d8B2gFaSxUw/CPJxTTebmGHyY3MZl4OhyMD/Q/UtgXiXzpShpVT2sk
fqcyeKPHoInuvI5VD0COjAjNTFK5vn0izP5af7uuuJkVlHvkDcGWDMf2nrrRHjiFRvBW7C6EGRF+
On2ioiw8JPo49EU7A+AypTY/fRDJBTlcBIbhRBbwRa2CUf5F72725AkhOVrtpDQj+s3h8fo9oRUm
GI4WT1HSGJlCNJgWg83EFrQodndQ65/garL01jPBg7UN/2oQAq9sDkR5x6lvXzfJuvHXUX+kFcMC
6X6iMLMDlQOQZL17JEPOx92rQR0xPWDkpPllEOahJyMPzT/Pjqp1JQc34rXvLMX+b226vDwEUVKc
4Z3a9jLTRZWlXli5boVoq68LRbgHdaTweTaiFbFkQ+GPP8/0pWqXjk7EI2zDl89zlC19gKkwHP44
lX4w6zYYyiE9lUSx2n/FGlFWe4k267/AQjwvdTkGSlPxIRC4ZbBxKX4OvW3whRF14hl45tcoVZTl
bMNTG/pTKLW0g+y5iiWMbm1GRXouJRFQO12bNeUSuJOO8O31HvWobylNt5dCg2TkgUS2hrFYFuPc
O9zfcR77WaHq37KpTCht+cW7vy4zkiTq/ROCdcsUNvLxFC7T9yXw+tNGQZ0THUFw1hHOQw33NFe9
sf2hzNxfXu3YYTNXTpTRf7arINDebFfGKBkIupEmkVdYrWffDhfhBauKcMseUftUo3BBjdmtpiE9
EFdW8fDw/bcIhPpCgspZq/scFfaOTYsg5TLBaqUsnfQfvonopAa6XuV7hp71YubcM1aN5ZJ35IBb
PDOWOHIbRaQ6I1t5zU94r/7EFrdfedXho5cCvzQuCJmWbx2eii5Z/m1sYwu2HMQukEM+vTqm3Jt1
NrY3esTogUmqR4Z9w8jNInlI1W9hd6BQP0O2fLA1Zzj56ljNnzDeNbbmrM4S6yuQn9HK6G3Ld8ec
nl1U/gHjd5+r6UXw/1RYBrFI6tg4fxCJcze6IT6hG2CgUtXABtJY4zrjo/BugrbnPNqZ0z/M3y5z
1Pvad1LwUZuJZiVBicVFl/EHrKIFov9RUaNRYN0YSdhRIS/QK+Trk1j45aD3n9+v6uo13+YhVU+W
1AINnXC/Yukid8l7TmWPH6p79YFUTt2VzAVhjNvyxrqXVhi9I6yfjPVM/Hn1LIiRIpLv9baZCKgk
ZDhlwWKLBqMuJpc/CQjvUSZFTF+R+Qrs+1zd8Q1NQJ+ptsqA8OmShU/r4xjDZj8O5ySaUIeR5X/U
TzSJSuoxPUgM8GAO+3cjj2cANHw9EvUqxZW6PQke+BOEkWn8iGxys4EekHOJHJJFi/7Ge5afUYJi
XjsuLE/u2kXJcWhaWpf2hkTLZKfDcLILnrZfTOeWnRhB6nQZ6VmQBHhH0KxTWfd2VJvn9j/TKPS8
J5yglhCOFPNMZzHe/DQKams24Sl3QTMzuMYEW/2atACW/JLR2cGThP3FA8PH9KdPkuAj6es91pof
fb1RudtdZes21LuKnCQ2+z3sr4W90NhFBhvv3LaI4OFoHJ0k+2rM/Iuzih7weMtgX6oqF6esWqbc
6Vu3IMD1DeumNzZmXxLu8r/+oYvWazWgrWNM96zk/zgxqGInV8jwTkEsQXoxjK9MJ8NvPv2+D+5d
0B5qb5tC8i1T+g6srO9uD+3GWdaTGFTMreABUR4oNm8rjFzpc7wMAoRTy59JqMb3Yt5zlc2FmU6Q
CpcFjUxuVHRC5mHcm9B1DdXMbRxDLzAB6y4LNuRM0dkHnpnNu5fRrn0KaxGW/iOke7VK+TOCvwY9
u286BhtbsaZIK5hdi/mKZdKV3oUeDBXw0YKf0CA1x+edmsheIPFpNFofGiyERWC+81/i4IPiPcG3
iK3n3+dMXutls+PpjYd0s9LheR7JvPz1MARR/Lr4PjvZ2tnPbf86eshg0RUAeYQSOkFKwoMW9EmK
Ud/SYdtOzt76rhM6xjd3vOvtBos2iVj5yQBTAdp8Ypar/LOp9x6+sB253aOGEi9KtXagtvMqDsNR
4tUr76THgSbmuBhLyONREezAjVK/5pTTvCcYj+bFIDSb5nQKp1coBUcBqQ5hrVS2arqOnRw+S4sU
vwMDosHiOHHeLorKUfWmeh7pIQXccofP8pG/fZMaahs3GCFQCVWyR5uX0cadGq6y95q/KY+O41dn
XGnJdnMXsMHCUsa+NER90GxCQQj7S/LU8brP132kdvoqXwxxaZkAZAodHvRMVWDqjN9SY9BxTMmE
ZhrCWcAfG8uOdVE16faMUREMXCHt9gLmuUwmtzMFa1tFUll6LfCz2knfK8pc1NXMwGs/kZIu5ZJy
cOnZDlsfRPEbBtI8tyy3jk+5L9s7fFsRHOinY8gbz8FEu0g60f1mzcUfIUXJ6gd5X8+mprWIt/Ux
GJ379C7XyYtbX1bXU7LUSgQKCkvW/DI8DW/xSF7EApm3V5HQP/MSkg9jznc1SQgxhjQgJ4ZTZAOy
ZPGpqUyaUaa/PsKbd+6OLyAi7eTr86odJigpv9viLhFKNrr+G5nBVVbiDY6H58H22426KH9A+HpR
MWxibft1cDfPqgtvVL9rszJJO0k9v452lRALRlL+F/SVfgRuQ5lPQAUEUm9fJNyUfUANhncA0rs7
8rUZoKYvn7PMyOwgeqYU7MecQcCuvHkgvArZKP0auc5Zv5WrGrAleZXQVpXiRBL9zs1MLl3oUbSP
OLDilnjP5iTuCsBoKZAKr1joj13N9f4SLDe7FyhvuAZbDvtO3daHgUbnfO6RqeL71D6lUO6K3A+V
pA4ksQglQZBYVj6av701rUiVF7CRHAwi2wJpgdsakJdja0u/Saaj3cZtgWcKVwBAYRHSJbKax5F4
mReZ1PrFXPseNCeicavAK0Vd3G/cNbABtBMZ9voI35/o4yIi3+0DqDKO5gHURS6wocC3gi8+UH6V
hXEkabLRQFol3F7A6DzhMQvMqxBibIAp8+It1aJn/ZNgR9L4KU9aH8Wshss1MziwABKA72GrPAP7
yljHFfmpB3VDxPz5U/FKz4DEAlGKNNtenl3mX6TPaRscYGOAzXtGmnikXoUjc7s/TacF4nMPMWEH
PmJNWrRSwmrfjgK9X3chBqMRYxjr3EcFRV8xrcOGVfFLJlj9SnLcIPGKm9hHthERC5fsREIEPrPt
isrQoYySzm/988ccge4zB175fkADBnl4mWObmfM5AfHvne5do8s+WKpv4LCKw2A/v7VH5GTx79tG
XCMektPkco2JZ60sUBAtUBpnzJ7PwkHyMmUVh22ym0cqMV+54HUV/whp+ld+e2HsDWA1zXqDSWIO
oYLGmbT3CBecTGIuoodMz8+borAmwQaXjJ9Jtj+QSlmGnOtoMfr0NT8Oyst+f7Val5s5Ue4Is+qN
Y6Lg/JZWNriyR1/+6q8b7luk5OnM/AFV+wEFgJ2l4JhGOPSAWQsBYjGSHWR4gtZk1ppOyGPBqQHN
Tp2Jhj0Dx8z6xb9SMAUlLsx9KdxgJj3R/awvd+52u1rkiNSs56Z2EIXOi6vlHGY5NOod04qN+xtB
+P+U56fcBEU9EPW3mmgkeyiYKqwfaL6aOtOWr2jIexZOWpd+NWde1PLDYSsTAV9iaC0NQo4kMOMv
918m3tPFkLGOr7c+yGJ7bfnnlbvMsHMcMXFEVubnX4cZ8AAaK2k9DkUGu7/NBI769wSdEGjboglK
IJnjIQa7OENMGprmD4Ng5W0I/pywHUwWyYJe3pvhEgNWDmD5SE0rnVYdUkiHyC5TDwZZ7rIufzPy
xgj2j8FyjCr5r5xm/CJkm/fkeqTVhAwJ8nsqpIzFslmgQdNZSr51XzGeHPsyxoVYrNN1zntxf9i2
SHQ89Wm85vwjs0sW5+0H9QlFfinou6dMUR5d+n4ozJogonzIMpya0kTKPogrtqj3KfW7k/OABobe
XYUJ2+bfJ1xILJb58xkl1iJnolMhaYys+Pk9tOpdk0k7Jkb8I47d/QnA4vaBgFQrvuL8rBjMPwt7
1+SHKKHiapwzr9ja6g0SetvNXf19ymOqLNW08Cs/nbOgdwkfhb77i8YG205LSEk9wBZy1TSYy1K9
vQZd0XagnCSZFIZpK4+ZtTT5+Mj7UxaLgzqAW5bQyS1mTeL26CLTM4bks5vZZSkUsBR2rLnuJlCl
nrOUSz5L1BFl487L7oFNryFRhC8oaboascX5rxNAaPEkSPH4hqu9OqfP7Dw/T4TLIjw3zd+TQkSO
H7pEZ0S6tmW3ARHAxioCW+Tm1t5xq/fGsSMtjwzoltz58Zdrlyh5xeQCgeRbzoBghdxz8PdLkOkO
tWFD5JMDa80emJlCk0L9sahu5S/VbDAHEdo9lfgoZtvc2IHNC3615bqvQ6qBmleQWxUXKqtQSnoJ
gj+UFnCJBqG2w7r+HGQ706LR1SYPGqLmH8qfdavNDtQVUr4vovkYnVRx9U/cMMpe5MvACBFiP1t0
ui/vli2Ao3KTrEsuJKsiV/6ncRe9y/tgWbWdy0K/m2c9czDUUuR8YgcntP/ka3pduzj7hnOWioGf
U4joUP+me/EpCCl73KCp8zHirmdW6MEs1+kh+ZirWTPU8JQFzJVLVcjHo7274HpBWWMC4ufkbhzZ
zkto7sdu58kb8m3bqC/VMi0xRVVgWOqES8JR3hISsnRKb2qZvfTiebgELYUhuL5jo5og8Bt+UOTk
RxvWWgBie1uFwR6CXMAinai0rnOCNWWr2/DjGehg6n+bhdGtbM/lwRephv3ryhTmzndt5vMHI9Yv
DhcMZL+Cl7UOY8Qv8aQ6Lay/ZS+E4lmLtdS5FjZp2KCWHk116lpaXkWYcE4NOwOhiNbbIO+M9Zyv
qMWVt1qR4cVljnxgtFPSYIBBWy2fG4og5f9BlBJ2J1BKptO7ixNGc21/x5QTxsO3GXstWnNNrBVt
GyUPlU3bMdyh5asSxJcdCIOtmyHZ6j0LT6NY20dVJgUaWuV5Qa+tjCl8O907H+/WD30+9KNA2C0e
UiHLP1FZZFTVOaVuBAdADlBR9I+m8fDDd51zPjisEPm20hSQGwiFIwz1EX9ESPaXS92AeRHVmkgg
nz0qBH5kwN7hqwLkN2mWSe1MSpso5UoDbG0Yfm8y/NlWYmKkcNFHuuNb4I8Ugbk4W2wDsRG8pHCn
llWc7DN+WDyWHokkP8HtjhT5nl0W8ASmPV8vnFTYN3CfsY0DEuWCJYGg8VwXUL7JmA67R1whsNSE
UhclCFcVrQ1aMGpkBRqlRrOpl/V3m5s2G8C0qAHhylbak1Bw2p0U6PpITj7s3nJkhsFATbTZg0Pa
YVOdZtTjXKBX2xJuABg6hOwZb8Vi3LTZxAFzSAB4cQjux6nStQJKwJDMaAVZO++hYZH4+0nR7CMY
xXknDplxNSDWPOaOx93djE4ggh1cy68MaciBlVpVFsPmV2VA4NbnXqGeThRW45JZGg1HnkrBMAQw
BznvoUStxAA14BIHoWrYNSqzeccNB3yuLzjzKr1/pVDMWp2fm8F0cr3v4J23d3xqB7CXL86eHKen
iV3ub2mAcXniBA/qWZSBlOAcU3VOVLo5y+69pBcRx3UcQDsV2RSWmPa+NiLn7TW5EcFIvdSle311
28H/Tn/bs6si1Z4WAyzs8peJJ6PTCeAcIkWQ0XT6F5fS4wEiakgFxYhrcFyylXIhJHgbMGHmbhZ/
RU60naWR9jH/KXYJ/3DLwfftB1aWekdm9wiCJtEQgNVaeknThks1ZsXKJ6uUiyivl0MagiaPGtih
E0fIswbLTiUlIyGqpMZ1jMxG1qTU+hwyzM4dn/ZGVDEiJOZ4Rf2TdmI1X3/wm29ycBbsyoehz7Gu
mhLyBYV3+ga52Z3PvdG4sqvZAW8sww6orTBSRM/wyc8m76HqShO8Hsp11z2pQwd6Xt1k+plt7Neu
t+zGKPHbAbA+rFj4lHdkG1mahNifyvFlLFuldr8xX26GVi5+c1rWgQO/Jor+xawNzDOdD72qsEuU
QXcXKoN8IlZh4YDzawhk4058CdjAiLJ1sitXlEkZuJAZOvOqAZF2VcV/9u17/6TzM4IuNNOvVHkr
nGE2Zm5zrHpmi6qx1vN2fylEui5Vx/deUq8aGxRBiNaGX3oE9raAMaDWcrMIsZrQ/VcpGUWN4+4d
7ar/Fq/W/e/Nqf+BG3M4+CvStK1rVmcsCD+Wb9g6EWqZEi237ccvtwMd2EflOjP55Ba+UMykK7xZ
zKxtM2aGIzQg4j5hQ+tF5SkaKL1KPwJs/aKIbamJfJq1AYMGTQlzbs/jLNPHTx5JuJzrhYox/BKh
z7CVfHWnJ3X96+0J+vKuSBh+SuOQ9PIjGuzQOipGLXOWE7w+mejpT080l2qnhVHSRAB8Xpc2Jnuk
Bsn8HXg+aUvpKuH0QNwsQBDDqlFFEHC8CWaPyS12FlpDWEc2W8qRLjLLC5Ean+O9Vc6cyMNgxRgY
cRVjD2IYuVqxq97oTE5Q90Pn+eNZr3KXyRSa/FKye3pVKNVJy1ZIWnAqGD/Nw7Or0AfU/RYQWTaA
6zxIebs9HtpD4434n2DGCkdVdmXm6loukTA6K+62AA7PSacM6N3bUeTI+vCI7rRvVyGWYf52efIz
NqfaLKdP771iJdDrvcDFEktZYhe5oVG+K642fvoL0QYvfXjUrxiSmZDu8jiwMeq+VI+Wipl7fSe2
+L/vSLyCT8fpYNc/tFT21vjaazZaM91r9zuXu4fghPGnvxG8XrOnZN9LkrhAHzNTnLE+b4h7ncDC
jONkAoHT0JVjXwibtGIXYXH5hmNZbeTzAWElzDxvJo1bB8s5ddGrfWleIQfXqXPrtSYLK507FD8a
IanSCMdHZEp/G2SIgjL4yjaQKmE8RxbSV4xF9EwmoqPqzQWvdABzaGqDCh+bd3vK5oqIIUSIMKSC
rc2i0SYY4GIY09mh9dq0ufH9l66ilab0YLhrphOhyfDOhl+rPYWZdH0b3h4mB0oKi6LAZKjjfw68
F+xmKje9HWAZcN3WrDcoM3HEwo966QZCgpAd7xLm9y890xDMAg5YLlpcCtjOxmyWknIh/mwnACms
uqfQ/8w2mFK9QN+8roIb032ZgPxxY3rSmoAs5JcAsn6Psp2+QcwhKvN/MQ6i7E1HLOEo4riqocJC
Aq9+X0FcYG3kofugUdM0VNoLXrE31dQfQ79ViBfY/bkEdiXtxyREq/FDI2JZMXlaGOp/Fa4Y6Me1
CZqa/GC8afKKemdGFpXc7LaYvbPXtWxz4XiBs76MX2saavdZ3xkN6u7NEp/BDC4sM1sleCxjmWsO
vhPzUTf94cEImgtz91g1ujOqT7MMJKR8fccWvIoiMPfHfwwH3FCVIIVBDlUKqurvf6aK3a28B665
If4Ebd52Ii+/8NagErBKmHWl1dSYFxPIeJ8YHGPHkJDv6kPfM/9odcG3N3YpKujGQsG7vgqVoE8Q
jKA3HZhMCWCSJsNJr0GgY8BJKbbwan5DGnfymj0fYLOIw9haylCS4YTntSNcIsRV0mf/AD8PpvcY
K2WVz5J9pVSAP+BUMZagFOkD7Ns/bkfpoTRdeNwankh9GdEyy+xjeMJudfUcO6QLodHn37niSsXe
6zWFjY1JgJIMknZeDon3Ofz0ZNI+brhRbGemPgG7AgbyxnIOBMekMn2VbnwehV7NfzPEdZcFU/r4
QFrE/S+mfPBZW+bCbUW6P30xHkqm8lQTdSU1DJbegMXYOFILHEN5wajd8x53Ixujd9MdoijJy/Y2
7YsNOnsH3RrXwrOLxtuQWRn1dRcF4+g6hplmnK90Je7iHgdGPfC7+3eJECHH1TqVtyIMMQ4FG31U
3KDa8tgeBuQFdenDV+c3LRSo1UJTBrrB+eq4Uhew/HHo1qGwnM2NTL4lwJOnHG2zNzJgZ3GzSpdw
GzTXFLVfysxvY0hpQ7lAyWkB8gT/gteD8CnpAEm6/C4+Rf3RamQjcAWwPvqO+PF3f6l5E/LKVC4C
HgvS27J1AKfz/fWrtMzf0FouRCg7sn0do4Dz4kd9e30gRy2nnDHHgAkdc60kodDWqw/hnkv2zGzb
g26cpm1whLB5yncw1mg/T33pCTjyhpXpsZi3PwDbxEk6IpeH5Ik2nENHic4/kwKqK5biBsqq/3dT
ZRhwiz1KlIqp58PAayUmJV1sI61+V9ZmRCQyYGv2O5TsXkDv9MLJzZhyuzAm5nQkUxyJ+U28z0W5
y2UPT4Jyts67NGcjvWlRHQCT5HPuZVd8KDeTuZS9Vt2s79ZIh2w8HlKg7vsYteZHumwad2Pptjaq
4vmDkEp2v3+EzvSxaFsJAA/0sF23cYlDszqDRUOlmKhRHiuuqdsH0rjZ0/nRQCLnczh02e/wYQsQ
5cTf6Am9VXElXHUHiEa5NlikxXFq8ZBhOR7lbxrOChvUCZX3qR5zepjyRtW6d2S49rPrnyC/92lA
2EERFii0VNzmuNHZw3L3p3lrDA+wblFN2jgRJyXaV065ucXd+3zntT+ad0hPSkKSa9oqjnXB46fT
wvcJtqMJefMEn0B5x+qeByTkiYwO4adx2NimqIPf9hN9ZtDM9QYc/xWI4yGEnQr0cl3mr2+uRyiO
J9mARYw/w7LLx+tNxYaPb3/NL43R9R/PAI0HDyUh79uO5UP6qsjGileeb8jFCb5JKoApvinRL4QJ
rMBisyjL9VnhzHSQBld71qRvqS5Hjn/IX4p/ImX1PyphvpMqe3KrCUUDo6GAdxDZc22LWGQ7bJBy
MnrZckOZs0eFTurHdAWVr34Js1XF2H3LHK5Li2KmZW2AREXlO2K2p3ZpVl+/mHZ36FGxyyWDQveZ
YkEGbftrRPIWqgvpng1MSOMcQFXNgKp1ZfA4oQznnoUvzv0NwMv+4X25TPyeTWGM8ecHFhWdzRDI
ij5Nfj8FCHEAnI8VWTkrK+tU34E+Ahg3vFqaFV5oPsw29FfqKwpWzR+S3cOV6JSwbo5ApEqPklUI
yLMNZcgSP9copwhomIkk7YwQAE/tnbOC2Qar3tyEPa1RQJdLWFNVPCdNbvz6XSFXyhpkP+V5r8CK
PslFXAxflPDgr+z+BjJGkSC7kMaYhS0F83/NF9rIR7BkTQFLlpIzak8o70JlVxjiAtGAxZIRjQMi
FChLCfDyZH6mDPqKiCprkM6/fLkF2Kd7fDWSMTkhuEI/kXhNKoOp9QgTCGFpsYnsoQ/o5LyUcx0e
bev5rJ3jyJtSMzPk8hRphkkYWMfj8mYZffjEdqhFYxpNM3oTVbF62LBYB1GRO9GM0w3y4viKY98V
xfgypYk3qir9RMZNZpsq4aJ5yfR6hiW8ZqY8QXe2OouWfUsalv310+YwJdPH/Wha/FVh93tZyNp6
YmRE7nuCNMeMfCvoPS8kb76etSiKDEBWW5alZ3BIjbCgfBlgXp4Yzu0Zfh/lxoadjx5qCHL6i4Q4
hDcO8jLoyhXpuPgdgs7WHSD+P3FxCPLgiXAM4ffJNCaV0XftdzkPCiILScPYW9n2q87F/o0F+ATP
n6MY9T0oKp7aQ8aXQoELYbwJNzvRnIxH8RG9BL8TJ/NgJLFbqWRevpz1XP3thItZ4m/Vi65cDKpj
rXoKnPP4VUaw8IePHseBE2mCp/GGFN6BXhdlhG4h4vI78eW87Hh6IeEwX1cf7dWH8oNdznICQmN/
Ye22ahl1Pwh5rzEfzlMt/upOWLqHrNmykvWBt4nJabO8ibjw5XVAG1U9NIuIUdtDBlVnj60WYivw
Wi22AG1Uw60Hb9za6H47whggTPBVOBAIpOwCkfKd0W0A21kvp6xhwF5eftS9o+7QcXaWoqpVQ5oW
8OSL3z9fiae0OcbNUrwHI0Yl57HXXBmbPRUkvAYA1241DnhYweR1O9M7evR7xqTkek16mlJsdLzB
54afAVPlhnXYiCIp57HQasrEOt6irmaE8/rYBDB9OD0FOeVNThZj9NuDkPDqyYyYXL1FoqqSKQKr
doVzu/xTK+y2mnjPRLDzGKekJmxqmUN4UuMPjJj/3EaSL2C6DAGtAaEkUN6CWkEJKceOL/IozUHu
NtPrI/DovWtEqVWSRybNtnEQTqYQ+fgjz9QD2GJHmzapQWNQADNpPRU58m71B4G70qUn6SQ8ot7+
KikkhWaoEix/AKF1mkQNkseFwaRRljms7JN/AYX4oUHcSm87HHLgFLN0yStbhR+Grz+D54YqS00P
REVKEOPA6QE5aP0YVTjd76ryhU3nMOZetJLTx9v4g3jmt92UtPl2UIXlRv3w8I944gRhCS7lNs+a
lKOMZhW2irpPfVBEgkNBmvpXD3wFWKTYjjlA8QqB+1mqJmXY8GQcOXhn56N4WC76A5mpWAL338Nn
7AZYIq6AEptjhISQEXG+MmR+BP+esca7jZvjCauzyrkOSbMuRY5NhNV+Y9wUKS9el8NP3ubQxusC
tyud7k7BVdpkyKw7mflwCnt+PjsZmsuoAIMKfNfQgjEoRUEMaROtWjWWmPNRIDNdm2eT1lJciXnY
8+sdAz9O4aWMvpC7HVHd2qQhAAiLfOAhLGfN2Ekv+I0ofUAPwcTeHcuMhaUudexGZBTLHyjXMUlO
HowxqTqmoqggTT6cecw1YAmJrlg47q3DOxjg/UyFxuA5qsjLgzy1gDN5jTm6dhFIVi7ScruPOa1u
Ug5w2iU2rwSCb31GsZ0rEcrSfZP2UPyBo7e4CHDEH4fQmFHA4XS3LvRk4ItOc7elL0td+g2vTxI0
ATlV5tXnqDvMLwd3QxhiE4Y5r91EJCAkbkfuyoheFXy9hbVhj3HBFOXXT7HxTrjSQ0xo/6mO5bYR
H446CinjMkf94RFaIcwGkMJLrB18foqe2MoLKO8dNccuFjT28FhRhDLWHh/lx7prR0JLI5fntew9
3NYzI3fsHZ8JwuWXVw0tJQobIPZFx57gb79mdOQDGWW3PXUEwNyJ3//+NIRuwRJ4S1VdohrshtXK
zfrhdnkzwboGbpb3wnshah8uuC13yP+mpe/quzgWNayivK9CSaY8bGsYWIrgq8kg8xncYU3MJacR
jky8lU+tDkYTjjps+J51vClV1rZfSAn0cWaczxggwCWHJph+L5dmkne9kOkpP1kcgRbULllmz8qr
bTmSvZmKe12tahQ966zOwxFkAbtk+IxQJ7y1Jj8u8YVA1+uGF5awhfxvkCyJNaNe59wmOvPaIXRf
MLnd9lGH0lQmvejVlOxafO6EEArulOI6CKRlU2UpJ/k0Ub8tb9I/zW57SLKMCKqks1zPUdmr1I/q
+LjFFoiRILG6xDPw7tUwfav/rm/6GEY4uI5NH+NtIm23WDAC8FRW4Pwz7uFRuKU0SPVIFKJpSG4q
cmcjHzISHl/tqPcwA1fw3yqlDMMH7hyohAk87SoknJ0B+LHrXawRrX5kocKGbgqqaxkRefExBpsy
6sRFdGYbrB/EPFGeJYqHXq7a0aCjjhtImf066zbo83ns7WDd9KxPo9HYwts+4qEXECSmnwz2NkG0
m6sa1YLSk3Ke8EH5/y7p51B7JaJppHw1Njp8gr6BkvTrpVXwFMBkmhm1AQrTh4mdHq3nwuSkTUbs
91a3EH0rspRkdAx+1bUwlRhf5R4+IYTSKmJZxTn4V5YzVFh+N3/SFMKeAMjfe1tT4g8EJnsTNDaC
dIMhvEai0rbRTHXlf2xC7TbO5VZ5HlV78QHEJYgWghq3OJmNnlDDFi/FuRMGQGCX5SGYqT2G4Yzb
4jzXRkLjAOWH63UE6EEtZUck/oDiiuDbXNj9eIbxspK/x5oe1TFogz5gcSEzu/tNTf0DixjLGv1d
wbozh2ZZBlKDHynmeX+AQ8W94D27mRozgf19de63W4ArrPqmrwW7sGsCyhlG54cPKqcdakESx75J
BTNh0d+TnckHVxZa2ITjTjILKEjibMwc6xy3XGF8QzaW8Wx5TkUSv43fuxKGTNo/9HlkCORjmusj
ITkoRa+oIyifPUHZWZFFYeOX/4Gj3yLuyKGcLw2yO0BdAHEZHODI1y+ZB+0VUf1G0SK/5Z5wE/me
+zho+vhZ18LZQnryjbCLpg7OmeLDh3ypIRCHWFVlHmKrylKlf539PxC4E/X2XugQ8SCt0a8MCb+V
TdkzsA5ZiCrfRhR5V/0SWT8pyJn9tAvzZakvWNYTfdMoV7liKNlXU41H7m6WArsQJj/F6F9u8POA
wpjEDiWNFqqTVaM50Ee4+GzRsRXFofcXk6Hz5qdfSx+VOIcyNdd7zFfWXSvcJxHhcfG8xekUqywn
4JRMkzdwYSf0Yi1mk+N/mLu7dyemkFFCQed6Yfr/bPi7B4t6LP+oTHqmsVD7tQrCZGygaaRw1WQc
rBPK2uiHKL1QVeHd7QREH4WFhddHPHdUJN+0DJto1gQgiBB4yw/Ia1g3/XXoHb1C/zaL5aQBJKDA
mW666WdmPuxawJdb1nMxdcUPSwnoDmM2wHDYt8T3JqOfghkkPqHxbxeQcEZzhoUXjFaO/WyL78Ah
btFcKQJBIVP1KwKi+ZZcg4gqpWSHNo6Yaa5p55cgTSMq+j6ZWxDVR2cVmaTDLI3JjF90sxlKQ6vt
LRyNRmPq4Y2+nI5X22RXw4Cp4nOGFr4OKhL06ZCNDBzf9AMF9su47ityeuO9z7YG2a9aNewktlpE
HDecSHD2nJSmzQve2spJc5RgUBVgRDZ6oZxYHmicb2jj499YVB+1NIA2TXJWmURUqYOfVgOgVmJt
2lQmVGEjsjxCGQCeEIm826fCaAQGHZcdrY1f+Y7gl/V7gQ9mu4i5Zb9uECudZ6Lheu/IgeZSqtWb
KhvQyB+3i+W6zKleJtjZDniG5ThS35nnmDIB3dpZj6zlqP4sT8Yg1QQvi9/UCCYoB/k4dagdyB9D
v5HZC1M7cTzvqpmGQJDdsd3Z+/DpPCK1koMNL36Vffk1HnP2iWb2Oa3Xt2B52hAXD/fZVWiRM/Zv
CJ4+y8KwXOTlucguTNMMJtlYTJI4QmpMT/M5uFAcgeHc+VFHQagDqoNd4wQaE2XSMY9dRRZl65C0
1jwNxoaDpoT2X36MshVzWtHGEe7/Ap3YLHrtJO90YYW455SbDUoXN8PdqwXKNOJBIhUNz2LCFvP5
qKUVIbPDequezgEHfn6sR1N0cHIQ4jryT7VHO39Tg2Ws0FqoIDd5RA2nisyXOxAbtbi+BxmNA91W
QUlqzeUyNxZwrLRndt1EV3hlPJgXvSbpRYEeRj+W2qff8SiuWqLDDKEN+xAodsrAZUlKO9KiWcLt
r9A6fwgeshGYcu2lKgwMa/ciL9CrCBVn6ayYG4DMPfGFm+VzazrGu3nt2QUewpkfjLq5X7oO9Sga
GDVgkIw6RovZo+hbHy2Jn95OnQcbjuan/+ezY9fv2tjLwAzqGT0y4ANTB+TT0LNmkpw9zPOhadY2
4lnpqrwmvuyFWFYotGHrMgJO35o187qMX1Z5oB4xRhbGLt+EWhXL0EclNjZo4dKgksqQ+yKzM2TY
ZPOEhNrmfcpVmSj0a4gj2yy8+s2O0oXxfn5WgLMvz4I8Qu6/7FuUi42/pCztbPg/aCtlBjg74rFQ
wiewNQY8LCB1JmADGDxvsd99e43uNx0ixdA/IjvLr783Vmv8SEKvaT5lYejtWv6pE+RCNShva0ox
X0ngJ47wmUdGLwvafkGMRFpdMyZDjv3JmHpNrDRYqRjZ4gs/gzh0Up9NszgRl9kwYq2pDsZ6rWpG
DkYjwwyRYPPSah3xD8gT4b/uTvm5Mwm68JAjYX8feqwEctSxOMPIZvNKo1FnmARCrEA57YlVMXum
kWqNusq+MhbGXV6/2/sDc7Q1z8gFeutZLZ/xH5UNHjLd89HoxIRlPdgEDepa7Lpp6B+MML7pnMyA
cAASglgNSuqcKSLuGFGJ8ds/YfnA2h418cmXyaDBtSFATFuFQH4rUwiIWXFKYRT7ul3rDMabyhqC
8xYPu3GNWxxs7VdDlGzwfNqzQ91+iYIEIQg3VJv4DbDshy32PVjlbn1r38+7BbwLhMb6lHoem1sM
NoI5yWGuxHqxcNg7ePP9tUyMT+J/+eH0VMEyCSkQcFXDm89ZDC13syWy1PSUImdzOnKjTx1UHvVi
boCNW1i15Y2bIUF9VaYdkNZuoq+b+nfo6s7/ibBqvHCeRRVaQ/tLzshN9Q87DCzti7aRkAhd9LyX
9NK+a2OX/18U5TziKhEjbQrCVhbPeSAj5V7AUBLl1V+ChqRDl9WRyiXhUHbrE6VYESHAxnhhHKSp
4s1X7dzjvFAJqCP+2t9xUsie35kwgHH1zKKQylOc0areoY6h19cJovxO9jvm3gkIg0V3NLnTyeff
H+AeDLQcQ6bmybrbetY6CUhKPm8IvlwSCDjh9M8tSuLHyM2t6sNatQZYAfOCs6rDOdfsxVcapMdb
daecJvwcQapRvDLlF0zQOVDnHf8EsBmAds8uYaM081i4/7V/9PciOo+cqeFpKFwC5hpfOW9I+ePe
mdWgDT7CbtSCjjdqjqKKLuKstq/C2Seq0tkyVMxPqwHndlEF23eWfHt2f2uxI17Rhmhg0wl3F8KC
rWEIf36rE2YugVOIwdwH4J7baU5C1pg0gMRvNh4xm/IOP0/UvsdVP7WEpb8i9wxX6AJBDSb9ma5/
83BL5wOkFksy+7hCUpPHW97Y+B9R4/YARJDVa9N0jmMvfh0Gr+QEnE7gpIoznT3cRLW+58FNC+ZM
CaoNMMeDRWzQA57dhmMV9oPYPPoOKBReLKDd0tDY8aCgFdcTr0L90azeIfEQNAF5Ukm5Q+GVt/w7
OXuQ9tEcpMNLdrEcH+MU+jSsPLO9Q240zt+83ziP6FrsEKDHYgp7pXNiDLycQKGXgvAX7WZUDW8I
OWwPvLxhWTfTN7J3Yi5lNUaHqcui/kEoWLBiUGZ8jXlXVOhEfXwc4TzEJ0gxJF59HCg+neRl+KXf
PcY+9q6kc0lOAWVrlOy5+2NqGNbkFYFMhwBvV7cClF44QSrAjGKfc9EhmhBvDleJsGdiJjtVPJzd
Ks1mpIwAzTUh/wUAn1PQOOpeuWtWzEFiVsJh8bg6Yyvc4j44xf5Dyfx9w5pQoum66/YlaDq7skQg
VtU0tEohNfmamaGhIuHyi9LEZbSeKBF50PCndAlKKz5rrf/cXBTkXwhBpU7jEppdkzV6WWZn3yvr
O+ZI01EW92YTB58I2DnOZECmENtRhP5F/hi9hOrOzvidzqV1R0rotFZXOLOlVU2xD1rY4EHgwpfV
iTqbEzscrGh7MqKCnxQmZjQww6B8ZN7PIFvYaycowXRP2mELKb4Tk1yLS4I0wyeVFaZdLlC8DsP6
c27W1Ei1OGpEpzYxd2zK6CvqkLgfxSGmlKPu+wutbGreAw1p30BEvpOnCR0WK/0pyz9PBk3ZFeTB
K0nARk1gq69k8Rb93Ni6ZTdXtXwQyi8EPYuz1LhRt62CSPouTNkU/03r/S+OAW2DUYfsbANDojbw
slJVE14hkTeArLTE+1e2E7A5wcnYxkB/77qYmEYgro4wvLiVgQlcY2Cz1+rsJyl2u97Z1i7HhRP2
hhFbRkaAH1Xgljxn6MPzmUNNTiAsX+a+Tt97zR9EIf7D7PDxND8VzEp3xfxHbBEdnUAAmbPSXqBq
zCCX5eEu0khjuhtBBFmLcz0audbz/yzgV/js4cuDwV7x2ONSeHDz6obwMscapXvxMmyutq2t88y7
zuOVx49EeF2da3TCWtqWt9eYdNuLSNWppd08njoo5qgkd/ERYBH1CdV5DXprxVB04gUOo9/R/tVE
ojRDfwCE8tbqAgA9Z14QziZ86X9GXVTZGRdt5TpoH5gN3f/iubeEoo51k9ICfDIVPMwdE7rZrJX5
VjEurRtTp8iw9MQGl5VmByGCqp/un8blxERRhF2lhi3YZQ1MAL5/EtVJ9YtIhFegr3Jrk4LNOgiC
Ifaa7ren5r7CJAwfagwemqyDXaT9WG+LJ3u8ZF+Hxw/WQsIVEOD7ZGzcwkycZB75dZfPSXHfhDuv
RLZqjSDu8rssgDE4KfNrxWB8Wq3Xzjd59K8rv5MF6d7gtXnD/ConNja4kihrLwwANqtAYn4glPbQ
n1MaebZbK2w1okx59i0sDJT+30UbtFW2FSn8Obcj5/b4LmrRst8Rmb2cXJ6qVS/BsHHqsXSy8CFe
7yIVZY7XJenI++zg341q6t6sKdTTVB3tKJZfAxOOY+WOHQsZILv4QTlwwnWXLxWZKdQOpULOGdJr
UJo1GWIGZAYu3N1GuL1hvh0feWwrYyosxFF+yMznJ/4mhNXi4oCYVGsFdi31V3PjFT/8xYCCEBk3
MVIkvHmzTNoXdHqERq1fgMIDy0B/vbFVybyzPNNET7/6iJS1Z5+QfI/rJHR7My2qGufTjj1AKcQj
3ZjuP2vt/iOgBug9r91U1h1eTPEENRi98m1vUviNSZmscFiBb8EiOTv5VSdD5uMa3/dGkxia1IzK
HLpyinvG9yncdhdEZODYiSnfMDdfgQGbjdgxv3BqGxa9u2U42Kf+ymi9WkPTCVLWzKiWmPH76EFY
FYmlOLzOVRvS/2ik6dUab0VRjMz0gBgJkaANX7ADO/l0yv6hVcXx1pmNIQzX8OKwn8h3uyILeRCp
4P5HZBcCw++WCDDq8n5PjojVyYvzKokUGW28ENVL6MsJAGHdtVMHJWHTE2fRIppjV6EO6eaW/jyA
CUI74fRUPvOWFeIQhCgm/69oaPrigr/sxBy/X7coXOzMJjQtMIFODxd/2ZqMRqitttr/xVg2HENl
bMg7t8meq5gLOe9aL5N6exCZ0gb4jSSwLI/rKKm+YdlfoKwXx9xQxsuI8PrcuGQXmf7kDuiU8CE0
oKfR/NKOiKQlhvizYidB0ETzQqsqApv4odg2X/YvXHpKDDvpLkm9Nft/FNgoFSQzdfiMO9tOC76V
I975JtR9DeQaOo1vJJzzB5xAHQdRxr96ElF/TNX1vy2lUr8pEXL2zFc9EDSatT6IzPmdAHfijWlr
a1+99jKPbNQup8x9A8+6ADxugU2NNr5U6n62SO8atqy84TJzx/XnmQJxhww8rJ3tn36n6y4k6XIY
KJEI5wGVT50C+Fkcvzo0+hEGtDox1sBcuMpC4gGYeOSVkxcTFqvimBefrxzlK+egRkq3oS+RK8Ne
moKu22uNGc5Ksjr9eyeE58BzFGp5m+yAWCRqhxbJ+XLu+OiO6jzDR95ijkZihxfcMnYYQnWdaheC
xlGTOMQ/nw9BmNWEXdYCgLkL1ZipUP8a9eWqsnn9hJZJwr2noAR+Z63YJo7inf0oeFbLL94Giavv
xdces33hwKNaaERkEmVw3o5gB/iKLsM3zq8AtgFJOFBMBQPxQBfHxjbg5FEK3QMOf+7zvm9VzW9R
tTXzpoTs8oA9ydxIUFXwOvTEH8VjScXxg65xOjaH5cRQMi0AXKboIo8DtKqMzvDAAFFHDLOok6Sh
kgIFFY7AsaeXMBnK++OwLVNHsUSy0uPnaQJ2weI4KDpWQYoakDgCWPT0wwEoBplnaUyTGzh8EcjG
RAVYNbsWRLSmoGxEuobGl7li9AvtwcGu1i5Tjp+urtE60DQF4rJqzqzMCUK++bhS7lFY7YAPsAoB
Bj4uyyaDRJ2XzgkfzIfwzn4l94kSNXQ8/Y7k1UQ0eNzOajq+JCKlixSX8kinupDEM+c+JxlSZV6/
YhS3LgYX4Jv4p/ITyM8yPjbtqpRZcH0O85ZRnKGlF7JWXas/kOG1I2qaiYTTE1zvPEu/PQuNpUwj
6BBT9OguGgRZ5jYjAr09JUt9R+cHzymfqRPno4988v1gxZKsA7wt+iqyFBNTB4axy2MXpE1LEOnW
gFP9QcgBZwF9JZGLbdrH3Ip2QvMw07r3RMzZYHTjC7m/xB8/0fhlMQeFZeD71+3wFAOC2RG9LAnN
7AY75WDnHOvp0n2d5srVLEUK1CW/VDx/T69eMtZxC3ZqqaQQbfD0XPwEHsKmp9CgH3PPn/Khc5pY
CvUMI4wCh366YscBvmXkrK9EKS80gfDnSt4JoersxU2WlAy85t8A1ztaxnxWRnK/ncPx4Eaeb2ms
y0KZ3II3vY7yLRvfSUK9dRHGxny3g9R/y8rKlDmgcjo2uFu86Kw2ftHpY4Ot5o65v7TFIXKMQ/ag
fKOywQcdpMQi9yiYh7Byg86Es0FE2xbWrLKhy3IBd1khLjd4vAKCKnJ23yzji+g/bpymkzvaaHdl
ZxlO/mmBSo+GHlzSXrIUSzf5k0B3cqswTyvTcMRY3iWIp7HffhhiHIKad15NrsCYnHdtcBfihAzj
oChDSgjXj8+tB5FSh8WNDN62P19RRlNTILZ97K2c44mG/Bj34lJp9kQFD78lrYQGr7TL3LTegyjs
nhuKgdQyIJh8pEVcDAnNHrJS8CdbEW16r+G3AGdtdNNrDheFQlGuLlxvWAJIR4BH96JJWP/mgZnR
U8FK+KVALK6kHLEP0sAeg1czNaGtz96R1S3xj0KPcqo4tBKr7V7LUtbJ5105iLeVi7bUm2uQyp+3
75SX9RCtUuAwU9P2wnjt9W80W36frg+27O7kS07h3xzw6JyIC//Mc7ZiP+Y9Aheo7INvAeekYYVF
DhfZeDmMNblTQN8bYfleYBsGHwFvGMaTQFHkYgc1J+et0M454B3dc50FizEolWeOaJSd3766l8kT
vuK0AA+UgfSKVh1RHh74Kwzi5eLu81VILem0Ps5PpDyUQVw59lu8dQkPNr4LIJDdMRAX3uk+76BN
e4WR5TURtgBbiSWGMDPbf5y+wJwSBUKYY69MAotO6VYOKMZ7sF4DGhoamzLMSrA/fz0k6Jr4a4Qh
ri4RTRJlNfH7W/6CfO3Adb8CkkiVAFEfEt4uEZDfZ3nzc44+vmuqXgSbwEF/FLMwOxVUMKZkwqXJ
IKzPzXYjp8PuiKYhE8ZwWYO+tynjoVbXHd6ea09AKn8Kmze6RRUlepELv5V9L3da5wS+pZlGjigo
sEooGIP84BLoMkklBONqOykI9hb/IkKGceEdEOp4+rDn9DeNL50N/2DQ2NBojmVltYjTWvojIJ+c
0EJhS+DCYZ7k7UufjqsVIRi7r+wlbcMkBNxfF+btiH8m2EqPTpIu5Y1RmklGTPU19Kd/4jHZPrRb
/zi1vrxm0xq8gUAIPIVKjuuh5vH/DkDWFrpq26yo+5kGpW/VWS1+TsahWcQHs9C1xaWnQ82rYaXO
3+y+8gMUc2VticL3vScWUMJ1C/kX9k1YiTJ7fcsp8KvWCn9nn+I8uxIydJCpYm/wDMlt8GqrZjWn
60eVHLwA0cW1vrUM+BnySy1hlo7pYZZoxDssOT9PP1f7lHegrgavIkN3i05YmncaQW3tfVXRphY8
NEqfgaVXuFqcPM9R4AfF5a2rCC7iiFPQK0zB8fizOO2gd37coD3+euZL9wN+LesGcchGUpqHysAR
9byX2Air0OAbrcRgwqKgyQcmH0g4lZHDxagzrPfSKcSp1q9aRuiKkrPBULiB/UE4LX8Zv/JdTM4c
2hi/NQNv4odvEebQBZGVq8NRYjtVl8noQALxeNsJjY+mfFZyucbKFbAmqDsAWC4EV6gg3TQE5Mc3
ju8K1Ep6Tjl/ZOuru64WlaKs3wS94NiatRjRmvpNPEUbuuDml1DDaa4x49xps6PEhCH4kGTll+26
W76ztn3seYQ8ZskgD117NHBO+oamMut5Bdvn/Xb1qQrpExBocRwh0aCUiSbeel51KvnxHWxT+uAV
zGDG1YKggXhqPdkXlBBnDqoVANddZ4DEU33oD+fiwzp+wK8Embdd+s5/ZjKtFR5K7g1X/zzBpNv2
EcR0sn7taacp3Opj3fXgWf4MqLftKnLPcnAqZcrjEDq1TVjRsCVsl+J98KZMMB3BkGGqh4G942t+
dvUfB72z8FeoWBx87OtruehKEX65D+D5mlbXnY4dqJhlFPS0Ru+9gggWS0SSui7c2ePaabOYPLIO
59Y33r1u2mD0bA8D9zWEXJuvn7nfXQje/aJIlbHY1j/MoK1Vj0mbOQfcsqStW3QyEf5/rEpF0dEJ
yFZ2uFn8CfqL6UZmpymSFVDHMLXP8ISrps39gyxakpzgkqNculWYlRb8FVot2a74l6rUCSH3slaI
4QGcniKAZ1U2rKoh4jc/W3KaqyoaNsAS3e3/1ueVZflcFuuDLYBW4GO4aVmpqi473cc/QUWDor0B
DjKKvxJhAVg5otA0NVj+RLVbGLs/NE0KLbujJB7nm32XTC74a+HHxG0QKDMsZtuBw7g0oT7tRifm
u6e+B1wXEahPIqpeBOSevODGUJhpeWsfpbTlfY5ZO98Tf3Fdgn38HS+rVyxsFUtiyKloJooHHhNZ
G//8yz37rc/wogSmrHiBnPhnXeYEGG7xYI8VMQZ+NMTjqnO8pfvqxwOakeEdMLc0He78Gg7Emo1f
OZDGYyG4b3vt3tSoZRYgeCiTUqODD1kjy+IUiFPIMqG7kPysONZ46B+JjznH0rn6qU8BK8hGVR6q
7769C+n4brlvvFGq2SWtFL8/iMGH8RtU1PSLhrCEaMwoCCGIT8hGA2MQBkEy40VCD92fuoywNCmV
jg+UCd9miccekEiApfDp4cNCHAKWdQrhnlKesKUYPMo/QyAt9OO8HH2z2DEFt5P3YmMMDdL4o7D/
fGko4uLrKJEjjW6WtZIIk3+yqRFK8gKeW1hcm8NTrcwcoFgPgw4wN3REMqaITG70y1gf4XvAAlqY
lAXa4B4prC8i74QemLmoRSfZ/6x/GQFAMIEmWnrSxxQ6B9BDZ5C/GSDKyOS0y1TxZR5OV73EGEnm
6dPmB/P38VnRtApjJyQQgg08KoJOAuNSmtyAyC+dXA4nh3RQ22pn1MvV+L+r7cMAnq1i5kDoGgMb
k3IjH2YjW4fEzOFHOgpHFhPF+DL2EVQq2AXR3VpfkAxe7m64sQ1pCA344QoI5Q/R9jdLgmwc1x6c
oy30deTTSZXCI0PoveGxNlRAYOu8HegJJHTjRQeRXCasC3E3H3BIL77S6tgdxZIOVo84jv3Q4McX
vZyuBeWOtmaErUsbW8e7mzNI3k0/9hiZ+7tx4Fw6X6T5tDjmAaV1CSll3qOjiPSyptnyYRr4oBRf
ilPr3plM6LTe2/WGjhblMnsb/8SnNLKFWiTYXW9ookQfobaonAYJ8GlLzTKj/KGFKjv8bIXd/uZy
RQ1MqX+B29scL2ZduTxT+1Q9WUQoSKD14gHfxwIx3IhdtWtifrbs+URkvUzuriwJJnJ8w4zCC69s
SWcBjRyeQhFYfHWjPmZq0sJXtkOi7lRJEDmDKZ0eQ4WSYWr/d6q6v687tsENEy7zbrqS4nVLb6mU
e78i70qwg3fumhb3eFfw7FGULoKtb5IPFDaZ1kS6EZ4cS0zlmjkXpB8Bd6n74mRroEm8YvgRNbMT
7wcBxPViqfcwOSlG099Cu0dO0e46xpkwX+Vw0F5QvAdhB7PqWCkAThmrsVcqQ4CmAQss+tCKT/wk
shcLeAl4ktH1dGBWTCwIyyjPfkOysK+fUNhXD+bE6d8veSHVqPgJJbN5j0SoyZWWjo8AqjgnCWLz
iiK8iyTooxj7xvX3H38W4Wx4N3d3CsnWmQFR10S0lUT1ex63Haw0FhNrYfyvH7kWzQTutwI4n6jh
c7/Ghn4qFtMNBxrGU2ZpHd3ZT+fMSr7oYB4Oo/WDrKzzLvq0y+eLhvzMMfNJpzs9wPkPqvghdh/Z
WDG43qqc/uhD/yGqGytbec5pNuXkiGVo95cDNVJFtVJ3BqHegIdXOk+/NUZmOsRHjjedX7A2IcKU
JwUgf6EKc5oo81NDMf8v8/VTvPPWu6+ixSy2ZDMw4JxCaP6dTuJBrqVfmhGQgD//l0w1VKQMqdJG
urwGD/et/2hH4jp2LkbYnw/yLGOjzYEOSy+fecCk1taNwB8/iKHMdpJtkXt8QoKNp52GqjCjoIvA
lvX0gy0yW5P+PFsuRRYvz/yz6flrFW1Y2uUGVBCjUUy+19t9dwA4QeuodvjEMf+UwGKVcfk+DiS9
OJ5AFxGIjZePBH1Ykoo5guLqUyc6+RyMM3zWT5kwvemBfxjt6cL5hE5HItZA0wBsWiKfcNp72iRx
6r6ixQheTp9T9kawUIu6H5jfCoaJLDMuF91/1Uvr8znd2P+bLEJdZGDYk3zsn6D6PpilqzgfjgRp
VvzNSorj8Br3v6Jc1NDrVSSA1dYY0bP1C5WGhSD/eUcokuf3ehUk9N9akS8bl0V+M/wOydoSnr00
5R9su6KuGTWBIUNqLQau12yidpB4NlCXuh9o3rTmiSIlAhxONVK1Dua2qnUuiowaaSFlBhrzLOz2
dqVLMurJ9QSZpc+pr9pSrKJYjgRXoz7IFBJxJTq3PBH66KHg1B46w09PpSHuDP/J+Hu0i+hzkxVU
kajGa2lCwZspGb9AF9mbbFMWz759J8jaKNYsXAMbhwMpBrQZIz2QHlQGHdiyAiWvL+hv/jVZQRDM
AuglTPbDZy3LpWZQzKXyqIlOTk80ZVOm4OwhhSdlfVhoWwVDN79t46iu7HUyURodY/M3/yzL6zyi
NZnL++R5Y5ZpHRRE/H/yDQkqJMeaAf3E4HEpJwWSAjMUPoqGOyEcHyQPSEoZdNhzWjjhEiMiyEWn
SAaqHHJYJdzVSrGfpHz2/r1+11BkZEMR7kc6JodRiq8nZq1I1GLlhV+E8r4RaU8Q1GX5YUcH0bMy
xJMmaeCuiOVbR3+ONuom1uqwXduECH5rH0qYYN5NsPeNQds1YqDtvXsD4ukuxY1GIk/eBz90FYTk
mN6V4+36Y1Pb7R+6sCOOp4LHqad1mcOOS+OhcDRZ/k61ppCow7pYy2v6K7FfLQdliAAqLwzIuzkP
HxZyP8aa+pGioF3OkRchG/Tveu20xxDJ7eAlKfr//gWL5srtP5VMJ3FoGzvKG82sViUfhyGhSTWb
2JbLQ17DcUSyHqfEj+Y5SdhDvyNMiGZqsNhQUi4f0qGfKKluuJTUatILdORg/Uhwt2GnW3oQZ28u
J7zQsc07Tc722sfJkFA1cd89zZGikuu3VXWYkH1vLGzqBzbJs2XW0jcaxDBHpPfKrHAobOVr8o5l
HJoRXxDtP3/+Uwj7piyjT3VkWawGkremwBTvmRzrDexJvRgOl9o8oPrhSs6eqKHr0/PgwrWeaCGL
YWVBIP61931tk4aqd36Qj+oJm6EBsr7Q9mHNx5RpctrZ9o70aVHcIDQ7wyj76bsQBV6oGfvcA2hL
DnGrWwMDarvjB3RlvVDZHxkN2tLyeC63vnaKnuM+Oc755aNPdKlsC/V3g3nlgdtu6Y/XtLPwnVud
ZRbtvFxxW0c/TwOUxseJpLshmVTpY/voz+E1KBAgYnJ00Y2GHA9g1nRNyYJWXhvp0oB2y2Hu+UPa
Jop+hprlN0YkakhBOpryWHBQMQsCNc5hOjcz/oCPe+9u++F7FDYi9OwT9LErhcQq1gTRWrQZhNXg
p/hNUo56pPGPBX0DXE3Y1+X9SckXxuti2L+1nemYTIBI4BEzrP972q4pqvZM5v9kW/ESHor9cDIP
pXIU4hM6T/i7P9rVNFsXUOb2OAVYHhEw2uYBBUyXYP78jSgwWFOTJTzvNQJ2c40HmG7BaLboHjfx
mQJif5HsBMOBSxLJsmrpWH4YaM9v4KilL0VTX4WoBy6xZvx1V/f7S3oHHw8fL7jQuX8haw6X4iik
B+pwUt9ybN5PmdVHgEAwmGwDFCDYde88huYs7FXaARgKTzmmLxdumraMNsWFMNj/QmYB31mfoIJO
7jWNQphtK1J7uaeNpwty94lVnQDNSDsiJKd8kO49sVxDa4BCyy6NUS/+XzL79ydDT+T5oB9YIpxc
/23FZ5aEvSNFI9/G3Ygev9xd51gkWesgzK0A0KIQQsykFsdSorntIjuu0i7eZMBWtle/wTE5sTRI
vn9rE8RhvFIpMY2g6FDI+xZ5ETKvjD8yYBCCqqrKTRSXKALcTsGsaGBbTBl3kRMzKXBVzKY69mDw
w1u9yyH9BkdIJ2f74A0Yvjev2ghcOtBnt2EKdM8lnx+3n9FSfBnaY3Qf4vjxrHEPfSubf7UTaD5K
kkD/lIo0u+zGlzds5sFy2mLIaEu0KAIxe4Tes9Ckpq0aPKOLrvR2twzPlQH2RB/JLz++A9bajLaE
FXCLu9CD5Y0WJXu52Ps6VoF25K7RPjL2AlF5xQSMIbuggZ/gxX01bey7DDejgwOzxzgoZ7gSLu9P
jnBVuWzzxvNjeJVLXwhoWrTY+HshX/2cj+vDk+CqToq1IksQzihnH0WMynkoWHGRbA0CF6Aa0QCZ
1j7JJNlUNfcZwiuGhFUbC+u+q2+k9Df8ZviRzVkW8rhD3MpYO3TQtYU1iTOMe6OEaL5/tsCxkBw/
P0mSjSE8lodkXlkV4Okoma03BXcaiENs1q1JC+4Ek6VU5FUxytoBGJRoCnfgg0Nb/PnTJl9dJLl4
fAsEDEYY0ZgcLq56QuB7ecjN3jXb5QQ/nKwJ9e6ruD0+mVAlebi8XI6FjM+OdO8pPl3WVCxcoU0L
/hsHWqPRxisi/4mEjz7dm8FlgVdREF8dAw0lmERm9WCMjHMRLrXsxdA5cMruL+h6/Xily3Z2VvTp
ZqAxQ24mW4aN8hC8j/CwAVndBwulxiZRdgrxgDGm2MgN4775QKD6t8DFf+ickUk0sJ4wymJ4Xdhg
wa69TMkwMR4dsCrbjx9dp7EOqtKzhA4/Y3qs1dCKjsa1XW3mDip82Ag6FmWIPlaGk6yr+1J6mIVg
cGL0Fn8UGwVbk80QLlskptL4rtCFX6XWSxSAEJ6B10cRjI5e8xbBHJaJ4soIaofYSmkUDhbNf+dA
7BuylIxJI6OXYfCMHD5AMw06mL/V9raApnbK5jR2N0TDq6sBCVSO/dKQWYotbIrbh0skfPaotv6I
BmPl1N0eLJqf+Z74xGGRgfBQJOcjTUcKnZWg2xyAhB7Cv8zkgvDkw1p9ZcM5vIUxnA5ERIR0LFiN
5JK4pZkijaYqx0Eq10QuHtc+2mJUwgBVB62/12cOyq4JCe8ZG6zQd8vXLk/CMG6Z1cfJcZxxe/7b
nYKh0zPKGXYUYYcaBGJsk7vma+cz9YnoCp3eolDVVnQPL3hZPoA4plmNvIZAVAe9+CaswkF+zAsa
N9EnY+XOnUxcxxxzh3tUlpNidVwCY+ANU3fIUFAL3m/LX9GWst4Z1ehro4hf8S3zHOQhFEbn036D
Mh2WthB7trQ/QkQeeTxdrX5JmpLzSDMu0PnWZKoiTkZjh074yEsnUUfafB1V1Rq7xJ7TKE5zRJBP
amB7jasGtndni2MhgYNJoH+6R4mvnzVs/1VEVT01tZBY1qz4rWoQmef0Ifz8RxLY4wZJIPliQa+/
GwP6d/+oIUQ320xjUYKn+exFcNlx3RnhlQe7qut2MwkHZinQxNhAGNFiW/HdnILB9lkZDXgrGhb8
R9GJ0i0d09f3g45D6zIGYqO2fuoU6bq0JdkXl6zKBOakGJCK8g6TlluhAFTBfz+dvKzwLg7ZMRsP
tKTc6Q6kse1+d24gqOksx6piaFIzCvSPT5qaQ3g0HyQaOCAja/KDPosZ9qp99VYepA/BBU56h9sh
p/dyCpD2oFWKXKwZExPwBwllMWHIavkSs/yIpxd/hwQF5WnBNPKCYCxdeKDJF1O8x7oapbazeII7
bi/92J0zCVYghVj3MdBwrA1JXXgQL8LtIx3rE70r9YIVvT/dHBiSZVpCLyTKUEnS0tD93zHIZq4C
wzIXiIM7jNWADAuCqyn6J1QUi0f4Q+rocPasJQ8PGazCHZl5xCG6AGWY1+eu8qsv+JI2wqTkIIwW
8RsEYE9Bb4iG1aiiBwwiTNRCI77EZKfSVg2cowoU2uwgtwCMAzrSy8Jv2oiDHxPyPnkMwFS/Hpa5
UBuYngxdGGGH3Xx7cnZPslp40P8X5lBrZwbLoe5l5PiLcGngPMqiL/dVZZkBEWLnvaXgSYQsuGm/
oJQV1Ux8ZLwXu3Prh3+XTukDwHkyOBFNddScBm1fJmFTM5jj7Fb08DGPt9u5Cp2t77J/5wOnM0fu
DebtDC3ubVoTpCYuX0nXgM4an87ccDHujeFjHfxVR3NWHy3w/dF+Ho39CO1eSPbEW3HoBLYT2lBb
jVcwb1vdRBY182Ey0eEAtebIJe7n3ZdQ8A/bULr1q8zJ/ZJn+yRchceamSumJlR0iJAXRgI0Udsh
reKErT+IZjcwWAqFMuX6c3cnhFJcn9KmJsGq9a56TkDNUVqnzBT8OQqcjjKwJLqcR3+zWOnhGOlT
tKJ9gUjnisTwPg611dmigRDyZf5XdGKiUV5W/va70yt7/LRavY09DLW01AQ99QjHTKtuSj6+g+7Q
FOOonxmvHYBHtkNkpJaT4cDpwVmZkEswgrda2yVYYSsaRBZygDBsB5Va+lhTV3UGuE8KaZ1M7aeV
rZMYMVUqXWX14kYpFpN4ywej2REqSl1V/LQznsUByTYzgH6NtEeFjhGSPXA91D3r3f2gkXTkLY2e
4IqwGfo+6p+9+5ELGPsJ/7QHXK4CLoTTKiY1D2WvvdyPmd5fjtRpTFkzBpLMA+MlPV03m6XW0xXu
RGeThx8GQ2mYU8z6us1diFTcWtEEQkNbwhUfldx3AnfyUXVgeUE/77m8PfkudlIzgxME7cbmQbrz
EF6xfbir/KtfGo5biIkM1F5OVu8Dbi0Y+CakRpp/P794efOUz5ya9QUCkmwCt+PtJmSqMbj0hHfT
j9dVqsrz0AQEKQPNM/BaNgLR7KI118FAlzyq7RwHTocpbhovMSs/LXW584tubkMfmcJjNJoPTMJw
EzanEB3E4f+n29ycHjRf5DiopufCF2PX7EV2fFj5w7e8ybC4kQ11aBAM1pGcnKjm4EUPFrvo6hT4
Se8Xe6tCq0LqeLLkns6Ul7rhj6GvQKnu3AqPkENplR6K49hqtB5AGtTrqx/1+b1akjPZGkd137ms
lZBdIe5gjySBHE8LMddI/JUbt97rpCPMNZPRy3DY1ubart7TjE6tYHL9XaGEQyICXRROzbesDeIG
Yb9DtX8PTAGK6JeTp+euXgM58sfs1vWxUWjs0xrZ48qcjuxe78qy52DW8aJZbu6+ck6PZkS2NgIS
sKsFnvOxSFMuZJtCtZByqTEkY+hRrMNdXYzw3chVrmhkPEjSsTpR3XZWUu0RjElksQDwRJf02ocA
zKHHy/sJxMilwDI6m/8suIjqXZbbd1YxlsCiHlsHAUZ/D7ksg6hSwGQhlJ3WsJaCRf+KUZoxsrMX
4Ei4lPxb00Ak9O+DDK96uyff+kult5FDugDLPSYcl/4eQHB+rE8TDhO0jJCNSKAtZcyt/Thd2UPi
auYLSE1WYnSK7ynsxysY/Qe5j8o2zPDEW1jrYXyGYojSw+ZiJ+7+wXxUVJPvTiSjfuCO9z5BGamu
chu441xoIls9y8+SpOIRRPv6Jlx+lBV/ymmDR85H8zmBkmd1zfzcNKHz5Y9ZQVHnQOf/r0ZlSX3Q
xTYpudzMd5Hu55sx8bA8J1qHH5Mj+iiolkW1ZzjEkZeQhFf0ZFLxuLtcp+vDDn0vIh3LmxkwBM4x
Y2fOfY7iNjglSOyEfJc2vHlc3LTvxkcng8dCrIntSPVSbXQK8TSax89NBLE3P5EtnY8LXYKOf+MY
I48Y+bj0m5rmJ74k1PK4icGJFgMy9rCQj1I5RwQb1ximiwqzA7VRPC754R0iF3Si8iE3kI8U/tmG
Rr4Y1L3PS7oFLrx90roBCobrae43dHaAh+eyrexPcj2ZWYQtJKscWNeNFFlT4NX3vXuMmu+cYC+7
/xu8Kt69thGUZrxjAiiUTqSv0+QztmMFcfHngItJEwmeAFjwtrilYYP/3sCaqN3Ri9gSC07LAyNX
ILkTpp8cpxTD/mmHt2fHeYp81yCxbTkkABG+sC/gRD6BvqB/vRSq900V8Q5JTbh+4A6xhQzvvsCE
cRojGV1TBoqeDn115s4/cEdc1vx93qCWCilO6chFjtuAMbkuq7gLDrYbfOkX4fUtVb27p0LasmQN
3EtxSlJzxOMJ+jVIuQcpTGufKBU2VG6ut8g/+wXM3jCnDeEPzZgYNPY89H+UjLzyglhTisi4DsVj
kbh790Q6C9HkbLIxpF7QH4SlwI4Fkk+Rm7FoqrvWxxHEN6bJVnbHBoB3LhVusTyqrZbO2Oh6XKUA
qaSLq/Xs8GX5RSKQ/RtAEEXj7c1el7/LPJX9Xk5g0y6kOOJwyriHfFPODajSdcwfAMR8nAHewr1a
XswYjLZWSLbsLEJ4ZGzFy7NixMAQG7fNcVlz99o2ePrKrFwl7mJeAH4LtqDM1S8d4xT/tzXptKDf
X0/0m7tU3Sj0nK9awZM3RXS6gNJje2CO37CmxXp6kl2Ot87PxzXcIIdg9Cx7tcuAMKfnqzH9+QJV
jY0TfkrBFJGX9IFV6QcR971mnUyEz0tECNTzLGHXUe0VZic9r+AUD3xK2QyF8FNJAtvJVuWM7dGc
hXxdi/2RPLSNegkbdzc4otVHyEAS9GBVYVbWZDAlEjT4i4UN1Y+1oOwk7Eyu5UwtsY4V6eAD+ezb
FO3fDmKFVqyrUXLcwpxWff5lbEC5aACUosAW0W9ClRcx67r/dhvpuA0oo2qYNduJfAdD2ok72sxX
acBdak5ABNOC4S6JMbjuqRWoKQMY2v9mLv5x5LIQOz9siEg/SYtp/Hu1vzJKz905vM5NYU7Mzq0Z
dnSF+iVaX6eIfx5eyKi7LGNA98kKcMZrFA2z1RYRnrjSDaBx6r6uHW6bYDQmk1qO2Y7mv7pkxmoF
mAfOqr/tMYAJDHPsqHVamsJ0nlp2eJAx2eHL1uz+uMGM5KqoTvihSCJuAVfsZlBzNV8PP6OXTcI6
gkSwsGnwS5pckgj90kBjDMlSLtAWtPiiWrYgc99j9v0E9qoFsF6n4leE08Dx60S6t3n53UJDpfjz
NBUkRZaB1KOD0r6IFZmSYGEH/3L4YJUSQGj9zq5+h1eEfngV6f2kZp1XbS7e4FTLZ/T1Vd7eFoDW
sQ81aedDWZ7mzWRDCz8JxNtQtD2NfZKgPVRjBODSYjeSYVMFmBgnjjMV+Frw6Awhc5LG8gzGOsn9
cnTbpbgO56Ji2BuvyUaJSZlWNngoMH8JPZOt3RqJrGbSyE0Jp/ah+SKr/Mg7qpIRoqgTnRNmwPfk
QEUYhxbYAuwP+E4aVLlhLKDPKgwUEt18gOC++DKpZQUFXsKBv/C3OxaUBIMQ6o6q1mvbn/Kh5O71
Xb6yTKoNcl4GhTXRgWRtw8/zlxsFXXB0VFeLv6GzeRH9UHs9Zqx7+6Opf+BMmVkkKBUWhJFys+Vp
VA+wY6WqrTZc5it7eJqLC/ab+v96IuORTwvhloc/EqGksR2fPFj6RuDU1RpGiGBahnNcaoAmEKlO
oSAsqb24elkVnwebW6bgxoUVG6X84UXx/ddZL3zkbLzUdTWw5mtUJ5nnvqRbrOtAP+qCqSrfeX07
46JRxvSI30vWWiY2krMDe0nmCDWsvC7rTifwOqYBNJldfMN7Oh48pgwvWszDkiGKFyHll8CtmgaX
LCgGzllgb2kudnvCCbnWfqbrop5eyKVfF203aNIwpUUAikCpInTl+F3SLgcaBxKHDKDsc9QsFWm3
Y3pMtN6MZ+7BR9ag1lhuzyrR4BOGo0C5Bkaa+1ZjbRUgsqfdnty8TU+T+Q4ke5j2w5QXcgnnbaql
gtb/hTARtT15doEvQ9dIeEYnsNIGzBp9JsAeQqawkza1KWLpTfBBMc2Cwsiqo00fm1RYfyLK+pfg
n1zVw9TLD3e1dzMsRM0eGCXnkXh0H9ovOwPY4eviz1Nxg4sObCdluk4WPhg2Ii4vrAG+M+SfgsEw
DN5MYUTuuOaXZjInhGwIEWL7VmvMWrElccn1Fp/7AvU9kvw7kHwZijOp9ifz8er5yAl6Y7tIyKUA
GDR+3YWSGbpEL4EH7b1REajdH+CB54evPHNscqHOSHyILsj3UPxZTH9FoNP9it0yTfM0+h3TJZoW
cY11jhCezhzvoTqbSnqmq7SQP0249Hvk72c8k4XaLeHGPqC+aCHlzIYCHA6QVDCKu19EPvl3dfk7
zqqhkuCOWcB3l/NbSgkc3Yl2LU9PjKUNKHhiZadFCG1uMu9ndE5P+HBhNDZ42fdiiNNGuWAtpV7b
Fa8Phw/r4/hdPa5Vc7OEqej1PH8md6TvGPNA/LeZVsAWuNmn+FjlRfzogAxWEvp+/kRcCFIOyyRh
URLSkNe7FLeSaBoxcvePtN2AdJ+k1M02XZ2cvB5RI/LMzo3Q71nVfNtOi0IBcmqdGVIlVRiMuHSN
XeCQHLVJgGOJIuKqwgrJTmFhZVM2ZDgmW1JDOheOgIKY9+PY4CZyeg/NgxqlKL5FvdDYzOEzQDUx
4oPJGJtN414EQ/tuR2iqert7wsWQpVn3968xba3OpKT4BWn8Dh/XiVMd7hObP2/NWXayyTkWEXQb
uZnWYZcsmV4Hpa8VXUVix6R7zYeLT+XQCh8TjRLzeVDm55fL9YfkUAThnSag9TK0DyCmeSBXozFv
HnP0fOVgWP94iIpWJGvev9y4omzAjjgWKWyZHYb2swSYvKOa0gOF1JsW7dUuq4RX7ev/ojKyePyd
eNDt62OKgTDfv0p/ep2XnmSI1c0kmtVLJ84liVsqfkltlsE1Jbgp/dlcWhjaJ7mMUutqSDkUAEbg
2OCrkH3DZt7Pv5of6E6kfE0z9Iri3ec3Mw5ZJdJVIlohovEjk3hfOEiCfSEooxnx8ywIRHEkeq+o
1HCgZ7i6JrIJKjd536JNLSPbvDt+uBFSm7PV0P5SZbNE1lWJRMFB6VGAuwYcRp7rliTrZ5KPFQsM
e75IZPVj6WS95fBspZY/kk3mAFVZ/E3wJgvxKim0HPgLmwKA2tO7JjvU4vx+7U0VxwuQ2uWD0Ir6
Yo9L0BhpWL+oQoUF0AXsbGA9V4oM96sQH+SkNT8Dxzv08HfbwB5cw6Wie/4mZY6tyzaPO6LQDf9J
AG72h84E0fhuyVf+ZbqKYxTPvdI5qMeU+Jn0c4oM6TaFfANnzvh8ALrhfSum+bMfMsCaHkYlH5HQ
CZ64p77KCJE8LXXwxVjAICdmWrS+3hdiNepAhDvLIGJ29PMNtGHOR1B0mcr2HjOeH6f9M+HT6Udx
a8l/IJzO4bbDjtVlAxw3KJuDKOd+XtEpLk5nY34/q+EqKIq2bhDvAMfkHzqaNZ1xHQ/h/T3Uc8lO
fUYUvFN9Nm6B43kfmIgmm1uRQSMK98yf66PSudJxBU6vbNv/N+PPmCAEjNX/TvO3DZbdeNJzV4cx
ejYXm6GeOi2UYpPCFZM1zo+jJ1u/Xfvbl6OYa0PObd20maNTIl4lIaI95vX52XgTY40B35YY3Ipt
KReMM/YIuL5sUQU8oCLSXeb4RC1AvsV8W7RS8liQbAoL8vfa3bNM2RoUpcyRP+agvVt5x+z5BJ79
mCQuWlD+ok4cFQ6zllhDFUlumPpETre7A7AFt5YvOqYWa2QYoyArnkP6ISXg3vgRXJY4uyb8RvNL
Nyp8z4mErgOrvEU3A0GTAAfnG1ALmZc8xXF+UvK0uikSM8Sv3aWckp+uHvORjH2ZXgbD2cWvOAVY
JvB4mGJ6XjMpOpa9T4Z1xskD02Y7r8L+NTo3CF67bLjxZBQglzGLHYNE8WtAuCw/yLpWop1fjElA
tjWRVTczofUfSH3DWoCvZnsT5LKt4fJtEOWpCwcSlZSrhA2sRe6WtP4KOV6rUWAi+yjVdiPyWsi1
gMTJSlse2WvbsWjws+QPtUi14ClKSvSU7IVIPkwTToG5yeORpxiH/N4BDPgZPmNwuxuJ90G9Zu8L
29lc0mmgTVnAfL8snAhTR41WRurbBtpibdOet4AhAwZFZiQ4s2n10LCevrd5gUZ1HojEI1kZR6Fs
ILK0xHSc337OUwJHoMmjezDbLsc67+yhMH3o02eRCQZb0aGlW3n/1n8rIpGJLMF8eAvhmYez0BGd
d2Uek76k9sjBjbj/DMvGfbSfL4h/c8J+pnYatcKkuv+LryCcpMTqSjeHGJDjlssxB61a2nGE9yhe
H+R/h02KtuL1kljNBXCWOerx6G2iNJ+0WQ5/WtWb4V40YJmCoBN370+V/w6pF9ue4WcTal20Cn08
YGcvS3ct3ya1RH/ogBdefazYGyZazkyFQnPlctn2uhfQxus1taqLRsZVEvN4khJhtCdfWb1WO8RB
icEAD6hhjSzs9+4xyzccdKctslY02FhCJZ4FPkvNTEUcChkOxPLD3rLPafwZtqncyB85wz+HnAvW
r8Y6n4hynEfc3HJ2qQYCHaoX5s+ri3bRyWvslI1wfdbQOb8+4QEmO/WKEfOHzVVACLAgYTB27Wa7
gVPsn4bIvNuFbgMoIAM2RNrwvSUWOw/OP8cpnDK4zQP7UW3TkemkW1zBRtLc+MuFSLrL3SO0steN
BE5diFWADcof+Ob1luFdo+PStdStmU7BZBTrw7JP9yENXLtEV7vrO9xhYWu6ykwWgV9gATxL3Oct
RuGo7np5kKfj7uDb3/kaADgA6DNuELm/IU6PGCQV8CMDF9SDAlqQhUjZQgLCRT8D9fkEDMG1ZszB
/sQKa4jD9Lh3vBcCpiDo5VerYfwb+xDGfaOZTbLqIDX30Kf9ffNxfBe0VQC/440RX2qXd6VZST96
KQs/IpHJh5Kf8RU/Ss4yj6vZ8ui1AVrn4PhZp3DfyhHPpBooFUymdO1bfHR0AIgRYCkTY9XY5p66
u0Nh6oHEvKn8eW2W8v1+Ow4xIw4zEr3uXruGFKPGCv9COhpX3asrx8XyPR+xDVJ4K/pao8WJMpcf
foKwjxEhXLNQaO5+ZAq4PCff1gj1bz7VvYLCyidRl8pCPSAQJd3wtTN71yvcrV2AQnpQ9ya+mK0F
Ri9gkmFMA89Cl/XGlwvJsFhTiXy38zpdTXUFUhaenjI1s1Xxqq+scj3jjRQTBWkC/sJ/WZqX19D4
i+ppXIzG2mWzXNbDZD9Ca75VbIL3MrqFt2QXkwdeRWIiTrrmP5pLnN1nRxNzYJV9wtDNfTemTZwe
NIVdxOqBbF3cYNGW8BOpRfDjb6DCz9DxSWEh8k/VBcfbldFaJxxev3FVU4RELyXYfinFLIfITqoI
B2bxnw94nL4IxaGyacnJwS5Xv4HKa9ViN5gYPxeaw/37KEgrJvxbRz1hK8n6Uvnw6pzauCRd5tgB
Wng5dckHWPC2gfmpdk+FhPTMGFRnnZaqpPc1WJl2OogowKBGj8nsLXZj/8e55AwaoQE481uD1K6B
sH6OlCTJMCaK6EBuZ/yU5Wc92Kd3qRd9DmLLtI3RyKjQfrbYNrAaQLAGD7ju2HS55BdwErHMXtPC
iyQ9uWihdhq8phfTh2odLf7H9rxVMz9x+o926jCqestbSN4IYKqukpufg4otmG9qMRuPFdkUynaT
k9OarqAzFmwDR409Mp2GTcIS0dO3eAMtgiq/vVH99xJ20oTsoX5ruKfHcl4RahjUIIckZ5imy//Y
8HZ4w2kZL+1pKm631umfTByM5AL57kQRE3ymQYDCvBMj+NMOjZBQU0Allwzfjf75Tyleoi2e5JZ6
c9zKK2u1FQJNyRNzou/t6vVKOBUXj2ilAFohidPjwl+8MSIQFHfcJvUTvSQO7FEInnZPlX3awjbC
Mf7zu9V2hrjZo8kPF/h3uFfAfawvVUAU6uC98Fqp/Eul0NRmm14tnoDVzPiE3YVUkDzFZdeZC61V
4umX17sLRKde7SjKlRn5onRDyrKLAarjgTN9CyF6OAxvRk84HFK/MRVzfF5HfFsgpyVH8TWU9z2p
sk89us47X288+DozwT4S9IwAvoK3Rggez5X9U7j5UVSLJ70VsnEefX5c9TqNmttBO6xbf9PYBkDs
7Q+fcwEyQT606KzW64h+w5PY1sGsbmBd3Vw/oD7Nt1iEnDExig1e3+MkjglmlgsuyvXL7I8sdc1s
Q2gXYCMjXSDEWLaWcCLaIN8dQ2VX9gXjIdipU2kccNoe26J/8/NZgZf7m7/SlwSUvgqAdbBBYNiR
RjFBhJmetGnBbrpdU/lPTVrUKC4YngKatgRDM9aqudn91WGWM0LrpAqY8DoyatznO9HKsocQxDLb
q/EeHuC/Asx7f+izRfL2EQfKvaSEtAA5U5exwI9/KJKprs0np796831HkcZtOWNJLid6W2rZdKOg
PJfNjUo/jeUPpc4hxiqWZulyVoWH0IHOxBvJAYzqD0lirXR2qf84r5DjDVNj/ZD6/0AElWUkqv3D
SvRHSo+2stq16+S4rVYuTpL7F3bfajsnrixF2hWtmzScm29nCAVc3fYeIXqhH8SD/0FyHtcIDHnD
2J4OOEv88knaFplmiNa5OpfteYXq44f5mEQbJyulPGcRWFu/PAbxC9lGqWr9KvAQtQruP+K/IUOQ
A1NseE69Z3Sv7u/hK0KWqvfvL10mrTJZPq6bk/+9i0aX1XGkNbxEQVdTOZAXma6qaJFZ6UbQ1Hkd
qrVqroyOQZsH9cU7ovx8ZnIcLspZePdAL2kXFbtOOmUTHwip4/sJsr5jRfsF9lqcENFZOKaFSSH9
vXHm5td5cNMtc2fjQnf4GaEkZACJLTxuLQSrppBUBxTjNAzN1eCv4T3TybFIdmS35HtdVurkitud
w0batClSHYh9ETYW1VF/FwBQ/yovjsXZpesJXU9hMDTj4BciU941JeFaNFjpSnyvMxzMSIFM5VoK
xWQLa7MzzKJfdQYD35v3SQ9iXJRXs7TKGEoQlXsxTAitNAWDH6gd7Q2HVaIgS3qsy7lpEML4sT9B
VqFoa54L1HP2oivSuf2xkxMgEMYTbyOIIee/D3E86UMqGGxql248s/p6odf62gYuerqrdFPK0eWU
RvdwsRFVvwyV+EkBZ4bvusd0JV4bt2ekN9E6Q89eu+8r9+21Xe2qD+c0gmMXTm2aHAu54AFbPqOw
WLhN2icxbGfxH+ExWz70wkJt34H8lwFYAmj6galCxwWFjwa1dXlBBB20e8fDwSRcS3R4nk02v6pT
kHtFT5oLB92BZ/zc/v/N+ZCvtPeyg68bJ4Y6PIoNowA0s/4pYFLm/qB7azJyY3e7mMixVhWebkJe
q8saoOytY0TOS//6O8VNoSI5B0zXacKPx2dtJXacEqRMAJ5AvwmVBRLwYpwpoNblqIgseWzdccAF
C/Q5opcQfgKRTb7Hp5trrz+cXpQegzBQKzRtas9t8m/u12hzy8mdLL4NY+8IgV9n01EEnPFc17gF
4zOy6G87iwKky/UUmKKbSGG2ifFqNIU9qCBiquP2RBDMqIZr3q+aO23tUDTDjHs4gI0RKg60KCwe
7r/XgLXK7XMTpXy+2pBZ11Cis6Lg8OEh3cG29xKgcJlTJikhlo5F871cidCzrKfcElR1XOG9WgHe
opZyx3jmCsMlM2Klo5NE/jEDFZTzAUmWw4zHZ1+cxlVNmVT0Jst6YhtZbklAoHPnQ3w6bEv7s8zm
2C0M+v9hA+2ldemoC1JAm/IoHIU8Slhg6CdvPRed1x/FadczDyP6XGssCmWXaSAjsPE5uXrzQ84J
v9kdih0MbxEgkgX23Q2zHI3MDzMAsOQGvCdIWAIOleQqPL987TeLvuFfG2/vJL6R45RnEOQa+zTx
YB9EBInRtH8iaQNGUxnbFbFQKREALkqkctjJK+MKiTULG76RP1QiJhxaEgIDKG9Sa0CltdGjSPLi
a0QxgEI7g0BR+bjG+WCaJZgErJwJ/oRUtJmY+ueSfF1Vfc/ZAzGIfNdOxZMcViF5yY7ORoZYh02Q
R+CRWLOA7ABGgYGn+4UMpzZu6KI5sav1qpNjy3ehRagQVYkrlIXU4YQ4GQvd5/gV5bsLh/nEEzii
bD/BcrSk/Xtpx8PPlB95rIrsxNuLX/RvcTJwYuXEP6zIm6gYXyuZEktnBOjuRCA1zaY2kmjzpSWJ
IrkSV0cV+9+Umz1VTjxY1jyiLop8ZRAl2XYLcCnVtFKntusp6RepSPtDMwHuYD2BQaJoexxqM4c+
uu8fEBz3t/snn1JAWv57PMrt+6XgmxzOBemU/vwVpnJDsLVXJM1/DofIJ1Kn/VoNWgrFy4ReM+hS
efz3ogZ2ZiDxqpWm6FMWPjBPqavqcBy3OzNnOj66/zN53LiHBai2BAP5pS2NOvyYCHNQGUwETm15
UrnwR3FBJNOHUdEOWjvCC7dIDvUsmAN9KxIDn6RUkNhX+W9OfkGP3LQAEiRUD8aQzelXL1RZjBVd
BIe96NUs0f2bNGRaacxpfJLl4BRFQZvrIZPs0gZMg6DcsIpG49KTEgA0X+ShcRxBXmGzS5BAuSQy
ZeyoLCNrcIcx+LF2X3ImQXXhdRlXxBTuzuL8JuoO/CYliXSF74UrBJ74V7vXvZDOxO8h073rd0W3
g7c5yrw91lPkRBJK2+gQPoup0q+NyUTJ+3FPaRoNzb7VCNX5p99y4U9163X86LD3qsBkIYhL4h/V
ZD0L+TE7SY1w02jk7fZ6OzoOZignSfBuvhk6OgVurjEwH65omjRfuIE9YLbzD/PM3mtw2q/ZPFsr
yawTwzBIKkl+5gh1RWWybd5wHu0fvjiVmRScTbWG+ewYD3uUXQze0i/n/CLhoKvbL5O244absxtj
JDhTIw/Z3kcEd6fTDUZotRvwvvsS647xE99PzEhnfCwrVAtv8XwriJXlOOtTnp//nJbQjYOSswl0
2zTlIrHkUXxmuMYhePb17NVhDI+4CMbkgixgaZi8K5fy80SVOkngY4LwKLP/94okgZYT23bNqhfl
FZSiCmQVCM4Tx6S8Wpqmr5gr19bwkEYcChVe3UucDm/Yp/CXwtsJOaFCKvkED8lUQnF0IpYMZyhz
gqUwvu2C0eKWgonlSq4SAu4cFW2NCu/Z1j3m2n0ycLUjWneWKZB9ZtcmMN+6mmv/RUYnnMjuhlzY
ug11ZfXzcPE7FOj2jCi65FvWZ9cSw2IVr+T5hHmIo+h9MZAwcgGDH2IlkcjuUzfd5mNzKtbTsC7o
h2ep/tM3+tJ5qoss1boEPWWa/Ri/e4pcDdctFXAZgjt8MyCdrBe03wPvA1ZexISddfckyzeEuDkF
/mYSmaJqsyFyeWxubE5pSIIZHny6OkOtTUTpiu4T+lP35KbUkJB24FsodWpICB1+saWarx4dKBL/
FCa17X75mQIoAZZ8HjhzCNSUqRxo2vpoXlBD2ToRAJBzNxlvaKzSgcCK6IvKQOUCQJSKpa/g8hYC
GP0RGQFNFCQG1e0PfOapCZGzUVNrAI05M8mqbv7CQNtiN7efEWBKKttH89HveHbCAuQn0+HPxZFd
FI2uMze0anipZX6AkUrPBPZeQHSGB6XJZ1kP/nkIlNHMWNAc73o0fp1zfuc+wnU83Ig0AKCYLAHN
Ka+GA8ly+/gYFPlJM18/Etr2qLmjhnpLdd/2rPd2zdM7JRS9VU6BfvBdQyfPpd1rdXYPAPg4QoI1
KulxMpACwptX3jTK2LakbStxndn/1fBkDit197nK4GN+yEuQdhwIlz6mbH1brhU+wGjenB+26/HX
kdUA9Q2YkDKwd6uIU4pSSKBApCqBy024csCmS0BZ0qA+/LqfcJOKT28POPXNHDgRduICTuO3fIo0
ZIeMoQlVNkXXu7M37GRIBr1HyWdD8bWoArRjuPnLfKF4zbRoopN/qkOAiS4OMe463ynce9LXEcDz
pr7Hs1zNoYppAMxha5T+R8w4Fhg04IdrZzgiNpzoLrRRwmrqAwY5QYD6TL2WUvh4VGrLW54rHwMR
gvbP85OpDsk8u9N00K4+JcGprKOvzr0YL2t66W4Rf3riavqjR9EPPiNUAqBcbRcD6i9aymLr9s31
FBda4MtqR5OQogAvYU5DmHfdjYoUmU02esAII/10JIQXnplOETlXnA/4XemH013GoZI3NAthBt3o
4HiTEbEMls4UGo5Wnc9FUgHH+6gA4OyqiH4enhVqcSEBuxMDazXt4/z9rsC28sWgbZsUfeoJm932
R7BOOJh+Xc8OGrxYL2KS9hlzGsU9nr6BzEZNOMzZKy+uu5i2RfXP/78o8VKRo2V+kxRDo6ON3OTE
K4pEmPY7IOi/G6B7jAQUFfTCpbNTFsRtZWpUXti41ZbJbejA6LS0jaiXut3HZ0Cd4EQCx+u+i793
pkxAKRrO2QOfEplIML6bBZOYUWthgiDY+qJV+Drma4TsyYL6u7j8+K3bci7gB7qPeVziMouY+xtf
ub0bfNUFkScCqfG1DTeQxPLpvYWDXVsJt3tzB0sgAuDbBzy/VymQVbgfxkpwrXO7RCDNkOlU2o6U
ESYmQfO44YPWQz7I0wGI7rSg1Cc2t5QcxkytFAYiaRfSCZpRpz7z4PxkUaBTL8PIcdgymbAqi0D1
htZHGpj/oHfTl5U8u0RDzNIUx1G0syexwsAI18cEEkB89Zz0bq2Ypy560wMIkmwW4C82f1k4r9vm
sLiU7KlOjB+Q3Q+e5aflr4qvd+j/covlysHZlFSwnNA6hkJkj0JmoCmIBkVvOwQJXIQxb2Zi915r
q0jdMQNiuRphmXqOSFBOFPdl0SJHjuGKgn7nzcGTq9fx3M6pOvaVJmcLiXH1Q5vq/67RsxL00G83
z75I5CJe5baOaCbI5XEs1zHnCQcldIq3KyNtmV1ATodaMlRS9kepG9VeUKg0Yw8MDrjkQmEHUong
KNkZelSIzIpnZ2CEAWG5qFNVqsN70ftvszZRYZgMvNJ+68CYX1QeEIDRzxnFHW/r+2JcWD55i5fF
FpbBE9pSOOfnufJjfMr/645MagBhNMDpUgvMEkgBE1Dk96JSKBhvnTyfDSZycj23pgBdsqnaQX5p
jfTazhbk4KX2Yvtm1RSJ3qJ0LSOlfQDHKXP9nxu2iwlVcNdwOs6eWoXhR01deWp0GDthp27SrAL3
ie+fIOHV35UgGjVqR5XdQM2VpagI8ZrC2C7OQeqYrEAegH83n/jGH+mCbrWgs06ipXJTEkWMNwBU
/IbQleg7BWQrvwjgA73qY12UhsQAe0sNW/WJjRTqYvHPJAsSB+lGDL1nGC6oaeX38pAfpLCQskIP
eCUnbBzP3Mxs0B+EfjLg+Rjc5xlWArsSRngsBwHbfeho3xP4/DID/Emvjsk4szT/huYmc6nQl6PE
RDRdH66OWILiwtBW3mbhsAch9sQUNO7B27hOPZBPD7An3WAeTvi7+bHWKQodcZeMK++wdKwzcG9S
N1YILqfB/zGb48IHIYAu7ZydrlFxSsboXtgjm2T3R0PsZ25r8a/T/ctfO9/s2rQwUb6crt77sIeO
UCBzYv6R9FZwMmzVJ77ASH3JvBgBVi2TpHlTSM48ord6UwGBtsk7Uj0EarmsQgGbh0BUfRT5ekVy
S0Agz5kGaY6Yi7Agr8I/DRt4vhVFZYlQFtwP/sWBNPPQUHrC8AJMzPvgIJei2i2mFFxnlnuOdfQA
M8h9BCoz6n9hNcBZkgrRaIaiHbSqlNWVXe+DcSqqkh+aDP9SNfF8EbqG2S5mAGkNF/dJuJfbcsJv
1ivP/zry7YsG7Ru0w3Y0AzDn5M5ECQAHjqhUZ3f+gs2Z/xWMe+TJpVuaf3g3r0IBhtJ/la5Jv8Fp
XgDS4JpJ5b9FbDs/rVMnHSRblxEbTZRB+AIaw6yWADn8A7STBx1iBqJAE5M6SPPxqoLBwjoP+1MM
6YSFEhx4twne0nXvDxwRhtr7jWw9GnAsCpO0mEnqwluUXYZKaysYk4aayB3oMWBENqtxVVBW+s0o
v7kzvIwMaB+HjA26dXLLFIr/evfO28KQBulDI3yQZMsynh3SCeVx4VMp7TVpP2a7gSNYRRX94WNy
plyMQvF8wb1yWoQXF9aftK9pEpAWOPEhIthxzGTho6ED5GlLmOyblx3zCCu4gqlVXulj7UsI1I29
sUjLpVgzAXceI8Se8yF0CP0x4p1pc4zRSYaSoCwL4behL8NqMtnImwcOBeDTd2qj2cpbAYMy6W8M
AWVftLoICY2NPcHC2+wNijP/jMPdzZoPjbeYhU0QPVFNjzhzffFn1CKsCxpQecFbATz0aAAns5nD
Vdg47pAR2G7fXp4eIThkgxoF+YgDTIH7lM9pQ991sfriGzX37B1ItaW6hX9oSydfV1yoL7zOPzPu
dXBR4ylRfhL0rfxLzAo2/B/RXDuewnynr9MDNNlYlvo7hsbrK7ibc3cwdeqOtTTubvg6aahlDSw5
y5fa9MR9XBuk4ETPA1mO/PIEr8S/uTOVpLujIursPPLpvYvYFl3WBDd3H0IDYCOV6/QwbEE+FbuP
8qCdlTf0/bqjxcJHKWtLKGa90+PoumkUCEA5rcv8erxgJEgFy8kQ6y+t0YPIMJj1AuGYH0/Y6zI9
RrKiokT8ig02ZOfbT8nf9SYwuJ5gKSk+r96HzlEebJf6OBsnAJo2igcYeTEGTBFst8eypZ61pCzh
n59Kp4vTxIIlW5q0pqg8fz1BgrV9fszr2Gqu28oWzoOFzhzsoU/JG5pNivZdq5A/BhgqywMe8SxI
4AAGx9ZLbmp7ZS+kai4/hvOPZces+WE/SFKyGDsXw3++8qhR+VYt0CeDt7uKyZwljcnjdIxTqrdX
wxsFHcnTPtYdKKx2g5ECtx7LColgOGoT4XGTzWsLfsdTr4nOkW4uqf556dTokGAOqnloPNAxaSEG
CeEXL2TBly/Dh2dEGK6WbdJnMvv5HgnNsKqEL3D1f4gSVmChtNhAGo+rZn8XHKEwbvpXzteeoxzv
MkwgUT7xvCQ3s1h48eWxwayDJgtfPLwf2YjonJiE5KJ/nlCy8tYX/sKiLY7+uiAe5mdS+3HDO00X
YVsd0uvIQFhgO9amuhFnpJMC4Wf8xDreA2AaAuiimDuHxNqVgmNKj3Tn5zUko4IaPVoYqLJs8Xa3
0bQ8LS2OdKzEIXSYPE3p4yyBGrGMSDSwrqG5TAWIi78mHzCQPoF0iVPAmnaX4jo7IvgCxBH13Iu0
yqjkZrQeZA1R59giqVntoLyb01X25S5IVfH6fiQpgXk16O8MQ5cSKBkCB0TWTHAfOoUbrEYtD81J
Pbt+X+/MW0G8KcFhI2oRcVx97/sVpCc3Fcyo9XHkuP+2nu1PEdUcGYp29hyc2Nh03aUP9n5SAAGl
lynbW6Ymtlt89DTTyYDhmAwafBZNgDf91hd/CgwSLCHkyUcYhgUlvzJ84EmoyfRSOZxJ1CrkqCpx
pAAZmwVcPnmJXYFafx96ie7HB8dXNEwGhBGlIsI+pUMULfeTBKMlOA10+blAZSJ5+JWd4tecjaHb
8H0T/RZ0sNqxHhgHqDvURWTUWB/zAzzcvVevGt8II5MkmO/RakMTGv0JL0Jf+DoFsvCpt5EFzq4/
YjAif4zPeWumHfJHdPW8ghmpAPBsb0lvoiMq6lrxbNqVfwN9HIXW1tW37WOkHgC3AbBw/r1T4R5Y
vDeejnA0Fe1wxl6a/1iaSaM68M2vukYubScGdSXHiHaocKG9D+nrZwiAfmFZSUdvgGKsvi2tmsyM
flvARVwOZyQ2Q9XV7ERPuO1Uh5IJPc/r87Dzy71cBcQSh7y4ZlZAM/jv92pqaTRaci49Xn1UIdUW
KlffsYowWa1bLCnpw0SJd85F7RsrWFfk02vqxEdN7JZhIDg3R/5soREo5EkaMr6nkauhcblFBqMY
63Ol1Mp0nL3MnO24m8PRmZU8oab60C2cpfvX9+xfLq5SszbdxN8LTDm9ZiORa8Ej/Qeqz0BpL7BA
zFkX5mt3X+w2QssIb3l9GEBNWyUOXQakvEoXarlbHNwqpOHQFjwTy2yKf69LBNTh+hPV2EYiccnU
6z/jo8mrntN5b0dti/Z5bFKapdOM/9/lNNTHDQXkfuzzxsFdyDJddK4sY65VGqzE+ME2UO1hS7Ru
huISwWQXuB76TYI5/20tg+/Hpw7khPbu5KxBAwP6rdhmH5iJjlzC167b1/0kPH6g77Mb1TMciQeP
gtqNce/ZMIUCuaGHrgJgeZkTkfy1iA+COHNwUTeZcvmWBsEcwg429xqzrNnC7+FpbbBLfqyxUw65
FoZMOYzIUqpfUHfDVA4mUaa6HIc6NEbnswCa1R+hsbgN/mY8QzFV/ccWUgT3Qfx2iXOoCojIXKc9
IQNR6Im3JjGF/vdL8OpMBMKnXGLA+NVeO9N2MDVyzc5px6CqMev0losujuW45BTZ5bXJ8Ng7zZh+
Ebz0LakGbMDg58dab8B7neh59ngOIJO6n9mJEm/J5inF3D/LuKNqNXHGsMcxQBs7rvObcBTQyjz8
jDkebGzlWrcmkYocihCvgEvNiEuZGsu0O3n6AUshFbLWxfMqb/Z7CnjzurBjdzWFuj35MOgFyvi8
26/6tWw/z4ZqLybKmQkDQwOXOxyQh384eqjaMy8pnOjXBw5oUeIbGebpBbYFYdaDI94KRQNUdDUt
ckmF4KHfKyxp7pqZ+mgrfGUsY6WxGYe7x45QMCbUcgsL+VfvmBFNUrarLxb6WMQdXwLH+OE8KnQu
4ZOwo+1GCbpUHdujtrwx5+8d+pvErryrDHyRg/9E3D0k+C/DRwuLOCnYCL8E4zZb4M5PeJ/Y5NXX
Pg67An/mCiPKeyqRdOyh3aYetFbS2m9AWWCy+obSQG+k+r/BCFAC9QzPYequHsHSob2XBUOfNVme
MdIhhxAOCbHBEHWw4+07YrHyn6rB9Dp1dP9k7lei/k5A+TIlVI/UbfAe8M4mog8NbaPMHe3ZYBzY
tgyJhN7WDLsKip6oDYJGYnPU+Ka6gHGb4An5KMXTm5yFlwPQ7gygbf1YPeuYEh1GdeoBcE+QgVnv
eb1qxDHvPbQ3td6FbEyylXQIwLbr0PJgfuSK8rQyJd4wOnv3bL1aCjRNmjyK40ah0DrFNQJSk+ZZ
VM/vQGPb2hlWpVfxSKEajfX3ox9y7Gm3hHYXEatTq/4fHyGzDQoBEMcFDMJjjRoLLWsq8FgCrKkp
CAti1UUOdmLVzp9V3MGPJfDwxAMCKOSnG4+xOJ67oZDuaf4tkOeTMwzx1jhalSwTll8jXzz2zhBA
rVKkGTrJl5K0beDEjXKBIPaPBMAt5KUb3qwIbmuYxSF2j37H8b8K46Bdyszuyi74vAoCAihOsTjC
p31dE8xvhUmQ4xLNls1sAkCmYcl5uAwjAdP0dLtwVR1uL52W/AU+lAVRvqDA3ojn3xZMtgwceQPp
G5sd/0/eCdAo8bKBE5wSO1Al7P6Yo0LLTUpF6PXC+0oThsjP8+YUp75Nyd7Q57Z0JzPy5he2Ju3d
o5OIzUMAB7H4rzzCXOg9nWh/6Z9aEqDJmZcKCYI9w+w86mgB8jAKHaYnrjE7iBvpv3jK5sUSZif8
2pTf9kzLMTnlaGCJ8VdK9QrKkpQApiwNdISfuN7SbX1q9/lZFp7cCufA4//UzibCzs7jZE3y863b
qEIZtrjlzl72Wf23MSCi6z0h8NLJBpJ1CivfXuEnZXaZ3A1I+YgM8fo72L3R14LtLbw8CV/y2kpA
ZvcDXBRs9xFfQ7ucuPuEKy9z6U9K+eYz5XLLUdfCcWCXSKo+ymGr5+exEga4YbXMNf8i4BPz5QnT
p5DbihY6qRaq8KTtksFYxkrEL+tlRTgkIJ8AlZlobO1IBgXvXtSdhdNQmgpWZeMzLo7tqKGONRHo
nVfXa62TKBXAo2nuN/E4OfIunckd1emlN8H3Pa71FIHPhIIZyuI2YL9nz6ir7S+CYNFHg8ZCwfKL
zJUb1lGW7yAFtSkeczW9WOTo5UlJYHPLasDMjztIrVhVGCNM3d7O4ghNYQ/CIMakqn9U6i58gSj5
/FBu+DVzzkyHt0D8UudPztfOjU90xlxZTkujI2SVoTeWfW5INwnfsj6CPcE4NuWKbZ28MlsenK0R
frry+WV1s9oMmbjd3WlckQHAa+ffY3gZxUcDFBAJoHKpMfs3zYGzmjGcyVGRswd36tcMK6y8LDp9
WjZiUpqLDhn0l++V1z+z/C4DUoo90mBIWME094fNl6ATTUu0Z1RN8pPhoZt6uice/hHNFdVMJKWH
LiQ7ao1JcNoFwzvCpI2NtBp4wdHF4jNEovOUdaHF9l8E3D0ZYZ+g/g2bSznwvXtzpkRilUuY9xHB
Rm9FMd2Gto5X5UuFi3SN5OIn7+lGZ1JeKRjgoG6r7azzOdpVfyfYhwr/XptHI+o/1AuSQrqTboJ0
6W0YuahlCeWzLTSCkAdYqLIIHeZsZHxKVFODqMJlR6/qXChjqmNqe6i5D1Ju+4oOgOz4VN/OJGyS
Y+0Td8P4zcN+YOXReWwJ7CdhiW1WF7S5qsUsfzTQj7p/Ee9VmY9RLF8Z2B4y6EdsnWM5nuiN6/cW
v3TI0CKvBBKJ5bReDxgoiyNrC1Hc6ELx5ppwmXZaaY8jbgksd662N4YPC03TfRxmqHrgql0vy489
YUAm0mfp1nySc6PlyH/oSekF2SklvHVdh/hWDVeLXtrIrUEsDLTuY/sos/GoUoW60RGUQDFAQuHc
svkGbq4YxnOFR98ToJwgWcq+TGHrwyhlccb//qYeJPEzV0ExVWCPmWbPTxJPN6axc03ct+aOErhw
IDcOxFmWn3CtsWzMmdSfaGkIb7tMFc0SGhUePemTPGvOublKUBKpXivjt7tj3Cf8DWCBTs647qyS
D1BBtEUnd6S7Cm/wfgTdpFjZ5kWDlB+V2urgiWvg20IU2fRQrhfgLyj2NxcXpA3xsUfWqy4O7NhV
KdEPYzFq5Az8c64XKPEYxMBV58A7iFqVmqtD99p4Q0DCQEC8f9JOgiikjQ+9hDD6YW6vrhd9i4HV
zCKHDz0jIGOb5qwdR+fFyClvwJZiOT9erwAo37R9D2uWhsGONAnbNN2gfGOyU0YbUr2a1qm2nv39
UJK2myUdSS38RZ/VWlxGFCy/DudHzOIV2HHZIdcogKILcoWQfAh63Zg/hJJoimXx74YhHdr0erbb
IQqAlALt0Bbx+IEadW2dVHuCwQORB0S6cnl8bVbfMaZOv/T+pfIoyrhc/qVRseE8aLid/MHcejT6
hybVH7lfXwjAa1NUWheLKyNIA0kFJhoT58srRdSJ/uNSsmlU9OwPapphAZ5XVrIHWBSFU/295ZLZ
j/b1uWv0hUN5dOl2K8aeriidEirwjF8w1w7C0QXyIK0140nEYX04Dk9FLfV67QhIHSrH3xSKFnaq
tvrRphkNqxbUmlYvjhS/BkERAxZOwF9F5I1SaOu+L3OynBMix20C4EHkZnorQOTSaTwlsMplwLlI
3MMM4ZPrOZc7lVTGIIAj9FNvhZ50v8XCdai9UzL/fd/sNDgsciYeQnIXibdP+C24yEQCxJ+yoLuR
fKZcyTnDqM6BN8qfNsYZ2Eh0MlRfqUxj6icN6ZHONfGRCRgWkXwixrR0EBqmLH4ZQc0ALaarJOCB
R73Bgvn73pWmlRf5YLCR/suXt+W5t16CxH2ju+YdS5+u/PvQ0D2h5JgHrSGmCf09IxgrSI1gNuvN
WPF/wzTNkdfnp5BzC0Um0Zzpzj88mzb+SxUNYF/rg+o4SLhCZYi8AzV4CKWRahhhJ1mAcA+wmL+9
qof+AyFobeL/u/qgBNbwdOHpvpyWWSvCUr5cg/MyUOpJtnlSEtPhO+nIjDN220Vp41EWGpwWWdMH
MOQ50KN7IzLH1jubowr6g6H2gVeqfBnplV/Yt8sact9k6VNb1olyA7GyBFuzzup+ucMBa+mHzGtA
PO0to5VCLRBVU1x5MmDv0+Au87R12M6zCkEVjTd5EZAfpkQ9utCHzd1Db6Epd67EuIeMXbdDRGy0
KYFWp8ukO+n/beCFxfWPvSJwHE69gvIrJFRjkEehYQBgBHjnbhD/LwFWXURv/AjzUj6YQOIoEAfU
fmj2GxOqSf2QF7YKddACC0+XpALqaWxEJcgn4OGH6IQ8hUnOBDsN63y4ZT7eyGhNOqLYRuB585Sj
Dtq5jbg72CWlwaTGCEkJ+bOfBPQqCpq1e3Q0bxvWvZm7FlHof3IroQUJ4lX74Y1sRyTF63MUey9n
JpbF6A0+L1eqAVMBOSvQgwrgo+97iydGm2WJNDN/HINN3dRznEc6C8kP8sT8oQOVzC7OGG0aU8L5
R7RYJ9ODsmzAMImJr7r+1NYJL1xpJYf4h1RCI1OV2Y0kj/M1t5GX1NaGvTzzNMlNrXq0c+Fijynd
goQRGSoxiqVSVO8wNJ9KoEBUSOgklgmHX+Zl8h2Mq39GVA8Lp7TsvEzI3USgN0IDhp5PzOlvZLxX
9mAXLgQ/vil8KrDuo/6qCAyBXW4B0ykNwRTXsIrP3xsYmQBJMoskAByf186ZEi4BJn+XErRCx/hX
dj3r9GxToIiCiPLKHrEINvXS5ZK5lu4UWm5BzLToWbROCOQ61nzaIRnP0g7tF13hZCecsHdNPWgB
DUF2aOTYOMJX73UaHvVDtoUccIzC1hPhSz7ctGz6oRbBNd+RtWT6c/IR8bDb7LruFQ5jI5EVSPbz
vGrzQh4mOOEVPOdLaiXQ1bqnWxvBtA2z2411EBRLzaoY3SfIGSIOnSQkyA9GildSTBSI8jm5B8Rx
MQlHN4HGkTAIwmeiv+J21miOCHUWKOde/DZ/q0Dhx0pPDisTZUJCnc8FAQPeUW7v7UIFwJp50ND2
i4MTunyucz/F22Oqv1EYjSv1aCQ5LHL2yS3wV0D7Utw9q3cEwOC+oDNDTLL+J9E4EpMJEV+vqN7x
3AroG0fvVxYR/nNINRe7WFgcZ6nPuH0fw9Anf2ZL7BGcqXKjaDZx8JpaVB0DKln8koF/APcwtL1A
WmhLrFjI469bKO1BBZmtHH4jwB3rev9kmQ5xc5xZgk3+4yWASxsvi48Nkf4ggIVTObPr0w3UzMsU
Fo325LwVL3K7cdKPb8172eiv9Aw1ABpQGdcgHPCIOJBn1uQnt1dtFneTioqQGUD+Lbv2v9MdO/M5
tgt/PvccdKEEN55oz0vQ6B2Wpxh5gZ6P4Fq0sVkcwZ4cQNNqW9prwFx+THNbGiI6runFadxsXHvU
s1NucYX4paDMMSbH3dy5EWj9VN5sF7WGXKp4tjIViFK7cF9kxgepx0Ik0DJZzfmthx/Zj6uljfKz
5zTJkauUQ9GtbPJxomuJN5iOZ2SQR+lLVTi1GzNEfoYT2rWtsFDEh4Qb8NEbDh/hIg7598A/c8sY
/MnimvSxkMG32XxwKoTTie2NLJFOhOcrZBtg2grCuQVHHRuRiNbgs20cSqmBpo/a6O1SzWUn4gBm
CaU/IbG5mcUCWWi3P8i6PUJhQPAyXGbsapn0TC5o9LYaVAD0+UaLNU5E1j97m43zoOXBbuMoQkjH
n2SqjdZionxfCiYi6cZmTc6UQ6RsQpyZz7XJnAbjTVZ8x9cEmwCCast2VqD+/v6nyPCkOXAncHHh
vI9b3ywf+g2bC1TcyATOJ+PTLG7lMWLzfYQnaQkhLb1Iho/pHiCHbPYKxhLjWxgTQNl4IZuSTBAP
8XD70ZfgpodpfRXGWfiqvBsLssbBkYgUiOiucubtrZ0efS6cwgXndq3+rTGGQ9S7nOJkCY8mYLAV
SfrBKAMRQQjvg7Ij9i1odDQJjDGjZVZcumcvMGxul9TEdvfd2rr2vd4SFJWMLh1FLHqi9urolCET
eFNRof+PYemSIkd1NtVxj01i6hP1tuWG3WwYvjI99Kcm7CSUNW0SUts31GfxDtcLANYT7R5N6Gfw
l5SXkzovvYBBX/0XI/hDbS33P5f2VAh6sUo1ttzl9881QpL1+8ZOSGehdbhP1aESz8Xo+xCeLBgF
0eKq2/bqLAGm/X3YWCQ6fFY3aQl1MuHzHbS/TD4WHmvMYS06nheWXbGcyuyT8gsvroEhAO6+5LcA
UtQwVW4LxqmNQLKoGKFeox1LOiJSJZHQYZbAHkFf5Anxitm2RBFjXHlt7gul2KrM4Ru+UaFfpNyu
9Pp30F0FFIAN7afrL1RMDMWd8dRrNn1W62z0qlkUQfUezwzMf7gwT37Fixj8K5HbbZAS4AxeJSm8
NreMl3VHBih4mt7G9CgyYmvLm6VSyHH8wsgkz+Rtq0TPvUX+k3wGrLsGTI9tRrxLTpyFcZPW7kbz
iBQKej1EYd/8t07xZQemhq32inEl2PRpzk8AXt2USb4BGd1UXJPjr1bU9UCGRDuIMOq1ftofISXk
j3ES5+VfSTxDWhWViE43CbpgjKFhKw8ioYKhuqh+aTM6tpWVgkmJziPOfnadJqw4rtYRnCMqrSOP
uAPsLZr+qOMxICCCZuPWNF6CkAZq7x3Mi121rfAMfyIeQjPn9tmj79VXbHq19SNi/TIuXcEpIwLu
hmkO2Cm8lWwDo2lmdc1ijsF3dQD2KPcucgkvjoQOGyzL4LSoS1vyPhcuJSBXVRnenLw77FLSiHDZ
byrYUW3CmZUaGG6CoMs/JUJkSQLewIptgLWE0Yn32qPmYfHI1gzakSgYVME2OFdKVAi2IXlqELOv
w4hVA1xUOt1B0lVAPEn0sSwYYYBpX+jfiuuBVuGDqUK/nZX/TRNRYJmy8IPCr+HwO0HYyGYVSJJ3
o7C+S4gFT5MZ+Bqg7P5wL7lPB8K6ljdzH+VyPkTy8LVJJGnzQAfMX2906NOQoZtU++0QTtLPYzB7
Y32RITTqr4VpzHzOkzUHC+GEMTAJGOq7SgG5slTQuDbAnbjjcxSXpMnCaSJcvgWx1HJ+omFa6GRj
QqfKGlqZH7m977qTazFdJgNEeFz5dwdg7TbMcyctfziMADhQyL6xZFK6OhKlbqvteNzgLlBENofY
Crkt2gugZuqzR4PxRDzNI9inVAAbHdaWcOjjHsaZvKA3cXjxasWaM9rsCMu2Cek4faRUmkrs8Nay
5/gmB1Em42kXjiR5hM9NRFCrCMnwognxmu6NX9Rw/Kxyis632egBicPLlbesRc39jX49ApiDHVjE
RqFls3cv4bLWinoTeZJf4uZCWtkY3ZiPAQPWXdP1cMHra7ev/2AR55p4CHDeN4baUZ4XI5AZMbJv
H3MGKMo6rztqDZxgGkvuFnWwgTb4LE7exZLPZZeM054xC3zf8HSZ68ytGiFis9AaUDqZRHatKFvx
qbrSf9wA9N3rXva4IgoMkYZPu69+pA1Oy36lMNXuqAQwgxwmQ4aC2zLdh9JGIpVTBVB9ZfJOGDF0
t17CHW+tDXix7Kpn62sI+pE8DQjiXbjBYcrigAeci7PjHRTLOSYYtK5qh0zyX2LvKiHWlbwqo40S
DTOlrnSbh6rTE6bSEdcyUZyxxdii5szDJ99A8hfPmNVeVNIZUbh8TlMKJWrejrb8mfTOXWXxZuad
23GhtvjnrBMG/7DHss5rALEqa+fFaAijdTW8APpUDmH6OSetydlKzad9aSO3fJ1PUCSqI8ZqWbiq
S6AsE36r/3scggvZ5xTu3FDD69KObOuuzBQ1q+rfAYyAdP5vUgAC06ZhfZ39iVCx+mKeuWznnQgR
oyhtDT/iMgXarB8j3Zt3HnuzkN6FN4iCyfI9gNsO+hxDKZeFfjNt8p6+wmmLJkuytv1AhFKBDVHn
7KAg/c3I0xnc8rHtFnZzf5lh8E5yB/2/3Z0n54Aru7KdRMNX9EYSvfshkktAb7UQCP6VnKGWOAcL
pOWGpVGOL658hM1wZH5RPja4ojK6blrZMDfmQDud3qRU3KQks9p8lsy9ZTtKkkeoM7bf5mqJj8wb
IghwaiuuI9S585fnafJUnktiabQu7asleJyJi8rrFpHLxrBxnL2FS5ILpROJ02iIgF6SzqNGeXk5
u5uNc4dcfftXjpFkc7ChMGTdGywvmQdT7uvY4A6ELDhaLaFWGAYn7n4temPmjKpYhJGGsrcfWKuE
fO5cHJ/VPLAKGfQmkcpmjqBw4cYQbHh2XdCFn06RBh11b5Ofh9DYEHS0kQWhBNJK5mVPD5D5Afq9
K0hKt2dUb8Fssy5PaHwO+RwtxVWgp7JJYqZmZPwwjmRT2vHUQALt+c8lSHLg4JV+LjI04EJR/dIU
ti5LtVHIs2Cl8M0m0XY/ybYfJ4oqlZmgEXWzcEdqLE5TL8B1cch+lqPQjJ1iYGDaAgJ4PJeBo5rE
5EsJBqSGGkXFEKMvL5SOFca72bi+BmUQrbkcJHeax2ZrTXnbJdnC4lPaFTYs+r7aCdMUUUzitqzp
2u4GDYdT3uw00XAWgIZrIVAXn5wx5I76ZYZ7M+Th+jGwOlMUTOSDveM5kQKvj836j9xhl5rVusrF
CA5adpHzD7hnqqAApvwjY+yq32ccVdLquhAxvJUGMxZnAFcWoIHH0cU1rCFdDD7BItdRkkA7uzbv
uxDitWV4wTLjzItjvHCqj+j722qYWyjUm7zBkWQtzh82qj2fhx+lo8TWc2nE6uy/+755AlezgGjZ
U0ztaDV7tqk2uY7294rWUJgssr6Qfg3b5+IQWZAMiFwoLkSJ5pWAJZ/2QqOLOm/7lH8T+cFnYwtN
5/fPv54wD07kHuwkfw+edvDQhShocClZKXlDctaWKsOLz1uM+zXkVxjNcGvzNkBs/FoG5Sh+UauK
C7qAb16/eZb5GE36BIdReFMWLeX8emOmUEyTawQzXdG4AQFc/w+KIeIgFSonf/2Gzyoj8OgJA8b8
peb1sWPqs9lK3aKWwUdEA+mVftjCEE8N8oMABnnSgfpH7ZUA6ymz8XHw9f9AzrqHkKk5+BcXj/p1
4Nq1i+MMGvw5vog88Q+EI9jXXJG+uq3cGojJTahhtQoWcih59V9lf3iWQGXEWBJMWqk3DhcoQOUi
cxsGQfHZIxo/RCUcM3ygC9jMf8l9/jIADafmQjaIkOQKki239JgbzZI+qLd3xZIjOxEDsu9Xwkl/
I2iHQS3AOSKwOXMXvSuCVnQvFTDxzGxQysllJ9sHxKivG+tTzzMMt8ykFFlNe2d8OpUqfzMzSIYd
GqQjuy5QLN3wiX9pHX2+DdttqfewY2G9Y3ipJxyCH9R6/XAYPCMCwKReXXm46Jw1sq9tYQyLuYYu
RZ8e3Pwk3gZrYViynbUJH418Gbz7GOYX4YwfgP3oB0/uHlz2QGTEejB2IX+blgdInXwoNHOjG120
E+0wcOwetk4VANgyNHEPg0F/HGz2HdrnJzEdxzQFMwEXYTFiaPR/Nc/K5GXoJb3Ps6U+TWa3cvJI
oV7nLIHoRN/e1vNp37hwu0cDVwpCGA59quG93YTeWRIFfbpE+GDW234ZcYm3JkdhI+yYlsCKrXHb
emDyJJYdexuEe4HrwLO9l5lNkpB+htjQyDSLzhJCZ6CqMVdbjgWsqoGc+62F/qF2bdnUvCdHKAoU
wJJXVKUGEhkqZrqjLFFJ4TbWl3KQ5CegQBY7jiWGs93YPWcr9EzMRHlYlrPRmxxVUhkCrfDOi3UX
LuuUkLs83qhp7yeqiRzBsDzJbmiDOxqNRVNLYzsKPVW2DvOdU+xwvq0Y/p0/tQIJYlWHfkd1N15s
tkXZNAPnT4dwFU2sPs14Asers6Sd+BiG4StJ0VStrZxh49Quc1lB8iwYJTEgEdfcPf6zLgoku0nC
+jduj9dHeO9Np+jKeMzIy7Gs4afo5ndsyWOeIR5FRhSYjU2qLDtwckTAH9DfRSTDzpNzLEbXXFGB
YLz9NEeFcZv0KW5m2XUPjFYVw/AQLPGcx5NO5IbEnbjxMHVBJ+bnqXt5+2mTUs86E+/FqESTxchr
7u/rCo45L258pK7ECPRgRyUicBRwQ53u7bXTCFgi17iw3DkrGjQLjPfRh3B6UvwOKV+CXchM6b5a
TciRxZAeQRI3awNpm96axjyKawFytVIEIawpH2I1rG9N197uJIWzt0FF0I6g7TpOomvT2H2mLjU1
OUAPfY2KkkJbnFfK7SkpLzlCt1VkU7EwVOxboTTuYR8cQUnbt302Sq3+CMA3dCLLTa9g9ggi2OIz
GfLMruX6I4ryXwqUjHKEYCoSlBI148XMA4ORgWHtHyyBspwo3qYYaMZzg8Z6q+/N8CaQIg6+AHUl
si1VEzERTdx5nMQkdbAyCZ1c0mRQey+/8l561LAO3NUUL2D3cUPqYUVJnqQSVokz5uGAuth4aTub
anMr7soV4JOU+MpGSYULwD7kb0iNDS0bw7g+lx1p9lIeJrS/YLWdo5BajIbo0e56CObFnEph3FLr
eQ7dhqHLZ85CO77ycPTd2lFqW4hNPB8aEGK/bmu5RO9eu5357dn4OPP3qq1Vj4MrRHipfABNId6C
WCP7b76PjDa6zvKfCzKMaS4AiAfyR4AFgmDzwKARnZK57cEv/gMc23cRsDEWpOFKxHYyVpwbsy1L
ay/SWz8n8FwsKCed+bAhqDJvtvl1XSfJzIX4o+r4DoxFhm11XLGICCY0s/A0BHt/o9COrGr22inO
GYdE9PF9Iy8pJLfRC6vb5KJ4UYIpcuFw48ySeaB3XgUHlf1WNuJJ9jmA8g/kcTAD9YvS0QN4oO31
JydzKkdGmwqkNODxzSq6nd8O0tG1hXoXIXAR7KJDDSm2LUSPGHFHotMpQFipQueQaaxHJVbczeKZ
3nAT+zu+8STV0duwJmW865dxnwzgfKjaySxDTQZeSRLa2ViHsGqHHBiyY2rV/+e31d0e1ZWiR0wb
Dxqjmxe/0JHdBhczYU4lHfVqdAax1mNZEfzDYfJ6V1Gas6dOjSrIWEqo6luJNI7KFK671oxc0xzE
lH8NrAoqN32sObQiqkQBgtBgp1QYz0rR4Dtv0pyM/pT85Sk7XAk3jtDlIXQjkGo/+72H1ZKH0SnF
9k6xhTLGLh6AO8kC1Nk5ebiYagrS87sg48T2ZkhZInnc0o3xEsz0XMTFAwXvdKu+yMPRN1LPgQUc
cHfWTwcRzLxEWl7U6IyexsWT+4mhWlAH9ryY/ApMHSf+NxU7q0p/Qrpd0gaYH/ikHRXVw1z/cb6W
IrbhquF9OfAhgTsK2nGDUljg+1T8fOCEMf4vxHj7eB050dHT4dr8rfRS7mSI4vnJvXH4z40yx3fa
OvDNGv7GugRK3XkCi2AI/2rxrFmVdDuK02lHWafCvWiCrxHPghfsS0IQBzXZ8aAPw8M2VyY8Kqa6
ty3oS6QZBOuBgbrAz02hckDXFe3e+dRCncgTLIIgwaTpFaYgIND2sZ+ZecaTlLXJQSJEZ1YXsVo/
vdpv25Ha2tSXJZypnQLsdom8LwIf+pEaItO6PDcF5En3CZpYYrMeS2CqUAg6wk80k17ysCp8Av0d
YiUBwYCQzQQPsK7Pv0B6IC1pB7Qx1gmbZ0wE6+ESS5lPHTKN6+UhT7H27gATepABKw3BFOTwu17Z
h6gS78SBPnJhYOLkXt24LHhgdOZ1a9JWvaThJ97OOVvzA/tlmEALO8voCTi9KPXMJuA0RrNH7jeZ
FMN91syUHn0c6hJ19SRObAogyxIvL/QtNpoY99/1oobKF01fQDypyQdSmHoO3cObTQ8SPQjTNTSq
NdBMSSqqiyS6G5vT963woke+GxguKL35CNp6rNeAJ3YW9GJeqjUPLvLXYJez0AWL9lAeXHRweez7
TQVJmj17gWBUeuCYBIqLRa2OA44dnZ6LTpxLQBWnBBnLzafVH5Luko/juPKJtIaLAIZRW9sjXmgM
eLOnkZMmOZS1Ks2qrecDRRmg1Agak0VWPxxZuoKwMnOsZ3qqodhF5ePEpnxwXfz5tU3L7RBq2vxP
V+mrHIs4EjFSbyLxASCOausHOLPEcDDsVoS55xfZ6ivAbkzIaYhVnsFp9mzWzJPU9jn6w1y1k8WL
1tpm4H4RDCzPyuqnbvkiNsGU+ELVexIDslVsXm4OA9D9hXDrKkSfWTc3IBlne/PbTgbJt6ZA8s9K
8p74spzl7ihVxNQ5thZnGJ6a0gfnXPTTN4buWeP+n/1CTJ3sjty6PRyOGJoNXt4rtzigh8SrkhtX
ubRij9zHwF+a+TQYv170h+jfIBCVazeDvQYj1g+np2iCeceFUtMKqUmyDhZ/o4jMKcZtjrpoTc7C
bCxZckaOmzcdePLBs+XaJg3WqQRMRHZTFAkmDzCoYJXPm/ZxXjb3rweASKGMe54SgI4W/+fSjYtO
ES9jEDPQR+3b7+rXchyWtGWK1FnHo3lKSzazsWdNOqXNVS2x8vP8M9/zZPpV44RjJnOTTswM7675
rn2OYtQX3d7N563QvYX62xHNb7//JhiJE8KB7Nk2PCliYk5EhgVNTRBAZ/VT/suukPsjlIq6AZ4k
emMNGtZZjtpvXZDpkwQ9K5OIVTQOhCRpYef1A5T+vjiy6UVK2840Heibl6o88GhXNkakH09Yme/w
QAXdxRCkcIOBOU9eqzU0DE4TSI3s/U+Xw9CTtcGKiM7pkq2iRvLF/82YWc97SU5spq26TmSGgzb3
0bhSjtMy6tZG6Sspdo5oRQ5FyZzLwob9pGZRPgYsQImCkVjCrYpRmxSygwJQlEbJHLvrMfKt/Y8w
wxGBw9ZjlUtXJ8fPHQS2b1rabk1oCbOr9EVTa3P4OO5kQMVNerHol1+4NpIXgyqCwX4J3tedwCil
dotlf6rS67kIZBOVDit0Sxcs6YtKrI/H9wbpQLUrAxOnnm2bP7MWYHVh4CMnsUREiAzJ1c0b1O5D
MH1r8WuF6TR05J6qn59kbCf7pGQR8wX958t+h1YUe4F97aKHVzW2GlqVUSs4N3dRWEgYbnB5WVZE
/mXtqKTB1rzlFAQOEI7LxWkcRBqkW33WPP2p9ugi0QpCCiRm2+Ovj5l5lNJfs2of+ae6dE0hJuHA
dkRyxaX8l5mzrXbWu4l3AeIeCbYBT3hM3YMHDUUv4oEdfY8yMH5CH63Y1qT7f+OxxtqXGOwfSOCa
LE56l9y+HtmcfinZ51XaD2LXMBZDPRFjuD7pmV/etAp+jOpxWNcDKM0n0akVYwRj1ALrgYhaE0pI
tf/RJK5GgrtBEOpQPjI2IVyGiw5sI/KumGIX8vG8XoZJTQ6gSRMlJbw1flTAiJ01O19zSvLLAGn0
qRjXhQCKUnF+t35MSGeqaFk9sCt2hHR+fVccGyQwV49iy59OJAMwQ/hHLKJHtq0deSnjiiPvEpa/
pjyvB7LRDurGr4leIXMdnkyU6c8Dfmx0MnvGSQQVMNl3R5Nd/uadRMgSYnk4w/YgkZNFW9iZ3sdh
g6OqvuRcUtlKdLC+6jFhjHoD8NSgyB/NWqO+URS448zk3fhQne8ZHGM6yMOYHPd6YQACbHIuFiRA
4WWxXgXe6o+Rx9m+4Lhj3YGu/ratsLdJGk/z+cODdCDvKwe8PLZigGoePn+WdymA9mqMYAxpI437
j2KSqzEvhAOkkHXaXM+0+zWjdHC9wUkwFWxdTc3b7ftbT2o1VHQicaQgNnXH5I4FJ7FPi0lABZD1
gQ2f1FSnQuwy9XPnlhTz+TzV7gryGukLuOzp3+LEvtlXhnw5fGNSywd+cAIFXNlRNBU9AYjV3NLs
EceJ804bIrL6GLV3RZt6LHCRIyDyoddmTwnWzu7MMOHbpGH61cRhtzTRQfhsG3Pbymx3ra/Z0uru
uMWPIBAotN0fAt2ITyYRVVTzYd8CFzEkFSX6XWjc4s0NADJEDhRs09HejV6VGvwWL8q6cOGR8Z8y
0/0xHHDQiEqUHCzBfDhBbJOaSX73dACtUk3gplmXy3LiL9MF0JENGYDd4VmSb01DBz0650E9cHXX
3EhLm+lS5XuxmJyaSX3sZT2Jl4CepRN0YJ5yWxY2c+V3uH9Z0PgKhs45d1W2HA5jJOGtB1kQFm+w
+Eww1rmroshKkUSnzjm55D5gMfc4CNF8A+eLVQPLWlH6AvuKX4yn6TlRKVgK/FscbF680YhEWqp1
XJPGHZ5ZMH98XKWihH3lTK706aou6YhunrjQ2ZrFl+WT7+/1ObppZc1OaEy9QKANLWo3gTSDMPWX
RmjJWvO6zd4GQhrR2+VE2tJwHb04i8eH7ISYElRg4naBuxAF08FJfKsWmVd2Ihsx22JXffQ+0ClM
7woo7mfbuoFH52q1OAxNF25ZvXRe/0m8oViNc1X1xPQFeqGDZLUDwLt+fT20aHI+a+SxXV/HmKKX
WQf+Rb3FXFMbg2i6SFKWqAwDIrIwo+t3K/JPszHITKge/YvGx8K8uwcB/4DYitf+UVHzFrgLSZsR
v/KnPnwUep4itHX2eblcs0Gl4gtpE8uwQ90m5oBCi9q3mGXcdo9aX8mVh75VT3y2OiAHwkHagTEd
m0EXFhU3u5Q8X3zGDdkZ1uUQrDDbZnz5+qY4wNyiqCjsHALehNVjusYVvb2GY5h5iUR+dx/i5n1t
td2UfLcQ9mdtW3fyWjUk8X7w3Ysbl/TV5fzrAVm3XkEPHgJMEho78kcuwiqslooWUE4GMLWmwakW
ULUjKLDY6ZJZYmNAxFko+zg8u0+bzTqGa0MV4900Oi/1yEGHgQahbBhoGy+y57BgCrFHFoFLL+aa
cF/acnwyZX+YYFsYpnMxW/TfZWZ0Riq3cSiQiVQLyh1aJs8zaSU1TBS179jzXWk4G1/yOea5kDUV
IGpTuUdgru/MGbyolUz6BLn+UO8wDh4X9T5l7CWQjrKRl3D8ljCiQ/Iqv94bV4hZYAd7HgbQl+tq
WfOK4O+Bi/S1dSolf6VYiLF2UuA5/A+JMuB/j5cN+zjthVK+a0Ysc42dnPF2DwrOJDASpiEu+8HC
rrXth8XP+ACoGS+Hnbpfw1UrpV5RVSx9UgbpbPpzGNcxSKwMC615urnCq7VZXeO8UmZlqA1ILSIy
vYI4Xf5ZBgGxV76YGyOf4Be7TFWYbR9T2FhucaDfriSnsWsVFhAGQOPjiGQMQXHojuLJYZcrA+za
FzdWsrzKQhf8F+EyUydB/w2Eh/DQoS3e3++7IKDH754iqgPdnORRsmuHlr4qaW12KKuQ3kXIy4ey
OTNtqNCz83/m36rIefOMd1DnSlrBvdOwoSGMV6UhA63NLVcjsKLhW/BwEvV58BzH9pWlQq6fcA0R
eUZlYy+PGvX5qI2QL+o64Wsuc0zevgcAKrFk4bgSOBSMOP3A9y7Drq6/9xAH5uAwLazoeNgxs2ET
G1iBvNplSI5Si9kwtNM/nF0QS18PZDZsT1LxFi+u5p02948PM+iwqrMhtSvtgp1EbU0Qk6veMqR4
oZRSxjG5ZclIGmrRbPD4z1KTbmWUZYmGjp9mWGtrq0lHh3cLvr3Anda6S0u4sH/HHCHrOB4WbGmm
QOD9OO6SPyhW1NZvnT6WnMD6tCntvIPAhlBJ6REgN95qc7RU1DeR5/fsB7LYyj/kn3rXRGONYGha
yy3gZL+mv8hUfgNyq2YTHj3flKW9mt7OHvji5sV2ujqMCgjX+4kQuaOMzYypR9tTsD8GEVASemMV
ZMhx+fkoXXRzTTiWojxi/0vxOlTILL8KAGcSpguGFSDlCbWNTMP+NJUcetz9id3cel3WmTyKOudp
UrFQo9le9PN692k5wBxz2Uf/gQnHQf8HPENpXs3ULrNOyuQ5SnM6wHOPLw4IqIdt0T1JmpCrhr0Z
F+3Kz4RqQSf1OPtoLhl59MYCFYhqNjJsD8ITEJpzGEaN8wt44eDlRf+BuiMM6gmMnsBjQrMIg7rn
cC2AcCU2OHnoTt94q0uE4+6fMPdMcWT6A4pVKVrfy+iUN18n3zwV30/jzNmTTPJkjlW8yTULTWf5
x9HZdyrpKZsWDvpKL7IvxW0WzJcSgYGASqCTkWPczrq3ySlTuA7fO3PgjmaXkk6CISCOf0cBhCcU
9Yc9yfn0HtWM7GBTMxxfiqLkbdWvouW0WMx1QKDM5rgkqeqdOtMHIB98ST9e3urj/dkPKrHjYtV9
r4+TW7XFqdSH5h0aKU0lwtLzJdXwoXRrP11zmkmn87IzPuZ4ouYK5J8FdMVYkPe8Kv7oMs9fuZns
pP87PnjcY44Y1ls8t8DGvxw3i8F9IoShd08DWEELgZ1Dp1cCtk3GSuVLMDaWCoKKqF9AtMwDA7kA
hmX2FgMMzWMlbk1zfYw+EPhkbrLEteO1Bb1Ty2kN0Qn892N48La6pOZpKA4hIDDkyImu60T9TNiE
Vcgw3GEgdGPY6F9AMbL2OETwkKLpKl8ak+mLLiQbZnExgds+phMmjU+bsVxoL5wvR3WvjVVYFYUm
A/yZw87wGTWarAakj5jdHAFcESxudKkI/58+CKUlCquzpMifi9nX0HBebzwVGMzCtWO9dYqM7SkZ
c6GOOEJOEalOzdnY0Gk8p5gaXQ1Ix494q/p5dHufCvPFky83U1fOu90Rvv7byw0dv53sjiK8woPV
OsXGRX1fRMD4WWXURyGiBOMWkXogiAF1580leToGq8NaOirRTOGeZChRLbUw5JemtBC7P76jlMsz
ktlPIL8Mp9jqgbJRpRBb9Bt0/n3ccE1wBod48OWCOIwqc6R334t1upkFgL7WxC39TgjV2AJ2CjSr
l2YjUGc1OHPa7DaAHjJmCW/Uw7I36J0Rk4jrnrA7bwka8lkMQx4pXRVFT2RPrfFKtBiJ1ayWdL8o
nSpwGZKE8767hJW4wBz0epvOb7HV++fGEJ+6GTi60VOFjJIpY9ykwrPEkG1aa4Z9i8l56LWxFDfg
nBhPG4cb/1SxEVN+kEEN+VnqnN3lukGHq52xyW60g/z73IuLrpCMVhL3xj2ehKe6JpbcGT9pn3MD
PMKUJcWxPDwnFKdUfGMiciI+Fsy3KJKiXrmCZ36Kpveqp1nJ/pcNHJQXH6TqYQqCzMi7/WmjPHhK
r4QPX6WbiXNeySXVU7DuWgpKA+J+096edpiFAwnm+AKBOwfz60U51PKHgNarnQ1eN3oDsXh9VKnF
ey0naHVoDSajdaNDhTn7PboAS2uzPXQay9eo6iHGlR5wk+waaywWlm1mMQRMxZlz0t8qDs9+WgUM
lKCqzbap0rnS0Ryst2son+wdcVthRX1ZO/+s5Q8k5VqrrzCtbzZHTHx68BbCyWTjOSRAA2yPIfSN
4ccF72OoNUBYw1XIy0roHty9y/1p2GVNuNgE2w7mWY0xAW3EOsF+iWsyx1zyKfFauJz//oGHDX3Y
k+p6Kf/e98+/13LedVYEPcuDfpSBQOZdqJXwggdp1NXiYeHfptNetMfwdEm5gvTkoMjKr7Jky6tx
UpaesJTHLxT+CYk//LUEJCIfm2SnA8vKJnQ66aU987cYLriiaGmaWyKJ++khKG/6cpPlpGrUN9k5
5Ipk0JAxdM6Ncj05/7k4KqJmQlD+1/i5+gFniKUMozjkVXeMnLgtwFat8b8vmJTHAYlq19LQGcyC
YVgelWRkNJPg4qX3CQPxffnGUth3fMVusshT4jhzffkLcovZLacEh14wc6sfvwwPZSc6vk5aCGcf
pfHlB+j+8H9zpJry5r942G/Nvi8Lv+eUrqCioN5Oxgg4Zq4uIlGXbhDV3o4E7cOkCIJw9/IEq67B
c89KepXGPW22llcoXNxBRHi2TvJ7GaZV433urwB9O872or6kLm+4O3TTz2yDTIMa4Ah+GKep7D16
Wi5gl/AYeEouR5iL4Ot7cB2v3+dBj4CktAOXfWPcJe+VJkieoQzPVJw3w84JowWAVNvVvStKauGn
jZcC/nRSMQ2kUVeVKMV3QFg4NNpdtCitE0dNaugv5rri7zTL/xwK43SPm6GyzTobWFgvkObUufXh
tPEKHZ/k0LDKidL+8ENVWszUD3sUCKN7GpAVfmJPVQZbSQz/mimpIjn2cygvyepFar6SAD91zUM1
V3W5ABCbsiEyy5A6pMYXdPHMmMRfUnk8GwGXkgPqmNJvyamhq4+4IY9WIh54Pt/t6WJuRd3imVWl
DF5WXuMJGntxmVVQCmZM88O18SCPIhuVm9QC4ysc3XL/Ep1656IfC1EtL2E7BnZYHvtpMhlzEDyT
i15p1QmoUtKwRvRFgdqt/rKTaDWpJVQgI0UzQ9w0t4U6Zj4LKSGOMxiJOMwNs2HAoK7fp31WAB3I
0EqScRgzFrvxMPd7vJZJY0a8q6UnpmoARmgG3OgnLdvGruyL77uJJ1VHULautiYyUAphEHUYK52D
ABZaZ2G+HUlgOSyjC8vI6Ok7RRqd2LywgphAyPw57bVwP9nMbadBsg2e+AlQGsz85AlVT7WDIntA
F+l4It6LJB8LsbQbkeDaq/hoAlg+vycqULBPDyHlu32GxH5HITyupwIPjeLatN+oSLfUMMujS2h2
FP2gbe+SM7xIGViCZklNR4p+CwX4EU1KzpSHZNNMc4MBu5jQG8AQOoXTl8iWKqz1taUIx7jXuwVo
gap9tjgH/9L4qxsJ7YyPv7s2Q5AsjJK1mqiwcT63QsJNjzQ+0QuThXLxp7+c48Ua3T8bp13j8fnR
Rne/hguOQpz32RPUz/Bb2bki/lRwMoOOPNKpg5jgv1tYDQrbKgz/AfzSWXzOfdBwifmw4RMX54gU
9nb5YrjUmi100OXeglwZX+SQvS3y85S5mx3D0dOAB909/RIkk45NER+w7r0JL7Nixb1dAgNQZtpd
94+65m8P8UAwGC50a5x7fuVjbuncCVY3Sly2W6s4cpTEkZJXHPQckbnrZk4a/150zpmuVaXSLUvh
CQ9whH8swfP+lPRXZwUUx6/WwhkooAxVVVjdwkLiuZLResvfsF7UWKoxYN52w/OVtp2YSFO1YcEt
ZAM8g/+E/W89Kb4u+sKPELcRbw52cAUctVZDlVE7iNDhaO8LsNBG+7ys76WByrXjs22Yhqr0cv3E
1quahE4S9YAsK2G8UcAHNVw3+htg0c2CmARtFIh8sIx7G+Pwcad9nfrXEDxH58J1kLiuYc9fkSwe
UHjs9t+8moosy8ZX1O5/XyVuqxSaHiW6V9ni1AIglVfoQeD6KEa3g05QF8IStv49Hm9mIq6B+QVp
AMGmlZNGFZZ5yLiJjPcIoFVDmsXIv9LTnnCh4IpMb6tJNpGm12RWBCorLkbDr0vUH6fKam305FlO
xypWaSjgc1eZx9cijRpsdXmfPtA884urzWWJtkyjxF8Qtw4CsRT7a20m2N/TxVuwo8DYGttcWXb/
QW/CUlGrL8lRo8z9UfxESwl/OxNk5ukQV8Hg4wTSGbmwfa98U5/CgkPI5i2Jx/yDjk/pjvQw0VSS
ZD+BNYT2CSAuBAXAd/zkGbOIeAYffrU4OojoXiTcFSU00+/Ac7eL2nEEdGLXGewdmMHTWvH8+M4/
TE0HzBg1t3QhJixdB9mgfi+gSZXNsGzCxiCKXj/ISpnFh2adpJR5GucsTu0Y8qfupmQafSumKH5Z
WkEmo1OEIOjzvC0qAoHADRYxIMvjbf7ugOmx2leakcZJZaKrOTB5lPJvjQ1JM5XGAX7YY/SRAGys
UEBgjeU3Oo42+bWiYAOGcInTo1bloCg9fq0Ps0ZZcfRAU4XEtYpNDMRgZeKyULMc5n4xOrUpGEWY
ElDw4yBleOl2sT2Kn+SEjchFwqKU5viShRygWjqeOQBX9m2mKmrOtGwSCNNTykuj8GSC/GMgUKnK
WHHUATIX+v2Hm+Kn0AgcdlO30rNAJsxw1oT/YBizCsjp/Nfm3pQQG5MQ/si22W6F8SA2XF6oKvGv
QpAZbZ9+k0Bj8/+b/Dpo5r2bSzENG6j1Lvjks7w2NyQNy25jWCWGz2ovGW2rjgwl69tJFOIvOqca
r5M61cWwh57xyhjBduho4hpNL1oXJSiykxAy32rb55f9G61wGsvF7xDS+qoSSGtG7oQs3XB0b8VR
ZVZF1cfQlj+ffqcXoN8QZS/Fzu+Nvfin/P6E4WNfqk0i0IFbkt50f+vSyWoxTaTfHtWswLpTPBVv
0iW9SlqlDENxdhbo80oCuXi1rpwodCrSzOe0a1+EQ8K4MwVZbrQAAtyIaup8gz/FDRn1DurhsEhj
7UkdZJ1EVYCbr4i0hSZJwekA6aPWfDPjO/jCgloBgygEgxM7itFfyhmQLPOVVBMOhaqrAtgE5ByD
Tl5IAPZHAGpEY4FmgKgVIkAwhzp4FWgL6Ll07ikC1vFZazlDRLe6XsllGesSx7j6XdoxiZWrCiMe
eaKBNT6DVe69DT+hRKSh9aJBYWZlbnXTBnWUe3srFBrUVUdH+gRP9mwOGJCmccpeA3/FhBsfclDc
xtZlP/+i1u+xM7lziAfv8EZDlfCZeiQ/8JFO6vRBqDtT/RbojCNT8yAeWTp8sD8khl5mm+wsyPJ2
EYuTZZTTQJhoyxRx2OCFXveXuJ4g8uf4EU+rurjk29jKG+WuPBSZU6CREvwFahaCJwRPO/v/sHwj
WUW75EaIc4yoyOhveaXYuQnmPLO0nbsfDv0HrPsajBC+FSmKdA1YfuM74ZQgXCJ4CJ7kOvhxaKPQ
ZA+ahWPiBFZPtqxOGcbzoSDi/TbLQGZhPEM1NBT0ayBlxopQvEzTA65pdgA+iC+zYE0FTIZYPREq
HV1sFGEsyRN9JgsBlIMRYQPxoPrMSzUqdYBE/FJ33qyvwONMtqq9IxpZHQ1gfGLujNJnE/RanOsO
QG9a+n2qe/+obzAwPPpLUoXwzfq4K75d295rAkBN71+MBMylRTsJZOjV/QM1kxfajZTv6EU7eptF
JLZjW8+l/SCC1ehwhRow1RAOBNvbQD1QEV2Idcz6w9W0TzHPJmo1fb5OgUlA3kF8ahP1fCWtcnoh
TbgFWPXMvlpNDrM8Jt8yxY2IwwchkAUhA0gle6oz2J8jqMRvwP4mX/Qmj4GtyY8LoeNFKQOErBpc
kmvQpueMI/G+MTllIM8l6m6F6m2Xl3bRsa9C8pCLmrjFsxL4fBRQ8Pa0vuP2WbS08un7EnGL7ZRN
KMccwa1EgZBOhcmBPQIUZW7Aryxc9fc05LSCileGTEMur2/hzpyzftAAzxtk7/hzZCVsLquSo2Mv
/IF3O3V0nC1a9mhcLBJ71u3LrJPhk15HcstZx3Ghykf7fTu408iUizsdxIHUj/JwRIHs4QGnCgjg
M+UxyPYNRtS+rEUiXuBlp6S3v/QvB6jzLVt28a1MLf6ns1roPqg5sP/66QaVwCZQUOant1znMKkY
CkYSivwi/6fZ2e0Spfe6j7XErkbS+SmcWJwHYVtD0Dko9QYyRDAzlUjRkUeFyvQe1HPDs6nHdspC
LnPBA8ECo8FGcvrl7UukbtSELbcKtsCfrRX2AgyiPaY/IuLvlQVN06/TKJ+bmk64KVxf+iN0kUX2
BqHjvyFnbjDrNsDkebwMCUF5rUvitWdhbmafxuZ5jKEY64xGzS2AJny9Eh2eKHX0mrD9cbkrzOxA
Fs1clkXEqTiOfJiHv6Y8Hn+Rilpz1YXU1PKcTT/HfPru/y4TiJgMvSBS6oknH2VafJzQAoifE35Z
O0vPA3lWeujeCxhfod7cd5i2GUgOVrJ8mLpbowUlWjweSVxw1eugrDV2BqKXM+KZ0lySYZcWYEb5
dcK8/A2ASp2cYsSqjVYxcVKMuBaiHYkqlXYHxciihu3BhvRVppMZYWS7cPi4LFqm3mAehEpgSyG4
qXztuoIyUJyhdxFV6wQNx3oABbkqadzxhAbxbLoJxc95lBZYoL8wUXmiAU36vXff1jgr+kFdAddz
2Fjef6evG0mTIyaPOxCXwCYkrOPDXKaxYMtZPgTAYsPfa/Vb4pjVCwJE+cgGAGY7KlbNdN4570t+
xD3nVRhDZnohqfrcVTiAbhHWdL6Zk22hlBWRQ85jdhMoWJUJISRAL/FneyR1ogde4C7mg/tD/N0z
ioqJj9+zyAYlzVzKpBdlXXjDFPtmmv+ZLLCGQdDhk9LO3ecUOBSFIjv2UogPQWtmQ30folnz7x4W
AHfeOtzow5KiVVjNSIxxxSZpCg6y0baG9MsZgnFw+Dn0a4MWlrtFvfksqGD1iq5tyxgpG3vxtWH/
KYtfRrDSotdR5xy3Yn5K9xDC1FV+/87sh46fbXba1sur6PjDXFyKawCcvir8wOFo8F/U90ESm0CS
SqMYzWLSZxnlySatkRTflePYL8576sW1SfXqxKkNaNeMzfCzrT8EBKK4fDklUG2b/JZ4iBZIgb4R
Ljp3H21fMtKygvOSBkOP4fXsZhI6yXasgWX+45H3uT6+RRb24lCe9Fq4LnoIgDKnbFJ6Qu2SDaRh
5qxwKyzKMNejxecG80yPXJO0hODL0OB+iyaJmYoKF9yEsCTzmRJhf6cQmLZ37VHapz22fOTkzKnU
q5r9H3fiWZ03kUvV3HRpsh/KfaavrMj5JMoXUUfrrKxfgfyMc+9oJBS2OUZbTHktzfI7Am68wKpk
0Sliu14xT8a79ZEarzhziCo9uaVoAf+ZP9zEXeWUnf0cj+a1GvvX8zGNW7+ijqpnmlrFhOm+6dOx
rRlS3pxsYbjlBeelAaZEQf8eX0I37L+7u7j3LoiwLpqWf2HHEu4+N+dAVx08A4PlpBN/WTH9UELj
u48guVbjA+BfgPm8w4XIU1b/Lg+LpYFlE2Q0ez5l4CX8nLoOVUGw67z//FYIJKFYLfdtgjI4/4gS
1WdhFY+Z+h5J56eXksPfZjd+9Vov3Xtg8OnnYBe9/QMLapKjY3nQ7MJTZB1pqg0jZC/4ehUIWziw
2dRX67Dhdjt8zstBTxQkDTh3bxEq9lwCLxt0XN8w9fdhT1VipFRExeA+Ep50igxn4m0oy//ei313
iS/AlqqLfZyhHeczm1aNvIra5xQEwflalgGW1pskqSb1hznpXcPdva7HfjZdP3vdXKJYJQSVALrN
wJeM4pHpF0v7DCZREeVSqVWnIpD4N341XajTv7XfeipLMl9pYNL+xvkvBG0riqzEdSKYCWDmVMEU
lNgKyFiOWF+F+8cKagLmz73SpxdHD58uNlDQ8JZlORqOvpD40BFLWg9xSQ1uU7vgQ9Hiu2o1jGSe
4857gCZl295UWJhKmpbBTVyNHxoeWDRIBLxa6zEWxB5hCKhVYQu3bbbLexB7eE1p60hWODPiqlDv
zvG35GlNhMADvJrP0L6upOGDxh3Oy6X2d32x3RlKyqlk0TFmXYeBupJQCYuoFagqY+E5QGj6Zg6q
mFShzLOz/rq3PvxsvZYgu59zzB7yqUpDgzesTzt8mxNuh4n+IyVnh3AxIbOqagfpE/xZE44Bolnc
fjbGTzrOOKGTEhVN2Af/Vz0u1XtUT38mErIn8uRgqx+Ft5tlR2SYPMW7WbELuEE8ezU7TvBJ6+V7
4Q4wNj1hUseTvtV6KAUl1Cj41hbLQl8RcjIINQoQjX2KKf1JOIO0DC9CyCYfcsgY0OWsO0qLuBgA
L2faa4zDt+jxY/LUjMvS8TbT/VfklEx9Vl4OnJe3gH8/9NWzs2iRe36igzccfODAbzqovvpzwcuf
i9gd1A7lvqWfDTKYzJQZTgOuJvAISXnf/93CoSW6jc1CQSW2bao3KgsWk2kmV/N9mlRENQA8SxlZ
qECrKrVNDBlsqZ2isPZm7RB9+3kC/WJCZElY9rpRouj2ejWno8Zz8PBv7QcirXWQ+QXzFGU7wz8H
yD6DWgT7aGdWOK6U8mdPSFpKPaPNS9Fjt/CBi/nYLtRzUdKbS6f1Ya214MhREIdQMNUYwXsy3LEc
z2U1lNCffI//9qdLAA57HTl49h6BsNhZ4NXBW+26nt3qHviHFOCSTyhZRaVQBwpoIrmLA3G1Z48n
y1wYRDdEeql3Tf7CupaJj0B8GluZNPC3CxL/A7QdtpilW2EBVBqw3ZwLxwX3yCta04QlwoLB9/Lz
MKldaITpcXEZK+Lw7SxlCKnSEUqsDu/V0Dc/xhJR3nkjHdmjsl9+iGoHJvkZKlI5QAsiPyRR/Sry
o1tiJbmlTjXSeRJSWpRjgSGPREE1WSEEJ7so+VEYjFrZkpxKkZte1NF/L6e0vkq4ZY2j5KcU51Ut
NYDo9+v1u3hsVRwMtzdDeQZ7bIBm7ZmZ2Kn81hvfopOPt2jUOEoBUl3yjqnkuhKrJC+udKL9R0du
bfLEQ4m9nKW0XTzqMO1AP56YWInxNQ0gsRKjuHnW+LzpFq328IQ5XGlmg/o9yabDk3UnnQhwgflh
Q9t/VaivGv4ACMmNYTzbq/wzYwol+IK0ifzFeNv/jcUxPU2cx/A75b/wLtVMQk2KeEpnMA33WoSh
ivMyFwl8cC0amWu5ICWcytSlarApnYqP/8vmCU+kZVs+AfZyGrLor8kmIKsWH+Ln7VsIJzF7v03C
nsyN5G7sdzE8rFanfjlFJE6DS7ADgxqN1kjHlRRzp+GkJ4duyJtXiCHR2vO6lYgWORbeqwjnUNPc
sBhz1GhEuitZmHDCltP/iYvQRUiXlHKxrbplmrpnw+0iUBRq6OUh5aTs32fwKi5rPS5c5RKqhLEy
UHhLuQjMdc9vD3HMgxfO2CUCsOol4j8DpX9f2UCiXYtch50tgO2ue8MtOiAsSSJUXW1tLFuWI/uZ
ADZgflCXA9pWjNcc97dN1lmVeoa7j6RNyj5R07AL389gQ5VBMqWv/kMLb/k8BrkKc60M+BQ/z3Fv
6uMNIfTDyJny+RvCa3fUGZZyegWdT16euCWH0L0b+RFedEy/08abx/7ZzXXEH4LFOUAuLLT773Zs
XGSJKtl/DOJTsxFFYJWGoZs0P++uCY4LRIBtjv3y8zCAozyqh4JPlMTQFA78GA+D8dpwgDS5oLRz
WTOveS7CJepwoIrsnoXOpE05kfsecmpScEgAejnKNspSybh0G9d3Vwx+eOEFo67qnd2eL4/UvQRt
in0u1pdvck1KScoRthrLEfy3Xw36fWCzqAWSi1Gj7m/9gVsYqyeI//uXtYAuXXYOr9kZqRL+ah3A
RQvh781CChAGQ7MnOQV9cvYe5RnGvz61jH3+FiZ1qciGe+TePjYUjCd5+8hoh5y8JW24O9KhE846
xd2RUrissQDUaUvGH4jACB2igDlMgEqvrqEdTKgSh4gYUQbRacRByp+vBPz6mcVse/dAQa9HqMqy
WjFB+Q5i60UVupoKh4npTH7fPAEgm1I+5NNArshtawGbJCyqx1XPS/KZ3XzhYT5EP1BiciRdJe3O
FVJUegmsWBUx/beuC1aVPeXUwEJYlY4gft7kIXY8EiJb19mjjRCUiealp4kJVetuxCU2vUwheDuz
Y002LOL96ahI+ijMiIZeBWg3jTnKNagkzMNvhQCMbL73sdvtbc54Ijct4v+rnn+WunKY+6eRV3xO
3jyzjdjxNEafNLacT4M7MFigDfYZBOFgkTDusjQcuv56yoTsLwCdQKWYo3MYwLRu03RgZodLclIT
ICpQgoRk41dsl+6XjdEzcWF6KmQJy2EmYrf4+NsPYBG0/TptPVUwP6r+R+Vhi/7Mhx53JSfhVMBm
BnnH3rdZjLQyL65IWPjACNqBWAVAVXoiirZAMf7YAzm1SwaXekxQNzNDoQnwp6NxEGBOkVt0Cudo
Z5QNBX7KJH3WZl+ehSB6zO9ftPWN2QCcXH1vG+Wbh8WvLUx0DtraI/lS39M3ERKr0Pugk6I1iBB5
hn4upLOPSnWdHgXLrYzYoL/aVVcU2T3ewvx0pchIU5IjwpHUKgPP5/wZRId0YAYwIvR6L4p4cZQq
/5DAYu65Ue4T+qejxvgpvGs7CwBblDV3dr6EBb+mwPjAIKzcMZ1U/ot/qqXvIAydmXxNOe0ACJwW
eSHCHKOAk5NpzuE0DP6eOfzHyRd0pDe1FNQlBTdYC0AWRgLvBbfSiFFTH+qscAZ6MUcWpeSdkGH9
bh+g+/wBtc3TW1SXw73PKJILzI3pLrTknPnVf+UFIj+oKGZa3W/Mrauqm/UjK2uiGF90B/SyisxN
cuNSFePT/Ry65XMcd1HQbT0/KKHhQpI/V7s4NTDn/i+lyqQFVYjxNNWFNHXzjPnTFPqCZLCmwjJa
UrGL7cHteDerN9k9+qfke6X6RCsu0OJ35nmeqi81IedWLC4BjM9zS8JkBXivBvpwkVY6hWZ3cSWt
xfj1IilZXeElqQNsQVyUfX1VwbpJy6ztkzQ4mibZTBX42AJWOYyyJoAbJgjwNiOc4K9CwFRYPHAK
zySFABAPJpLlYE14KRaCaBTK8l4NrsYSSrD+2YjyXPHmOe+dB63Q6KyxKF5LrSgd+OiIb6bFRbVW
3ph+vAkuTGPBVPDhG/fQpm1Qaq4LA18VSYfkt1EVkWEMl9QaUsuKVBufIevxq6ByiwHxhdyPO+O1
MZg004sAZL6uwL2ckUEzPWr2/oujtBfngnqJfhyDrz+ZlfDKGxHjrCTt70T+9OcDpcb+NZb7QjDP
sItjnNaFWtCoQ+ldO+qHFIUBFrKnooNu3SRL62oT/QnIEABcZfh+0E03Ask30kOfNyXVHIxpoSRc
l19/PY1Cj8sBMEV/MDCx1NvODjjYdyjybsA51w9BdsyfMLLOvi39rHez6msFFsXq6gNI8yBAn5qB
trKT6PeLWSwatJOUAhFHqDXbESS2/FYAZFCaR64ajK78YHMIpD3+pM97wa0wETz1GDR9f/p8+GNp
JalfLF/S3p4iFYnk07d9DBp9sKamNViJdqUgW5O41f95bNEK1Jx23aOUXb+hxZvN3FKOvEGEV3jD
+gLaQ/IbCwcOmo21RiaPLOVZ+6pdS0CaGfmg/KiIfSpgbdByxSE3sKYbiSukNnPTFxwPZiXffLb+
kA6TCVMpjiObJptBTgzdQBKTKZP/kEKUdt46YenmAP2IraUO6txbu5lx7fxeISfk9UEUr8t58X1c
taukqu+OR3K5KCMFqaohr+fThaA4DgLiggFqcj19l0l7TyDqlCLWADAggsZAZBqpgwqJTSSaNMTZ
lL/tBZqTRL0EpHBrxCfmt6Da7edjuCS1gLiF7/dHOF7U5kMnZy0TN+099ZDoz4lLz2q+muGHuKkU
7QhkjEH9Vhc4vyVjs+hxb+6AX5TjWRebwy8YIWdaH5DMxBuaGWUlHcJhoxXdTFg0xXpeSe+zLKQs
cDlx0kQ+uX47r2rrCeEWsnF5UtDCb5NUoOCaQQFO7OCexSUieK3Xq2ih8qRQSurFHE7ukVF+rEcW
U5B7/7XwflAYAkJv0hjgIMKQCKEvGVGADhH/D+zXafAiqEPkgMOaUgaxm2oRb7AyR+kvKuqrZFva
asKiZs4EZZAvgklTKcGtTTyjYGhfgG5ixy2+8mc4kjyHKDugq9ObcH2Qve/bYiDbMTBMDpOA/gne
jEECEmo+9UnKsLwiejiFRL6x/LuohFNqcPHX+UjOVqVT/Z4NAgNHiejpBNFPbFv5MkT6/yHTPAqM
2bNojgBx0NLDlyVl0+e7BOuIzsO9nQaqx/vxEcBofobVQl/Ct5JvIS+QzDucUXy/X8I7NuAfF1NJ
ne7CZSyV/9aDo7SVFiT/8D3+DLKZq4NfxVnaznAKXaVCtbLN2peDpYhcp9v5R4mB8kWvkX2O0BK4
ezkft5vxsuzRuoGmNs/OMG4uqRhkG+gtRiTpqinKDhrNBnTRDE8WuHe976p2lgbgyluTBsyeiK1r
SXZo59bJrZrPoJ4M32UHHB8jfQlDiZpkj17snfgiuCYdjUZ0JqK80FvCH2NuWtG/t4FaUmjp68jK
PjQruGBWMi+pa7nZFlbbApJWG6v0IARJB7heOkVU2u4i8V0mg1C+l+zANC6aeoQ5ljn08ElXQyjV
7imq//8DvZfld1koY3v70vHpM7Sed2AZmX+2DRMW3NEH0+B5NcUS0L9gxm/6FmBMDAxtXXOmrOF6
vPxB3HwUiEDKjJ+vuAzs7oKYXA/at/0gZXbC7AfnbnI5a3r9U6IOsHlk19s7XCUBE5l3xZA+S72w
WWCw1U7gJYT2wJZuPGp7TZV9QniZm4BZNYIdZzzZZj932wmSG/dtD78Zui3/f0Kd/5WAeikxHxhx
oG9LQc+0oBzY8AQi9gMiSW5JZoC1wVTqPY0Ls9aREBXjFY2uoWJRvQms9UrgzfMDCzfXr13F2cYx
CZzARXn808FQphyu9Em010pegWJGd3wVmNxbUPvx/tPUKjMSZDnAdxI3GirD70S4VVO+Yk2n+DWD
IYt5Ipfzi/Uc15KBuM433BW17zy4UcedpP+Hg0zCtactLJbPnRYrm8hkWuD7YyrpJVFt/mTWH5CO
j0sB/9h9dOor/8hSSS2TgNIJXE2S70mfkOsJdhBJDScBOaoRn+EKwQMgM2+zFssDYNI1FNXtp/ab
wDks+Bnpx3hSIeUlVt/SyKh31WmOG0AzQgmQCIUf2qaY4GlxZanDX2kA0UrNinxHRa3aSkCTy9UP
NWHFn2KZ/Wq00XkUhex9ADlN3M2AUxF17rfZ2AD8H8TyuVTI4Wk8EgWZh0reBTK8e+jdtstfWSiY
p/wtQUe8v8DJ6pvVZ35JFg10IcipUleT4j3TZ7juHrHRqd7cZftqndLqCfvAlLulHnnXmbsKPuqx
WIa2FhxhwHXOXckGlS1MerspZzIMFBVnwMwWUKpk8ZmqC5Q3mf1+8KYVQm2PUXxyTfUPqQJFO1hE
bZn8SxcgL0R6XmU8OkZ6fyu9AlWzZB8MiK2omzrq9USCYXp6R6rfN51tM12ELlDQoxbo7ctMplf7
Z0Mw56hWL9xhedw/FsRtKyBSGm7jUXhNmQz1aE4ZKxeYkO09bNGIkDuzfiZAw1lJuMY8Elh68+Z3
JqIoGi2YgRqCH6DB9MbcVLPSX5NT3eu5gXYW3g10KaaL5xgbYyZfjN1CrcZ7jG1a+lp2lP2v7aay
Wqo0+K8HyqwrIMe+jBa3EoNzGtkk8dvQQ9HH/M3PwOIG49Cohffr7omHG6xyU5zZuD/qhGS0D9Rn
9I8pDXAEO0XW9Q9ncLmyG99tONAQkfo4n2xDXFA33C9dlc+vdiOhsdPIBkkb5y2y5nwpbpAaMKCs
IcwUkCnA8/wILVlfzm0bob59PINK6Am6SeSiNhqU+k+HKW9faO7OuUfcrbu71I8Ssk4U1pwMksl0
nO+e9jq1I4hzNHrUe060N50YZZyCutGY7qlxWRoLVwMjQCQXVeRxsz9XcGYVAWQ8S0TStXKjaD5n
JUq6aTgHYr5ElwsGFcwjtMANdNtbJISpL6bTDfVSZiatiwKCsdvpbm5J78rKFvIzI1Vc6wJNm5qy
wEuNUnL0DfyP+dWUcc9wcyzsm25YkQlOeDJHl40yx6xUgeY4qWDqdKyKVLKOwITibdCboE6Jsye4
JzpW/FUgUoBy82TgjqNZzAh+nW6m2EXZ3Fue/XJl2meL2R/rvYNDhjlegL+Bx9vO8QQPkGd/RVE+
zrtG1TEiQ2PGzq5zD/Ti2FLrKr/reg0LDjGWFJec7SVExsE22gIFAcuc3SIMvwfdsnlvJU1xLy0w
w9gqgUMwvlw7qIsTXmINeVk2xqBn4aIpwbtr4jv2Dxmq1/pO22z5H8WjdlUNxeHWkvmIS7IDtCZb
uQxgMd9sJl1kMjg3tEAudd6LMk6jZMAphg8BEu5njTA9tW2OE5ZsMxSCheM+i4NPiLeeBI9Xl4H1
P2xEQTQaJRPscj94mpiBPS4VnErkSBNoUoW9l/CQmceQGiY/y2x4nJS4mb4UCpMddStMG+ipAOSG
VdT8Rq2mgDzdyz3bZacDrJxcc30XodiyUAvwXoJkW1bqvBaqyk22uoY9y42aJWsEh+9av6+eVRa9
Rs1cjuVMCneMEUuFiO9k4xUrcGyTxZ/SVXLTuGeH6DZzvqiPrziLgCVcil/7ulqTImOL+BnqT+dr
L0Dk2oAYQs5XTPLH5EUzIkGBj/d8uJp3Utq6mq0hdIfMm3nUxQgnEPDohswvHjUnGJa72zE2RA3V
rMou1p1Xh/2Blg4cHM9iWHshBmC6S5l1suyWAq7T+Lw5LqtduGt2y/tU6eJNREAVNqSFMsyft8zL
U98wrhR58e7SEIkP1DnyHTJTqw7xNoVYb7LE3reRRpoXka223ZieDIs+QadI29heoJldulxoIBDV
XWi/kHPyrg5aDgxVmH6qF1xoyaAZf5GaVS84Xqq0a8m2WoQ3rzVckeppNhMgt4cPwtDngFkWc998
d1IuSe5ky70piFoelJkhFB9qOVEPXsYKj8S8EdpKgxR5Dmmc8eZVyaCite6GiqkXxGefOWPX1YPm
QBypFstz+aGzVzuXWdonLOCRfNPLMnBKO5425JvbIqfJEIECMtx+tFjzpu0+xd4dnXpsp1nW+N5v
WXrFOFUyL01Bcq5gB9PcmL4Ty8fL6Wpby1WT4C4aI1QukjJaYMkSh3WYyLNq9HSlABMVwXwZJgtG
cfR4lQnlxpkbuf5uM0JzSGjFHF+In5R+izoAOQC+/IhQCD5gVWUyPgGK2TUOPq/O5QPzhgwAnX9d
sAVWH8fK17GfwHLKjFFqMGtLxFfmrQEsAROeyVEyUO+xzwJH4mxwg6lLTyiXkboV3KjWjhjR+brD
bomXu3V187WuavWWhBbejA3JdfAcaoxli1Xor9ELMEHvKe56UBe86Xh0qWyuCOO5aLC9vtUU8DBV
W/5fZ9neo7LYm8auZd9ry8hWslMya/VPCuB3DPEBweV8PmWsLUOgUIvgE4+eArYT6MNwLAi3oRaw
vJCNuIscB2b2kaWYP51lR5QRHdGlydu1BKmbFyp1P04U864beioPMBMuWUO9XQBmi8GxDEc55Eg9
8vsuHYZ2pIiMf8NtmXL8ETSaHMX/otpDgrlJDtpqqN6+NjqkhMUE+gLjEkurmU5PyqRkS8vzdOU9
YYbgcnwwtZjW833zadGFVE6ZgtcDcLkcGBSgbs2u3agnqSsFybEqUyakBOh8dFmMCVy6qF1f2USZ
HL/HIgTrMYK+OKSWEktjlRBFTIGSYViLUctsYwrf6dP++fGnpcpPihxmowHofyz5uwrHJNFFKyYo
+QGpSZ9EeJev3zOMZc3ivzwF4ldaiLMC5HRJLt+oklo7ad58lTXNZC7j0DsBQedrSkuTx5RP6caj
w96iH2SGn/MX5ftDGIlfCOVrqKbZsubdIP0nxYYMUfJJ8XwZZD1P67kt0L7M9zA4JGxpcwvhzWBR
oY72+evDUKqJ0WLzeuG5rPWHXqXw5BiiIIlbchlBNFWCj/Ua6JvUkm2lHbYv519hqTL8gdz6+/5v
5+euC1+6csyot+N1rQ+ugXVTWbIFbqSy1xzXZrkBnwgNe1lmy0G30y0v3POpPGBwQnCaAJwoPyUL
iEQLshjAPkmYOGF09uMgJNtJLi709SmDrjKoeI3Cj7ELJ647k/PklCVFWr8H3hk/48uLWoTtex0e
/cVY6TKDPGfwaE8yx1zuhxsdy7Jw7Ly6fl53j8wgEvrwuJDPHwEPkxVuzr37OlnV5NXu8dOO8h+p
CF+LIKd6Grqz4YJ8rjGe8vGRjFVfVTvlD0ePSsTKuR5CyqXQ9V7zrdBaGLa/CowjueKjfPD7485y
YGMHlTB6KKFExrFFWxu9QrAYfnutjdQbX3H/NQiOPSNTCqWv0eqDhHB+FbYVz7Fiyfw8nUtuvFFC
dk0wQ7HPHBZJfguxqRGcnZDXw6J3cDeu3HQEOx90bwhePDvBkns1n3OYgIzKnG87SZsJUu64YIOB
o1sdl/+/sDeasKDcC58EWr8w3mZ4unJ4fT3XeCqTcy/sBhQ9/yhgOoGvWlYOT3nprkHeLVWv7ZI4
tM5zmXgFspxWE89agtJl8cgGKTsrI50nawj6KH2GheSlx0DJ3LfBibn2UUsJeXTsBof7Fumw9yQx
J3kgyRIIewgj5uGvCUAfPbAsMJKF4adyOCKtoqqtvLtvWhvqM+aKukR55ExxLceeRndn+fyuLj9o
GuGind4fbS6bZuQnOKjveCv/4uGlvDHDGRPeqkIAdQFN/618RQmYWyL8uxWGBtAIYQ0nvwE7SnJB
UrK79VNPNGDdBr0tMsozHIK4veAsmpzbOSXOe+myQH/xNkQUY2KzdgrugGfX0DENihR8Wp+ysaHS
d5vxrZMCCfj3MsRb5K82AXvt1nqROUpyJkLyeZSEc1nSIWyF7nhhsUb7e9uXu7T7+pf+/pdW21i/
sh2g9nlR7sCzQ0+bQUuZsoAzmwg+SlmaASCjtjqH4gYpcgHrgSpwUifOcFaRVsEky8wwE5eSEtF7
ztpc1scqFVPb0bIiSokf9/LV8VibXXTVs7CsnyW1edCU4OTOzZBlM/3R17W1CPylmsny9C6IeZk4
lEqkmE5h5hz+pFObuzgR0Tcx/VZpT+v9ii4AHL81UhpJZqZ3OBI53ZuuruytatT2rZx99Me/fXsW
CFGSEjtvofKIGyeBgIO34CL8XrRiWbmk9Vfh7vipLlkTU9QR+VrWJSm6TlTp8sB5N8aVyLCYAYQr
NreyfSnpePHUvXLzY5YO+J2c3gFcljragGF69J/pj+XUMkxfsQyN1AYA9Zc6lHoRoFF/r+SANZBZ
xky99jzifT6inElCJe3s5sDUmlIWFQ5OFkjicry4volInkOoE5gOurJwuT49kgvcnhDPIgrDD/UY
d1o/ihRojK3TcqJ5m2u8M0LYJDJtFcS+VGypF3uHO81bT+FxRsIhpUGKLB6eUVOKt30jzj+dmVZI
xJQaqVRXwdX4BDHeIogycGsI8oHbj8hLTubuGM7eYrM9ncj/YfvW702U58frLG1ynl7h8YY0WfpG
8MAVFLle7IsWiesykDBTHrnqhXaggXgjtcxdco48t+um/Apl4CvuFEKLvluofDUbsyaCprIwSgFR
vE/WX425f9GgeztmjzT4svx+e1QxTEoCdlJhlMqodlR3OiPeQLCWw5USoJhxu3LY7hYEv8Ur0zRF
DlSmstUoORe/+vXO1L4ubZAli7uiKWpvE1w7JamKLowf3idUQgWS0RDK7aZtEYPyUqK3IyCKC8sD
qCtuFk6xi/NJ0ADpK771fKffU4UgmQNd4VjDsxfbD3V+Y1iPE4Yz/e3dK6f38jqyYz9QevlW/MFB
r//yIRGumSVIM9eWGNEPuc7cRkZKcM42CkMXaAaMlQURMn7UEo1Q+VrKn2Ycy11kJd8bMrtANUV/
WK0rTTMBahcRSEqhD4l6vsxcTRygKkCsjyKHLerbjjU8oiorxBW7zQ26yspCSfcmOeLhbguoK/QU
HmT8OMeuQ/VyXVOrIkcZgy7+ZenLdYObPFKeWg3L5tunKJJHQWQah1RPWUrkJzxC1cDzyoTvF/Ol
rT2XmH4/RBQAj7QUSF+NiqR9CQ7MiS4t+jyP+9eD81wSh0z04dOB1w3FZcaxwiMYj3ooIt30lxoZ
o7zGGLPXhbI03f2Hl8pr4mv7H0X9KaSVnsxn+M0eoGDdOCFTm3oZ/Ya9OMCV9yetx7+0+RauSASX
/9jZRYtPwa0JbwNgG0PvwWxxJfB5XFeyUPqSOVIrhzhC9kAsDfuUJAKpm0ks21z6rM9oJvNN4HzP
qgmxBnV37h/zM1GLns/v/noBF5LyHRZ6f135u933oUftYjC1Wvia2fHp2m61RtyhbEiYfsjUYON6
1/2M41LMhYWnh5EJDOkGXjZjzJrJ/BQDmURGy/bP46MtsOq0KZXnfFaHpiSxNCW3MTJL649EOmVc
iBNT06I3Uoo1ODOIeJb5dnhBaTOT6yoXAzmtD+2dD26gaE2if2xFC7HKklaBRBOB8cDkzlADCVrw
bfKBMA8HtYj5byCAtFwNfGIj0H8xU//6jwgtCL1IclS69tWJIp8WB0neewKe/U2BVQrRWhx3fxiq
msow6N4KFFCGCrx3rlOEO0ldkFPp++IJ4GgfBfkloGmz+97KfWdvWtmPC6Mingj5R0qTqX4SVmn9
hqFmDhuGQu6jp/lXtikeh9XM6F8X/ZtxSYDta4IP75BCE9o9cVIHzvZap/XOGouUi/dLnhLFhNHr
FvnwHvneaNcu/y8Jhv6Ema78qe5PeWUDOsH+VPpaTJzMLz2iNy+rESl8/0Gb4zAjYxNXug0Lgba/
RuZTrc4Odq56hzEh0vyUc0Ry8RygHfWc4/weEnZ/MPb6NjkortBslbkZMCfKj2Ri1RHOXigqADZW
deBTySiurPZ4v9PEM1gCj6wVZtnrkVLle2ttCKXqICKD/w+SKlsSW0yXdd4yuG138ElpALVPmN9I
eehN1oK6fB6jxX9INsm/0L3im30GNur4dQzt99pVaCa1N0LKbtGJcmKn+vxdKz2VEzjD4wqQ2kw4
OichORlb7fFH8hw4gby+WXmmqj1pr2/oWt2Zzq1TxKVj/DIArZQi01uaFeJ0N1cqGtMxqJCu4KIb
Sl/YvOLbFsI+mu6dxXVu/9p5TIh1BCw/ydagcLWov6XAjvL2ECmNvyrFh9hfU7kDQ7wlzcqNIfxJ
oDhqP7+wnWUjYhjS7cRYewf7Ryj3ZIN6S1atqHL4K/YCxTVFUqHL0E1FbyfxSsmRIU6pz++9nWXX
jqLorW87t5+Z65Ua1P9KfIW7HP4Y7YKkLFgitWStxUFR5cK8L216adzVy140Yhb45xwJmLf6hJ8K
PgLaEeq/PTMqwtKFRN0tj8bZdngDp2+nj0rKR7rdOZPdRLJfx0gEbtfZ2Mr63szSdyvS6jGi0PgH
GP0LKrFyCw5jOGoHUxMqV2aBDTMKMWY5Xn8vAvu4FEh6RyUl8kSIVXd97wTrZULF4h35jeqxbxXZ
CRsAzNNlHgc/0oCucotyJPkSspSWhcdD9Rl9hfKDoS3BT/Gttc7EwVnti+vGFZ+aIZm0+upFUPR5
NksmGi8taIEwfqyHtXmU1NWFawMJA5cPfBaGmKWaW8W9S539qY3h0WhkSSPNhYF8P8v2XZTnlHAP
JyzcWhi+BhYY7WVkX04yGUJ8XX5gB2Rou1EoQQop0buB+ZFQOevpLZD30EDKUnXwu7fXIinftrqJ
TR+d6h1Go08lWCWO/IBiCA2JwYtCG2i7OG31vczVvQZSL5dJNVEH+jHXUTk2QZU/mxP5lHOBS/We
ye8fE+lwQw/sUYpINJ7MO7FXOeSDKPD/HqmhGg8YRMM+infu/mxqiNXHMs8s74LQe4LYEyQ5BeEK
SZmxeMXaME2c+u7ZbR519a4MQCsOhjeslTMlFk9HOJ7S71FXuIYfiVgD5WEHSx395ImKf9IPsaHx
cwQ7lge6j5GwvWhV1VuYBvyJWT1Ay4/P169XJjv3stH1mZSP4tiHAo81w5YHmDNpq2xPrx/0NbG5
cxQ03qGHXy5IK0K0LIEpxHD1oi/jvynIhyiR5ITTN+Vh8xz7PTKNZotdcK+gLSDpnY4gSBTGxfvM
75OgEPkX8l57LONzhQQs85sr5pdy4Xa0RUPcU5/4zMGH9kTVOfynbTWXJDmgHHLa9Npgwu+Fvqqa
lytDVSq8haxl2Zmh+0h0AwJd1vFBMngu20oW1x2VuIqUxcMdCcgqiIrD18CBEJCg+bt5qLiMk8ae
MQQRRYb4Vk60dNp3Yn2JAkib/wBIJiKPP4S/kmBPSWJDudU2ax6YoBdqJgD6SZXG+DBMJ9SQFtmv
eoX/2c74cFCxd28nV2rosCxREmYI98iwVekZ8QX/BlbqpyR5QzDssJjlbgZiYa2ZirNHK79G6LBq
DYq9xN44f+9jcdI39V6yWKIjsgM5yxBemlKDDbkmbN+5WG1wk1r80DstjYy+ZXFItSG0MLuZGBE6
fheTSRa0e23S9W/AvDSmHDZM5zM30BmDv711ikMwdLc7wmJ5a7BA0d81otvtLBSZYKyyKvn9sNn4
QJPbN2TcSMRpAghDulCkM+LiM7aqgik4yrTksgDCrd9P7UVQjs7C3E23kdzQd9yj+v5qPKzhTTmm
8jJsQ/i9ckygxrWdCtvl/KJcHxUOaeNjsiuX+QmBlCv9JK4ww6+g3hCEs06D8NOh5oX+ZRkfC4dB
mw4HLMeFZCnmg+z9rhwRxTZsNM7PqJPa4yMJUlQVVWxI+EJSXJ2VyozUGLP6k3+sjP7cDPl2G4v3
Z4T29hbBlTN3iNexnwRow0xrVsrr0R/Rx7b8HcFUmmsAhFCMyWt7MCctsFb3haT01SD94wLjAUDV
eQ0TFDHjqmRgaqQ+UNs93oPhu4lCrMeS+C80gwKMFH9/SGKJJ/mezAjVrez9gIEoJX+QEdF/hbwn
CmzGvr2OMibpKbiDav8W5IzQOWrGSYf4LIapSN9aGEg+ZkwML49SlJsXzgSpluyIpA6W9Dd3gKcf
iCKoBlcPRBOB/0NPzv0zHtxhB0aKyeG8ITxfkmkH6DwckM0pbClkT6iL95z8zJkhiZJVPDLsw8JW
SDoCVmz0NkM85xt4+ELtj4+5gAPK/PpyJxcp/5Uo+9ZAHKM/dL18jCvTIeylODkHPje7NTUlA46k
RkajAfKJvWUHBzfYXb3JvtyPd4K2vJlDmvluDe5jpfpgnFydLiPv7Ch/MrM2CNQq45YUCYiXX+Fa
0dluXqG+kn34PZ5qdbU7oLirn+MjjruEEiH/UgTptOiksjPr//pME4qef5HljPdnP37LAj1MWl67
6rwKZ256H9d1Xyo6SpfGT6vPwXUohVyUgNKJBnOJiXRve5iFoN+b/vxYaXCqd1yOX/jUl8zM5KAT
EqijZ5uRhp4qj1nUUUZQenC+k67Nc9JLcY542bb/qshu/DvubEoDEluH2jZVQBf+n/gQW1uKean5
XrTCo3RueYGXPDIP1P7/13caHKiey9ulxER7lQt7pq63miIL5iH8w976K4Gz4qjMWZWs9U0jBO/k
+fY/r3NDvbgES9d4r88cFBOxqxFhIx6o6MWnIq0ZeuE9odIkz6cdslrgfSW2efrCx6xYCRUAJNeG
hq+XNZNlu4gnSENnjZxR4LPR9MTWL2cVsklskjcL9/uxaWaCfgFrXABfendbo/Ud4+R1c3r3L1Ae
4kHe2wPha61y1wur8IceF9f1RC5bsAAwWV9EAprh1ddOMq75QTr4DygTOrFw1AaEQhf4oFkyqKqT
RWEqgLv7gEGpqrZ8ikxtSsC/UDl8psW8l/zttDzuLaLoHkxVK+72drmHSN8wICEI9D3T1lC7xN7o
5nDO5zaU7uY3IoXKdWHz+wokYfjnA7gVx8CYkX0tS5juEbn7lIgMJs8A5lIE4PZV0vYZtJWI9p9w
tkylRsK/7NKlACUYb08drmFCIfmcYx8q3s0tz+EisgmHVrAB6NfeDOcH8m1Ud3QPwZBsyOnvcRmw
2FBnmZ2gJZaJ/MCi/DiVI3gScTgDyxz1bzdQelfUQq2CE14JHxWRd5gzoII/04rRxl3Vgka0lTg+
BBqN45RkKK71J4d8t/aUpXFcbJlRlexnEXAQvdmANZHPJTuIfRk/y5KIV3XVKWKq2X2ZZvtLeVir
rnZ5Hwwz/6H1FzsGS3RSZnrobciVTo01O6yWpygYWchdocq9kcC6yz/XV4sVpjp5shwqzc4WTLFi
ZLg7SmqQ94RhOq1ydaPCA+0tpUhcWLxjdkMwAP9JkuuhGZDl3ANc8/Xf8ChUnruFMWQxSAhfe/Nz
3ufBwVU1vqrvRowbQY8kiWnPdCruSTS7eVSAD6Vby1GxPsalOu7BBDQWQvuaF1Mp2viiwV+x45BE
HoYqjqVZa7ouaeOKnytD69Tj3xNnp4e7w4EF9Tx+D0tma+tp2pin3sTBurJgO03z7G6pDMNG8hxT
3z63V6+6elb0U2ENydSKKzPggmBOP+WqGtG/sYv//LB10VlpknctmxUv98FbGpvaGbWw6rhjgjqn
3RoZhvoWJgCDuoXBWomlaALfAoya479kPNA/c8ietswpHr+BPFOhNF1HixE9hlPijodufwoCIijI
pZYtmdPUeKELqa56eUp8UuAqkG94/HYqQijM5L6XlVMgfOengAvYG6WQR/b/s1Cls9Fk9mFhdJrR
SR+LcTktvyZ5RjvJWAdkzaBtk5dM80vWUoOwu+vCcddCG5bL6GZm89e7z3IzpmUsgALj4vnkkMPw
cBFclTtGDvllE2qxIOP2BxcTVJgQRs/LFpcYQb0DECm/HgPlflnd3/50ubqmCVQsWHnrCCMvYpSJ
0ThICWAl/Qc2Ed4YVklqbnizI6rKZHkUA1koTX5DEFCd1TUgROsMQMAL0Xt7ywVBDzN1uZpuFd0q
vmhlw2xYHw+vYCoPeTUrQzcRNtoROC3dlZmtSLSWSs/Lo1c2MWOgo8qWd/MQaeEEcVcZud9HVlK6
XOsvvdBa/H3KcItM2XXUynqpG9gqxonyZfCn3OXTV0w6wWsiqEnlnMedZwiicjfb7JV3Tsr5taHf
PJ5juvMFDPv9xIKaVEN+5PA5p2qsccK52ug0YHlKkGQaUB8w1EwWem4R+f9L3ZBIeBN1dHJi2Mv3
2qWz+r6L8oX980GLm02eAMmbOmBZD1mdQ1jNHJFYrXMFTOIB2d2sFNGGA9jBMR2ErGMN/wNgr0NI
sUoNArv0jQb+M+S2EA5qQDYluUUo30QySrgy/NzfFrLUhPI8lQJxkVVQX1zlKJ6RCq25lgpQPQUE
z/EAe96FCAV1m556kKQz4bmNV0ZUvS/6tT8q0FQwLUFK/zZpdiTCFXrOasakH9Pkx5ImQcxrAuaj
sI77KK8pkOKw7jTbe+3fQEm/4vkI3JJmTCwVxNzbSS14mXnf3FVqzscj47cLzXSspZqMfalZ+UVV
yj6AotRh1FU/RoCXj+OpIOoj/qF/1bj/5U5smXhzwVeikZm6Esp4HlbujXNE2Vj+Ue6qBiiXItaT
AkqH+9BoT7Btx2lePG+1uULu2tly6fqXA4LqRvKdkoSt6bUyXIUwPVGLzx4UjGLsSLesVdxxPLkU
ETLwlrualpw8t4p8Np4xtH7JtECGu/gkxT4ItcxAPY8v3FSLfkJcEmHrHa1Z+vtxPOdRJYjJGDld
MdI0jbAnlI0tFCHWsAJdyAL+msHYveM1f1PQponSURKB7CDr6iZEmVAKBE6hjmae/g0eaezunke9
8fMRfB/3sOAFLipyyHwzOIXuzlf7uxXM79K/9OPkeehXBHbS5aqn4iRo+hB16b18fCKsz69vC0uf
vFRbGjDeSlbd1aBckMhqW9aYj/JIcJ1V4BGQUa3/9ErYUxlmlUuyQZPEhuH5Ob8PhrL5Yk6fHQM6
vz4V9bgoPiUUiQXfMK/OOH1G9KwGQ6pPNGlpee9WERThcwX5eiHOLnuFj5WaGJMOH5mNsGesRc7M
ate7NPcwPS4U4YCloDHrWDOmD7Uyx6I8gJ+4Qhv60NsJ3cAeULyA4lLBnbb3fpbR5xyHsLsEylv/
STe2f9KhwxJMekVUQNm8yry9768ttmGxKfYHbfE7KuC5ExkaRUracOopNsXl4nYG1NTHPFkavH5k
9BLBpxBvyyWFUPL4wTe6qZlxMDf+0/ynjDTVsAWsSRmtkYjyHiUu1sARqBko/XIP2PIDbeEiwqRl
4aGBfLPsXC2+aCqMTebbcFiMr6dltnGGHjky2Vp3BznSskG6sH3MFia8nMK+QwGIrk9obyFVPh7f
GydkZ/ngKr5NgHoooxfj6G1sMHSL118tjTNDTMWxsPBgYe/sU7AGL09NHIzAzuhmdaxbBPnSDBQE
jo52c0e3hgi5out9CE9jK+DKBsufk+Eq5khd/6IjIeJFBrov9TJW0sy8dxW1KvGlHWdlyGa8Pvkz
VNov3mnx5SFb9aS7b6VYbvukIQO3YxAvqawa/K0ikRUf0zxkvhFqGOjaTvnizXaGHh/zZbLOysxw
rLgQE7l5EI0tovtCorV8v27fBhDD6pR3n3kZSkv1RYcgfSPhnGdPskic3v+eMSHhw8bEQic0MyCM
K/OTIbR7GUWg5tLcd+RzsKFhphB8xXtieuWywUJzexkDwbQUklyVlwFePGuOnQC9diXQOtuEfSXW
Fz/Yl9YKx8/zoRAyM5WSd0PPk/5uwofdf7USRzgbVE09X1sO8OjSlkObt1EyLUgh1J0QiO+9nqam
mmHUMNDg1F97FPj7zRF6s4RFLTDEbfx/Ji6qPxDCKb4oGgXDqadAeYftf1yvvmazMb3LhBMetzuV
flGzkDeuqCVY0586rPV3F7wxOD6EnyroNpiyOmc8y/reJheY0yqi7iCyo8K0uyWVSYcmOI0bgr9Z
AZQ63yP3Qgm+UG4YR6wUDG3Nq2lyWJS801eUG+qVTpdLRXSZBG8MyuWSaQuResHI/0docyxw9+nd
e0qybGO/DHpt7XWQcWI0kFf0QnvGGwACgopjIDLNKbpuMMgbIWN1jsouP2bTzrsZaycpyhjfIQ0i
9uDSvQsNok4pCItBN3Kpq1Zq4Gqv+sR+CmRru22imNhGOSu+oFfTtIONJc10WBJyD6xss1ILxv2o
6CKiPDgGrjPl+Gv9rH9itRfasjvJ0V6yF/1dVlH85aHMOs7QGSxhiiW8TwwF4bOqVxIdUGNftv1g
02xgdKQXuPWJnz0YpdiyL10dzpLQOVeQN2I73ADbtFAMVTX3CE7jM4Ujd9muIU4ZlhBIV2CUnN7i
DOsqnTCJk4h2tve/pdI65fPOXhy62T6PabH+ATyP0B1irY1cMaAWFEsDQ0Njbh4/sHLjPHk1iDOw
X/DfVc8FAAebUN52eWFDc2mC0mITZQIQRCu7vw7XJSA2IwXmHiR1Udow/qUwf+Me79H2sAGlrlBD
xyzIaFLF9bg0MAhEepkUngqMW4MQVU5m7cD2nfJmsBtugXqbWAfuINTgDyr81qJCS1Jkc50M/3fC
iPE0UwIxXP/0aVXyQGfgSo5fA55Pf65I+ukbPo1tJc/abiB5L07sn6BMnw68IA61SgbFp12Nmm9y
WFriN9aruHxX2aJDkxX4z+LeyiDsAmSETqSQaZZ+FdHKjUJXNGMs6VETf2zYf4258i6dyzfhNkKg
dYiTjID6K7pvm0MbZl2q5ZB28lvxqTgUrwsLUwlYHlSVM1/4eqP6tsApYno2oRj1sNwtUCzIQxV3
34cAffe1L8A1cbPLhzx0sJk4WgzL6LKV70UmONgbFq3IT0AN9VStaVhiLya+r+ZReFxtOGowOXzC
/DxtpomdYoJB3aEGW3zfJp5NnqFIOvbXgjaG7vRSQrlsdVLfL3GgASoo9ZmR8WFPU6iGGNbL0a7v
iw0f1em7ldAPC4ABaRLyo14hjU3sTyTG92arx1DFIBOhvrd8NTqLJwXZ8QKSU8AXJHx/lv+NO4WJ
IEXKhYecPzh+O6JiZwelInubL8xDYJLdc5tPiQQ6Hzt8/nEfQ1NILDPlXUjvz5oN7VJyQMNpisjY
TlLOuf7XIWpZj0t24nhf4i0Ul0tnicAlWz/F2kjEOwaTQeUmhKYOyRFmuprZdFhqOseZv+vFDrU1
ss7/8P/tTUr7nmehbkJtK2qw7qoBwL7IcK0VHaV95FaYBNy3dLvSSf7+KYx88ja/GJQg2Rl5xVPm
Rvxah3qe21ctlXjvnw2L3x73mvsfEaUQJAQzHJjk+gT5R5j6ja+pGC+5H/rC7rQ+BN8SjZCDHK5K
WL/6gQMMjv8AfRnfjg+q33ZSt4hu2cR6c9p8nY84asjtgksWnT1qJ+ZWx66QpV1eg50k3S93Sr8t
8PT4GrmCPP7Jzl2TmdaZzce9G2G2z/DDLFA3cWoN1Ml/3XYLaVVvpzve9uCXKBnrKnphn4mcfXyt
DRszuavaIQGuTWpSrJDPWA8vvrxRhHgCaAFi1jRtV6qma+Hsf+fnlJ62sZF2axGksYW/dk+YBQ4e
o7mYUQ1K57WnaqIfH4JoxPHQws2uzMnPbXF7BJ9IyT+wF74GuHwaHL6Ov3sLYrLPj1BeTA18xzaA
omX+/y3ObzWCqz1Ls4SQ5xBXLYIXD/589IJLnnl9fAIaUoXwmH55Z2tshDw3wMGo0K+KOoOi6z/i
D9+bGmizwBgMEQZFrHU65rzMAKq+7sDanDlEQmqxU79u/b9egc7oO6RCJgPQtmnn78NI0Q2n8wA5
lIqsRPBnVtoIbk9+3egkn1eMxZsjJJLxCsFaIrsobuLHppZzlexx/PM/4F21QsfhUhaPuSXrlFZI
qoiNTG52EToYErvki+aXfcAUsG1IcB9TiBPCfqePZ6o42RC54Ub0FwEhBXYr2rZNPOsOqiRUxFmZ
dFUmUnS42ln83lYwhPDfNBDsfC0gxc4bIsUOyfJgk39alNKvIDV+CRu4k68tMpWc+wHpdG/wFDfl
LnTBQ2iyYD9sfgO0snYhfXuJ6LnNjr4LEE47WFC9Oqn9UI9tHpMY4Ic2e1VM6e9YCxMe55+Yd7vU
1chhsxZuKfSX5Eiyrzwchkc5B6iUPECbUCmDHrFvWgt0zTHKDc5eHA/isIslHgIeRn0iovGhuuJi
Ld4dIY0bvKYsXGh1XCCIh5GLNYGEpfbiDPy7VWJ0velc1Wz4CCFZRnFqpqq6BXzwpPYF68w18/06
LCQJBDQcL63caAOMPkeDGjnOrNkG72htRVI2irKo0epKmf55a8qnATZA32r6xzzoBvPHEWABSDwB
t/pxzz5ocZUk17SjYbPRE4oJ8njvybd4sGo0I/BuFR9BpMwM2IYI9uwUDtrYPuaJZrmq3xt8DPFL
nLcFcXczybHvUQRWMwtR+4Bb3MOI+6Cz8M/Im+64XHm9oH0qWiZ+H01cCsCnHzQ/mGXwIUM73p9o
4Wdj3xefyhfug+X634aQD+YRNKQ/VzOk7JbpMAgJW4YC4St09yLetlJ8nnRIj5wbth+9LRA4Ya8H
PYgUXEeA72LqSZ9uDZVpJUBvDbPuJKz8oGlccHYiADr5jh24hJGQ7naJ+vigA+mxWKrmd4YgdSML
sbSUmtwtrhDb7d/GcgLWjac9eoFdruwGTz3cK24UjB7Wr+czE+LGxqK1Hs/QP0/MMaOiR/VvNXTm
BV6tZgW+1gqlVymxC4S8oUaDpS01+eFdmt1FNpVy0X7VHeA2K5YuM72zxUt8um3oASy76KhagXx3
ktmn73DSa2ZsBB4IMFcsXLehK2HYM2rqHJgLhbub1cUXdtn9pvRZZwwKbG4FKmCJRoF4NDDpDR/z
9RGB3oC+7au52LhP8eTxNafs8C/0gjsBxSzRsDp7ay4FRitX52Xd+W/Z4LiZwfCc4kjx8BDyfRnG
qoxsfuKQ4rkYOG07NdPCasWtelD8M0XUbDlEA53F21cwoyRZ0h44OyCZlSgDgoaAW9zTpDn6+a1H
2W4JhgM9NFLX0cJKcI4rXMxGHSIZ0aTDc2LcsQB/LCI+yGkoScRqmqEFT7KtbRlZhL+c85m05Wdf
RZAewdxyLMAc1Ni/dmRstcb9Um4FpFM+7wQWqmFqjMgf8+I0bu4VbeBajPu69W/5x7grfKgt/uKk
8xudoc3pJiguidnCbtKbVPPGpg/f0hvKwvwYWh7DKhAcEQzBwi8WT/m99xaXdcXdo+vGvzcuRAyt
ZKaHZGXB04aeX6+3ut+FSBXn5bwXlROcIvZzYWDYjTSZhs7wJ/Qu1KAKz3whn1mvnjkj3qeFRqq+
cDbRoEMkOO7piBSqKt5lI1BCAk/v/C1N6F6SXLCYe0lipX/L9LGyJt5FUWKh1LpEUUYI5AMI+7Tj
oVvrZB/JecgXgOwMo1FPYYwCoGajbOmY6HbRXJJR0tWWHtpaK1pgkq0qoEcrltPVH2qCK3haX7xO
qFZwomy8fYdmxGaXizLNnO5fD52qafuTQBaWMnb1X0I0mkNqq40FVlAVif1Zn8RI0CMMO92Kmx1n
DVc/ijnEWvXDXaulI1N9EHZYMEyeNnZO7mylW9HRQUdF+mnMXagjWr2UDRYD6vMjPM26QlyF4yWw
H7W6INJUkUBSXENIkOi0sESG1Nv4M8+gqiidPqrr/PxVvYwf2eX/31EN9AZwPZnLpI4eyUoUtruR
LkwNX2c74fX5uoeVUNXlDBe2eFhE+KuXTVzW7uAdrNsxGl6oMtJdzSi0QV4UPPYvUlYdjdBwoP9K
AKiddReTcbua15q0N3MWL08jtJNgli1DXqfi9ogdd6jVPBp+Z00+mG5+6ejqsxLuyhIqnBy4aMk7
DlqdSPikT8XS/RsKPEJ6Ajc2Cw9zSMc6wLWXMkYJYL/TG/tzH3QU2ctrpm+fJjEL4g3Z4YF+nGqU
Rm8eEGaN7t0vSHcL5BcRonanp8gH4V7fhYbJEHYA/rtQuFOKi9XeGMmgWoi7gxyb+CuboC4FVnv+
EDY3H41Lnk7weoFmfjYK6EzNReWXdlv0UcT5q/Qf1H5NHDDDnGn3o6xFxfJlXj6T4R5U5q1DrN5N
f1S5heh/U3OESUbq0oi5gPbJ7Feo/QN4YqECVyYBPFVH1b5LKYx78LH9FInfJljpfzUqjnGgbBmh
qUxvvrEDjYF5Ny7X9gxunrjBS7MTFHZMjz9Cg7yYw3AbTQsYL2d37I1oQxgOMMsoo+m05XP9YhxA
HOlL0DKYmGuh8gU1C2gaLv+06r7Lob41HV+oabzDeStJzwfP1xO2G+CAurxx9Oez11UWX3vFe9kH
aku691VZkIsElRWIItMmGUe4rQn/gMNmnwsehq77ru8VgPWmBcXhwrfLSAGTqeSN1Fqlslup0FCF
ZmJ2DfF5HpUl+dbhtJI0G798yMsYSjnkyiwTSmsxAnH5ldvib1gRYnOaW+sDm7jvlZQ5bm7UzD83
FHks4tFCdYRYpgB1ZuFIiHiEsDklvKTNQf85PYB6mz75AtaYJZt/Y6u0zx8Xu8Wy3EtmkjBTyVS8
9jnY6RkwIH0b2Yc/uaJN2bK7cMszsLe/vkIV58Cj7fGj3C5sw4pa+mQ/mYhzMZI+D6d9FFL1X3Q6
9PJ1m22Om1sC6DfoFUPf92IRFd6WGiL7kk/htI33dArx3mAjHqnJxYbIcSX+7d1lzxSTHkzp5Cmx
FLiJY6rShnOyJgHUSAEEMfuLiW63yB3L22caXP5xfnLQHO7gyvUACXpSUnFvrayCXjDD69s3bzQG
8VHSGbGzJA5fxaneO1u/dGa2uNYLGp/PPCJ+jRz0KFM+mu73Qwf7fiB1QcQjk1g2xEQt9RitGCyZ
Um226fjY1OgHPfMvNTmx+hnx6srLmf8kt8ZPTy2vuXUiLk+Zlf5XhuUNySRF69U7VcKR2HPLJPGy
McH/Am04PTDMwFy/I67ocCX3nPgiRAzXWMRovtbMG2ofZF5lAJLALF1AcnzikjFaNACX6ufBR6vh
Z+Rh3hyjBjkjGI/Z57e9cCkCukF6KAniUK+h6wXX6J/r2YF29s5JqmyNzl0QihnJx3xPxmzZapZV
TM0q4UtddZCtUjaOHmgFcOy/ytqkxCQmLx61Ut4pgGYTdYsNIzZY/nJQqev57FTiRbynOj/JC2wU
kzsxLVGF7YHU9h06GXm2WweGUebB7+sac/yl4D7Th0gvmpcFZUO7ZIZoe5gI93vXp4RpJegtzOZh
Vdg8FOs1iL8T2/U1RnPnAvMtULxzM0Rw3tPCJEi+6jaz2hMwIlXYOQNg6Mjt5/aF+ufDCCU60UUx
Kp78lId6sMEyx32XP4qXWJvm52VnXoxRQiXH1ObaONoN6lKRRJRcg8FaKQkwOE2RFuMg4052Utw9
dJiAswOroPLRYQlRI7xI+m4PQJCXNIDnukHQwrNsLIpc+E6kn2k3eHjQLn3crMq9ggWQU7wkRKgH
KdfwdTIhqdHVNKoulvz0+ba6gogxUjcKLBo0cZoMmRLgKb6YDpMOtLZlI59dW55Peg+pgJVo1uGj
AzI9r/GTQ1L9LfBsCcZNAOwesxZ6agUm1ixhbBptkKqVZSpO+wHxw94qGzl8V2igSX4xCZG4/YBI
oGj1s0M0v9HkBHEPrXpY/qOBtEoHmJ8P1I3vbADq0W9+0UOXUUnPiYbYypCogsitU06WGC8VISpK
0vN8WtV6UW274Vum7YZrsF5m6Vd/sWz2Nvt9srHn1FHcmxHLihW76Tlfd+JANL747KUJZ7/6PDoJ
mMth/q8QZ7WOWGInSECUT5vZiBGcXaPDbyMSksmqSOmXzJENekJRYfoNu7/FXmqx4YqbaLT3CbcF
Gll/U5Q/rZ+LS/8tef5t4TC66svP7IlTuBSWLau8x312mA1SUZOA/iOtnTc37tgDyTeoEXDL//Xk
es9TK4fKdmw4Al03P8QgbsoYj4x3k/kXnmZzu0oAdP50nrDJopogC6lFbS1A2GVpsB2JHXmcyY79
ZApcNLOovr9/RQiBC2V+pwsqmW81wz3VG4aRclme7+dmMjI1bzaYniIyNYlIKm6Pkul5GSoRH7Jx
xgz+dA+6jD6cI5KthiFietUzuvc8CE83CkR52TEEP7/wSRwvkbhy7URRpIjR/dq8GIBQEq/va+HC
pIdzMay5EIe/QZwvCVmXOHhQfO+kCKwatmCweaBLL4Zs2ZzhFQbg8rgU3G+9Ua4+y1Qo6tLPM+4G
lVtgPM2c3d2+Fsd/7wKrWiXym74rw1WUKM69qjqPrcxbjodCp0hIvDYf0N/HdBdtwffT3bcuRWR9
x9duHO/Rfe+1s0GrdaBWDgCpC4eW17HxD/8Oohawy0fQKlZNFAQiZv2q8bTiKUQetkvhTYqcE/Y+
yfkbodh8Byj9fd2xEX8ZIKHVMNo2tPS1MqCi0JQYs6E2gfVjCe0RyFMyNwlu91GGTjWuZGZUnw9N
YxxhH/K/3dlMJACBgt1fejfemsEIetvTTKV2jx94TSjfoVC1Q2pl91cWU2QePNtX10Q3QcaUYo0C
5EU+Hu5jNCcWrztUh4foMeWDUrviM8mSSPa3Vc6zwBCUqWnbmXXfCOgKW1daaq0iKmKphDkNMIif
wmQUqkd3ZddlzTPF0SazUEW0QLFnb5F2/TgELcstfkWqFdyFF+ILVdsQjwYnwgnl1IJQ+Lao3zEU
UCaXlK8hIZ4WsIv4N8mHRArVByEJmaFHukEUuW3a5LKN6Cdyo7YAt00DdKXA8q91nAQBHCxEIai0
GFfl3gcdR6++CsFebty1ETItzidc/2OA153nE9VmTb7TAhMRmyNkI6G2ev6DBKyBe4+3CsjVNT+m
ZreTBlxyexONsDxzsS5oECkJ1nEkjwOssY1FqPLpPPoL80yn1KI+TRrOQPkozG7GP+kW06I+xpNP
wj0H4vIhI2iYbXpMNpt/fkCv9kULICpHaFPXDsr7wFTxOudiafVhqGGUxoCssrhzzDUkIbAqajmP
BaJgS+StU4HaJxzrVqaa7G/YWJnZz7t/GB9JLK/U6h0VGCYEwKdnpJ5+z4KCwzxZn1myfunpZ5h3
ujPiDYS3ATjzhXTsNtJDXzLlCULiDm6sKurLxmYCZnQN+iMNmeFfjrodI2IknnJN7mm4oeeO3qcv
7p4tQ9wF3EmPs11Wy6VVeU92fB2G0v4WEIUp3ljKz5sIlJ7cbjOXcVWIEco7g0PLu8tV9C4TV38h
+M0TeoOoXGZbvbp5ivTCOcdI2gXvowZoYHGuIoUVhmD9VRBV0X9OR8yjdY+INOzh4KuWjfw6R12u
kpHV9sH0jcO/dvxuPtBetYveefnh1opRW76PfXPRaf0RXR3xNMaueId3GeWES3td3oJktYn6CWj6
x4pyX0UG05hKPqbyAtQF74F85XtJ7jhVqbxRAAyTr3jnebfD6vbdsq6mL5egKINkDbH5cj5V9SI5
GnHTg84+4GJEUr+U0T/2n/YWfWXJpRVqiiHTCZeqYbQh8eT1kldKZONswHFCnT7SRWp6E2BxizCj
2x4JSXmB3EvoUx45Uhu6doRgid0rsc2HnFj94vQanSgqBdPBCXdM5Sea7t57UvWIpcg5F/C88Dzq
P4lPKuLs/fdqtdgSHSVMzcKIsA2zvt3InNv4OUBGbOcv9a1J9tWsSwxLEMNAZU1CgO/bHZPkd9Ox
3iUU6BiZdCHF2No0/EyKKQ9WHZu9w1ZZgARKdftFLeVrEpvFFaH8UPyVsxidN8Eu4fp9ohHC0zxI
SPiMdhbLGdpJtC6PBsP8ibNEKVH3X+cfCSQY7HRRFrWR8WBtTex0sBw2mGNijXtag0BmXEPy/386
4ydIJR7h8f1nDU7X504R34PSjf3i8Rlo5pxerT0ImJYOp3RwdelWcf2Spt/UIRomCXGyDvFL4Be/
vwFaOs8DTyAHP//b84zpLUyVJ7sQlKux63wYUQhqNy6ERrceKZRvtNa2qutrNw9AFR6Q6F+ZYOeC
py8G0usYWpd52aFPUJdQsZ3oPKWuxpIM/feqHXH+5wO818+K2IvBzE0G1BTTlbXonurZYDrCSLvn
Jfp5VZRY+tTiFDguhTB6TJwceqlNS5oZY1/LpbiNHngeSlkF7YNvDYg70acyNjKbQPnVNn99WpL2
CRE7iUkjD8HXaWo85UcUb74wvZ4Jq+ok/BcN2jhYlgetAzzfoN55hIxnqQG/FiFDB3nHKMdfnzWc
qCeglA4U2+a1+A/ntCF3nM4Nw9liuymApxcyMHlCiIZAnNaF58VH+iWvR4UpcxoKnued7QohzC+A
14cdBuO3AKkgOC9bSXovjqTf8i3UJ8hww2/XYMUKzmnXwZMGwsGKaHEiuiJT98I47sLVbvhSLHDV
XFeXK8x/K8c4gnCIXN34smLU8blRU09HDteggTrVDfKG+Vkahru30n3RwVwgmMW05CA9yolyfFfk
+FOJqtp3N3poUpLc9b2LUg79NnOUbzJjdJ08QPmZ/nXznUxjRWTwXNIAqSO/d1O4lNnyNOEI0cxw
zYXXoNkFyZRqEmYF4TpycMD2bqDfgfjr+LXAjgjacngMMtp9fY1zL/zSkBkuYADDsZtEydQiMoY/
XN3Ib2mIHxLqwM/SZAY1fh6UkoYHi6xr0Gy0TahmB0UyjWBxOoJVVGXRBfcFIGiga3Gs8Fn1roEq
D4u7R3mlhlFDhQEPnyUJuUggjS9Oe+RBIvXvvqbAwe/f/JdwhUXgzTXIFnBf0poFiELrLtbbgNkR
HoJDOAQCznVTHyfInirtxBNcP2AFz1CHUJJAUfaIGOm1wjcaAYqb+ec6SqxcjxmUyQPr/sikLaE+
bTPOmTDKc45kX+wqSD2Cmb4zHwsdbvJgHc61w9hRteCjcev5VniuC6EJAdTigd9OfA6hCOEiFr6b
xFA/fc0XLIsqlO9108B76Jfm3LO/SSDT0E7P6WRF7dJ3X9mS1iJG4/0qheglSpZLJlw5Y364/NIF
1/+tXxlYRC2JFZa4uUUn05vMX7ZvAoh+UWuIVIkBrsrFrpEkeg5xoeWGEFgQs9BLWucduFNddzZK
oizB6rbCrN0rPRSGM2Rjdsq/PRiLIxLKn/CsEmaXiqXqQVNH3+cYGaGk1phBzuov9DCof2s7FMXv
MU52BLAItW2rwM7puC91aT3tBoNXeo7nGbgydUWE+Cdep9Y/OryVgfJmyNZXfisdOAY2V08QwJwx
swhFIdRTARuczDrDXVBB4qhTZONF5SkWzSfuBifS8d3ivxIQ0TP/IInrXnzpvwtWdR0OQbvXYrX/
vZoEeEIUYeM6g7xnIZe7bfPqxG+xIC6XDL7dEQxwWDcKXQC2dejmwCzxtILAZkC57uc86EvVX06F
yOYphLmPHkNn2MdoDF+I1YzsbMd35LuFlGTEr6xfcML9pXkbpLrN2VgO0y9WlxoijCnHIgnc3CC5
z+jeCRGBGsyn7SlOrXAFeZqUx0ny2/sdpL6Dzls6fVu7/pKV2wsp2ZSZT//s82wzPxcrqmuWtqh1
pC9T6AculhhwBzpCFColtkBUL3BSlHVlJKv79dk54C+/tFYbb8soynPjKaM8Xjc2KcSpRQBgzm0O
TFVSOw00ya+AxS4uysGT57g6AucHW7bPzIWUILCz/dQDyYWC58DNIdSSRLHs32pHN8aNZe1ukdBs
zxoEF4JlHEyC40Tu84PywtGL2qESblZCbmNenTOgtC7G6vqA/pJQl1+lmvExfazAfoMya0y6qOQ6
vR5ODKQeo1LjHvZh82sAAf3Cv4bswo9osTg1mV/3z8DSXz3mHAHjfdxJ72ovF2l1C48lPllrsskE
7u4OYUHIzoOQ9vR0Y8lf1lCAa0STpAaM0kBQc94OFRJACzCrPapn6aEKELH8m7pVkBR63GxQ4UjZ
Ze9FJKvB94HziVxShU0MpoXoTcA7joZikuoSL/ZuB1M+9q/53T4CHtsuWuKxzSCOTRr/xp8q0CCL
QGKuZiF5e/NTbPAHuUZV+a0XKDTPd7MEWSOaf2G05mIzVZNP4wxyYAgG9nGl4evKezjvOHjaIBs9
oyUFevp+cVuDib7qbN6YhQ/1Uc6hlRo++HsbOTh03UxyOu/FIT0EfxiyJmg2LjADFg7kagbQ5SdJ
qygMplqifLtBcZDH/6lTOtstOqjBwXHTm9JLx7J+b1IVefEbukjt8AYtM7ejhXhgCzMBiJiWMvJG
a0P2dJo1mgaN7HQlcN43dCL2HzpA8GtNJrUJ7kgYDQWh+rnEVJIBxbNRhYa1jh1N5gncW91x5u8V
FcuyCETLoikoff9bjo480LWtFjrebme9bYFXwfu3QdlJrMZgtBeW5EIePd6L3Ygvshkey7Q+o/Rp
+qo4AHJlREGuS5ihE2VVAUpKBAPKIv+AcUetGpaR/SPNCuVWcCN0OjlhGsRRdnCV8Ju0j0T03t4M
OeWI0wsTG540BP+r0pYQwCLhI29e4WmjmbybqGW6Cl9TS0L4c+Oq96fdx6tQJF6/QEwzMFqQ1Wta
DnRHr9Nra88r8hA38vKsp7R51m9tfGX0TLNcQDd4eI9Hz47TUnpuoBTvVBDP4nfUGWeAKqa/ShVN
SWWp4IEGyISaqlh/T3ZhJFuniYvcdunAE77IzJjA0Pj09k3EoA2hLdw9a0MQy6NWPJXOAgaK6wzA
jVT0XnFsvs+LFo/1WhjjvNlU15NQ6nJMelRNKnGZZ6UTVIJzThML6eNW8kVwDTvksJki2zXchk6g
xujkE64+GLeoYSrksx0GifA4PB+MN97R71hdfcS07T4BvgmRff0Tg+lnmC+FaWqufdayj+pUd4Zk
srBsc9/4SqAsAKQKH5oe/TiRry0Igy6+YatC0YCqYRpcPplETgNSdP88fKNZKe5O3HI84xQa8XOF
YVyH+WGjA5tNidc/Ys3pLpj01OYf92TPC2ValLHrnZfCKW+lvAF1YRwuYhc/03WtE2qEsIz1S0ca
jDoHv5PCiJOWdUK8PxhXHMkoeGkqRNa8lsEEeYKUK+KqtlhJ/tXjpSRcVsTFYn6x2AWZyqOEp7oo
iZCq1GUOT3SUumG+E5dYBm6qlRtPbAVUYFRGisJxY6wTh5wG+lNq/dJSEN9IWs9AZatxyiCwWo8s
wzIloJPiS1NJKZO9kxM6wDcq5d8tletRWbkm74Fddmyc6FhuYWXgCGMrn4C0bggyxUxZQUZtn9Qp
f1zbTTIu7ksfDFQIIT6V3//+fBcSmDWZIvyjlNwKx7N9neT7XMXvP4muhEmgp6CFEQTM7enhWGAZ
uLtvjfnK7+wBaXAjjYnxDj/x+NdrEFOkCJopVy2PXD99sLHxIacTHoxmVtTQA5dQJLj/3w5eXf4S
tc1Rfy78pkz53IWd6xg3UtL3iawFZTclM+vmNMgKFuTKBx6XBknX2yVVeock3LesBzaMt309cImy
bjKcth/o8bsvVXXNOV7tM+xgOGt1tZGTLkavd7NxMaGjkwXJ22zqvIbXkaYGpnNG8vEDSZAZ2eE+
xON8l1vguvYYimboD9v1+ukC4G3jEPWykRX8o6AzWaSIZZjlNJeash9UpFwwJOiwchuKc0ud8rvK
zEdt53tY1zVJyyELtrEoVdwJnqqt8L33+KxPaQWrZW60jFxp1qIYbzMByKVq95h0bd5j+PJMAu23
vDyyVKksK3ziWOWFg0TdBGQOgWwDbymbAzOaI1Lk9D4cCLr2DfN0JpwhLDM+6e8Qbc2gbDyUF007
fcNTRg96A7QeTDWhnRHt1dH8ecBNWm3AisFMaPnKhSZThUKciVYV72yejvohpElsRaDWeAW3ovhy
0koY8OlYJCm8W0At7cbX4jEL0gMc8ivsT+G24Xd2bCVROsY09GRwa6Qff2H1ImkrkowiECzIIl2z
DLG7XvCX4QAJtNIjJWqqlqiPNh0xmCm2EjZtqNwJ0/wh2G2uSWpoJJ1URrLjOaIMtPLyAZDVpfRx
sLFnASboI/mNGBW1WzADIAP/BHVyxRgFc84LZmrmdzoSHUTpTFQTO+CgOgKen+rqzMQoR6kjr7kX
uVxSQoEtnRtt9jx6mwSN7K2+PWzwqtmrShjYOyWbc8syIB++hyMWtQgCz7NiuKB0M/y3OmlMQVN3
uMSqVWzoEjSZVkbowmqKxllL9ds6f0HP+rveyYrMfuJGk61iZuMYerls24LPgk/fVU+NyIjeJ0Xk
kW6G3oW7EQMN7hW1/p6KG9Ipql8zuPahMeH/T9i5ek9Rbr4+I51NKti5NoepFRS7qL+ouz3es66A
Ms0awGDBlw0qEH1GMkRRS+/eV77BJjRSMK3+/AcCQkmVWfyTNJk6uBdk3GaipcQOyeqdr1KuA4ER
6b5NLgW7wedmsXIc/6kqskLnwosmbTRQsJWxehgrLRSPN+NdIBLTs9GdUcA0xroOsjKZy0N5iUdf
apz1L30VPy8qQyo/xDcfGNcy6Fkq232kmwCtELzYln3WbXobkJkStyMorl1rhk93VLIHioydrHAT
4R2N4fJmx+oYye8B8dSCJ6bs/EUu+61CrvevSwAWWk0sb5G9L0TWY2GVp0MVOxhu6ygZEcfkhHMx
nCsSGJFKBFsqvNxnZKrxp8D0dbtrmd6ZOGkz0VmXsLL34zp8snTNpzNqHBCer4ZK9RNb3qKYR+CW
ZwXn+I766aoWB0Fc8m/zI1wIUn99RaI/4Ntx/gL154VhK1+Zfbm1/hZunqgCxHfnI4oRCYiwdWKV
Cfua8seCO/9QlZgWtdpjDk4Xg35awg7R1t3nJazol5vgCl2tOvoLd/YcJqli9EWB3Dr7be+83S3+
Q9IXC4MqRTlScndJU9u2OrDAuBPC0tZMsQEJ07B4c/Dquf3qmPTqLFrZQpEEQzm5ZlhLMDR/620e
x0qIQKMt88szjVktF/7voZYFYIf20LV6KuCG4IwGAG/3gNE4gtgggxDwzILp6BqOd77YzlQ305A0
T25105r+492hrBcoFhGv606kwcIBoqTA7Az71dGYqLc+N4DbeoFACvFb515iywk1nVohScKY+E4R
02PIpMnSvOZ3jI7fl/+098KYMfzuzNSD1rOmLiti0TQvaOvmjskTSahgZbg9laYgMeXC8FIIx9v+
cjSo9GL9A92tYJlFFoQk9BHL7mz3aVXobfhs5FG/F68DalNX+o7/aZEqQpAIUTqCPI4A8TbbqApS
/ESqogtWLaGQI7cJ317YHAPX8qkpK3285hWFvy9wB/7gjUwtKDXzQYNaPISb3IwjyePHKZc1fcfy
2E02SKuMYgXA4sKRQl1+eeU3j3n0L7knJi+BLFM+ipfUkp/JinW8IUVCa6OEtwkkJftKooHysTw7
2ld6uvwHd62BTXR5pKrgDTJzQna8DIM77NDfLvVXWjwENbg/9egjuj0hFy+bC94QdQiOTB/UY4sy
EOhn1RgpSpm0tW17jlfG/GIutDrO0P93eRCW5JlJpAyrpRiz+nqM43ZevdK4sLIy1tZoCOvQj26y
dzVaXM0QAWldSrBIW6ENwDae0EBXk5PeQApU3e9muoWsC+e1yVC2jMLOyBQ6o9zMh6MeZuCCiKvo
ChBachwXMPrc3JiSAybXQ+Nizfz1X8d+b0uDWcPu6lF+FU3wB/mmzsUS3+b6xgXdUyvkc7J7IsQj
JEF2ATzZxindcNFctynTwr38L1UJMbhgCBIWIp6rkn4qcc0tenUlsdjdRqtXbJnQ1hvFxOkE0nft
rv9he6KV4AFspP0n0Xarn5mfeCH77WYrqTB4aMaOYAynLxxs4Z95wexwfPEVRel1VTpUAwAf9465
ImE7w5V31wHe9dc4N6UG0KAnTtAcnCcSfiC0ZP4y+FNkEE3pTw3s3ZQWKf4MDP8cKdAGNYiow28A
qhBE94pqVkO8u7yz+m7kBIxXoRKXrvZvmZ7FI+uihcFWssD2LYb7EFg8MehGpsY+pk1O4sciiz5h
gAKKntgTp9jo0SHU56WTRdAPNIOKaLLKmVF/t/vggHEgmu/9wEaG/jIQGyCdxMaHgLLNIvXdY86Z
WS3XN65fRV2YG7bE8bYfnTWZkgbsEv0YVeDkC4Ony+sYS/ecuMeVSQckojmXLXXk2K2X3EXJbi78
zHeDX8bG9DO8t5XLr6kE36kxiTrmozGT95MFVZWH2ugyrfYMaLUD9OjMtCtqjQPATz7k0l8KarWP
mc2KT25vBsWryjP8fA7zg45H8G5c+elefRlpCiD2JV1Q+6aMN/OI+z/3lJPTI2sJ9r6eHa77TO/g
EnTdyhXeO7EGZEfAGGkZIM9BmsEGMyIcSd7bPDFymICM1wc7H4XCIX2ScXV+GpTnG5TIUk3DLC7m
dTZYD0hvlCU7HClOUhWM7g32cskM74qp6HY1S8gItYdCmlCP3HgAIsVVanLjBpiFNaU/nivK9nRo
xF3LSh/Ny0Bro4B7lvANBJHLTMdXO4xY2f5aAAGPEKl5G/y57uPuOM1ok0jT4Ddd/nICGkxlmgPF
bJwJsIGLb+xIT9vxYsWq4vKU7Khy/1Z8hCJqtXNPIW9h/EBnKIAQY8HURUtxeRnU9CUlbXDtim3Z
8lGf966P57ENbyUiMFUjQHG30MYeq4IioouJGZet+9mj6F0eVK7acPC9xJpNZLaRfElPSC57nuJR
3YP3B2yDq9Ef3WcJVNOtBIW88BRBb4pGkUWQTI26tXF/ASayJxSaVOoEWA7HhomYFQK5ag7Ed5VN
uml3eXkbeys27QYD/JSJjDhkfLXkpHNIuvmOyEjVBhHrIJI8ALVAyCKhJWjdwcV95upqf3Ki1bm1
sAOE6XVCWjj9HbcJNRBnlY25/NMwoQkL4sqp946vNhxqTMvmdtq7TcXy7x+WyfHAVc/fQfT4tFtM
4GKEe2axIxbn11YDZGDa0LS+D3Hdw7A86tGOU/MnZtodL0mP12MOTlgYUSxchbLYc556RjPf8aSy
NefXesAa5uUf+7jQcdAc+LyuHgrF/DLsj0bXAGQ48O8Eu3wLy6xpSpTECRsACj0zOh5goOiR9Lm2
byEeG3zUJ7kgwRFkAXRk/03BPBWA/lNbRq8o8NjmXUOUI6t4TxIIb8cup3zVvlipJF/Uub3PjZHi
se91isVgVjkSmc2+TebMKQvHfqQDm4nTE1VF7wlabMS66yZMeRhIQqzYE8kAj9ggrvX2drlYxfuZ
69PkkfJwsgu/NikZSDYtPc7BD+WXGsv8qpkljzyNP7bleDKHo7BNcbYpPkJ1tqQF0QqosboCWY6X
s50mj63pb7vsS5Utmin2+bRuYxAqHW3hwf5muP2fVgs1J41+rJH7Dd148HJY0SsSEFByfIRoC7Ln
8BRFCkm/sNwNZQisf9xPtpgUDRLkOv9wh3/PLcSh3J4dG4JTvtijB7o2hMnr5cNXS9zJuR3e0Yfe
4pUoX1xYqKU0dnzAP9v0e7hfuXTFF2LUcL1a2Wy9jXIs2WpuuLo/JvnYg2OO/iJez3oVMD5J/KMx
D0QWZZ4o3u8Ota0ZCX1jB+Ayz8bKF8xSiWwKPhIJEei0dAzwOVXfS6fJS/e9nZBl+liQqvRu5Yie
Qu1Wpy2D7Qnf6VtSYPLGGOz3DQpWTRErdLv2MAjiBkncz88WCNhWQVUIs49anzW+P1F5FkrkTphj
+nDiRUcpMFHcNRDm3nVNSgMfT6Z5FZZpdKBJXffpPZuQbu8o0xIckq20kxG+YucMf+pDbFwqx5vX
5cSKkngiqKBerrDuhvIsMNrI8hP6ZRCSaR+/WsnKBqJYDqV3UAVMINlOIfRH8+pXuHqIzRq/eh+5
6NGXyYGoddBzeoWAJpN6xMCSVSagAAzuW/Gq0RZwRHFV2No2riurzoiChNI7uEvrfti9WsMriF7u
HsVrvmNmex1qTLFyCCO0c2sGSjtX8mQy2gCn9DRgzjOhlI8l4tg6JZ+nAC/GGdSXiBB8Vf6YnGxZ
/gbo3qqfH6n11aGYcbMTuIeTkCmmm4KWI/WkTKMe4GwJEanUFUY+bqDpV5R7lUWVm0198eVBxT4F
whpv7Rd6h6UmCprHIXCU4AWBjt9DV08e/u1u2g6tP3xDEHMpgYrYANqNZYtFa6QTlxu6JgA2twtX
3bCwWXjy1mxHcKY4EwAkbggnVlL0PyOHq9mhLiD06r+uv1qBU0tUZ7CVc89qaJ6ErRpykvpj8ajC
yVkwvKArt4rMIPFQNV2mAQqDSPqXGqjTbVbaIkF+bOL89lb0QrIgqHWhpdcKi9SOEYm1Qvr3xPhb
cLBEVENbDqpU00jenq01w39e2K5i1s/KTQj01EaJo9Fn1KxR7krBfq6X98ekIQWHS1WlhvkITliw
FdAw0/QO+0rztU7zB83nkrgADN6sm/gACuVLCsH5lSV6T1ivvD3ma8VKd34GWEQyb425mKil7kkE
WePIlSe3TNLBM2Bi/7Pkwj4MRALuZifoTR22+0R2dX/kOxs1kk/2frciVVVPX906fAmXzJZoFhcI
5SPev9jhuRqhao6ZG2FYSDOoVuWYezE2rqVtjCdq9LixSVxAWHUylRlgDeBELSgBQ56sQazAFClZ
CG5I3rH6HEb4Aoqkpstdp3NVzKtTsrXCxQJpElP/rxygj/KecsbsKH+SPFNCShvEDKzAIwXIFiKc
KRV+GM9EJ/RhTYuXylDeSdaG4K8hlID4DKU8V5V9JE5GgmwfjFx7DdFUxworkVNv5no3eC/FcsIo
4nRfiUkz1zQWeVvst56wqLlvCcRHLSJsuC5ak2pPG+ZUuHAynXVLNCTjBphH2wplb8EqB3kS8lGU
avsfdUtju2x2iPrS8qZS/wxaHrOeS9PJEwGJpsTwKcevBwgmohyLWU2vfORwTjvY3v1maFsGPTqU
1EX1Qoq4pUkr+VJGmTuxlB1oWOeokRVc+YkfDpI6bIpGRB0UuIzEh/JA0QXPdfuG6VDAUjofN993
UYi1cz+nHjKceDo502icHpNVfxCTx6sVzQvWI2vVC4WM/Ja09kjbBSREvrcAMbJzj8MLk0aNSSkz
gM8ki3E4M6PORZ3hDY2zUuaZiyPZkVY46banUgR8T8q38sBYNK5W0158J3UwadDpSstRUBEno/Ie
791SyEnWiALSSkzWdD9YlYPH00M2hIyqxEmgz2jBmV5e18jYZhYORe/+NJlWNbZ4ekRTvl1DXa26
NseSubdH10tDmJkPE9NWYdp1WpANHGv0AVp+VziSXtA6yuDuQgo5yOZBsXtZk+eCFqvyYAaUbQDG
dKa0HaHQKuu/oBdId63yZSEdvzeliEYFGasADBXhlw3BD+QaMHYp2x5xFXQCOgbg03abN/wXIRyy
TDeOPhbJUVkyO9IUaYdAuMmeY6IbUqe9RQIomsGuMy7e4PdtEYMUxBq2V8Ea6ft3+CVTChtBRTAP
fIRHjEkTZEphAC76e8IAwEwSOVc+5mEFqiD02Byet0d69hsP6iH34qT8qJZlMHwJWoWr+YHpedlz
vut/63tpxz8kUdSHKriDcY4fFO5l6i0+69ICrIE+sv0txrtYDkakCgszI4Y1uSpS4PnwtcKwxEWq
Ae8HhxvMjXF/Sw8Z5Cz/+ikDEnYYerhBR0AB6rhMWhNHaHpPqi5ytR8Fbo4e0Et+9nwjhdlQ1+sf
tvpDF6dgLX2bt72UqTSMQh9WxGHxKMVakL8xhp9Ed2ENqBlrK4jc4depRwrYEN6nYo+moItYsIL4
HA+CE2zpTmAPq2201ydNt8SaWMDm7/RRHPVJK8WFpGp8UjkJan3FqRuKtKWffLpCh0Q7ht5kq877
rUaReVCxaGAUIz9GAlo8DxBCD7t2j1KXpTzH6tw1mgq6RvSwTXo1L1XRMzRx5LasgRgYVUNBzUdb
AFy4tb9LdybxZ3FhG60fO9uxp1u9bbZkFQUD+66LtdKn6tAJoS0wqbkzez/ZnPwtLu5o+a0WUo1o
5YJry4U2tiTU2pntHZ4uQn9h5UkwGPIUPSvx/8jhxQmBW8Nrf0956Vo6qbYvicGe7fjGSmGDxF2M
0MN7F364DzTL1ZKESK6x+RWp3uNMV2Xss2avC3IIcFyMlfPIt2VlMkTKNNiZJo7lXyW8AYLeNeII
mkJlV2POyMvClhnQgqpPhmRXyTT65g1Tk8bmYITxphQ4xwkZQMPyoH8q8Czrd69p4EgQ0+SXyU95
DngxIaG7FmufDFrTbvGegB/YOq9cgrvymq+8qUZjsAlBH+C7IB3VVT/v+kSLNMlXetZqOSuOwLfb
rs5QstGKKJuXWr3ybDpn6g6OW0lEWrPZivdelD5ZvCSy6NEUvMMpKQI+pLFjegcJ9Hq3ifRJAXnO
akfoS0OobztddGPUqVpkI6kz+TqoSHAX5DpLhgHOxS7cqeID9jgfS/idsq06wujsrHR5+06j+WF4
clfVvy+5xb4rm2eXtQ0RiCQfxZiiEMRDYkcaA4nkwAS3iPhzjHF7YtjsRY7CCdhB5izUoKrefdWc
Z8O233x6toaIH1RecPOy7S8+lz4oqz/BhgVeXjd0/Jd+nDrc+kcxWDbkTsJJ83AwscmK+s1BSBJw
sM15FQQiHGAtTa8vxQj6pxojQd3GlkXjUeAZyt8dTthnc7XyQ3x1zRDQcj78ph+P8wYNSI8bZj5Q
zIoukg7rSMp3fSMniROp78Bd26Wex5DItyDKhjV8/8g7MrOUns+l4yKetl90UBRdtG8Ac07qB85q
2tpzs4wTCm1OcAjweqbgy7k4HvjleGLXRQj7S3iu9zOf132BgVN2pVKASRr9GcV3/JeKVw6d79n5
FQg7u/AHsGnMfqntxpV7gGqH47BWW3OJZudA1gi0Vad8VYMf0ApPOyOXjbOMpvC1IIjyo0Mzr7ig
aq4PSS9WuDpHlhv+NNQi7VrX1TaNaR5n5EbbR90TIeUEi/iOlmWv6/15aUKbZosqbdRHEbX49Rfs
HKcHSHyat/pqdpQSOo8wLdxXvDBAh3DBPZm4QM4XXptkq1N2iaj+SL6B9/AH2md1QtSN73+S37b/
fxFfBdfL5sfHAx1lfo/aaceXK9KQynIIUguX4mD+J+YpelLX0ZGGtcPn2czhiQCBdh2k7Ji9Btoe
8X9YbG5j1gf3LSr4yQGXOBctt+flXYvBK9RT8j5/90e3bb88Yh5rwPIXwtB/fhWJ44sTEHfK6fub
97BH9GbxFvC0gNg15rlERQBSHIAPrM7Ru1uAMJM9GesZFf3gs+zGHNeAS/KsjTKei0dVJeDTMFK9
jU+6VmCUFK4VraLcTyFgtsc0WuBsit0R7EZBRExGdEfiqtrf3Kxe65E5jcSP9V0r68MDROYhfpcS
aYfKWWMf1vGmC/wnpowTs8vkajplBj6i19ueXxgnRImXT34vMOUPOM3Qhhjt4ncbGr3ZngpdbVyI
FYCCLrQnWsjd42wQeCOx4dgPkWhZFQlkGuw+CKBGFunf7kRCe/ZT396ADN2C/wmgWcgUDRrl8Jyn
UcFUQqOEQa8q/l+szxqxpg//SXGVF/O/rPys6mUDJLjLmxh++YcfAL+s6fiiQ9CZHLSwGVOBHwsY
VGTMKVq4OhNGrjg6iS4rCkcNH4D1JltbkBaqZGfJM2TSAaFIvFCufpihUdty83E2dyZnITCZphei
AZHdG+fokXXNWlubRFE+S//bTBdUDqS6975XoiU1ONVJY8d+5gbJU8LVdV+iN2dSZ6gcc90u55Hz
LEoAZkH9FX0mbmo8IeKFOCWuNIkWMiWs/TiMEapryl8Tfp5wCHQof2QL7Py7QcmfGDGHikzNtCoA
2aGEZIp7QPssJv58AZZpAEm22UC6nOGh57yt943Qmy/Lhp16WVrXq9aff54vO7FQ5f1tKLYdl1PJ
9vPhnlXENuR6RIEqWNb2WhOvF0r+Kkp/bAQAynQ/Me+WcaD6aR/etGvj4VPyrfVmL5XE6x8Db3nx
In5DvpM5TNWDzspbdXGEvSETRKrPP1HZxlDo/rfafMLNq0tUp6IHQOKIwkz3NZPgTvj+eAyHuhAY
nlYkdP5/haHioDQji4Ox+fdLDrfjyU89oyvPL+gosW2tXmwDw/f4i0bGHjdPUOt07Xz9/53oRpzR
p+OLXR5qkzu+FUQoSHv0IOaVnm8WIEhjLexJv0ZwpiJ52tUPYyI3O7Nk2VUB8tJdUkeiZr/BovxL
WEiba+83bt6ceSimas/k1zJ7vK4t+WH6F9wjTfhgDurug7DSDoR2sBrUy4a7fPxvrX81ftNS+Mgm
JLtY0Zr9/nKLSuyxJmL/cm36sY0Mx0oEoVxlXk7EQ/XzV7OpYZ0OQc2jdGXQGYMYRsdvGm/75or6
Fls5HiOTxmmyY7wespf7kiTQ4FzoBx9DV8xB18fMKztMsmtMPYataYc1PNrrL2amaAhveoDXQH2V
I4dgNFG71xQ3FHuSWSHceNfLxF2nuInMMQQ6tl1vkkGvnLZQPhPUcYtEIqEeLFB6iMmbPcL5w9vQ
C0FfMdYEWDUXxQv72or9ldE7mWn+PvyrsZPJjkc+8uwkjZhHZpxEOwAjiQ1M7I9wS14U50u2a0mq
uu++Za2d9pKHwSM7Iw/z34yChJ7iPXbY30sp5Ljmt94IbYIesZQfNKb5nGWZsexeiuAXCWs6tSXt
7+JCVDd/5WbFAcr5Pl4qpQGuuVKEVmVA6LsNtZfde+29ee0fNv9VyUJ6n3Cj9+U0OPcLtFWZUMhn
mYYPfgKep4Vm0AzARsUK8oA3HcO99XFQei7CTw3AykvFsL1NowfFkzMoGOQanYu3unXSgkkmzBrB
/nKzeoZxkRIyNBW0aDegX6tLpUwNr/bWjnphsloj2lTh83CZl4mTdoOZBI98df/mpHLeJvmXceaR
LfDXCgmvo3zjHVdywQVNxf1SVZvJim+mfQAfM8w67lrQCXiXc/X7LU5LpUcR75bsfoFFKkCLGdUn
fzW2eELm34S0LDEK2NGLNCyJHkgihfJqF/MOsIwfHuFnKI03uOyDzc+0vCyguabawbRmwgr28W/T
Z3j24W0sOStO34bklpJz0gjuUVoR6vChL7hnmfsXIP5BROnlnuf+tVm23qOM4cDhSxDRCwbPpJx+
E3O0u68xEanWfWU9FeSQRD5ORHqQQIvzu0ms+zzpdxZ4POrD/HrFTjqPAsMRk04YJnnoMenc2bYW
8KuR6GM6cDw4ZpstEjJdP39C38HLAC5oRX04zSjJ9Y531FXhVDf5rfGK0QkCQV55zyub10GGlqtD
6X5LKbr5Bl8Xu7MpXsZEBtu3Zs+hN2x2mYffkEYXrDbwYYR7jl32arbGlAXsl3LFMWDYyUPJwPKl
zrOH/XQvE+250z6/qx7eyw7FIsH0D71wuhTR4EZSClAleb3dOYSbecpdp8xNn7cemgGxSudIh4n8
llZf4ZzuOd4/aY6crHcz3JsVj/dmDIXoWaPniI18oc87fs3jpVELvlOmU/xoRgBv+tk8wRM6+ZzO
8l5Z9bSLCHjAcgVB+fWKK7vSkZphk7Lci/vOoGbiAAL/iQhZFNYhisoScsJGEoKiXumea2TstMYU
T/6D0Rz+HjGPdCx3n7k6qrTIVbbLgbhloWcbvx0W8fk0g8ofRtMq5e+I2cEv0+2v7w1ciLNgtzWk
gm9breLQBy89iQ8gffs3Fabk9Gb6pR4nJN2kab+n1OCpjiLeDzCncuYfrptvJaCuV9Jqauge+aSY
ILx+JQweLNGMICxyUL3XHM2LZzHiSwS3lcd+T5I9sds+GM/7hSdqv5JQEUE3PW8WXbcFoyW6YgqQ
3fKtUHdnGYcWI3jKEIwFk3f/5Ebdp0Klz+5xu6d02hY/z2gziQMw/XWPNDZnPRTt0ENKKP/1uukH
1S8SB0yUjDq0GzU8SnaEyn6KEPf3tEwHWP2bSSCABe+9UMC1wLSQxdaHmDm8sDBZ5fGK95ciXhgq
O+sdIAqtOcvw7gM8GdDj6dT7DL/ETslSFFYleIyaKXTFMdUTiwkZ0kjrS1kJ5pf34v+tg/s9E+kt
pZlJRrcKdRkW+XCc13vpaEya2iq3mA9IvQEWuAT09KZJ5sqy06NI1zH4bSq2ubMmNa2vu3WDhfXo
0fWIXiwRSAIVFfR8xJRrDMFhpCaJiF5EHWVXFsD78HSagxKZBTuG20y06LqvsqaSW/e0FKN6nnCX
h5/OJ1BytZkH5yS+NQqzhJeSytsckm2NVmx2B7ATYpks2QgcBtIeW5YsISyJQcHh1+EcAoOELp0D
ejX4isM9rhym4EXAk/CoyubSFq2z+YTWnsVKiXEHxO4842O+uCLRKOjtVdjSz6zlrf4V+uyITcv3
pPTi18uwakSGaNTuCRhMeIb5RRUn7V2skLf6OxrbD3io6YYIZ52J98tN/F3d5E5kXY6lun6PryuI
Nolo8P4y/nQWvbYPOOXh9K4vWCTWM2UD26oiYj5/42pqJrdmwQaTXPQpT/qWjYlj3K7v0/1MujrH
DgerOg1unNbtdwHFTmoh/IV/E3V72A9y9LFgqcWHv62TYwIEvXnA9lBufpVc8c54Je7EjLB8mC6I
Gj2T32fy2DJXyyV2xHAyZP0l5K5VVZw6q0MIHBFOw8bR5sXXugTDxasNDFYaDXrQnKwhzK6O8I5z
n5kbuJ/7wyRoPAvRdx9ZcFrx3dhN5XRNBlcGdfPjs6jXyDfExqN2XKTrhiAywwsbIO7JfHQ6l+/f
bVk1llzDx79HxAt0Ox9cPhRHsJ0okGV25WCP2Xj+CvaG/0rO0Ybe9v/gWbHjYFEG636Atp7o7/Ic
A4cwvSgOcXiR8VVJrAdJiHykIsd7CpqqaCeJp9oGEvIljXDkFwDeJ4RUcHsY58sk7Prq/agL4Cc4
0mvhoAw4KwPDRqPBNl6om7djk2wTU7prxkYGPbd35w+B64vW74m6IaMjbx5XlMwrKGzWWYjWp6IO
t6NU0XGTv97B97hntmPps/FzwimpPgDdoUAnCM/XMbrRwyM51FpviLdq6Ciq4qmx7rkJhDdxWVcv
WulheqUZ7HLExtdEgxT8TfdRJDc/DGehJ/NdxuI3ieG8CXPrVipETck4hjE+T3ZDupl6B+5HRSh/
Y0MxPIgHBpMPoQOzbU5AKE1JKR4mVm+qFt4anWogXkwss9cAiTJn2HkiRAsONKNYb1G+3xQn7YMi
XVvT4OJJX30+UdNdRK4eUvnoI7Xyxjw+a2drY1K2vrd6y8erfYRf9t8HPRN3/L/gOR8RVXg0KXpc
1YGf/TtXcCL/RE8SQO10EpVgouJBFjRuvZVrB1dfWNd4AxxCsuceDBvZK82LA73mLLN9gLeR5TrD
gBnKVY62WiJfPSeSQH67jexBLGhx7E3M/A+SWmqcYzVpMtgS8/fm1EhsLHdFg4zYJ+mpyvjbycXw
Onx3aTnwfCi+TSWd+2SaixpqSDClGEXC6BPzlRH1W400QI7fXNH2QTJf7dEWtVjAHRyX6yZVtzjy
hyo6QhPLd4yLjN9GQ/qy7jR+G19GK1fIpZ0/pBjdSJR/Nu1m86+1C9Br8lieyxWQmXQHpEVd4BT8
EJKq9kIRa5PeAAFVDLoYj+0I5qLReF5ztWbp9Wuvb2Mx/RkOYrYlKaU1D3pZPCuMEcVOArFbKBLj
TuzcJAvkDhPQ0xdyg3QOM7m/vVcFPExZ9ZORPB16lp9n+CrXicQIaZBnJUX0Kmmn9dca/0z7t/zf
2XSCZZAK6bUUSr52vUgXGZ2CfAlrR8t9s3BWWVMVqAAWosQVNHDfPvnaZgPo9DzMzBhs83Zn712w
6SUaLwhnuQjc3U1zptoz5fZR2eqI8vMDIDEEONo+aL4rptoze1kXBjPuHwX7LtKY+fuXDTOqfDZN
TmjOndvESHDkn1K1lWojbfhlzFFADDlqJ/GjlRBX/u4hxUk5YlOC2kzv3WqYisxybqET0JHRljbR
INezD0ZqNdu7cEJzHqkVpAj48Lcz4GVA0mMHU4dF7HUsc2yobdUd2Bm3ndWUDn0GdVo+e9VG8t4+
Putwq9nyeF6WwaPg2v4JBMKfWv+gc+AB1OSGyG0MOmIkns+DT96DZ5wqMMdLgVA1yz0GsdsNDX6y
Xl4LtzCaVcF0pagoquJO5yPpRvKCwun+s/rXscXq4fsiVpgg0apWlIxGXOF1O7PBiiF7BWHwCf7W
c7OBSd3xC3AFgLWZhBgBAaworzagy/HJreC0VqsDKBDwsEMRTZhZYOMOPI6DAyef0j/cqBRvOpg4
vNUP//vVfvKiXB+uTjMKq3locNNzvyKzpdwHPtqZtkEFt5fG88NKWMER5DwKbNjIrL3Fn/okB7yu
DnJ2Cnv7V0u8Ssk1ftLD1P+uyCMK8dj9c+JgOjQ+3XgtpaLzSBGDXV8vFdodfALugXk+q63KFPZd
Gkfw1g0zQaP3lwr51Pdf6e/E6Q++HIXy4+oPutUXs97LtGxRD92+G0hlgsBTR4+cIsekgCvYYMmI
NN4wnqU8cSkgORqQMxmOTo7fsYJVSTAzISNdG6GiE1/OFwc5gZgOnQEKjTMzzhLn7pwpAwVXCuQP
nJIoichS7Ci17FlDC5FczYEOWL3VlT3Z0gyyCUrpdczh2qMHmRragNqEqU/4kl+ebi3k/cOxbtBt
PryKrCkIcwLewxQsmdiqxDiGt+q2geIMfyUznFyAvnxeB07fRVIWM+ciapwIIzeAFdwBjYjXbfF9
Jf0xLRa8dqFX+zw531xjh0z5LyIxm3SqoEhIOE0+v6sVPLaM82qP5f0Kd8S9zWuwlVOokANAvyFs
TS+AkWdf6pvwBtK8kmDoCF5UZcSNMVIYx88kRqMVqSvaxVi77pjGamCroxyFvlVA6jlivXWGzVnw
NrQmYlLh9L8oIGH0QFiz7HGaEXO7qMEIPaxbbM6XGFIw5Pr77ldlCfO3ioDoSE+4pcmnN69Od6y+
t1/f3BUE8GETrw73VhPOxR3Wim7djC5asxg9pvLMmJ79VYUXuepNy0oD5pilJ/Ewq9SN+DqTUrQw
GY/V0JBEl25KPrTk91nZzDWoIz5RU0v7X2SxrI6RPFNNelCpM48XHX7WqzfpyL+z1DlIOW7YeHCP
cr3+7/ZvrS5fmvpp54J52VLrlu5BpxePFpQRhvxv/ZnriYe7gzbFkFVUsxzh2Snoan48ZWElgLCo
JCbqcAyRWg0ELmIYNqBTA6RFlZVbZoZL2FWf8/MdtQpxLUv7TZ4E5CipN+MDbhwAHTzLEn/F4eFF
rlhHniF5T800c8iJ1KrvsXGpvg8E/yKDqtPJG++FYPmDZPR5AWnlgbV3FcQJceghrBCL39b+9hB3
ZWnvM3/xgccB5RcCauPIjaQS2d99T5FExho6oObFHtMKLmcdJnI8e8PmED0pJTvVf02iscOWD+uE
2UyjmKj9H4N2Ym5aPBiD4VtpJaM1ftJuW2Z00R2UDBgKC29EYMx+qRIpor6Sk6u7VP/+zoW6L1+W
wrVbCdHm6wOou9gdJHXDAo3MorPxCY8P2KHypm+OImga6zUKF7zOdOZPPrD/QULzD31qmnZG9B7I
ZZmzi3Q7ag5+tZNOWLjIUWab9WgFyoBJ2uZr8+6j87N/co6s6UGc1kl6bZ1mr0QS/1benFhSzTY3
my18k7X5/kC3zirQVSADiroSnz2BP6dYLMENslOc99+gz3BvROZ664k+cPLbA9FiKHE8xb0g1IDL
u/r8aqd74Qq6Fup+k/NJy/x6XZa5vdInyZV7yWSXnNLt51eHeopBiwIZQpPlxWNb/ptXt167DiNc
GkTM5V41MMpCK78P2zat+HYn/LT1BOUOo1H+rk+iy3PyT2w00/jFT8DbrdE/cG/t4fogqRs4JsZz
O9mVoUIAvhsOPDT2Rv1i4b7N/x+smE95ziRMFZX+Y60pzaHBxf8Q+soPkSTbvyCPgQSkLzTpo0tQ
wJN2VomtG0gMvbWl7RREmWPdRARrCXS2JKU2mFG2GzmI43fS2NPlEeFaLKN2ONZidjXuOR1xG1oT
ICepZfsxI8HmLyZHmv44pgk3zNOTSmnNtbXTFHTzSMpW0ksKrYLXHCbdq/hLk4IWIFuRKy4SEreq
3q1rpEhH4s2KTxiUtdVBOh+2EGs171BLQlQk9RCII/Jxq9jqc1rGRi5E7cALrL6ExMUnPcZ/5oSq
//k8zqvs1GcKMrgiFPJ6PjgIxkLJoCSiFeHRzaIZ7qYYcMwrNB9103dx+XpAknrwEGiP/z2lTpUF
Va1bAyeUJ6XxBHtrLoi1sLBN/KdX+EIPeweEt0RannQIQVPQaZia+toNyhyTYmczJO9oLZmsj2fI
xmHN3T3OgrkmCS0Y9MkEHiSzMuieGJVa612PHH50v6XYxPYHAsoCfXZ9JYU2qPGzra4K5vQqnfdi
nA2AqjijlKlU+maq9CT9vMiq+tPIHKZLqT6LvVo2+xMU+w1g9DPb6sQ8vfiWE041MgBvArIXDVF0
jUs6bfrqS11xC1+8jqzpyl4LXU5Xwg1YxWt4lbGUl0l+cVUNZRPr6oZrHRHqJrsnrCKxN6rNOkTM
WiV/vSsH1k+I1y5jNsM/0FgC8FVnScTI9lRHrMx6C+8tuqbAhumYMMvPnHPKaaBvZJzUcK2GPJZO
dc/8gWysUHIvrWHjwECQVL51jab5Kc4LE9hIG6lH8N76jluKEzAXSnuubI4nybmoON2sfFFlVwd6
CnjEHqunm6uwIKg6DaMH9NHMbkum4B9FdKkhq9pRGF/AtN0MYj/xuCByrHi8tdIrdpQAuuNSYBDc
SbyZA7llWP1AZbtaDgkPrXeyZpzk8sQ9HrvpeP+GIRIVjuXm6Vwc/OL7JbM6fYjBPwg6yhc7m2Oq
QHuVjUS3IaN2kA244pLGkVhAJM0IZ8O5ITt7zDftDgupQIlFOyE1c/ZzzXJKzTf/15zsjQE7xZiR
875LWrgSbqVVAPSj6XCmHV20iGJoKJb2vBjCXyiP5BNrNu+RQ1QsOo+jMYdhjX3CXSzdRPSk60xg
pSyBzX5WhaU5RMP1VVp6kJHL4AmwVM0x/kpnotyHzeGwDfABiyvUTPeNU2sgaS5tDgHYRPEAinxL
7BuaSulzzEYq4WQZk0++o3AikzvzjN7ScOxmMkfOSpKsr47Wuq0vZbkbeOATWtOrMalBnIb6n9Vy
hXeUSg6RT4+i+c2wnVSnPzKh0bYCLMgC+2U8duFwRo0X2xJJ2FpSN9ywxjb/WRAuqx9R7nO1qQXb
AzJ6Ai0VtlUTy9h4t4vbtppzfK2HmA3ZcSeLDKwkl/4F+nPVQtXOJMoh/vDMBg0ljJJudDbCBT3W
GWbXPIQSKD1r2rMos/Tde6LgM7aMHsQaytzJujeKBfcjqVJrt0wjQRiFC/kXOba/tit1TAN2avWj
hymIqI3tncH3HXb3CcRk+e/C9KnCK/o/UxHoReNMcpO7h0IvgUROPk0p0nukH0iXY5jnmJI1GeSK
hogtcFJDynRO1n2ZHDdFUph3JvtBMWYqdESKqa57I/beb2RdrsGSvaz804Zp9EUQZH9KINmUy3MW
A+Z2eHp0ycLT2uyjS2s6oD1doCBqkoBt45TF2+PXZf7hNXGdvmimvjuDz4vxrBvvqbszXUS77eM7
vvEA5sCLP/0ypo6jhrRJ4PSjgq7rEhPhufNyYuONb0YZ5uHdnyeEwepypJSD3ifQsQrmZwWkMUpD
W5G77GOeDAoDsqE4ycKtfIljPEeUZH+RYGHuJXUflr4AzN+bwfaMIL+3386aFD6B7h+C5n5pAb1/
49TxP0Cc1+36qIyp3fYMgt2cNAGbn/3ZMEb2QOwV5CaqsDEsQ6NjeFYMvx3REuAD+be8N/CqPJP/
e5zyLw4TXy2ahh3irD/5AaIGVMm3ilNvWk7fOvlXKYuZAZzMUQYY939ZYKG0uhHc0LNzt8IkD/Lu
uRIKpgXzLrIa5OxSQlvYWTh4vl+x404T/B+YPyMvxf2GtseFpDUoZ9U0S4nNPSaYgseUg6vGccRt
LhkLn+8zhM3ilLxufBMsuONZ/ifqyX8I8s9Z8GtadxaSMl3gexxE0LvDNL4Hs7CSMnN1Vje0G4ir
b48mPVd92V1r8nm3v2XRlU4PR3XgE/qT97dUH0ayTOhRr3YU9DvRnTs1ByQ7cr+E3MXmsRdlorR4
3+FDDVZUxA0+ZjvocsO/i4xgs6HBq2YiosgT15Z8FVRxkXhhPeJAd26kNCqEovZ6RZKxDZiAI7pA
0rboARnUlodpAGeKytLJ85BzqdkqKrH7YvtSiEZNqUl/FPIORH31EooBRxoeLyvlog8IF4xqWjkb
3Gu4/urmvDy+vPCAmNOlU47e/CHdZapOQmOAqUR1quFOYbN9+Wm1fMl3HJjkoPJINJxCuyA1o11y
Odd6JImicnHn9VWqgB+5sA6JhMoS7siMT7QszEPTELWFzib3CfmvsybfX3vIFZOfKY30Zgj9+Z7h
PJRrj5meeaPNmcK3fu0lGmmN0nS8xuKLwtHo2B2wM1KQL2plqqX6AvCKoKYQPhK7YgeWjnjuf4L8
3/nv+PfcpcItzSVSJNOD5XG43OoRCdAIPWRGYf2edPNOgcXkfE6v7GVowPpQM7usCCOSP5ewyqL1
9RyXMbBz0HPZilr1httlIXhuoo2YMS+dn1Lt9ivxuF+/tWUpzXWS/+kJH6wIagD8WU8sY+GzjK77
jQ+Cl7ttEyXSwomeIBlLWZ7sGI7fDjOuhluA69va5JmLT/TJcEGPctlQFLJUllAc7IaoQugoluIp
P021YZhVFx/6/NA/kDP4KhW014yL/vQS/6Yl2Axw9m2XVsIISH5wD5u1hvs6kPJf8TjTvSoPbzNB
UJGZBneOmkEeOwZDbOLNMbE7xC7ZMbFjWvJtuEVeV1ykJrd5891ysFPq4jZuHI5DCCtzM5EoNxJv
ynIkS5sBr6ucgPoGhq6TZDlnSLD8HgbnfYCBUdEE4KHx4qVNEt8xTS56MLSXcx3tJ4qyltV1P79U
GxdCDfnN0BlsgEh7gVF2CUXK+QPP7exHrGiWwksvomo1Dnx2QXjdHuFlJfQXeE9/JPNe7fPY5b9y
qNu23OmCjMuMq8Gnm9KPIr+qIWRWZTUqGdtZY1kCO57mCsZak41axA7lNZj/3FBBTbrVOFQvZLbQ
KvOGolqrRJzw5kQFCjMir6qft8KODelaORntO68kJV6eyMxbA7vxrRRKtQ8ciWNaMh/pfrHREVlM
lvwu1J08pCySkI9navx5a3W5IOEWgngiDNH+cw0giY8QowbG73YNq39/CFJCQYzLGWtC7kCLWBrN
Oe31X+1Y2zUqAyoYK3kwu5vEBNceZMJFJVJ90K8XX8g7AJGQkhI6eLVBU6n0jecC4zN+z8QafR5b
uVu7/qQd3LYcBj8IjgePrpzJQ94ujJEOxooKCnsiajW+HWTJyop+a2aCdQBRSAwwUvutrFlqNxTp
8j61XxpNC42g3huKvrHFgJgFfKS1u4+4ekS66lix1KG2XZGfxQqQ53hcoEb+yUSUpzpJSSbKVt19
LXIFJ+jlP3g0W+jQxOQF3fW7Ed64YUC4VYV1F41QMevi8+G/4/3wittM6h47Exc4ZyvjWVlG2yrs
DADcACon+wRHnI7VfKffIzNS0GMwZssJXPu7Dp+DNkioNtxs7pmssp44pTkDMhQQsPXJrVbuSu0+
7m1GPO73HQ5NfKRrz1oPFZ5A+5eyDtuYAypbmoW5hMTM0cJU2Vz2qgYuz4Y8po4h6B/Ot0X6m6Jl
M/xhfHQUrzRwsHcR49Q1H79Trx9lrhXWoRWvS5e/IrN6hZzSVd/icxRfzOVMlQo27HmKX7mv/U6Y
5aHt2s8pCoeFhFML7HPZfc3KA786ouHJ/Y+eQs65tj/IJdkfLSbhO3EconZUYD20+JYlZWZtFVFF
/dcBcJJwa34o0UXOZviPPSqCfhf9wkftNw9K1vTgHRjWYDWAGlFcnne1EGC2hz4wV6YtGC2fqJf9
aM9MxKEKaWVzXmNNFjkHITZ+HOefXQFjNsMC6oj2h9VGkdziHxOqt2EspCC5y1aFOREmOI23ATsp
0AU9RudVKydhsBPOn36ivO+sEhiGtH6UboSM3vRr8bLb3o5tqlqjVfxaCjtWmcJmri9t+6ouC5n4
nExgRo5gE+RsoiNZSKrrBUVZljcVSzNORFRqx6B35W0qpzClfQ3jPYi52Ot72boJprGG84pRbC5C
Xfj21ZFTIG29CRvstDskBz+kIa/azlNUfxI8B9Uw3iu6td7iD+qG7qISG0+9q+Uz7S14ffz2Jbcx
Myh0iFgbMlJeKGlmoFXjOhPpozwr+sa0datRqtSVOZcTCFD2rNqIFxiEOl62Mj6/RGHMbNWU9UfT
AAG8uGaeuDYgtd7Wl4F5f3uIK6Lrh1pgKBYNYhKGGAkLx/F4BsxQkeQcPEjzTDr88t203fOiofr7
qimRHEHz4aOLmZohSidCT0tOodyY/6KzjRzBMBZCnROvxjV94dvcFPDtbyZ9/vqQlKi1b5sqjMuK
B7FWZ+8LtXW7cIjzCpFOcX6/LtoeslGJhQ0laWHMk3NwHoMEQYt/24VYRoV61Btag3jwVY8Qvwm/
72fZ929XO0HzQjaIHuR5FKxNLgHSJVeDU1iUwHMQkpjAb4u1FNPOza3yBJ73mIpm8YeytnfXH4NN
OhBJTKDSRU14Datt5g2MvglA9zwXNTPEQib5eGO+NWSbG5XEx//Wge0fg1dNnZ8yMaNBQW8JX9xE
ub/zZb3XmdREz3zy2oi4hnAJTdDmQYzL4qcXqLwnub5qaaNpS3vqaNBTcg0nGT2GuiDA7mOs/oEU
9Lsd19qhVWGQ7bUQjfb9fCpUXYDKeKFhgFZUF83cX3kMMNnHx+vaepHxVMCZg7gqrS9pLJRmLTCO
zG5fLFhii9YoNVEZKhMbPSYgufpXrAJ/WbYcj/anvUkj2bR3fLX8Jxy+FXpRgNrL6e2PfOFtDFd8
XIc6/OR8qaFtpn/mPOzPmzDgIINJlKrEzppR2dmPqR6U4yOCuCSDFCDiAmFVL6JczPpwjmXQdrD/
y2mKHLaPczifvKF41fA3y6Kt/i7VGLOhp22p+1cER9+31fme5+qfNB2EEwoCNyPA3ZydYHRkxFBC
xKdZcwniya1eSvVWz413Ms4tkH62NacgWUEvefHfNY25lWF/34El5OURVAAihhwpACv5cTOWFkCz
PSwRsjnZNNKUurZwMQUqYJvYgPlYvbdrBR+9Tc8BOcxyPHDzIXoyEvkJMGDx6gFVyOFEKas1lQFb
sKSHadBQz4GXDci96oqdalNhpNbWXztfv8WPiBqaIKjH3dGSUf+ZsMU46JrAaO3/7L5uXPl20/Uy
R6+ud1tLu5ju287ehU8yTZNaclc4Tf73JysKON2Jh8oKtWO/6JqpH9SagaRiS5LIeiMfP9IlPwe3
BzxsPiHxO5xjXQ77IxsCpdaU3SQGiHW3beg9zXtCLo75H+8PNjQjxy6Qbmk2rJ38XrVY2wL/qMmV
8sU154vIwGo9SBfiBKntiKuyo4vWFFp711ZS4/2IxlxWHo7sZRKY+sYwXst31lbmuYS6Fe5G/zaJ
Hdj+QIVRL1rtn3gw+xFq2R5PumEO2tQByAUAzfCpZkImTyOEk/E5ca9+tCOimZwraskMWr7n+Gp8
GpFpgiAiLbsAtyDrtA9HmuU4ziAY3NPS4ZAn0+Vrx+KEYsT1xpWYyTd+JOCHg01QjaVwc4E7TPnf
Urn24SREF44piA7U1ax0/Snhy5n7LlPUMlePhvhFKAmsD691173Smynf6c1SRqrykh86KgZqPJ6d
bsgOfXxzfjmbQIqNIWzsrL7N2cFkbJsETw6kLPWP1x9Z+mFe+cIidAtUnDb+y9CtOfcOKsyBk1Tt
x73HzcrelhivytJm3ygw6j9UNU+ZlqRK7NRfDOPrTP4xyUV9KumYvljSLENCxCCY+hjM+2daC5hM
KT7Yb5C3pPyUojWJRjvrD/2hRxpZDo/JbzTllb8mOM4/5O/0Yj1rAvyBnjW+x36qpne/9CW5Q24O
el5Ou7km6gLBbioHBToRuETM2GvVs1ZFUk1nOf1y3aGiHr6++YQBaqjU76YFX0YvblWE3neTz8Q9
CoGvpKMx7Rnsjqfcg9GpMPBb8+O8cSuDS8dIlr+fpXg9nvGmbF9fXB65fal3tbu0+oPFHTEQTge7
DSUbGkKeeySMB8wN0PlX4t91GvUXMw0BAcFu/zA4DGZOVoD3ab/U6p+Akg4PNjJFxIFyg+LdlQ7R
uZWVYuGf4n0CQtFdQ7CC6F6wjEOTKD8WzfvSeTs90HS7VScrabbbyr/O0omvFe8XhSfaFaPpwCYk
qxFD76ZOy2PmpamV7rt4Funo1wTfDVPIPTovLAfUeFS3pEhUKTCvfJGC0IZtH0/sPiFnFk0XHGXw
RV76Qd96o9wLn5NLB31VlR4ZeSJNWml4MP9J4HYeagCA1R81vej6xca2eKkcerpDCExsZE7eI2yO
gVPzMpZGVsUgCYhUPDB+5rPf2nocEcShb56/BRV0zuOG7O2i/yInEOHqJIsdNDUUyQwYHuliOryA
jkkUeKVfhS5ENz7AYbkKbtXyYNh5xggWGYtOgXQT7M2oBuP0Fe86CKyYGG6ijk+jUHDU40gjI8IJ
j26OtDakSz/vyQwYANOq99e6uBW0BqW8RIMbjwbh1ItioTOz4QK5lhOsfsjrZLruBEWBkpc0wHSv
vyn0Ngldu0qFK2onjVO61wrnzbCIioWvGEeIFMmsVEPbZexC4qWUkLbbJ9g5q4tBlHhV+mT3uXjN
M2+oPA4b0Rx8hTcA/8uu35j+pf98LCs0iHgKoTNr0i3BLj90FAwxPXaC7eoKq2L3v5wODJx0GZse
GIhN0lFgE2qpeIRXfWlE/AnelISx0z2EtqpN/jI3S6gQEKX1ByRKAKP7DxdsTT6mabW7ITLyz3Dp
hDxPyf6iw7zdYcC18aQNxouJvKDE5KuzYCHaiyaQFOhs4qgqemhXQjIL0bX+fBrSq/s0xljjn0K8
Dx7BCxjLbTsMIXHsbaqCg3T6TSteqWQXES+SZPDNSrivbu6lklUdWxvgRkVZoFufE4Y4N+IHvs/+
RAm7UlxMt+VjXdIc65dKaqM4zvGlPr1bZeO+Q4WFiFcUsjTzjOgtU4n04gtNKJfDuggLAS4om43p
8LG6/qwzE7HveVQfiqctOwVI75o+T7icz2p02bPV+LolAAHw56l08rWR1YSxGxk5+ThegvoTpkCr
iKkgBkqltemwwhqdI76fl8TOEOeigN8BTJltQ4Dnuet4hADbb9k2fLmtzy1tbIm9JySokSFcAmaF
bqjjXjw5YV5QTzzPIw8O3f59Vg0zH7bw0KEwZrtQ3WK2eU7mGyy1L4fmGnGRaoIbmMWzjoOvwiqY
oyqFHKO/PX4Sl7uTkWhw6kTvNug3WLSZfxe5a2yeMn3LwjCg0DUHgW9mdG35rp45RcNOtLTIdd2x
TOPkubx3k0mQc/rtuafoimBma+T258VvQqWCrnMoBpc859XqIhbOUE7gW8+bNsJtNCZUabAjFneR
q/z21+5n+hSCLVEhRHX7AymjeMd21UwXa8c8Sdt4jOouRLxMjL4Z3D/K/FuAtxaEtmQN5uhOHmiI
wRJF7L8DR8AcPn8bb8nI5+0kuO/AVmi+0jIyzOZzOYkiNmG+WDHLz7P3KPye2IF+3sGpazejNQXO
QaD/uDsgxpgXhCf7UQAD73rW0XOGbqfclvsRvgodiqxF481uhJY3QVfOu9CuGGrYJFb/P4gx8bg7
g2IWCJCu2t05yTrIhUsxXDqONUajjCvnDOLHBt1Q7t8U0BDKP6vtE8hC+LJxaop7n/mRee4yvYpe
67JUCGeVTIhEAy9/s+7w3cI25L3SA9kdazPo+m//xPysUGJFl+e9EIoPZNJ87Zs8PTUOClxp2yjn
np5G66nj5tenhNvPx23xS1G5gdZvb2+26f1LqZNgbDdjHZqR4AWdYZe2jMAaJbsCghIArUxuRrR2
kbycG9e3Aagmk95vprTxVZXjwGkoMTIkDpKYDdKSz9T7+jewj5G/Q4SDP6J9AfSSMgTIfG1MEJ6q
wtewEFZvaH94t6+h66/toCeEQQfFsxWv/v84rpn66raf1feZyxegviLVLapt/mm5iqqIwymPpjgx
owyAbxzfjQ8QAdTx45Mm4J4vc4wNx/eMenDQT+VE+39Shko2DQnokTcO5eumSnOyBrtDO9eY8VP9
KEBfRyDgoLrD18f+Muffa8jriDcUfVjkJEukTgucuXy9z1VvKfiyyl9dWkSnYb9BaeunBuurp1Cy
Mb+qlO0OOqIDjW924NSrePcdtQt0oaE5pWby+FF/lNWLKXht0yTVw+FXWF68bh5Gb1hN0JWo0A4L
LWS5y81vy+MvYEyluMJeJPUa//uUqPmeJxR5TqD4m2upTrGgB7dWWDOPSngncLy3Nvbm68xi3V9F
yUBS5uK2S/0liAM/qIf4srtMD9I2XYIebhoGYX1HGKrATBQ4O/jHdK9ZkLso7NbDN1HzYOz2gEFH
V32spaQlLGSPN4+ljNfDwNFHAJfmZ2DMpVkUiA9nKCwALqXS1dWUvnKkPTPa2TphaNZDFzT1Me0y
gSP+ixAPFK1GV2+Vc8IEYbDLFOQ5wVRBMdRVMNqQ7eZSuP5xdAI+4YvRhWhrRoG5xRgVszGzeuHc
FvG6HCQyO1pyD6Mwv6/uOdaXrhol6ayr73jdsC6yu1dtCjJ7CmStAXFu7/qb2QdFKT0KlilZzqg5
h6vpBDnHDwD2Qlf3glz6ByZyCdxRpj1vojWpkyr6wATIMAcrr4viKPIpQMQCkbPUm3j2FNTdZrAp
jSDWvNU/0zcIl9NpZjeUPR86ph+cMkyEZlrL4y33moSTtVHGgkPTBHD5W2nHe4PSMuUFlSLOrlZF
fyDI0//VrZYgdf8tcaKzF1Ppjq5f7C5cZ2voR9v5OI/JiSYeGMonaGBTo7pcBLSkKuUV67H3/B/4
VrppcDo+b+n6VASuTif9ArfM652W+k3/9NbGu8IbhbO+XVblxYanbPAiLmwTUorVwY1APAU8WYCy
y5B2E7akNR6PCygpgju+29XpeTiOljoN1Ojl+cC1k9cTSOe3azBqD1L65ljivi2cdYz9wDKqe1uy
ThhSab8k8WhGzXp0hAVXYHdEOGzQ+Vme89zEk7FjIXw6k4Bl8fsdSEuAf1jtQpabKMtF85dvgi0c
1HQnNmTUeoIkxhR1JOpktLzqni7e+JX8UQ+ZbsbLiuWVAjOHvAK6+D0UuA50ORXB4O101Ah4uVgG
tEFOwLXx1sz/A1gmoF+2AINYnKo3uBMgCL301gEd0BKBheAhbwJ70LtH7lqd2ERW3utVAWMZGWmA
WjjaK/5Ni0vIBbp/wJvq9nwpM+Gm2KGXhG0uJn2zJSO/F6OGtWAmzBS+RnArXp8Q8PJWycxD9zif
4akmvVo/amm4TP89QJMbC9B4pzlnXF8i0aJ5noz2Y94NqsAAkE0YuQpSYuBjBJmOrqastfzIsPpt
MyW7ktytKH+EMoibqboNV9/KvGM65xVUi8K6ouLKb5F8HEK69mkAv04gqZfgWi6w0mCvBiH4tgfi
KzZa+YcpWYx8RICW2SMNy5dY1poOFe5fik/BfwP4FtXpW/5aC/aE55FzAjd1bCluITl11zsvZBgz
aoRiHlvaZNREhO34SdOTbg0K1QH+mASO9qSYz3M+k8FIPn77xVn1UycbtwmwXntBj/KXIUMWqWLe
mpxJzVv8bbe5nt4ui79Lfq9G8r889cBh2pUx9W5Fj4VcSbhExlaIyuw7C6mzHsrnOV0WgsrkFyqD
jbntQvhyhMuaVW5lJLBYGSZ+L5FnOTb/7gEsRuOkmi8PreoWxAUBfgOK0KYctM+qBB3bC+0mCDre
SVBFT4Iq6AVT0JpDk+FQCZwb2Gv5fT3lw8z01S3OOc5qr6cYuRSJw1V3ea1jXsJWF+NerU1c6tDm
CzTo4no/c2vd4TTI5Vdz5l/ao/CzyKjXgtLmn4cfwfYgDGmsaOaOhBkCIrQXUmAp4RBTc+iuYYab
jJEExrYSirmrUnR27bMwmUYDFLji07x0Pmj2XAVndeaUGNckWsBODQV2D0UdasWYSPKj+sc2BLxs
t/AXE8JixBcNIrLFwN87cbRbbDAy4nv5uEN+oKFCSPuX3cqPiVd+vgF1aKQ7o44JStiZxTJxKSSx
WR6K5ysomxkMRY9PNmZ9lAuKxGMaGTli5MRTsgm5Zs2ki8uBoZNxLoCq/Dj4GWhlWUYZOZHAOwfz
jVVf3cKBxVSpCI9rkgcMqwXsaIbu7XG8jr36wbsanadjbftZQt1bZoS92HkLndXWT87MUvoDUEBR
1OFPtSx3Sh4tdrEXW5Du3vPLBxkfHREB9/XG4E8qCmCX9/4YhspbRLqemgbCdHRMhcXrVkz5j5LY
QcEBp59nzbrcYHAzJV7Ezvb7Olhu4JSDObda+Pez1emfiM4TrBw2fV9hDTgZeunCKMKTZbbQP1Am
raoOdy8rR7HIsTLd2WCJqljhu+QmdFE4qgf2EJLCY/b0smC48WENzutK3nczdhu6xevKC5u1EM/L
ZC0Y2hvVxWznD4XtAH91J5gZneBj5vfEXxMRFI3voQeAlEPn6xG6wj/T9avrzW6qQ9jjwBXw51Gq
06fksVY+L7IGBBzylyufQe5aa4O8NrVQ7TSV8916rTo4xhyzkiOJJDJYZabLScn8fUggTajTWm8/
KI3fXwaNi0Kdph+2K5d8SsGFVE98t0evJhy5LfXj8F3YCOn2accJlaQYALtZHasUE1oihqtbMBDr
Net1xh9xRyncNKvr0662QTmdvOlJAZ12rrOoSbPy2wirmFkVONF1qWj2YvtflkvJOJaWie33wAZU
pNWmWDySVWFPzhhDp6W5UE1LEjWnAdoi5o0drHB06fmKn8sBzEn0S0YyOFJIsBXey3r02kpmxiGv
S7GJErryOwhkGh1fopapCrmdcH9ngSTebO7d5T5jrp/kVqzkry3wRM4ppw24wazHRBKUJC4icVqo
WCHC9gUp5zPWInIceC/GUP3a+WlVX/VQNvLflWR0N4tcfNVQakC1gg7z4rKCz2uezpI8Ve2TXp0K
9dRTbJk6iIv/Ngp5jaxe36Yd45B40mPB8INUFo+YM4uf1nzZ5ZshzX4x2WHspxHYX+rDmagBcft/
vJDKrkgzYopk64sMzEJZ9E2bbeqZnBuvCvOkmKqh2H2Dwf7lY6Um7a5JkNeN4METGAbiJJDr+db9
XQrv0intbZkPRTOgU58LBz7pE16USAkxlFnrCmoA1s5knWP/M0GSRP/cD0dR8juyAO+ZSG/vgBsD
pz0nlK/PiO8LuhmHIfFQNXq5FerfERrdzfYqgBkAnyR2HHae0pj9XtFMDRlyfLGj8k4XivEb4tmc
jRWW2srJ2BB7akvjLaVP7/EsZLKJrL6MXtfHM0kwYTaNmodoFPpiyuy0Z8W8xk8W2oqmM2RaCnzj
DCH2pRje4i0VQiA6JbemnIo08xgOr1xNLqxHTueXedwBzFkptZYGW0wVppXXRcssc0u5m7YkAoAg
w7BbDyCe8nik5hFfyFbrMr9dN2W+Tu9hrJYRCB07o7cEtS2tihWOvZELLig9NiL/NLFBdLS+xxSd
qmh9Hp6yOoxbj11tjGzbavfOZKXqOXle+HNUTb5+ACxyS+WktxPkZnvOJeAh63yT36nBimJX6uDn
36gVmVae73zT0284S37nlnFCv8nOre8MvFnRJat3DOtiDKSca2l6uUXyl09kMaWLXa5f8B6zALri
FQSE/EL1N8tOTAWVj4UXaycSCbYEO29aunseF6beguZGlTv1yN30PqCYzTM8nYOtswMoYlmMaY+9
j54ioRTM8mHNKKshpJkaMjAPsKbqLjW5pWSGXnPSlU2vyjgp9q6+nNBj3+wZCHA6MloCqP7oggws
h9h3zrfqEhRKJQhsfgh/kx3tOTNPGIYQqmcXHPaCBX86hMo0JKKwrlIWDI08m/ONyjyHaOv9wohY
w8TARuXpScDLp4LIVWtxeJs69p259dLF+0Vd/GdXulPInQbUQGJg1JzEJu0aNj2rkfjvfL8F6VHZ
d7C+xm/6qOrz8Esyw79LA9LjZ2vsykqZT0kTn8KgpwfZ2rowxF/bZiWy3AzmJES10VKVDx7v0bd0
Ixa8tXsmTbYNhCaHHX0XZmBbRjFphLYxJHA5NiNOHZGvbEg09046x+cvckRKBipbovVqmY56HN+Q
/EiFpR5DO8C94OANGswhcq293iIEzV+6N5x6OMWsz+X9awtjUblNdV6YAaxX+w4o+k83UK1tOcGW
4BO0dbosBLXqTKNGm1WC+8FdtZW/MzZmbrJueosdJ77aR29EkO2dLU2/ig/+s1WY5MNaZDwf8Bo4
BgEo7a7iQWL/Y9LLc3NxMbGjq+HvO77AMYgDJ5nZm6aFhwd0KmmXUYjGIQ7L75jAujyTfoQW9pj/
o3QaWb5UCm/SfJTAg+0RWbG00YTCS63JIhi+cl8ca0yJTfhkRd1LVMEeF8Qb8e5xeJieVYFycRxp
v1cPBLdMWs1zcfsF5o3A7xmZg0QMHsvF591d2rrfwHhKmb0Ce59cJ9AvFrt1s5ToMLe7EYWstJBb
1gmGoeEOOGUJ/Xbd8EZHDLomsdyFzZde7ll6PbzDS8G0NW805GZf9YV1UT17FlJnt7dATkUjTjAH
KtgciWjao+zbWMFuDuQmoVL+8Rk5//q8KnPj6v/yT+XBdqVkQyDlecK29B5xw1sGHY3Dbba7ZSKv
Lqeubdp2i8x27f/r8V3hECuWiV8+LwUx+09X1xHjYHKrOtAi3fgU4+VwEtFkU3OTHeqVSUtCVfnw
pJV/6eHqLbgtEgpFQy2SyDPWzFpOYt4eW3DLl+tcDhhaZ9diIffkI9hmlWnDqqXHYAMveaYEjnY/
Cc2ENTCCquRRSJe41FCichHbaP6heXQtwcBEBjKdfqpn7tsFY42DSexzJLx5X2XyUakojrTqKPyq
8goBL+mllETZTjgNZjaqfQkVz2ktlGxqvsyTiikF8E1h1tZ7+lRV+37b3ww9wH1Wjtn60zXJM7we
wMhHRlsvd+F8j94w2UYUofeEZ+WAQgHqe8KTxVa5opDPV5iyRofBl474J9WrYxbtizMbVnOU8Wne
4LZZ+I0mKHJ++qVYsCLATtuQIKRTZSO2NrIjJC2PT+bsBSUG9JxNQCuvfbIzDRfxTwz9mFHTt+hI
aDVWqTZc4Y2O23oh5pG1U0+9Pj08LoV3xfP4SwlgfTdTegG8oZNGVzH7xkLf0HEVkjfWMoKyimlk
D3iGY5zS7NY9J5K4GGU6pYY4uIVB/93RLtisWmUPZJNwEqXbCrJmjJMoe4UvsS4d0U5apYNSO2gp
Q5zVOa7wnFdZFNSxSfTL+K2TW8b27UMKgv7HyRQkTWX3peZYalZICf5BXZbNQuo7mvu6mOaJy+QC
eLqTE7DOKBtkvgxE+yFhO3V3UuQbl+D26THCliK7Po+9bS06qCpnM4cKshBwWhSWcZokTJXKaYh0
SCPVi5Miq6N01OzP0VVB+DhIpKPpfoKsFubV4+sxCyKu8JRJT+5hCndUPyvd+wehrzqOwIKSV9lC
rh1UXjjVW5kOpWOkuBQuO/KKzbkljdGPVRLOCajWoewrRdjWTs3WYsvUPdKr7/C8QAHgkSqNWFBm
02Imq+oD2Goxw5HZcmOtv8UKKLKgFcoxZV0DAHMecVW66NJNV3CaAOJIdZcHHCv1xDsS7dMrIThO
wW+xi0v0D11ZTP446fPw7DHqviAAuoAM/2FdvQwQpn1cRgLinfS8lG7Uu0bh/6svP3PKqLp2TnZM
DyXUGLAw42ag8cfhTIuDBRzlpYOW9AStZ4Hep1IQlMQKOcmgO8E7MDdj+LXvPzK47uUVRlwlvGEa
g8xpf/6e+3nVkOXt0b1MnnAmct4eldwVt4/UB7NLqrtKRN5M9JDTfTOUVXk6kxnX53l1rM3gOcIP
h/k90MAbt+oXWtcet2Xb540toonoeLZTgvC0OMLi5hSGg9L7UXHiultQrppY2eGjq8Y6i4XL+kOm
//EZNYMmWeahtWRJulN7vYBDt5wyOcxRGwkv/NuX5OEStZ+SMM9JJeTCgBndArwSY1NSXmfYUY4s
AfAy3T2wWvpvaW2658kvXTDGK81pL0I5yfkJKKZXANMX2ZT4w5vfEhKBX5Qizo7nfg9OACpCNBBr
CrY4l4fHcHTWSwyoJ3SEARW9OXtf3heqvICwp8Geu/v2NcvfuU7URiAfoy5Pr+IJxX1R/PUgAVZM
e0Hi65YzrDRfeD1sv0TbKa9VnQSF4ruSXlk392WMBJALbg9FcLc1eqVJCmOBV+8ELuSJ8G/F9xC5
WGYHcri6rdGsO1iCbQS9TtE4DjclTerpZeGK0ViqkXPqebJh/piTfZd1Mgh7opVnipCOMMowefnK
2q70kdn2DFubTiMQp7mjj6ftMLQ0vXl75QGPF529RWJ7aW54E3VCAPTt7Fhj+UQyUhehvq6HU2vE
tqSjU1r2wN7B04TAM9R4x14n3UloRt/A+OHRiYwuMWaVn4yFIY3yWWt3ZodTga2Ek0Ujc3cvT504
bWuZT0C9YBxYgw82kCXTI0VDedtNqclL47MBTDysNuujGRM61aezSk6VR18SVTQYImd4ft/mnaOM
oV/aKPg9tDFC3GboJ2Mp2J2mbRtakUaunlqYoGobYXUggNAiK7cZyLxoNPvf4Xtivae8NNUjoGT9
YlavXRRAmg9MbqNbUBjebukjLrSVgUZ5IB44QD8uovxXgEaA0HST60KkYFLGlefWwBg8LVnsZb8Z
io8T/SnGReq2/SifmYZNuHHHlapLcVt2N7ADvy4Ih0vc2gkMTygWJXTb4D4KjXKfx4Md+Eyj/Q2K
L5Tw4SLhILsS8QrlpH8jzbvBgdw3vbVwCkzp7UHZ7zDoGJ4gTdVWDIMMLymElsHQ5BgdlmLxJ51e
gaUSiy/qKG4ufKZ8CXPSeOpGTC2V61pffcfWGqtLn9mmO/K8VqKjrRYvqYKRe1LcZK+v2alu5wXv
HJ8c5vFTrewv5vAXzyEijf8ZPUPbUw0Vvp0KyV2SKpxIL8IxZHN+bTHj/gftjHdw/6KCS0KHYsZn
ytxx5jgq9FeLUG2CSS1EwPAS7w/dx+ujGxrR6qnNriB79nu2zO/VtrocSFtNcpNrsSypDeBXad7z
XU6iv4LY3Mrtfe0ZNmrj0+nAm/nWsHWKvIBrLjMCbHqLghTS6XWaLXhUBpRz81m+hsHnP7ktrke8
nhnVGeI0C/cUzhWtYJncMoi62IO7X7uUN7MO46Rgy1UuD6xNuvz5geNApkJIoL16JhRwrDY7IfbX
yqt3NWT8zjpvbm7jOpPffPCm74XcJiUKyCxYJMwVFijG0lZgwcvA3sPTVRqoQIt5JaWVXp/qYNHD
cWyGPYd5oW6oqK07rVdJ8bZVVNFttyvbX3R8Ne6ATgCClZ1KIGGHiIAP2eFHf1AfAFMQWqIYk40j
Qw9KAM1m7ergLiQ4FRDNrejk8rS5pBrDS5U5mlh6CLlRLy5lSCt+oRjktxMcpymHC36rRETl6iZQ
sZ/6NVzSP5x14CdzaL2V46t6kmNGP+voxPfuEqs++oUjkDQcfEfoqxEUiArEn82WaWadKfR0aWxL
r+zLJ9kNcFueBuPMezYQatLRXwiWjGn7QQu7NVqxpSxGs09OOzctqg9hYv2dwOtOMV6GdHtJg3jj
FKrxXb2MRFnFZZZduZYHMAc9jX7m+gwTKYTq+Y7caeKQVLEBhsSaT7a3l/mxw+Rwe7Ya2XV2hRNm
1L25y76BkpKAS7F6rzBDHAsaIX46bE3Y+do19JT06je4asrguSJBZW14PVN+Vu24gdN4EOjE0JN8
nGvqgoNBo86OOsk0nsuTBJZoA1tOPopvsldXZIg5VkJP/JZZdrrlqUoThQgbD9NGWH8lpatvqAWF
QXJKJiyKtWojEkZVn1vQ7zC4RB2Sljeul6HFq0SkZqBCb08d3RwgQjyjS+can7cIrj6LIHKe0+Dk
3IPIeVtEAX3WYxzVyN+Pr/grQJejhnOWUhoHl0ZtyOt2VQCVKHJo4ToQGxHG14X8EHWdKcHWPVBw
O2ru3QpKFZa+lT8KGUivRE1Bp+fQVHsF8jLg+pcNm7XNHmF7QOX5JlHWIIpBJT+3e66nLuhnTzF9
RXDa32Dr0MJqqpEPamCxa05TSHHS/BGflKz3SG10wWT7KDfvIfUdDnl2zn1489N47ZYUdbq1R7Uw
6EAhN45zwmGqi/k1U9R+ZoVX7TS7X4gbdDJTuwLO3yJHv7wZkv9qfwHVj2MKQ5i5eY1g1mMjYYa0
AwcqizbNWjPu0CU0FGKidAb7vmBNZCvqogsaj5Bmu2bylvJzD7Y7Lg7HWEsRpVaF6m7zEwNPSyUb
+Znid9oyRyogn/RhwDZkOzRJIE/o0gZ2cajxeXuHOJ0vRm0DvlWDAPSzQlk52YyniDOAI9vxEMNY
QeUfzZ13w5ds8f0meDnjva1gb+ZGrIl0pwas011TUr+Z0eACAvfYbH3CmYl9wfZ0fJzgXR/nZuoE
qSiBElPYaWFQcyq0JwGMq9BAfePYpqfWEE4LM8GRDvT3cEY1Dm0lMVUeKXtD0nMvTIuSQ/0pkQJp
ZoFsrvc4WADfDrkcaF9sH3vuYChUzEZ8fGfeL3Ls6e/tSD0FWg2MXt2NCffVhhFu2TSddc9QDOHS
ZKj5yeR4FjLmbEIp1ggdmCN6UvELC+iM7A3PCIxBvqR4I2CjVmJ8PptljrCU/3ADnCEQOv3GUMqP
X834jzps1mXm5dii8ZYvcEOxBcUv1yeCKgG2QAA4nF01I6O60kWejdoBUeEJY/Vh7zQtwQUzG28w
oZtX3o3N9/33R5Mw5Mfmu1GWO4UZfnB5tDIdzlutx8kDST6AydGZeV573kPwejTiFVf2jSvKT2gx
zTziG3OdpQWarV29Ld0odEtO9WEivvXw66H4p9ZTihEyXp8AA9EiL9V/QhObIRWfksWVX79IEt2t
HdpHZzukvTiFXgO/X88H1/PGGP4L+zwy7Lg0TcYa0bYi4xculzkB2s5upoNXtlnAwX13l81Yo7an
8Lg/QDN5gp048NxBEerFA2baXdH94nWevGgwNEMs1oaGkxTeFVScreOaG6ke2TQ0cR8iZzkEuR3+
tP/5zaqQs9sQRntlk9/mWyk7AJm5psGOiyqSFZ4JvFBwzMNPoMUQQ17nbe29Dqm8ggiyWbqIxzhA
8mR6QmvqoRXX6drdoZ981zixEjFgMIyg3RY7/odd4DEpOsk77ezzUMGysD0mFBLPwbinXVwy21WV
fWeul9cUWF+fJ73NWwzefBNcIMeIMp2mhP4L5QDVjAfYmaoF04LoGFGFNS8OnEmZ46+H1kXYdZ9z
SGIudD2RPSyaCocroEHMENtsUfIUyetKXWonGPBNhA/QkwNIuGzdvoOJrDOHsz+cHX/zkP6Hkl7e
J09vmtDXj+ho1gqRIqFJTn63DlQxn+O1LF45h/eFQJ1Nw13TlR546kyOqpTImkTC8wfwSbGDzXUt
1AqV+p6RIaFR47ts9fhmaes6t/lqYEIb9lu+mGVrhxrA2nWG94okSRMpvFNhIfB9eqctZzMffjQj
QcMkzd0Ck9uJ+WerbEdiFNU9RVNb2eqIISlfasEMVRsyswpHWiXNsCXYLKQEBoxLiAFwgJfyD40V
WOlXPAj3HBcPkcMcYOZJDFLex3E1OFCWCJUDMfDaeug7i0rA240p2PtlUAuMS1P5lQxgdoe501R0
q6fOTR036YA6j3d/w+lnyRzykToqzcKZYtBbTiQdFVCGbbvlvnOknW5CLtpr21Y7g4kmosN9PXos
zcXksSOcNzoVmn5SEIkN4e6G4KOxnMsmTalo39x+PN8Kr9DO1lhoQrq7LNcHdxEPtzJZADaZqhj/
yYiByLtvSCOQzbpzvd+8WwiN1rezi15fOf9zp4+cLbVG4zz/gYqdGey9Lezb+oCr+KaHDlCXpDUi
//gqsy8XnLV4hxthQStsBVEVoOsTghr6SR8L+/7vwmJ2HZPbXU6c5sfg6gImIoNf+fteYL2PcktA
EFH3817u1mFVZvlUHkNhGKDojJmKMniq1wiq4G34aIwN1RFQeip56X62hztWOc6oto74jEKi5gxB
e4LnQYg0Be0iyKXeb9vQLnytFBa2Xc2I7apeyeC2CJ6BYjeKGNCK/UpXpPbFGFgvNbOkSZww4ZQk
rdW91rcqVTLJrj7PsQkXV4lh17DRbUSD82WwDyzFMZKxQgf6WBxgMkXWVIyiJZiYxt6YK6Dw8MTE
13h8udKZPMbdsTRzzKpbNlxkv1JyXAmarrZgB0B6YEnxrMJqVfeUARJVIvZzVx4frU7xILIZ7U1h
mWYvTaZoKGqNYrcmdqF+tdka7tnbrDeYt4mT9DMk52wvWEmxH6oIqwZ31wMskWWpbOMl7+/YWoxQ
Q3MqAZ8YDNBuqDtsXDre1RNd4ACy2PXxHmX05G7Pcid91DuperKsj+2IXJwH0MdaABth0J6EJkAn
ht5qaXXgBFpiHEV/UH2fA+ndUdFPfj/JRrSGmaCtbmzqfGyVqitK1C9dMPmtP4Fq9JjdY4SO3D5B
TnvUR1eWGRmgMWb/37ENHxBdJPP8tZ1sDBwYC0QYdi3M7supDIeyv2c3rUmkhb1bv85wpPMZmHF+
yBAg37o6EKGQwx61N8VXI6f6k8D2/SQXQIDn81sJ2jYROtiIWcV2MS0Kyv+qzOhfVfPKgfu435J+
l6zoTn9LP09Z2Vnzv3HeUhB3xJtoKr+i5zaGSbXEHlrs1eeDgqov8/kCi5c/s8AfSyp1/xY1qe9A
HooLmfLbeQ677QjxghXwbakGv1ys3tdt2LJLol4N5wdFDZ/GYHEd7bP0hgpWZ+dufiYK0y1WbcGa
7DI4oEPsSjUdnlc3kxnL4elL4DG4z9EedC4B3Tn4vyFSEX7WW8NvR5eCurPUKv5gURHS5pkPG/fy
eGcVP8dVHymea0v+aTcHMxwubRkaZjhQkCx7NrXPo/tPF18AL3b4oMLC0ghuh4/HAzjbbjLVhEGY
YROlczynH55OwQxGynsmpjdXLsQ2CuezgBMwZJqsTQlawWQNjJdhki0MAAMip33jwseaTO/xbfQF
vgHc0gp6Z09BuixL1wytWC+Dj9W/ekmSB3SYb8NW0cP82ie9V9lqoRXqYhYrkDxeKhnUXXXkhlPM
Flz/eZGIFf+QAPxmT2ztLugU6pUZTSoo/tLszMkjdEyQqRAsFcG47j97PTv+YnFCpJdkiOXnJgrk
z4NYNwNezLaVK2MoOGYmmC1nl+s+mcNvhjRxSusqjCUOZE4S+yDGJgtwe+SWVP2o7xmFGiRFwJIB
q98IyXpCwBACsk2AZGbUBksHkty2SE+kK6+kwQDf+viGE1S17dxgdqPt98nIMX+rb6K8jV/qq3Qa
9jwXNPZgs3PnWIBf/8JrXt5bRBGBW1Gr4ykVpdcx0z+I3T0S+rSZA1iEjdrsoT9aDfChOMylLPSH
+FZyrRELFB/uGe+s6rLm8kkRhyh0lY6Q4HUctEvQXbWQX8fLIyDNzPdSVvHvANiS2x6xnEZ4/TAX
qD3fjn7DZS8OyJxkirsxiYxFxTcCSf7UoTRmuaMUBnL1E4p6jkrw5ARtNE465ZIbl/pVDKem9TAu
RM74pK7HGT30gaHhegwxEyTvlVCZSubI059xOB3UxXOty89EZlNZZokm/0I64hbXLaqhJjL84HLy
1nf+4a/g42dprepSDln/wJpOmgBMXLjLILyPBeXpIXsfILxHZL2+2sojD4Cot8ErSn/1g0z+kxoH
Tdxuf/EZb0xPWIA2ZhroO56AyTZxGr0SDBzFkH7cWWflHXbEDAywYMxEUehKMThfk2mpGK0xzOdl
TMbZYz+yDfAFLCLsEh/UsnW2HBkweAimEdx/0I+39lyiGJ+roV4GG9B1f95i8PCaLcrgGGe4rl0+
IS4eP6co+tXqKsb6IwKVxkWdu0exAqyACx+/egeW/BAdxpDUHj9AqPAbCF2r3lpHBkqRj5R1vTE3
gyRsofkCHpBmx54RKhRyFGRG8/lk8YW0xlhsYNiKqHQvxt1RPMDbDyLt8Gi1q777dEtFlBqTy38c
dFCFRc+R2BeXXTgEHXnktEPNWqzfLjWvJV2iODED0G0SzPFKNxRsha7zSgyuCq/JhtnPq/+prZLD
F66iUDyg5ycOD713aEAQx33qOLOtcep1FksxAdCywwCbPirntBFOrANmyFycXIv9LfUCgTC1TMn/
U6kWVRLc+bB6hDDBLoh3RbRc7ar2mc78yGIel/WRsea/rOsoaEUpGzI09xt7Fydp/+c+yjed358A
lbKPT/DIaQSnPGQxNT7qZpEJ5UhcppKnqW/xT2FfOpMrRd3aQD8YCO/13yPN6kE5cRbaQHcd/Y/U
WGYRYh+bBuT2dImCMXifcR6aHIOOwjOid1g9S3d9Ysk+X+zVuBZTpVRNeiM4YqxMHBbK9O+T3e7G
zUGvCU08ysZ3XajXwzdvinbkvORGzsLddmq8WXJn1eZ488dSIl0078kx7EptU47FntFyyVrQ5KTz
hSRmEATm/AlgUEv8KEDT1Lj+5lt758wPlycgdtU77/Z088cffV7inic0P2L8TtviNQh8JPM+2GfV
qbEWOG+air+tls7DwYhrbBTtJsoOPRCEOMnhNeAuT4sEcSG1MtRy2UpTNJM++FUd6ztH557/S+EY
ksHbZ/eY1ZSAMe0qvLIW968U1KofwPVT9Va/+uURG3+KazNsiM4UWtE1UI9CZ7m0YqxiMirgj7M5
pWmOVctYWKsmkB5ctT+JwKx//X7sSKiPX9kptnrIlbFaq4mOkJpPZwD5Q8pGkzw3JRnqow/0wBfn
R4yO4nLeazx/f6okS2+4vdHktJu+JfewH+V/EeW358oDU2KdPwHzLK/v0YbuPOMD7vTMPgN9eX1k
Y9PmvMEnRK3bd9mOWZZ4C6txeO7VQ+U2XyZXIEjz7fxMSHsD3U4FiYHpFXNyXRn9ml5zRiz37HDd
tw5oy7UJgYHc2CweLMpH+ZHmsY66p/RzJ7+ToJD1igBlBBovTMSSCFj9ZxrMQMaepUndHq1uRgze
VHhK7P+PaXNwDzu4Q0uy3J++yO9bQheH5L7HebI/kCUPOEbTl6EnMQQQpDts+9KHs+swoOmvebZb
PN1b6VAfL1Ap7s/AwMDb3QFgTwoXj/qxmwnlA0BWtAO8GA0pqo2H0zk9zzBngquiv5JWi4c6GNBd
f0t4QcjCJmhnyZOLEHHWcg+WBjnMnaoVYVl0n2T74Pfd8UJyhsUDMYW2V1XIl7EaeC7lo8KH52wh
rHSlgxjIUwjkLuwJZuQqMpKI6RHO9tghJ32gKr+en6dd7xQjlP9mZZlKCjSfC7nmze1x9uHt7fRl
ZaAXrzStn2gVAGQgKlYZNLq1K9zUgVcZBekIYT1fs5kduA+Fi2G841phQxzWicvtDQJsl1cXPGcO
8YfGpOpGrSrH//SdSyBCr9LggS82a0tJTzK9TTyepQVB5LWLwuqjS9Gbgk8Qg+Gwg/2kQ0JgeNG3
86OIcrx2X8+vwFzvWGppYosXgDlrOBgphnjSMM211lS8xWuj8rYjGBBIzRvhJvkvDgxtxmmx5iKO
PTeJFJIdfeCIDKDm0rU+oYliUQEe1kQAeINehwEorkCuL4Pi7pa+JsYdkiSdJjabz76wsqDpqCJF
WjKBStcQIgxd8eeE/lkXb2t2j7/dI3jzYHLlcUGy4FN2YmR1e0cjeh8+v05ArW40QmzU/BU1abzY
NUAmiKK/b+PKEHoWP4W0aPQ7F9C/slbDsLjnVJ5yZK0Rrji/PXTxsb+/7a5FM0I0lIFFMIw7zIpP
OAI7nMm2D/8N/+8OJw+XQ8Bd8muNtgR+XPjnR6lXmz3O7NNEXQbGr32oTHsDCHJSsbawKDcA66yD
4ZfUuZshZRJWSNgBgiIKbk2axJYdsla3fmTCF+tcowFkCgwstBhvXfMttGRIPlI1TYOcCQ0tLAOi
1i3qYU0iRNLC+rSNgQtW8dFC2pmTb6MRikwNbiwlwGDFgmJ/bYIko7i1SUUo3bx/N4v/B+wNm0Tf
Y7HpDMd7Yt9oj9sMsXm6wUkU8HALeHDI7u7hwdZekQn/bkhzNOKTKLgP/QDcVtGKP0XO4MY7OXIt
/8vS+BjsrUm7itIlncGO3UCdTj6yucjKdKbrVADxG0U9RCXV5gl88ASPtAF+TV49BBxUaIAfrslq
MTmIn7ioqCFgMCGhvkaAIt1U0y+VaSvbsWlN9Ja8+NZWhx53h5BzD0vfCx6IcR/cTPRjNwliVMmm
rv6XnNb+ACXWOCYFGZzgTIW1A8cz9IIkn0fmebpNc0eYp+TX3v8/g4RLJPfpVMUG2xTV8YkypA+Q
ktSBqw883syoWP18jFZ1HUjBX4V5Nxjoh+/PGv1h3tDTe85uXcAz4hIUpHSWKb/rZdN7VBdtL7ul
fdLLPnPbl3tiJFtodZtMX8PMzyREaHjKKzUx7GyFiGg+7dxT3GTdLdtq/WjI5+0yNbdS6VifrdC5
c9Ha+WH+WVVQjmF/TwlIEMixfuUDjz9Xz0eDuLovow9w0OQDrCWjqli56+LrDCeP76w/dLuaY5tU
dZ9bVrF4jSLsfbOmDoEHN2Q+9SE3+wzmiE/D7thwbCivN5vS/0ljFgMWzBgI8p3mtrmC6n79+Fri
gFNog2NTB0r1MgVrmvXyfQ4zeDvONDnge4gVP+1j9MFhGiOISFJQzVi2N3P/1u45UXzkib+SJE4y
z3Od35Bg7paUrOlD8jqOyfb6KoemCbSjlWxXOzGDCSVLHhzQVT4jMfBJUf9159mx32rOb1BA3+FF
qq+zW8iQp/bQbkqiB3IjzB8IrsDGmYvsPRBXMY8Om06rIjyClBG2uMiHF0KwtQDB0eJwzwiFOSQu
scApGsNJfuUYs0UPaRfKgRhw2LP9wZ/N3aAfL0Qr/sOr9gbsIJzmVBZdt1ek/GA9Fk1kYQRdrUnK
craYBBox/8jWjQNx8ByT8BxRet/c0JzcNI2Zc5/0ZGX7lfLo2g1r71DqIzpNrvgkfdAkqb8rz6FF
Cjry1kZKICqyFhB/+pDbPpOmvHol+5dfWjE+wRAfGeLdJgxBR1wkscOvx6dpvpzQIQt3BGphdvkP
1WdDziV4PS13PsfDNn7cvkZJc9A54ZOcyvGTPgZIJ3f01PmdpJOBLKGT4yIFQ/ITEXleaedh03l6
6brZs9oEsxvOiGFMWVM+2BbN9qYxuMhJXdGoIib5qCLf4kpNtsD9S1h+ZIhmlniv8oKfrpqSbVPi
TS8AB2quQs5yYS028EYgRW4VNZ0jkgeTQX1fgFfgOhI2d9DhZXkVqy+XtQZ+3MPYZ5376IatD07i
4EV4Fsu0ZfKev7M0CA6d08Fh9VEkdIaIfOrA7OC4zJTGcb9hMVaSDQkCSqjFNUGlsieDvT45gfpN
tXlIVvQl8NFRz1BBXPXw4vlvMaK6X53VdxX5qeWB0J5gU3mL6bk7uSZaueZ1xbhaqPXUP7vS7oRr
28QT72oTXPD6NHpo2VZjttT8mVerF1RlnXkX9aEKzYbYYA/9lmGS+HdSTHGQu+/jhjhR9zeFJFRp
adPyH7qrc8LqMBOMNCbS+lE8OJsgoonb7//RP3bp2Qgy2ByIc4oF+GwHS7tbOjT/8Sa5A/b9pDdZ
Pr7sjsmb89zn6cjZ/g7g7taZh+zX5fpyQ3jf8S63qXrddOMT4wrojKBCmxIKmV9m8CXw8Mu8DXWl
nmjvmaXIfyM7tKlIt6ZPk6azt9cgU+xj0Mmev1h3cjnL5VglUFic7cyMt/4aRM8qaVelQYELedoX
rTvgXQArzFdj5J6PMgvQvn9dl7C9Y+AFIr8w3UrKMMSsaNp92tIZcMABh/S2AMYM1phMdjFwjmVH
UOl15TFji1QEYSEOxHSnAg0jk+fAkLzwUj4oRR3NmOtvpix1alTU14HlWdgrS7w3zuaZcL7AVYLB
k7ZLpDsLat0Wtli3DC75cxlfyYjqwvPoKHgGoclDfQX8hBXj+teH2BYqVo5JK/jAMKodyJ9TIdu5
DFAflTZh/m3NfeV/0xePwuQTb5qE89MJo7Mb8gS2KPSlgKYa98CyBQPaMiClGFenq6U3kuWx7Wjs
QRzA5zQo+GV+YJAXL7SF49sD4vvYbzFNMlDu21x+ckftpE+wwV5YgvcO7akXWKEVurmcKI/mP5Cd
WB4HLFdFW/q/qcopihSB5H3kP4h36b+jUoQbzGHDDZAuWzAR7aY/2SMazUfOrEhlWFY3YUa+2trZ
s5gl4xRTt5SJqwIBdLjDm7fziHudIL1dcDSVCVXl7cYV6XZ5c3+t0pN0rpnQvZHbJs9Ur7mDNUa+
TuV+SAw52tuNjo6CilbWcxu0flimKZykSSYmRhw3lZ6DxhsLyqXiuVs3S0RpQmmYDVOL0+m0kuMV
wgIP0V93J5+XH6+vQfmlaVOOsyLXU9/qx8QfMEpIo8VUPCG2zDlDY6IWPmXqYnsoBaTA19uDbxrz
uXunNHbysy4hYJm3bHv/pzdxHiy7/gZX01c4SMxZ2gpxSYpmN98QS0mx2Y93AO8vpxTZ4EHxPEhF
GXNm95lGZwJy6l2im8l3YJ8OycJHD8gAK8BcOcaQEwe4YPva2zZY9gv1BqgjO/Er633+RxlqJpuC
L/vuGmNsII+PaGxlHAT2rqe+rUQEudKWXxn1YnFLo75KUNhZ1eIzQ73SLLM1ZG6mM63/JLgMrMoF
nTKBcnrsBHj7Rhld8TcaTkmFb9qSBUFOVqy4lAmrW9nB1aOSEQGPnEwXhgUgX8brPkkHn9BY7IcP
zi2D7VuhMn32IImtRGW2V1XXMPOjsQarBoK0pn2oIcDji3kkRpgjRp44ue9srytflQazAf/QZu+V
RaJ+QsWpbKKwQsYyfumzarrXNMzbV32yGKMWaJm/HgGe0iS0ZltJULY/TNoz0MNVoCZIimYT+TD/
UbTgJpGmFDQCVCuJBT3yeIBgzh5Ebcp/Fhkmc2NB2H542WaYsOTkyEw/6VxlLdWkVfrelViXNcnf
5tmho0z4JRuKzj9wYb9inL3wI9dQkDjL9qnf0BFY0bNom+iXfdlQJKE/ApttJ2wLHpKYAI5KhL2M
mmt6s22XkEaDdRzqXqFO7iMQODVjuRgxv0lQ68681r9vDEou1NmC4TZKFszzT+SXDgbeQ0BoimU/
uk/OJodviDTurzzQhftUBT0uDyw/GDcxtW9OxtwXy4/spS00oy81ShCVMLlVki+ceoYaA0v2KmCM
IBlQCSMjYwn52OZNYvXMDKyhitP4VB3jqsOFK3wvFTXbH6PnxZ5ob1E3GTUWZAAZ1eCPpsadHnQB
xg6O+RWee6p3KxsSNErzRqQVm/zqEIrz8WROifiOgu9JJXskBaa+NIdDra6ZTRohPOtmiQaWp6D1
Psw27H1L/VKxKWdHfWAQKmkaEIgt996N5z95KUEp/e7xNkKkHCFpu4yod3I+xNnTjluJnxfKaqm1
trFV1EJWOjBmFLgJoZyMYFAYqk6rFA6eQ+AKBN3Scx1gRTeOGgl4IuQ+oSzSXLXnrK2MQ/H8qql7
C3kJW1LwPb48vF903mOIINMD/2PaSKMzd0drhNqc/vTBvSkNm+h1nijnpWOCJ2Hp7pg9mUTL3uM5
hpGInhYFyVFv8r5MtpDQJG5nXjm+9wPAqFwysLH5Qe8+S2NBRsRMUUpiujAau55YepEZVoNSRBX5
ata0qwlKTbqZnK15hwQVMCM1epcdldpfW9TfW/NEuqvCyWeEh0DefaonI+ltBdR/KJ1cq3rBXb1Y
MBDp4LBSCaWizrSxpEMi1m8L8iiRQCutFwbdP4MEbom06hrbOsGcgGyAPgemFbI4v4uGaVvqZwDY
7BEnLEC3Shh8WWkmS7sWOgFbJLjPy69NMFH5eFlovzmYDwqRSRa1c1KUHf+PdiVtjHY2DFlJ6drR
Ir+v1fVXPYsJ/UGQxIJuGIe2xE8ywUU+2jSZ9qJUGd1TVS8MZmAAdygjoE3TusMw6Z+DeizFspwT
QPOsLq+r4iVMoafmM6GEMmo27DI1wvHc9PybSFw0g6M80XU+8yohqfkOPa9lUdxiswcsY/lQh6vI
90sBuXQjU1+wg1QXv7FIbR+WhxTG4q5weoDFJ7vu97XOnVas/UBLfuyYluRpm08TptNIk2GX8DwL
vO+6x99BoXvqZkc79mT5LJtGb8IFXMe7HeEvZMOEVjvwUR0uFIOJcJdu/d4f6s8xnUG+YrDB3NZx
lQ2MoKcUj1L/poBT1eAvvRhcgWLNWAoDEawQSD+AK2FCY13No3zGXNXfiaAeSDShBUmlWn0zsHmN
hUVZhD1j8Q/68MORw+48aAzEJb93ZzOgNlJrBOW7iESuQfFPDAPrfbpSsD4q3Vp5TyWXh4LgUltr
QBuXYBBYN2C3XyjTN1PJSYiCN5jLdaRuHEPlO000fFn1VmrVOPmZc42eJpM5J6mF7YTXElsmWMzq
JpgjTxwZEHVRKpgedyphTKHsd1AyrvGLcYzgKqffSABdlzLITn7wa0JK36zqHlZXmkVnywLKVwF7
jl2rkunyAxmcvsTCkZSGkvGN+zYL4kTrXB2Li3HzzYwGJZhN7GJEyUyuLkOYfFU46tAe6rHmcJga
iw9rK/oFVcy1xpBAE/2152Ncj/TkBa8TUDWxFt0PQBcij0ESfiriyjorbGzbPWkd4xmXH4I5+Dnc
Aonsl1MxiCCkMOFyK1KWimqA+2fT/bMaFSuTjss97U8J+VUFETBbi840Q5an0mTo4RbNqBfJjNAM
7HsdduOgQgNcfjpzDc7VTYDgcVx+proWnVjrarGduRpnBlgD7eDy6AzwpjTcs7+oRfrzv+549vTz
NybzxTbwRFl22SF2I9udj05olysFgEz5LTyi91GYC6yfAU+6eM+epfQPC8gNQydGg64WAjM6PvSl
3ul+ZjLo5NbSMsChNrJPCKf5o1cm5zAnlab0QV05MPPWZ3oX/eO8QplYB5O1i/yNR7MFHKHcQLon
TvwRkxLAwUVdfYl0P4mpj4RO1JMDkPS0tEUTcQlzPS7hVFL4REcNjHKcsP5EbjlVd+WxOlq++BSn
5Egy8NBN5Nx5OOmcC+rnfBVAyN4CtfczfGmAPVyb2EoVPRYOJ1FT5h6DNoiatrRTdHR0C4PDXebF
0St8DAXFwf7/PO0CCMjoy9E8sNjHGXjb70o5APRVS5YlyPhuF7C+jnZ17o0hwnOKfWxV2eh20XGP
F6QXglzyMWoCNrcqfXXkVNMvUNgoBwrxJqiyswrtlUguaKE8Hsiiyje/bPwXD+Nl2vKclM9Aa/nj
4S15qzi6Q5Z+5Wc6f1JXaGqrzfqmVHFk7HqKtmHY4MR1vnPB6s663+xhA8vCAT4WucT3lBddl558
KQYU7uhLudj09Roy44LFB/rvYi80vBws+p0tOvVsIHty5VJMIFqjQltP5MahOP4PN8Rva+fvoHKQ
N5m6ml57rP5yprOz6YlI7wsVhjG87RK5IawaSgancAsp+rXgarqnuAhmFdgeFfqCHUBqMJq5zWxu
XrVFNHDFUshGSPgKeFzKFBzTeOREQMruje8zepExhNbwMnx3d5nvO+q6jDgpSwwpT3157e7QtZKv
Xz8vvA+u+KuPDbNoMXv1YELAM80k6gLdLcYB2xGt8kk8vj8V0ZYi083UKph4HbNn9ZUbe16s60PK
4ExJBKEwTjBSVdWUIUBi1AyyDOELwGTYHdda5vnyhOS3Q5wt3KPyTloLkpgWLORqxrlSAob8fuHj
zvrppNDjFpMmPosH0zpMM/5+DbVE6PzwHWzSZ/k4KBPVgH6BgVhtKnxxSv6VbHcIzRB6lZn4tjLu
kfkC8+NwPjbYlAcGB3qPb/ZaIoxi9xtyV32PhvvFEIwvENRNg7972AA/SAKizBBCTToDbOxkPfIV
6+ZRtZ0CW3kM3hhfkpMSh7/GoLc8Cc2he5JHWtdyczs8SleNXRsMGdPodKUVX1iA3eCPDAOdmIEt
v5mjoBQq7DucF07UCei1uPeZaGl3/QxmJ4lutpQQ4po+Xwl9tYolhJz/nNWy4gWXtXc4A8ycRmyO
HwRiQiUdxkkqLGA7YW0UPSzO6PgEz7AdDsHSnuN1SVV6EU8IVXVtxKa/C0LD5EsTLjSW7II49aKK
uavwkrHZE9aaKgAZAXIQm0uqKW9AX6edJncs2yhNLixcM6TpJwnDIqsm8K+trdhtGuxessQUkCIC
3KyS03b2unZSwdbo88kkSJZvdzwJ9BaeTrLVxA16jWRLN4erhNKjzt0qqJ3Eff0C1rbRYa75bDFG
4JXtqJ6WzQyYCID4N7cPSN2K4GQRDVB4iy1fXDfEXB/VeHyOuxyUaGrbDEMibl7yBclsjYl1Ndzg
y4EB/ypzOkDM71BrFXuJTYgiVdkaMXginHmQJEqc4SNvTAZAqP1wjzO95y0wGp+iKpaDbSzE9m5d
ERShvaSv0xWAxdmKccr/UEmorz0gY2p7z3sR1Uhrjst2/Sk+pNDvvDgN7E2jTFkhtQsvMsgq4zHK
Nk3P2veHYDdD2lYcnm6XvBV0Tt0Q3Yjuk83KPaix6rv+1bZ+GzGoBOGmRRWQ7bu4t0pYDEaiM4tC
TKFSeCd2gFtRyX3zs40p+dBLJcx5BsK2+KCJf/tptX1+3DmY0+I1HD+UbSkAy0+e0cY0iSNB1cQ2
QWPjKir2A3aEAl9uIEKXUTfHwYg4tRymJmHEb5zbnHi9JIvxO0GjWqyGhCzJSFqVJXOF4sjnGhlL
FusLHcC+Kmfo7JnBQI71rcKn7iFZpCYwE/P7Q3NG28s83iEty5SGY3TlihwW7VTbuyRGeJHJpDBi
796VK1/JwJkM9YwwP2MF3rRL9m0Pxa1OR4+00RzAldda0vTq+vOKP6L8EnBiY7BS2dAOEv1MFboF
tDKQ6IumFo7uBEgInsjdULha4frrAAOw9B1CTwt1aSn9RfJ5IdILs9hjj4MS+/R7HSk3IevcoGIp
86U2GjFsHWnzB/iv6C97Xtw56ZIYbfHB8Uelov3OV0R18ZeZcdUL5D8W8Xf9gDva5ZEpkLB0pICF
Nn52Ee7Zpdp4P62xhyKCk2Iz1nSVF2YP/9+wgLRieTnG57V48FgSWnha0H6egZHVbK+LWRWl+0AK
IF3rP5tplNtpSxP7Hdb+K2rlWdanYvuotzYt8v0HQZ+InDRfnwyaUacomE9g4brdAxedaItkalTg
O76zcQpqrYZ/8Afm9VntyTMoxmSX0OqFjOskW3u/e78LKgyNpiJUf3OncqidX0rslEoLGM1cvZ+i
dKQsm8JQ3ciZAj2LUtyVgPWWTLjNmok6+7BS2t9+b/g+FAm6/zRsabA/jx1Tzd1DXuO4NxTK4SWT
apcCn5WI10qc97J4c6lnVinSeSx/zn4XCRqGVkBQHSgYK/vK1gJiHpDrQRwiFrr7ok8V9SqOQRrt
xuvGPeywI/xA+mPaFgVUS38TFg+pmNGP46KHhAKaM0YSmdx+mwk/QPIhdFWdB7SjphM+RPTrf+ia
hwUzcxj50IWejNgQ8vwzg/XCinpUqAkk3EEjLwqIIaBgiidUumqjrU0DM647jRzrBK+OuWYMECCB
y5yEQYzRVY9FV3yJ+a5rrA7+rsgfbTNe/1mQTlHr5VRH5g+Kc6gvsjEgXjXGSjMznJikTVpdZVxo
4x0QUPJB9B1USf57WgtB2k5RTagO8rgyCbWyLeRzE9N9xpsob/CA4ZYjDEA4dCEcYH0Zzl2AZI4w
b4gbUoO5OoRfl8vnyEBmrjaP/StG27rnjCamzrqcViwrq6N3ViBFGjtrN/Gvi6HfywHA/vQ6Wy50
4DIZPMr+te8ny8cqB9bDM2d/fjS+FrJEQEvwQwDSron68UelW9SLfNhG0CGUXqm/0b2K/AwVQoEo
HYnKFHIDP2jFaCfgILl1GNDsoefsXG5yvjmDy04E4oCSNjQ/EZwvjG5nzcdWclGkNl+7k0SAroyv
jJclJRt81wTwu0k7pk5ufjahji/lXMEZEeBa4mnZ2Po2D9SbE7DXTqsJKbTA1Lcet3RuUpAA8dr+
qf+WKTsQdBhJAx1JMuyGQGtycS3ZZW9yZ72e9WHn4fOw0T3+TLut75T2o3O3fj/oXcdWObU+6IsL
vjHkf7n4+LG4kRU89n8AAu27yX0kcjNVr+n/PhQCpYrjp7CS7IY8VNYeynwT0pcIUVhXOGiPj2/j
0NyWk6i413csLlPUS0swo+RJJ8En1ydtUiRiTRq9iA7u6/FnvIz8OTN1iUnTaQReAPsjOlBf0x1/
Bs2Ukexhp/7eShvQb2IhXbC/IkKNU63jJQAEQUFYXVvQWeu3HCqMXiPP8BtK0uzDbrRWmRjuxtVG
UfkZ0HZrYZfAjgax08JPNcgzQm8rn1zFJ8bIS3u9PtPihxYTQVgYkg4cobt0sE+Nao5tliX4wD+a
BqJISveamPUrqcD/RchVX+mQ5CSXEAKgdTAu1/QPvhRdH0RJnXfULm0X1ofvR+xKOV9mLkXyBdBT
iPbH1eGrQJYVwADAZ04xqWSdRqdYKvGMoPWCKkdEf6UCKvaDgASb5kygjY2eHr5k8rbmc1mP3oAp
zrPDWI1TPM7/LjDy4VLKBL0lRUkOzfse2pgEF/1sJvzM6tAvrHrp2hYTAHfD9Uce2yL1aXomKhUo
Dcv2Ut1buy+hj4ZMOxRCvbbC3pK8okA/4XP/BWBGUvDxJElRp93+X4Cqc3LSEHmUDyntooZMZy23
rO6sIXL0+0F1L4keCQqUyLssqku9/oznkSjgBgUEcf7MWsEk/6hH3bnnTMj87iQ6PjzCTKsHVzfL
Hf06plTOtsYJUJ2437yVi2Im/qv1WXN19sef+lFAsqMznnSulcMuspw7v2a5Me4nVeu44ipcq4oP
B1pu3YOt3MYM0JmTPnXe2WvwY4yuANyTvL95Xa5mU+q8AQgineq3dyoVO39VXB5eJdPHaOYIV8pD
lJ9A816VCnVssa5pIzvMcatKin2eHXKlJmZJueSuHs1Ea4BxuagYpsFg73GHUKF8X6bUBD4sQ/pz
fY6AliSktjZY9m0/OCkfPqF/Feu3YYaUZ/OLAiZlJLGzYo3VW4CO2mZjPuTw4sqs696wAtr9ipW2
lfA/QSZZ//SZPNxXVHipLwDpM0oaiDhTTc2K7pAMtXUZhB/QUTtfwx/8NhYs2vwFWYrUBgwUwbD8
UqCgn13bmw2E2DBe0td1zXOrpMygNCPd1OO2xgPAfsNjxkbTUFeBgV0VsXWVVu+st/SQS5aaTawb
S6WpxxvbUPjawAc1K1ibVamWiJ7vWrVzYTsc2B2zT4VlyjQxQD5z2aiYFN+1WeLv9wDx+4r06k8A
yLXeeDQ0TxQ+ARWTiLqPmtSb6SuXuT/flCzM0pAfQpacwKY44HzANduT2Mhmwed1S37woq4xLGUy
bkcW7xLPKw85ISft0z6f7tE+wGVXKloa6iaul7OrXQHXpUdAjQLiHvPGUlP4gAIpTzUuuzhgekJn
CVfkvb3geD2z7T4+lxuoPo1FpOgnBbyqt2OOyYxv5xqwZONMSGNu28GTExCp3ihhpxvxK0IYCUJw
Ci+JqMi3NPRA10iANi2AFOlchL5hqD2htc0pyA3nN+8Dh0oMGFh/TtFf+WrSeoOJBgBgJbHw36gO
DdnI2e+7C5LnsyovNJQNHPHk8P/OsRKj0auIEaam7znMoLmnVQHSJW/JMoEAmVdUXEGGFkzyej2V
UvYje5eXIuttLOpN07gMsELXcjYkf2G9Oq/MHFhMzcipAdSXfswBEXDGsiPO0iB2xTRhcRzGo96D
8EFFcR2wDogt80f3aj/mnfiJ21bx3oDZeoxOLQdVP6DIo8aGNQWphig875rRMp0fSOejLrudhj93
7UwbTx7Z0bKPMRAvQXDqqvdY5wc/JFVn8O2rNK17xjCQXWi6Ygr+LXRuRI1e9LxD0i5xKfHCaTMJ
Bu/uKhiLwYrDf5+GLKdEsNvK6CYHHk2/X1O95rCdUxozcbrYzqNkm87vF0/AEtj1FAG+SzYnXrSE
UB7lcc1/sl56EuF1lo36GkbfZxnypyHwyOC/Rc8tMX8f93li53T8A+zMPquouJcI6DGYP3q0TqHz
AGTeeiGWOBz6Fn27IzHqtH9wR/L+nBI7WyNMv8ZdSiD8rVFywHTgsDyel7i627pkSacz3CXo2wXM
RViiaCKfq9ShHyxdeexC1Fj3f9V5A1GoyZNSBtY8ZcBYsW+rSdYObJZiA+HzmCyzFIS9gLNF6Y51
IKQ1MJU46H8olcRnbqaLYrKNVEijIhVM2Ye4pZcDcwdmS9GmmxPzqJ9m5fd2RNdbzBOeUvdxegrT
AV0RFEpqMJx48twq+gCtXVmi9qOGbmwzc5Z+Ighh6TZm7zb8fXBnJmGTjQpt8sPro6ubOgeTf3h7
LbvtkPNQXNspwidZqkSpan3lZ534/a3Pthc7m66D3hTSwBCE57VzeHXQ7U/OlXVHcMRuZ/AGYOVf
JWq/xTvtSS3iw/OyLWbHP5zDnQBsrkJADCvEV9XazrvbpQWclbnMStiXMd0X5+7M/vUV4f4EkELb
6XzViqGq+Jx9yfAUqU2eVB9U8WFv6mjm3WNGj4WsEKxHSv8rmo5H4CSRli1W+RLElTzPVtsles9D
v0m9gJRlVUmbucia2kMosqrLrQMtbnWXGuC/8YZwm5aPdgW+A871a2XuoJObqo8wPEv+OVW/i/pa
ZNsYUvIY2TfETp4xbvufkGw+BAMAYmuOXZYnOgrTFwLlfRV/A55TQI6RgbJfsF0zRZ329iWBkVqS
j6/I1cBGTlqJtkMIUCib90+OGL3XcCptMiS2jq9u3rji2axeYpCwPhhUTWm+Z5npG/DBP2it3VT+
ESfogH5vsQwvhvsYxzyNCMNJShEKe+9HWxJ5OKpV/RNZzhL04hqEw44CgRgsD9EunGlDIzxoW3/n
97fvgNnee0U7ybR3Dv5LhQY3qJFtMsh+h5CuQ7G27ZVzi8Od9x7wiWRck4b6UT14BgDQ0+0hs04r
V7JV1a2YpgdjcQYCxO6qsxSycK+7+4SL1SF287YnW4zobNKmsNTCz3I+KquFokF6nrUM6VlLfADP
3XsX3vPoQ5AIGLoZ0yepkw8XcXdLVAK//m7uOJkrs5N3zJgbxd5GuoVQbn+6DqhK0bgNuyHQeyQG
DrP2dde8i2qTiXQ0J12ehj+8wFIRmzbfLaRN543pa3d2r0UlCf8bmFUz0NcYYaDjiVnIv5Mkaixm
vIfy+DVhH0asChrwVHEFNsRXeq2q1g8Ea4x0yNua/16kOwDif8O6dP04AXqFOFGA9S24/wsK+rWk
nQtLXXCs+DCjSq0zlNIqmhN0+0KAMz1D83mvX17YgQW2WTM/GMBOJi/RR6kB3l8/o99Zylz/aRDj
nttQL5f0wrahB9ChJRvxbAMy+jCNfJMDJGEGslSjUw6Ye38KXR5CRZfKidmkMMqT0bYoEtJSbEWX
N8aqnU9vtvTpct3k1NGy7ILmnJwfxUvbaqeJAi/aqSP8CfKKoJUkUYL7wgafmdxweM9VUqMb/mkX
W/c5j7bZ/XyivgdbNt9kGKSKK4lq8rw+MowGUmdVMl10KVauTFeKWMZVpmbdeayHrdHdftESNT+D
B7awZj4ZrvwxU0JNfPj9gS5IfkECSXeg9E6lG+Jr2/v9IMJvW0g7X9MG08HrDkRQLYMX34JOe7jt
VLGUxII2ijRXtV/FqYIl1237H59vUyGNG1QfaU/GHLKVB0uDoU4meizlXQbFly0gplNXodi6+dII
rfawumEGxh2cVX69Ko5BYBNPrx0gJWrzeXxckLoijXTeXNIA0svdeSHIh2HI2r+49jBkgLhqGlcG
HWFZ4uXE9YWzyMJqcQu/02v39va02QDNkMWFw1orcJXkcoFogkoZkC69K7yqWA9uFSspLmtEuy5m
PDTaDscJtGDO/uA2uxfRrRccZ68q7Lb2j29UO1fL3I3098umylti8jrLvYfuBQGbouCVPKMKqgEt
Lm5u4NxhXgORHIbH3NjG0rQM8zh/uxyfsLCmL5GNTn+qyTeouzpqHlgtEqFCDUTHh/Nqcf3MdzaB
hoSg8wyFk+5nszOoeXEvrbNnZSecXca9QRSg/F3mxrw4MwmFGpJFJ3Js+/PHc0MhoWA5JlESVLVc
aa0ab/xR6mYHCgf+h9bGFT3Up6U6j9d2jYgW5VJPOG+vBRrmiwQ3t1BHEAKu4CmEInRma05uVt/p
k/qKyqxkLhgxw9Yl10CVlhY01pIIOsErpIqDoWOd/I5ALKcb0D78HrAZB6BIVFZ3jtcvD0zboc4p
ECiqqmOODZtDgalOHp8KZiduAvXyvg9qhuF6OotEsJVKv0XqTwxRhmuhTta0LLRMAPc8ufOdAju8
XYLNMJsHL/hvtiKekm9RLlo7ZVIldPMz+hwSFohYK8p+Nd0EhLIz37m2qHnssnYNV4hG071rNIBQ
Bw0lz316JBU4zncVRjC5AJtj6OgbxI1leqQJ55SnDH0XW3j03kzQ27kyJZUVfRQWMSEk0DdlUjDI
INmlHdroxoni7HDT4BRxQmceK1uUOFB0wuWPZUslPhSbK+53C4ke5JDnHdOtlHuY9++ayOkmisPy
m+v+Uv4m5rQFvY7nOcmGOdhvdv7vVSS2nlsbb1rKbzXnNJJnpe8M4cU4NC+ilBpt5ir3QyfDQDPR
J6gx5GPgngXX/o5F12iXtudAUeHtIomAZtC25ciIbDGQv+8Rg+yECfOZCyRp9ieHGmuGqQbG+mkn
cOE4MXDv39qjeHNBzvBVntl7wwVyIZvSvyGERTDSkbjhpH4VYoDs/KF3RnDPySbC9VypoLullJW7
GOESgBsL+YRiK1+XjcpRhxbSg64VepQClOwoPv5plUwAcG2XuYqu7gB6JI0ASwldOme3gacQ9GXK
jjR2v2Z8Da5jrBoYVNm74pVqvOb8Ej8e7qGhCQz3egC8dkLvtvys9yfZQECU3Ny8JSS04blJDekN
Cgisd/LXH49ztrqfBx67pAISDOXI/nR8d0Qe6KA9zAFZXlJ0Jrj2HAG79KqUszyxFazhG7Tuqohr
4Tv+dC810IZgGEBV7y/z7b2kiLea4mIlGs4aruLSI2RacvVBVKV8UM4ZNn9VAFhUmcDXtyrYttM8
I0o/Rz7JX/fS/DAbU572mwyK8hh3sShv77uOEsmwEUkVrDatFpKdZJ/DBJQHDzRHB43sEdU8KK+m
QSD+L6zB65nDAhPa/2kmQ3DX2SVpDpnHHr4rMn6Gjl05hj4rqaEibsJgHdoG7MEYYcyqMdAQBbGH
2g8zY5EAXcb9HJkqI46/A6VBewpLaAt2kFZr7e+lQ5WBbsJNGy6Kb78oCcknwUSbXIoi6s2txR0S
4AHYNqbPf/wBU0Jst95Lk+iJ4C0hDnqET/XhS2WhUZ2M7zTb7piFYl9XCOpVtcJS+lxv6wBBnLIi
4eIMsPz1pwjCdW1q3iAcoiRj4HQgrHoYYpRBLV2ViXe0hjR3ROrX2ur4FTTFkVacQ6SGwSg1PNSY
rfnDlVkzlWhMnjw+IuBlzdmjcYgtvKGR0lS1+JiWo8GIICLbRTVGFGmXV5xpdhG2eAKcqGnFgIP3
GxCydwMWQi57Vvcfutz8xhjM9n98pVmz5KkqjlG2WPZVeSAffbDuJMBLBG1m9o/zlz2iaPGL/2F4
VsMrWs8E/obCvpUWU8NVI0/Z1wDCVOLDIbXdBRoEcKGZW+a+xz3mnaWntxyX6Xl3shCa7Nb4W57P
CqhTnVsTgFmZfX9a4GriUyjFeS5oSw2b2AbW+ApbmuwoCcKxC3taGCJgJdNFZELCZBgyExOTRGE0
47EVZPW9sQzxPyoLYUeEJ6cZSrA9DS2yQYB+gqlv7T0PGNREVaGid9kF+F7HcSlGRScB7Fqggqzn
FaANam4QpB2M7dTUg/5MNFB7nb0Niye16N8lljtn4zJPtKcN12ToCW/0s03qsCba1vvc5XIFwAn4
9MYlU86OFJNLjrSuqJrWp1O1gyD053o7gWNIo79Zm4n1eMazb07qZr3HLyYk5j7XY7eqx18xL0H6
W1pjCcjU3lYfC1+PiYmGbp7kpVlnmLsjSWftutAzHz/+3Ua48TLE8qhrP+4AlDVRoe3rExlc+wpu
vVarbiPsBu+HjfoBMiqvQr6cCEAyoQLP2leTJw2lfw/hVf40NeLEK7Sc3kHozQRS02pgxAdbPgy8
IZERsa5pxP0ZBALIGUjrrb8XUdVOj2Is6KJBDAXXnK20Iuw99QKi3cUK2ka1qCpX7HCU7kpuvPGW
3l9JhnOlNz7cSh657XwxnlZgjHQIUhRJPYIF6AlWACXY9lJVyqZRpqN0F6Fv/QNy07PbCAjsBf93
kQ+s3Fc0NLaT/Yhfp8s4ycuJiW/sVMtDYFIDVSq0AKnKo9BBbMJo3hGUnB1lZOZJ+dZqEhdUbF1n
2TSMuWQyr+o9mwFQYcfddej1WKhMNXCIQnUt0q9g9EsdjaK8ZvugY6KeFI6gSb8Tdt6gzp9DMkY8
XxMLhXNG0RvnsBidwmEpQKc4dXH2KGg0HiO8rVK3UkAHd8qaUFiKBpHens9mIjH6L9JhJ0JKlV2U
i88r8jTkP1QgdPu9OBvpy4QS2mHaGWsALS/+XuSjYWb59CUiN8D5pelt5Sra+YPY7k1PqzUJCuQD
L83LdWUb1NsqjA2PTCID/HGBv4IgVwJHYSzfK/DACv9+kUlT/hIqa9S1FalmHUpyU2Ex1DApvi84
rlWRvKF/WAToC3gBVeSWEs2R1Ki2buFC273D1/FqNXhGEFJlt5bpB+jZ+w4vvvW+S3SyDDqptGiq
befk0cXB9wYcWB3GXaVbjT1woskhBS5K8WtRA4TLD1Jf7xaXMwyDWsEPjVmEwsKgJmxoQtUx2wka
042xs1I9zO5sMfEW+kPMQ0QtJj498oUaxqsp5sWt8jXB1I+ippDvQE+rgDONEMX1/98yLVYg3/rQ
oJuHQ9xLWyBo4/yI6lSYFowYYjczW4REOZrUn8LSIYac9enV8zr9t/oR2QtjoUsdKMSrJcCbciAe
TcKeQesVLmNJzyVe0V94/eQvwNOPNY3keKYF172PvF5l4Rj6IlNFUk07yY3kpl5RlnCwBgfmb0Cd
r/8yb74Z4oR22mJXptk6V7WdrUz4rvnt9q0ZUIMHdLhQliBGu97WMcUr+hRD4tRyrY83VdDKAwt7
5tOnPd3ZC81TKLgu9ZEalymmu3G/kj3scwshD4xCUyxEjhqJ+eBs6lNIKWVnfc3qdhI+yjXkyphK
GobUbLvIq0FNTmAfN7Wu3Rb1DR1AYvu6nALpO/1SPqQMWlzPZwJt2Hlc/Bo1WbdxlNwlXhg5UHXW
i9FtZ/Juq9GJUqmyYgalJC1wU1AhAXCjIef56xN5VwIAToWpZyp3VSW4P7+g2mVODFayRDyEOSt+
+bsUlP9fVtX4vLNOaq6POdM7ZiOSrrEqQyaCYTg76pfISE9Q4O5ZvAy5p3PegTf347GZ7Rp367fF
iqX+/kW6IgqDoq/rcDp135WBSIGsnS4UPwb4Ny4wdExC8Ouno42LqU5mR48lVnifnofFHxQDMylt
Qgt8x50CdD51hzq5f2KrtlNh/ijq9TAAoW7pg7kdWncxS0TqkSp5Szsjt5cmsje73eoCrtJSptxj
5j9f6OdV/1IZelOZPc5XGpNzGYdTcw3i13dcexeetXdRoKvZxAcIOLD+sgiGxINdkifnMmBbYUeW
CcANVGbVYUpOW392CEvTTBiihn5+EPGbtqlvTQR/qoeeSvFxRKOUclDp43Uafk/CRwP3FqPTxkb1
79YhthQMyf1n6DeTwR6Dv98Gg91ywqFbhE7EVCH4yXjJE8aFhGl6LJwwhb8ns3Ox2UBIhP9ZxyR/
PmC0BfOfwLk5shjqFnFHEzcGiHQQ9lj2lG5Zne3aJwnji8brK/36g51WPWiN4Uy3AixU1fN9O+zI
RguUJ8EKOZVXv2rHc2S48kvWtbLEX1ukl8ox4xDibEY1D81dLOPLZDOfM11DH+6Ou6Znb2qLUtbu
CtKCyOb++L7v7EWSA9MYr21aDUDOc+wXxm1ONL7dKX99a4P/9XbCnkj54hrXISEoH2oQLAl6mhp+
4t/n6G3c7UdsTrnba2t9v9P+PT/iU/n7SjcfN1b6DzYQc0QQFjGR8bTkDCWRkfPAceDZgcEigGv/
BO3mPg6/J415K6EXBIWN4GG5x30ZQcfF+K6Cxbwm2eKbnmwm3Hl+/PMWPDKyTOe64pzLd8bWbWLF
IKT7DdvgIFq8Z47z/+GUnDJTlakxPBhZ1ivxV7xeyBydIr+LMbW9dBY5/a8u9eg+53JM47wF9cty
acgBnlSYtPxan5oZCg5XNGxnzBs4O2TLZgsEPjoiEwzEpQ5bnIIIzG724JHrR7SM5cUUP9+WUvpB
sOvRvx6Aa8nybNaNhGsi24iOvuXc6YpwgwyHJRyO8IHVwzYtRkWgnfWkOHln8qEJxtfJ5FM1PjjL
rZDfuQclnYfuSWtt6q/qGeuCZiV3ajSe4x9d+m2zJNCFPlbZ+66rylcD04v7T3DJzuAjfhiAqm2U
lPQsWi8xNS9/di9iNyVp7Zu0rvLbIlxTktG0RC/CXxB9rcm43A105ej/p2x2SKvAD40RKPhfRKdP
Ec8t73eARb8i9lJiCuJWXea2cw2JW/hmgad6NIQ4xsKeMyu1fcyZBD2TIMtuSFjPyjyo0g0qXQT9
GVoWGAD9NVy6uCO5EhdaIxUSoJK+sYRAzeCvPMiwg3E7mLILV8b4g6taJEp67IqW+eYxmpsz0/V2
hl4xZMzehA53ZSwg/ZWqce5B/gxeHyowh60IUVTlt939ITNohf4Bl959SIqoOq+wwx2wN4xlQpPH
/0FrIbnHKInZjkNpvEenouWiTsj49kOpJ5b9G6zLFJiTewfv0C/jBMIHpaCC4iwkrapThPK6pW3y
zYKWLXWJfEV7CALCs7v1RWCDqIfW8IGsMraBrU8PL4iqEDkGxETAJwIOa+/DCxO9ZhR9Wtv2xe6e
4f3z/1J9TfFbKOFepZTCMNwa2bJggeN3clkTRxbTAxHW541v+utJd6vwsMgXtdWj6rOs4wdhZCHe
y28egfVKp5ilhHSnRaJpwW0PE/Jjt3HSxTfquu2aDGiBFV776gqjljoKrgHuGhJkO4NYDzmBxE4Q
ifbtbTN/9LZyrggjuwmM2ha01R+z7RPBst9sVrXXnsNBslUHa4ZBZMmBrZfH5Nq6VlNzPpwkAjay
1r+LUbh0TiEUa5Fq6X+0r270s7i3aqvKXT/8UdKgPAOxJQ3u43pKym8aSMHs0U3R2uwB8jNC/w33
XnUVvYKKeqI3Z1frwC/GCBSaBxIjik+1BXpxmsngz002CQyzD15IytiUe/OVWohJFf5+RKStDIRb
q9D9zwUXv5azMuyYWapcwztNdFM0YXMrK30sGPPlkfzQhm/FTwpBjf9cRC7Gcv4u6HdNsOyNxZ+d
NgqJXNQM/55vHxXNkj+lXvzQ9XKm5gUTq+eMzv6p1s23T8MRlvXRh71NDa9eATVM4CTV8eJl9G0+
SI6mNnTy4Qi5BnJH0iFw2dVUL0JNnjNg5bC1+pwWKZbCHZpNlJUgeMmSnN4tn1VH/c1hyrqZmf9d
F/x4adJgdAq2JHWc47EUms1qqbEsrpaLJlfAeN1PRgWPBiKEcl/sxvH1rHyPhzb5nF+XeAcNh1ZN
aPj8TOJGRll4MX5I3oPC9Ky4zXXwZt9EMaEGDvivwLtMUqTThrDkju9HOWFvX9ce0fnwv3mtMz83
W7pDqcKIm8ZfyywBwfGBMhtvNwvRBeWgs4MRxswE4h6M/VL99O3oZeGVUUBo1f6GdSf339YkdXEu
cAvOZxPoP0giH1VKtIV/HEA7kinw6KJS9jxYvNKD91PD/reJ2bxFsYrz7Z47B2lcKIefAiAK+6X7
a4JFu+c7FEpTCRGU1tvYGj/9Azaksj2yk9OgU5YfVYmzmUixvDmH9I3Zkt/lbEF/tuWokUq728X1
kyuDO/Avd3jWzYT/BtdVa/z0rLqFnrAZg0Nmax1y01aJ/Wj3FAUO8Wp1+hw3YwdGovu8/wMZEJqw
qF/BegxN7sOWL5Uw0/3Nn958TL23gV+B3eRcnudWapGstMXJ3EfatTdzARwLaUuCvCaAO1jLfmem
pCsfAptgQ1F2P/J5ibGfiuYkP5fHd8e60KrG6kRTN6lPgdGYqHGjdJui6jJbpSoU+XLVVbSQUv2W
mI4CVjVVfSuNGtU3QkeR+W5YyvxNZOe5U7aLPOSNIeoUtFCgUR3qNodsBfX3hy0m0AkVuvH6CrKQ
DstdJKTQMlu2R5rFmzbJg+4BxEZXK761W45ueHDT34VV0tEhqAyVGe3wnJmmmVoIfsNjymjb4fRL
KzzgfMs0wFB0j12kl6OrWmmisffeir6ElybjVU0VUMeYAWY/zDfi/usEMWyGTfQOaEQxvx3Kdyg1
b47gQ+4DDrWWBLfDU8lrbsJ64ZBj/HCeQZqF689hr05unTHS9rkNN+1PRExIcL+eI3kASBIUjDkq
uAYJO9d+mOlHopO8nX9cj8nvoOUYUrbdmTXyOLRofQEefXVxIhjacx4VbHgkL3ehwsSrt0fWVg2O
iKarH9vfbwYkEkdy3d3AnwUpsvnre/8K40kIXJ1HaEIby6xkFOQZqBUtOhS+iiOu72qBCsX4s/Yh
4vPjfJyj1Nu35ryKLPfisoAlan2hzhCcPwennTxcY8iZ5UEm2oP00LDcomSBDfocu0N9ESZ5dZvZ
zUguEFT5TAhZSGwHNPlYagJVeSwz8u8cm1wFv3FWJX4NtPt0+AhbdNPUJyfL802Xro3emdXksEqR
on1/CbHXx9RnYmKFBn9ZQ2A6eHUutMSpuyobD+2E7H/i7+K9M+21fHozfw8by/skvJ/LU9BAaYrz
/UCHHB/7BF3N9eGFGxTPq3iDiyFmpikjavp6mnA5CDp5bn8hNP6xtBWcyMwBXhDUs61IxdKcfdFV
nid/sDe8TYXWZAyh2RHyBSd8HI+BZVhe31tJpnNxggqnHHxzEHeEOdhZ0lDhfQb8/F8A8K/2aLAU
+fcfi96Ch0Ra5YR/U+INYMFTmV7Dy4jA98/LOfVIrzuBGXjdY0G9BFkTt1GHpWlB6LHV2Zmb1RbW
3drmPYYpLXbAWlf/67FMiAw6xpEdO7VYpZrw+qGtWCteVRXs5hUf1UciDAtMFbe/yXdrQvMnKHks
uI28+FOyk09nUUzgGZvsujyPtKVaelLsK2zL4M6T+Hp8OrSg1i7OMSR+LkbElGeRKTlOfSiiW0K9
qfslmsamC/fgmrSROKX6Cmn3k0QixNGIjecugUcplj3CE6L3jJzayADGBBMsFITlQggvMv7BcxhC
BH/YL/nQx0myQBehHElQwX2yqE8HgSwWJK/cgoFKXZg5eoEDL30R0OErgOtBUDv2ZcZ00KxjJBLJ
t0uUiLwFPAIhSqTvRgYlAhlhfm2K54rfJ0ai3i9UpV+9FR3aDDStOs6slAknY1Yc3oiznXO1+vxn
IYWoBUvuJZAlkNlDyHb8JfmEvLcVvTw/38nQazIoVG0P/izh1xCh6TeZdVyoLNVhR+JB2sXT+6hq
pimjARgKYYOSBfk4uZaxuRYOWLqHGXi8PrxoIOs9Fwobpxk9hodzRLlCRUZUq63sD9dkWgQmzTCY
pcYIhiMcZ4UQKDUMydQZGbAxRyJYjPDWjD67DbY+5Mp83aDYdUGvOuoFzxcJl/jkGt7OPu1nj1K5
alhK4WvgsVta3ztDHPQrVnVgGDD8WxvgI6I79a3mcA3WilpZEYn36iAXEnxxmrpqropseoI8B5Kp
yMcotjz8rsAKxxaXMN2GrcggHcIi08c3VPkng6zSej137gVbOxwO6AAcsAr5YSIwswpbD3lppyi0
u5tYi0TsDsH0BfrVWM8907ugjuKGpVxMdt87LBROdt/Ta0td7fAbDz87Nm7orLE/yL8btp1jqny0
qhrZDC5oajj8aKSw6Y2hcFATg5t0RVraoa152rO9jkaZJ1RUal7XXiZSifa1T5TOnDJtv2wXVKOf
or83kzp8wQrlVGME38fTpRhmZt24PaW0QIzyAD0JGiKpsnKgHGUgGzGo8OqHIHN63V4gMbPL7ZEK
X1Tp607LxE4ysXvklOKC9dyd2pYW1fFFHTaLO6nqdK3f88Gg/gjLvavzIGpB8afcByEjMZpGNr50
AOjkEVRf1NQeLzzl5f3hbTnZEGIy5yge8NxZ088CYmCOLAdN/bIXpKP+b6n+wYFgkPLbLIebl/L5
iRoH31dt8160atsfUwgIj+GUKul+nNAZbBm5nlV9ZqzC2uhTGGQn8NwPJ/d3eYG9dPFfpxuJQcvO
ZfSM6Fx8UQXd0XdtSuIOKsvmt3mX4qcvU5NU0DRBeshDUArOI7JCBZ3d5veyyEPgpS1rTmPE97qz
cuF4MwtLyUmA1bNHgz0znvBmc1P+ejnTXSGY8QaE438lWr73eoCCarlw5uWBh7lZuKDLUyVF4HbM
w63y2ZFtgF8q0PukKo0xWrYF1RK9aJl2/5SYb0oxBs2n8fwwojdwWYjsxtTrRTaUV4GSbTpdrpNK
4Cu0eRpW6dGyhDAYex81jA0XLt/0pZjq/fBaVa/eu+uqA04wrFhGediCtMNm+t/0+33EEuNB0A7y
uj9ZTZV0dG69OaNoE6TFzfZkzkMA2wz4/g/2XGKIwQf+BBckjCaShD7GBhdahst7v+7TRC8QoE0G
Kbu5OL+3i/wUu9VRTwge0nV+xruByCMWitsDlfiz/vYu9iEFSV805A19xaViggmK1POPCpPEe0gZ
SmMG3Lk0CXSQlcoiIvt06QzSEVlUB0nig1KTjNiuBJskvplOJUkhW6shkhgZuKQSmRYNw7TC0ULo
Y4cIikTwJsalpdyp7Ez4555zL3dcMj95nhGF/nbZXaSoPWI4h7G0In3VcODFjPNNoSLFaEqTMjj9
oQEKRgSfUFsIVvKv6KBWxI3INvE/mzXXW1zKGs4Y+QUEcB+dCx7IA9DkAiponSG66OqL/zbZS4YG
+m20vk0p67P7yeVc3JHhPw/AoMyNZKvwRBEvf5Ig4zCtrJujM4IWtjnqpr32jyLJZfkPPLW4gbhn
wwxO+enh2QzkJBBwuQ35BaHR1wM2mYfGVbvTY9WZpLRCcZhBb5tjUQzQ6m5Wn6w1CKr3+SySyeD3
5Har6+fQUuCMO2u5Zm1iG9+B18DBJczDER0UivC2mbTMo0eDf1Er/Ft8Jv4BFsl8BwcfjplAhm3i
4a/HpBEZLpsOYz4HR2CYiOSMo+D/NiE20ue3Qz2l3uo0gTy5QpizVoPqDjS7BAXiYh2zLGw2lYzE
JXlXPGm9K/31s7BfbRTUNV5HnFOoZ5aZA0APy6Iee4ZfI1HOHiUbJ/Z49BU+YlZLvhQ8q53VVrVE
aMOVZRhyt0uWXr+NFCi8ODtlDzKbzilIcU/oDvU9ETbNUAevEAwIkcK4JvIHGpI+4HJse/nryWk9
OB533JIvo771Wa+dIBdKZK/sPtdypfFUdzJVAGYsZ+xh06+grG52wjoGpBWDj0b31pmnW4r0/Qyk
2io8Yx9dr99XsOAitCIPfoR1QpGvKnJF4RwCzA0GfP9ibCOlAUHa/f/iN10p3SbeLB4ZsAtbs0a8
MUnZ2QvZl5haXzTPzcFwhJizxI+O+lOPD/m8hzwyTXf4dI/Xuns0vuroJZDZB5P+rCgpcvTXBKRH
AyFY0m6zgDwA/GRt0/RqqrPT00oUZJ1IRCWNDRnWd3+6Y2EqhojbyjaBXN2Rvf353LtwSPMP6D60
BJQX7UrVFxZf+Unpt9x98LEj/9KGbl42nsHQOYsss3BUQ9T0JQmnbG9qopQ2fDWBH90V0fWfc/Zu
Zw0eYAZg5yC6dHaywOPggp31M3MPpSqjeEHMMJgUewSwj46HKen4s5BIynegpX/QnLUpABRZxleY
o2HOqpQassOy6e3Rttrckacj9pvefpN6VJqsBuJDzqfRjAHiVbwkeVNIZnyatwSzXh7IM8/8s7YL
GUHESfR7a/g6HtTVvsv7UlvOpUaY6yfKlRIq1Rjsp1zL3vDQRT93u3x8ofC2+YC190NJzETTp6/A
McT32Dfjb4c/+sMAgSnRtJDDRFCOjKsAp/k0Xlp53iqWxWvo/tWKecBIltL/DZiKxogbRUahIdzj
zAByxvIPfl+KuARK55QbxCfEqfwYna5Zg+oCbDrTUJlZ0tmknJ7B0lJ4cBGC+yAehRmEHUgwFh6s
wcoS5tJ8AQ+iOdI9meCNK98Kne/RbNHoeYJB7v+tya+CmQ/euiCJj2LP5nF+31zgZlA+LgRJYWZH
7sFsg+OStICxk+Wj9rFyDS60Us3tvXk7yWJFm6TXnassOEjDON4yfWEIC/yutSDvpvYnjjivGADX
KnwRwK6jaamI3cHqFxSaplzd5JvGehHIP2SHlESMXmKvZhs5+UIZ1W7CUxDRFCvFcYq3pmgnoun7
M1PJdwBTiSBGTVxn9LJA5wGG8tkJA5jogRzx2taH/xc++B0OzVcoFZ5cwzYjRrVgSy7v8rQkltXy
qD80Eh3ta9A5ZbC1kG85d7efN1ON4vEKWbKqWIjKVoaChgsJNJqR44RTZMXLZlBPC5Ug36qMgZG2
c0AhovvzdIa2J4QFiCubJJ85OaAPWRM49T/0ZA+zInd48pseO9E090SYMneUbUCgsiCMeixAYcry
Gc21IU3hjAb5d0mWdhg5jTpD4n3Ydo7ueqe4TLHYJPvNyYdrfDlNDuROfKNB1Z8ebwzTYJEWyi5s
H2PYlQrXDRtcb3kDhVgxj9dumKmxZElpUDvpHmSoCc87axgS4xDcoikdBb7A46LCeaqFZG/AXCgR
J/qoqKC8Y49KI0Th5ebxxfxRDDQG3lmgYn3k4/jPa0IUmR0mnVFf38eHtMRpOLPEUscXQYz2Vywv
N+PvcwuBgza9PJbtJKWEabWXrYZWaduSnp+egabh7JVNi9rX8a3SrSy9eB0l2C55T+4GfeC80dS3
TUyzwQeV0jowJRvR9koUIUaMtx3aS91eR7BsFykyFKX+cGxpm4JgRpT+N/UVvGf8F9IRb+I/K15v
ZR/O0NYahOD0UuVOUngkS0taLvoN/pRqhcp3vlEmEg4L+GyyVAOSYwDICcRX98godYhUs7hrJxqd
uRHNl7BMG28o4yo4XHPqcaXpot4b9OTJ+ogBdx7kWL8QoeuYfHOWKqhhNyUw5AJi5i/2spSVklVV
BS1isJjEivjhVsKmRqAR3KqIiQZ4zaVofx/cWxCD8nVpEOG5eP9ZlR2TPjXlqHZRXQL8YwxfvmNa
cftWNohmvpKDuopQ2ag3eZrMh6Myzxz/TW194yjH74G0HPcMaQVLsqNCj/nUGzt4MyAqJLD/+hS2
laG2bzMZm9Rjq0PaaTZit0VmV1/CuvFsvU0drWXw8KM51aPBY8PP1AYnxpE7ZIpLGG1uxbXkx67v
o3oz6Og6FPyPgXgdT6aB2nnWt1byPWRhQld751CINLrg85gavtoC2TXgymSlCTlXRg5ouZWzshQH
uAQbTXlbweHT4djOyyNwqpmM+hqhihSMuDTC+EqwCgN+GLVIW4dVTJ6vSgJkzM5yjtiQD3dPJ664
kgakcF6RBfYjN3Jaaz3k/TnYNi0FFRPLXlH6+68iKjhNMFqJZ18N+BWubu3hkqYTUgVccgrhEg7X
1kLkcj08PjulJ9ncKoq0QwQOjHruODiPQgDv2n/oIbpY0Rex474nCsKSYm9c/YA7CGKGj+o3kBiH
t6YGC4ydeSoJ1SBOnBSvxlH1hJamyWAMrF00RpE9J5NB2Qmmh5DBgkM8iHpLZ4JLEuMHtIPBxBrh
fPVseOy2whXMb08c0IiN0YLPogP4sY5CixYPHV33eRJ5ZUBDTKe/lcLCQT1grvNV+4N5RPdxI4N+
6hYte/aKpS5wzFvflZ1eyv9yOYfGHfj8G+Kl8jWWGtLYiMhcSJLchvyG+9T4Qrjeq12mOsV4PMSv
obGB4TucKNrw2AeHkMBZwQ0fsV28/i5xjq5T9lkNAZRmX21QcwqCex2U9Yf3615bObbXb4NLoOzw
f5rfudcEKnuGmuvC8zJtm6rZMaO5tKAZ7VBLcBysYHxewhC1xxpFa7afwZXDQnNxrMbhN7e9V8wj
LLYa/xo2z8UDXxqloCy9QnLvjDQd6qMNBRPK6rRWTHX0fHegJ5288AijUDHtMvKmPGIFTnYNQZb1
d2+QSn/kEeC7sT1i5Wavt9gxzclNZDoFSvQ+RvvjXOf+CKyUTdiKX74CToeD/8IWML5iUAR+WtZE
R3lCoUOos33mP3ZW4aXVwnXoF2++w3+mAFYbNj9kips7rRNTcAFxavlfqY8xNc4hFU+E98Ox8Qwu
cgDBHlbKySGUNU1j/W5OyCYAlaDOXY70ur0PdmPry8suKXH20qZ0WXt2AuOTtq/FATn2MfkXll7g
iUShhPd9EjnKCWWUUFp/Jsx74QZijy4ulAj0AdH/BfNOgFts+D+EVZ+iNHNckPokY8cCfvWD6r4s
W+Yk8f47kJQ2UB9HM7jbYn9mIuJSrfACsJaqLsBp02pFhkiwFQcURGTlz/PRobJRE+qrAsLJXDdB
OFscTlWe5IBMnRPEwkPtjGgxmkmUOrG9adORCk1tcTowwpihzXCoc4wYCzpuut9S2qLv3Mn9s7AR
zKmlrVzzxwFdp6M7j3fpPL3OjPUjhsB4t062nNtmE6viLd+idAKAhl3fFUM+9ufNy1YvmkVZSHAK
Px4NcpCgOm1rTHs12VFqVuukpdPcCrxXoXjurANiTmhHY8/yBHovMa1AoNm/ezE+I1KPYYMfqFDl
DH+8lk1XMtTLv1KkFpUY0y8LVY/Wf2JJR2ll2Ox8T0aJ25qOjtY3ceBua0dFhyDJE9k9eCzYe0d+
Zw1tE0BWO4sT9XZHM6guz14nYrSMwhIjB51n7hjVUAQZG1BUROXkQlaiLo7R4VWe9LxvY5ViRZgk
4ubzgzp0sEHhG6rTMXG/q4nGpFrjqF7Ac9hsjYzo6XS10KGf4DL6iB3eWd7VgrBZWuMP8JXI/iox
a2PsfpN1m7aQRrO7GBDItw+aiaGm4Brynr61Fcnzr6nLbI/kZ1iFrPUQZEvBdbDTAn50DtKtF/4j
GKJvaNtQu+seuXVGVXjfsqw01rYhzSTad9DxMugdyMr8GS2qsuoP9XkgrR2taKAijmgnQxLtjbza
PDIG1p22aZ9z4hJagK55NRM++ecunq/EuN763BfCsUaKU4rPl+y5oldtHEjtFxMsGmZC7NxdeAZF
mcZO9VxohOkYooFFUoS7G7KNut5yyeCnSCG7zLJGANgaIPVUTEnyrLTJ2U/cW2KNPEK6I9FIRVuK
rB/KNOzCodFbNAdwiijdjwwVSvUJT2prKmvYrhHpMg+A9pIDm+mWeYrGZGmc9hocuhYzJjqikEnH
itnb1nS5X8S0NeNmRUjrUn+qWDUkp3udWcppujjMBtLF5YV+2JARchFTzyxQyJQ04eyEh76mnilb
HMLv7p/FAwE/csSEBaI/gPiNR7z9onTCGneFUjbZxKXNk8UnQPzGCa+mokxo+Ju7dTq1jOT/NSXf
6DGuXXswEL+wOvGEmXEtth3/Q36jGJt98+T57Oi2N+nc3GmlS51pYTnXPGVjLjJwB6nZIyOAo5Xr
Klv8Sd3j/JVZjOIOYCZYpSu+U9qyc631XTwR/X9lDSuotNfP4c2zjwqPLpgDLP7yejsZUyCOYhBm
wHZ2Q8ASgsgGK+6IQZJYLTPBZ/M82v/nHsktxHEOB5TBm/68LGFnBm8nSMDwSZfUrWXCPz9AyvZ8
TNjJpl96nLMaVVazQmlAr0Zu+Y9rMaq4XMAbVG+2jYuZpm5A3M4JIf2ZQVAYtEkJqGyur6B20AN+
ULM2Hj8j+gTE02FxSYNMDFDBb9JStAVMR0n/RTeJsQLGtQxaoRY2s1rbZTopds4UAK3sDD1tjCoK
xbAI/qwucSRxm3H87n3K+miTkdIzRPQOiz7yHsAfvQo9KvfjPdbl/DtsagLhgLzkICj6eTObQpCa
xAFjyCDQQhqMAV9T4jllXbAqCHbU1LuQyZ8JFtN+pI4lSuIDAVQq372rWGEnC+vcleDvoX+SpwJw
PTRznwScQUGEeTBILVAmlGprMs2+z4d7dXNIGv/PtOUFOPNFxyUQAmiMTjmZ863crRS/Dx3NLDca
4jh+2nfJtoRJZCyW4HlsLkd1JitBANF8taVm5yNHoWEJLyHP2qGcq6uGiFlepExjSdhq9W4il1J9
+BhtOiG0dQ6THJLT7MkQhG/5LI3AZfrEGBCtTYT/wcrCwT8WJ8PhtdIPy/pPJqV1te6v3Q30rYIy
Bh+CX0aAQSwJmb1BwIeKvnUFKxlNmScZBt3SuE4PEccqG5HHc54jvseyU+pwBqucKLzXcNojUwQz
uRZjeNZIQ/YI37pNuhkhpDJxqQEMMyg+R7iDfej8Sya2HIgoaUZgEigJhs7kb4w2eR9lHmMhfdoz
4x8pwN6RSMk5NpRfO0I6TfUJoRiv9EBba2nRwiWHO42HWMEr76pEUuMJOLVdD5vNyifklM9SLZDz
puNqd0Dtpa24bKeOmcuE1OdUJdbcJUTH3tm1yDP3b1rIN5p1ZK8Q/Yo91QfAUozRUkYF+rIj0sZs
4R2JnhAqSJ6iPYGQEcjuDfvM9nwmfUfwl7lEC9J1nupH+G/eaORMrOuWuPCwTyhH8j1WRF8Kur56
cVn1GE74NDTEz0amwt81VCRNH+IWBTJVAal8sc+D5RHExrxZVyFUnL5BpW6bhuCje6QfejdVPLw4
FQW3tba6gujW7KKq36iHraqK2iUytAHhTpqRy7b3yCF5kzSvLdKnwxEkFCle5isZBaSA8SttYL7Q
TvI2Sw1sQccAstnwQJEydRczIWSOtWXBcGSoGV07PyeOF9KshUG3twNVh813IBYpTlnbdN9xL1po
XXSmNo/BEORE2/NmPXeUpehY7ZgcWPzROjlVPZwkUIA7KDcUzI4as2Cc1P6eluMBCGPyJ2FMpwXq
3ZJ6Y3RcL0BcpYaLs1SC8XhhgwFtnruOgTNSn/EC2PL53pS5MqRo3zA/VQlusO0CGREscL7cRYxw
XjwW8OwHiWXqz1/ZnhnzaLJaPmhR0ZZ8R6oo3gpr023rUNDoADblzEgGUl4TZcfjZhMAatBtMSHn
9g1D5BzS+IWUQG+VIjPZthVkq2wRfKHB4UQ+wiAJMUZFKK559dBD4Km6VjYhA7Rn+73ek8zRIhWm
/3/tfigAQ2sCMkMF/bD856tC669i3Xsuw38giN+9V0+i3Drt1DGaG4cwaG/PZtpEpQ/K2JgHYY7u
PwvE0Ugp0BlyydS2z7kv9tZxE1ys42RuUJVtCYHeQYC2KGK4dGgLvmsmJb5GNgkgJLXD4NYmfEc2
BsUwJKdCq5LqVM4FnjXsNO8GZjHorMn7iGW/QaMHFLiIWD1GkoWrJz4eF0vw7w+vtNLxnzIEoPrH
uD0HTl0KUqD2UQFuPRlQpQSG06WHHaKR58ehtqvS6VYJ7L/CylFJ4018zuPjDWs+yd9zh/Bm3TAG
H0Txl5ZUmPz/KPPw/k5lzgtJehzmTNJkkXLhwFBDkCE1LFihqeUtoJLPhLgweLDg0plnJ7m9WZys
Nsw/eI9D45G7euJdhMV67ZkEXSFGVnYJq43K01u6taORtcgUe0AF0smGduHblHCWVGmjBAeGF/6/
ZCCrSS2t9ta9JRbuWBJ8agNGIkdAkSKdQ96pC+2QSN9oo6iKC8uUKOagr0te75ppGDjJCSB/GDc/
4Tw/QtLjSJlfT3loo+fqiULsDxnkcBrrGpR3xmtMDAou2/Mp+0dOAjVvsU1RjHWXAR3xcCuNyOQO
g3F4I1xtWGQ5QQc0y/RpUMKmAa+YrCloFyUp5QeEkKHnSwvlL0h6zRm4RVzaFusIOlc9LFtLpp1O
F3oZgSmjUsJupQw7DZ52jvkZVjhr+VKufKcskXnIOhkuUd94UvARuP3QCcPOgM/MgEsWAal/88DG
s2OhxiV4r3POaLNQwKQouYfjfKGXYFcYhiGM7m9lN2vzaMy+tbL1w1ymknkdJSecEdRda3D1pP0n
FXJGXh+JLMBzkI0cNXFcD0+9D0mI7Jk5F9VdRHMj4ojEY9hE0QfoOwrBQs2pK+7zRyJ7e7MlpImO
a6AR2PSlArLEuQyCU8JhYTb30RVMeuOzl7ma9PBuY9Y/iWghsSaF4iE/klEIQrRx3ou/M8pplblo
yfsNKgGlgcjnDENdtoiIBkSiqdf7g4LB+6ENt08TkOfs1oqKZv0atsBbf2yV32JBXA9JkFaXe4wm
DIWwUA0Cf9N66LRMJH7j0S20UTGLL1mlo2TeDPKM5U75arbgMWoZPfbhrXxvu2MTnsdYRpXEpbEq
B5S/MJWz6raNh4DGp/z7NSI2LrWyO1769d2v8Sl0UMUXiBgfcBMcV6Tm5wUEc8lBWfdcIxQ7BSVf
gHYECCeQ7q9Te4JErQRjOTx5udyXYwYQRyj1LfC0qvfIAM2X7oINieZIciiYRPAc06x2/FpFYu7q
6hZMD1bPfokneeh2F1PLnNm41v/SNNbY/G34+cf7KbhscwD5RTzTXdm4e3f9sIK0ZAK4nSLWGtWo
vkULLlJetXyjR57Ocsho4FB7MzpKERrGDlFZMQsJsnHtnBlttar6PRaY1UJ3mrAVGIM2qAyQEmV+
UlM91FKT4Me0gY52dxlS1GJRiHi6Ib0Dyf5IzuYsqsJTyPdxAeORhqKN9rPQKUfYZNmXpg2CoWKu
zXCul5L9T4zXkC5256tCJz8NzgArRI99LaSNRxwiJnc7e/UDCTXjp1YYmUokDQbLuXLDQPmSLLzy
LOo90UO6HNejZkipTob/9yv96S5hBFJ1hdVS1N9J68az6Af6QrMWHENINQagZRHRQiWZDmIaQBdt
pEwQ5ZSq+FjXa54i/tDefY+PlwLerHfGhv3FcDS8VatXONgya/YaZiUszR4lFU3yTAVWNAowY5Kp
PG4tryfYNQXmAwoumct07u0Ii8hxphSut51krLj5s6l4uaQp9oDBKed7kF7ix2Snvky0dtRnHaoE
cr/8qgMfBEL1L1tjiTZz76OuQAnevfiG53T4vV8S0TBN02vopkZW+UbYHNiUiTneO1Rzecb/x3/+
jnE//EzT70JWNsBvuH8vOKHDrGt5BANCLm/AI3RwOHbzQl9NJ7V3el4IJIQewDAeMshupXZ4CZsU
kK718RYuEtKICwFGIVN4nB9UCcN2zy27v+wPkfhJVuTaUFOzU0ZLq1pC3CQmFmkRLE0NaKSPNmp9
OBbmNYPV6WhtUY/mtxbOrZfqvHFnWL8w8jS6Rz0dOjDzwE0q9TtKnEjbkcfxuVfrvbbfGAd59JDE
GbK4tAI6WCOI08q9tIWdibdn+Jdb4TT4QOnM+Xnwq6+CDGFYZbnnI7xlJi1t7O1njCjP1uWpgh5i
T26YTS3vEuYn3MRvrrSX/v/3r6KJCv9mJa6Y04kQgqIZ+Fh7ong0am7YeGKvTnNRjLzYQRTotWX3
U0CIGtPy8oHpOKomxPLErSuhpnWfYMIMOh/bNwEQg9RyulgR0hY5YGze4TamGtqUr18T0z/p6Kuu
1UlcvYePvEj97e2n1GRwWhYV+RLTfbwgbhTGBDLzAkUYaU4qp6opq7LJvtSj5hW89P0OcYHLxZYa
RAcvzrr98ch0wn6FCvYBINkuvA3OOfgx2bFwmqzbrIFg7VmlVhZnCwhhbLD7O2EtrNPFa5dWjS5D
Ls4fcFX6vKTbF0lhorITzXu2ps82aklDLje2jfHBgZc32Pl53DlxSnw/ZAfQYWaCK09+sq/nKcR7
gHIPH25g9ZgvS413KO2kewTimfQXNilJxfdyT1y+BKBY/iKG69AiStg/4rq2aMn9Zx8X7xmpVZYv
vJQ76XARvKkhd/0S9ou5G2xgP3clxQaYoDXXdjx79bFUDiBGU3IbKTcpHZfe7hNRd45frmPO/JeI
boTrqVgjlWMKxkYuj1qXKNsX6CaxfoXElkyvdNBP3Ay75nx8kI7VTJZHs7AmFS+bEC/COLBW8N+0
tNZwoePAD2UdlNzerz/6nKMW6I6FbsFtlT4+opNHucgaNhjFmOUm+88gL8apRhmI4jKA+stp4utE
ZFDSHbLU2w7UdQ3STQa6s+NsiSM1NHfFe2EwE21SZMt9XTqtpnkf+qI9Kt2xj8bMq+UYes9b0OdW
TVDsCGzkjv2mhDbvMYOAEJ6+O4FH5mUxqWsJUwiWkMl2VXxUWB3Rg79+KXoEk+mqcRHpEJj0Gxb5
7k6t9HSxrdH86QS0afQ0S4nUGWG3TO+/m4qQWXZt9ODvPcwOzLtH0bMsgkNukcck8ZqoaQoRD/6k
rgcgab6iXRbsuV4WIXoTCRnfQf9N3gKK8U7HCHRtUuIetYxNVuGFSVCvvoGmVB/8xx7pZ1ZcBjbe
u9odWje9vXvhsjTEqoash5hRha+vaiHUl/Vvm/0qTqbooQrzFntfhiGrwOnhmYBwmBrCf71T61PK
HL1U8dTksz9VtBEGjWFKx98iFOOSwhwvlTjkWVxlzu83k4dY9HefTmC8XsaxSPTbP/7rEQYljjhg
vleJPmSmZofbVlKQZ0EISEO1z/8PLLMXNdNxbET5tavxrqTjAF5lSwWdWwIGJDaU7XIq1n9xWKn5
eKDWLSlevSUi/KJzhSswur5bJJgVQzzj7bQkAJOWkwE3fBD0tODmoJ+pC8mHv3ydwB5T98VBqiiS
4kKqVco+z5BRjLS5k473CwLcgisI5jnL+fnOCGegSGU3ZdEiurQUe13O6jrtmp0b6aiBAUcmaeZb
UFqiGddtuwjk9UKBntzx5gn81D+5VYvZBpYK/VgTbvr/4ILH2IjruKJMbpGLgH/rlofYjrS5XCwu
A9Qtw9+r5vb6TNUitNjvdMRsP3Ic2K+Q4ZdY7jsRogqCys7pG89p+0Fn3EsB9woUBRsz77SQ0Jd8
M4xv8uODULIUVMEvz6/2ThKTjqDnYXaLZOYvezA238gvosm9ocX1XVrjC5CGAM5kFEX+uG5Fx1Zw
AAmHAQuEiz1TyVm7d2A00RpbNGT/lGkfjr1kuBRmW4etKV8+H0IIAPDAaqDVSqgvO9IKRRfLuQR2
75aJycgA4kDmwQWO3sCahLaVfPhyMipV2VASmivEZAKlFGQj+om5+7ljT5albUtSckJ2GmLWyVYF
z2VzTMbaVpP4tG2JgiN28TSWzIxBhnVZkXrA0YSiYeUPIOksDn5Z4vitPa83JR+vByKyEAbV3nj+
mtOXRIoXJRvqaF+BfvCcLNjDHdXIC0F8BespcXHey57KPSLCMRenCWv5Z52tQXc3bLzEOgV9vUzP
UnYfEu3PwI9yA7Vrp/AHf0XCHGbdrK+ZnCpjuSRe22xml4XJHsd/rXqJVpLLPTCuNf2o9+mltCZb
ZXX5ia3NqQl7Ok/XrrsqZvvQin4tQHvj8i1qQX6y++yPwXhOWWGYCc7UJcKzrJu3qEAjAj+192JG
+R4139Sm+bsQKdyQdSq/gOeGuuMJRJeM6WKuetcQQ0jEuje0i4Qyo7NQRLiNMvdj+ZOQ61O8ce0T
42wgj9N+tlqsO5MW69Ss/j5bh+ywn8wjqmYgu3rv3vwSTRJEDyKfksyZRFHJhEeSCPgrlIq7i2zy
ZZP5RvVIobORdVfeSgftzZHVYmbGBL/MTaXHm24eGdGATi85XD43idU1qhiL9ph+Zd8PtwPfqmWw
xpHhJIp0WXCcJe/bvhdhjWehPdIT50oGP8FjFP7vB8wLo85KtyJoMy3s8fmolOK16XrtymQjF9eF
eD85DqtijWpwrJ1XYoGLEIdX6qu6yqOeHfDsSkKsk6KRlQ2APRxpQKCgZ/rxrxWbLOOBZBiaVKt3
dVAU4VMZha1lmluHQT6MDRjBfOw62zFWLdJ2f56yf5lhn1oW+vuh92wdDMsUp6xzvKr+KGK50LRV
gQeR4nQ+/X1VbQu7jC5ThLpmJzm2ZOaWRfFG+TIClUB99wOqjuj5cguG/ixuy5tpGCpXhAnlozJH
bU6Y9KYseHTi6aeu46xTlUXvMggIsZ9fwTHSWXENL8rp1LJu6AxznUSsd7+UdR4B/rCLvOPsq9PA
4P1RzYDRnvLRazCiRimtQw08iuObGGw+wha6V0RTl3x4YdQFu2p5aOO6YdmFHT2yeczVT+9EsKgk
B3+JMFYZ4s5XpE+UFmkfUe+HyCSCBnlR+i+1wOWzg5VauM1R4bGbCoiDlmUsHfxLRy6jWIXpyWAE
cotwn20jzo7SwOqPJ63kd81dhXpTWlRXZGuDVfqkbcvlcGtQLL0WfXgATFqV+2rI7xG0Yl+gcZ0d
15TNHn7tkO+pEaDhorI28C4hDpwNHPJeiUyk4tAvq72lrh1n/BR/FJ/i7NUB5yVnKG865YU1SgTq
DaLYX+SOdqYDLbri1x6w/BpFTOaFGb36POqDjXlNbQ9HnLq/OB6j2blj3/S6rUNy19u2q4dPVH9l
qahk56XwOalocxEzjI51lkCLgJ8daZf/ebYY5KmwBcebm3LtCLiF0lnZOV2qxJweTf3UQ+yQB+x8
Y2ekDKYcjLljBxFWe6O9VcdfdLPweiZELsS/J1Wt5846E1Zrrb/umyvufzXZ6D9/F2XA0BsL8/4L
civ5sjbk6WPDTlmfXl9Q7RW3ydzXRQVa4hkpBRhDrndzl11udZq15foHWTCPkx6Z851pBwOlQTLi
TnQMhWHDgY9Qskoa1dhubypWEUgnHqPLN432gbYwzWeuIqtlbDO8u9hER3WX015mqeeDfrjUiE8A
dc1oDueBXkapQAxTCB7czXYeVzZ5LxLLnX6qREd36LAZsxUlpRSQ3gkhNCI+XlHmhRRz5T4wgMkv
FTirudw4PaytJQo2d0odCCEAOmxk9O0LC+/OKQ8MP7hUTNFx4Y0xQHZe63Pdht65/d8gGbVCUkTI
OwKuBKnEJ8cYGFGuXAFnFdNWGEEM9pfMdoHK2mUX4rKnI1J0LIOXFXLLrE+9b3IAG3biDIoKV7hW
aNtSWV21gVeGFM/RVoCmmihLBNu3jTBmtsnW9RCc9rXpMS37lobHg3kLCl6GBB8wgdn2qDdatDtX
rbIsXnflI0BdNQuaNv+YR1UouE7x2J/u3FFnvC8dm31l2b5LsLe1zusbR3nIKr0rUokEN0mzwgcA
43YtJTR5huc6ROahEmtVwwmEsSm1T1zJM+oQSEDm3uJ9xKbVmJRI3+/PmdyAT6f0M4OIemkzkD9N
hXFBoOMZzjlR9AsR3e5Da14nQ6cR5cmh3lp/ESrL0ym7sqkyEEDuPVTMe208a1WRvEJjXaR8zH0z
CQzfs25l7rI+nCibNXoSkA34jQAQw+OS8ksEBOfBngSd1S+EA+9kUS6mQUFovKKyOZs+Hr3eWtoN
9BVJ8W2DL4kCqa91IeHBvJp7RST/D3l3B4lXY+fiLKveCBip1X1RHk0vRQBwqFHhNgqgni2pw0SJ
qSUBrkE1YYCTnYL2s3H2ksQKx8MJsJp6cRG5Ax1a2axHjh2Y2JITYar6akyCRw8RLn5SEpuTha3S
L89V6qiMKK09guwhl6Z9giHK+IvalLWrhdG8L/XgeO2DTXKOHFhnnmFf4Z3PhrQ2ykMbR4qfEI5x
w7yRtoceFLQZYZ8cYUUrc4L/g8FLX4TTDKZWZT8dffvSzaOA7QK3NO9gh9kHVmj6wO1Q88Mu4WgO
7F3oBLx4Rkuc8F38wOuHtZsX2oR3AF6Y4tbtAS43ft3gH3C6si6FKdfb84WvVVT2uwD2v9J3A4RH
Jv0ugnwLAGhCG+Z9TJbqRCIxwWY3FAYxZWPy7lhWCHJk4XOjXorOVAvmJT52xkcCRlO5gLvRcIpl
5Eh7BpOy6gW5jYHUISe5mOcTh6Q8WHSb7NP7OtzpZK/n2nODT4H8ztUBr6I4WFG+3CgDk0d0vPqp
/UQCd0oPXTeo4cD9Bl9CpPKfjkNLCX2Z8Tzn8aZJpy0Z959syvxPO6zU7EgAPPMijX0D/8AlmWDT
GfqwUi6WhDtGOncgyVLZL/kIpzvEIr7KRfKrpKkO6QoWeUpXKQR0YKA98+bAx7geqARe9/aS1O9d
M2pVe/bMTagsyvwqqeve5gx183xYVn8hPjlOkZIilTwfCIUDJaDYupiI28yxqo1yqPSMv7E91LHB
cktt88BL+AGbzkqwEn53mUhKe77qV9SytjkN8y05YUkG7rljvmDgM4stJNCT/8h3TW5WU9KgfZlp
RtXYyfoe61fM+mRIiAPin6vee14CV8H6AkKNfKCmf1qJBTAWWG7w5YArlABI5NCxVKS42GL3aNLw
IPyN51RNAyWzx9e6adI7KcoYPBCf4TwihLm2+aetDEEU1meSTXWxC9eepYPw7Dmw4uROLLZW+xt3
24t7j7mAtuhf8V+hvfjuuQS5d8rL52poJoNgNe37nYRylCb8ZK04iUX85Jwwvq58jrhs7K0DH2TI
HJXqUPHRJJbhv/6XyYpXg7LikTbhjZyCPXQPUoAjnm7JW+p2uMBL8Rw8GmcWxJWhf0aNG42bSxKr
lncnTnfCdgdnkq8dVpNm4txJvcbc9fbRhuVxHki+4aew0J0BQE9Pl+iRAyZJ5ZOIRD8TvIPphJUf
YT+CNeFgO4SGCe1BKCqhDsDo2rYB2yZmpr+2jzrcpb3XWB2Hjyy/JgQ+eOhVeA1qwaWxszdjzlIS
nVUT6Z2tUnHQQlAKSw875VB38Gvb/dLuXMg6YUIdc9yVnvmGfyVa2tgIESG3ci33uIJchl1qWvkb
3aRMY+IwfU5PZVe/nWtw1q73I86b13fsbahoyhuj5CWvf0SuUXD3yieb6USNKDECC7iC6Mcq0KWC
8rElZDfTSLBvezSw23N4P1FoKdoV4fK52wDN7s0MevUfa6eI4s/hs9DBu4vFvSMXT29dfhZ2gQ/c
3HU9pHWG6Swx1RbT2wk2c0cvkwmsKg4fzOvWbSgRrqMvpBCwZca8TzZZPl11Ama2Yw/pJW0BAUqh
iR72xTyGQDJOTL2UdE0b4fIZyCNWKT8wxPEd7Zh9iK6jzNBmZ5By6/zqHhbMT8cpkd8OEfmoO8lt
K5UXKarALBhiJkmOM+eC7bwSCNL9ISJg6JLzhldsSVZgRt7xbdfJ4Y8m5h/dbETwcyNI3O5Ao9S+
JosUVh7UGZTpI5RVmsYsh0LsEIa2q8NP09mosN6i6+mzCMJP0Yjt6tm6aZUpgdb89JQDVfPPbZUu
akc+0ltPW8wyPnW0bT2osg63guk3DLd7ihqcWgIgzP62HfwXRz+Qs0Iqex71cvj2i/GgzBkGnp7D
TbLdvVekXYa4kxQFxk8d8lBQzxF01FdaAGhb9/HF0x1yHVaQ95rdFZfit2LJCZ0E/+RpFKb+lgg8
OTnTCLZAAE7gUfPjegyoQhFHz4/V/cka8Hl+8n1w8Xt4dEULRRxQu0ofqi5DZopBiWkmKvZTzur9
YY6ZyocLouMjccXGvCDJu1wZYZgTxSMGzQ4Od7uIegaYAtXltENKPl9vbM35Fey0qowG9pSxKNcS
HyCDbngNI88/lm4OCZpx0NJibtQlmIVYVCWinInLC8YCMBHV587gCgnzf5q8jblcIl7zqZUorUeL
iEefqQ0z7K4+NWZcGGkWlZWlFx1wfgrkVUxmwIs8ppLJ+p/W26IyU03FKXZq726bqVPH3jLlMpbL
w0UolBJGQ1AjF5DKUYuXurAM7uQ8IGbhKj8KaJ9ndKGFsXLQreDMJK5Jyw9LJaIJBcM1UDNoC2GV
w7oJrQXPD1wCCIg8k0qHyU9HTJPrlyd9I8JOIN2NoVwpFvid26JCnrGUu+OyERE3S5lNXAALCzcG
D8UtvrGYWQk+HbqFtIPfatMGRpa0YFRT5KikttkJjD/AHMSm8AKRQMUcKRCQpC4i4oqk/1Z1P9KK
z67WYARQttlF34xlrytFu2AYArhpFYmwEk7yIQ/pVuckgJ2nqc6NXfsaNEvqkfJCKr62SiTff3ku
lx14iaD14awtHk9dy/D3mXOg+Rhv+KApzodyUjFuIOdGQ8W4kVOslzTCgiNIJ413LTnt2+esmxR9
m91IDempHH57dkLoPh2pNNGvJmpl/QZY9XlPCqh+zZvfUSAGz7Zesor+5W9/CRCJjvKoxfWJMD2B
bWRPyGeov9LjYn8U1TLfKy6P+E/cn5h+4+cSlITJAbJ38D84xp+JGJF4+yoIsiZdNpAmOx3cskd/
V7kO3sAs3jFmVHUebaq3BdlV6/4SF2U/AzNMjuLG3VhVVoH6IcILtBEmkh+kFNYSdgiHm5WMzl6B
aukENzh7uWBlvDfx5OXJbq/S1CR6KjX4VuD1MxakdMsCENNPoJdcQ3jpqHseaAaxEo173hIlIuwZ
QfaQ6eFwLLX8fo1FF0DtWVlWZ2lON+8eNq/svEs7ixPgtTdMZnRbZ4SqNDkSIn4eCPPZpqbHG/KX
lyZA3ZSMOIx2LSYQpbEzYdLfr0jKg0uqD5J4FZmWy6eItVoWQ8HbkiJz/sCZ9Jz2SFI1emP1jqCt
uQl8yHbCDn+FAT2Rnl4EoN18rxWFkhwd7gAN9f1aC3anSijT1W/h4TR84AT0OkpEadebZOnMiLzE
1RKeQInjXS60PczufUKOV0RkThE4hd2wzJ8W+9iM8e0BKpTCRtNodthlO+tkFqUoFiLrUmviwirL
saXEVHzlQ3/d9bKLDwp3Xia+LQ8gFEk9m2fi653q5pP4HWBhyzXBemJMlSwDsfXccskQFo4JHCSV
SzoBisRWN2Y5cfGRRNmtnjL0Nmm8S4W59xxuWCEERh+sTgedKxiKdUIhHsB7SWfKsHTEJLC1q7WJ
H6PjJ6QT3hLJ2nv89SwWB8aAovx6RgMPGYNm3vmYgl9WCO6uV7FMMyuZ3nA2O/Ldq57QdSfFfEd+
ePxTltBbWUHBUA0HEr0Ei/E8gEg5PlOVyXAn87AuC/bXXU5GRL1vH0XWPjZPrlIDR2oLIhB1nWQQ
EQwOi/uTiGZbGxtnED8CPML6IzBOXEX6XFTlEbY1cbZkXHxUvRraBUVsMVJixIGTDhDGf7xmKjSZ
mWhCFLdwURLL5LpAthkDpDNVjkzXc+d+TAScQYidNv85csfL3IDXldx5K0Ubcm83S/7zHxUfJtWu
HsMcEu5F+Raq0G07deJOxdmYH/d7jIi5ifDcVlzN0ech4MCXTmykyp5arqckSuUK7YNFeoheQxzh
CfcQSaXaP2p4k5+fHKuAH7U+glUFSjTiaGSfY35hJsfWKWnOIDfspZ5qLPs+Bd7cPuVuPszUUZXk
sQdE7bg2Tl1DarwLEmi03vMsDRE4Ce1j5ME8fIZp6js21yn4Uu5MKkq1EYAynNrZ4W9Mgbj5ud0G
3WQbEXLiYJ+ubhBI1BUH8GVID38lcTgjUKrapSx2zpdzXXJy1rJ6M3/rY1ATLdS0w3pZiK6Heqvc
1AmtH/Wwq+Rauvk6cO2g34kneqJBFfaBwq/4aFGbCzu1PwxObGeqhjYLFw/xWYQOZ4jgbvEZksdR
E54yN73Y16CmcWnFj/IW5jOOH1NSWMp7fzN+i8Bpx3mOgBEttlVK3rqVpZN0tywOHqSyWU+tdBNU
4omVBBIn6XmWr9TyPOvgtWAWRck3KH40W3aVAYNsGZgZ3+LB+seKwZiCdWYSJgl+scNdd9oBDe0Y
ZulFM5vf1fx5UxqaiEMWXSlZYk6bDUfo4XsJ/4wrVVwYmW5U9mzZ1MQNlegvK+ZeCx1N5EJdpTCZ
f6QxWjSucT5Nw4w6vQmgoPIDGOINL1THBmjzGrjdQjSZLSalIr/vPuERbHhs+fPzdZcarO+sXOQB
MKRc4VETOFlEUqnw8eQBn//jF6BQg8fnUSErgvEoBJTyN+e74/DQf9LYi1MMAPR1lYylsyaongHv
ewCmSyxRdsqbk21SJ/D4naSvEsFyKawrqr7gKCH7bjvj2blcIfZevrbfjgNstTZuM3PTUUSkwdqA
rj6o7XvQ1kzIBnaMQS+fKPkha7IF86ldd5OTjnjOrSV3sEWQZRI93gjES5Fl2WTIED/WvLhJrAIZ
mtFg5qwHDRwLq9kib1DjDL8eQx4f/MfFM4olVF6RZGXjEkqnLtkz0WfwxfbSqHp0PuT2meLBJckL
Sm2AMemjuDsldmSfZb+V4BYM+WmGvXQwYPCpYGe5dMcQ0mGZhULqk3DowEgHXiDWVXiHYDLhvoMy
+g6daXfT2TiMVAzT2KYzb/7+gPdYln3RMSPld2pBOWBaWrvE/TIAEJvaJ6OLYti+Lm7Z7WX/iQNr
3IAB4iuQfu1sNmiVR76oDz+EdrtbEU9lMb96G4IeZJ2jMFtlRdt3KIgI/0PZClSZj8X+4YhzHRAR
bO+XE3tpsoEXk42/bFXtNs/0WJ1C2o+S95v2wapfefiHCsKah3MLQMi9kuxCaVtt+eFXC+NwQy5Y
hLUFvOFW8xnSdwkSjzulZt7CmrFCw+SfQh7xawPLg6MImAFX59bZNY/d9t++OfoehAeUj50lKlUf
jCYRJ6B3TURZD3166nzuxYMvcYGLJPL26KeGMkqb075+/0z2Cz5BlDPjQxwpGccoJYiYDqJCVYzp
tlgq8Hi1dsqW/rJEq3m41dPdsl6pbP8NxCoKjfC0DGoU+lHv3GPXWHl41Qe9kTDcDtIF0ALpHQu4
k5RAfMsySU1ptLaBa4GD/TculljaJnQe+mHEK0J+H2mrA8l1sWrd0Xjvrr/bJetJYfZ2Slv3TUdF
60FrkZg1SDDRL+B/Gq8QCIgIxgn2dKyeIPdUyhckPB7LiV4GNVMeeSm8QQmLeG+2dpcz5rF2w4Os
GnXXMNcqVGIO/guif+XkzhIHRXB3X4TSmDgxilRpwZ4EzIw5C1mJ3ayL14Zp3YmCfvMvuruzkORC
/HyjD8dGd74hGED/FvzxPmwAFCu/xTdlPWhqWSvGWYvM9VWDLQi8f3ezTgCuChtJ00xvf0iRX/5M
HkCCiz4hiW0RZ/5OPQDtBco8tjMDiW48FM1eaDrer5+iPR/fQcprk9PQEJaOKnjE9xpUnyOl/9Jh
RVZmLKfYX9e8w3ejJQtsvFheuN2kzDiun+EKonSVnYis4FgkzTa4Ubn0Y3StI+tJ1n7xNOfW074M
Q19T5g8RE/zyFRaXe5BZEBHRNHy5xUgk5nSL4gBLnd0TJP4/cvgSKMRrOmYa8Paa5z+wL6P0xKBE
kS8UojRdIN4MzoYgTVKPKUhhqdfs1WqFMKA/TBd8z+fWQ8eFQVVTyyYwPlJgIxOReyI22dUPfDTp
DSd10EjK4xDcuOW6DACHxHAxqoqfr/6x/Z1MAieQg2bZ88X030qUbfvZoyDc8MBfMDu+HdZZF32Q
4co+htuL5gwBXmQCxHNj/Jfzr9OnzOsB7BdFCLwY+Yyefl3oxqQXDq/h2bqcLvgzUUkutIaXF1e7
XOHs0PQH+jAvC+azD4mC0ARpbuSUAsdcVASy0ihTjPVKtBMmJAtAKxsU5kzSDnq73XK/WxATo8wI
SMw22eGDDrqhy6B5MuNN6zzTT+qfYdoZwcydDv/+PunKft4JJEsThJa3yD6Bfun5XULoylNcY9Nx
/OigCs68P41vn6TBrumNIsDk5pHRJtRTxGyLEvLI4e+UXXsw7QLZyic6XqbAviK95M4XlvWK/OPE
aghx4S7YzxTSUAutzOAJhDCHwWhCfhimzo4h1Wbzx4wT0ypvvtIO81on89MQPiT67qV/2XVPOv0o
jlrG0V4wR6x1eJnzDAw5LcgcQmRFuvAEof41zIzvWvPjsw+owdetxXjm4tlEN4eiDZWPKdspXWC7
jvbyEInTy2tOm6ZGQJ4xVMwnnr9ihtsbvYPHOagIeQ6yXs9Glq6njZldc85BTkR7U6yQZtpFGIL7
GNBtz5WZ+19kFe9tsYe7oeO2wbt5Q8Ug8SIt1BV90cwQ7B887kpYz8MjgUhCo04N09euCuOmYQgp
cSTXvxv2et8ImqPAmkNEUcvGIxT/Vj25YibvGTyi5GpiX9FQUAl1OgogxhNiaWyEELshiSwSQQnJ
f/T0xyoikuJk8jpQ5RB6jzA++SOGT0bzoTmzEWWjYYe9TCz/wPADEC1jY/FibV7C+lxx35j1UUNJ
blTk+S1ANKnlbypx6z6J0B5hbzVsGMM2JBclVGPQGby3TeiZqUWHmH0LL5MiHn/mJYQU0Dn/P7gw
UYP6mSHeDTcpaVvvJXunTVH7eTgo/3WQP7A+/GktWA/nOjP+lz4a/hL4d7Z+NeVtcHht+DFGBb5O
7xlpE8N6fk50wWnjnwHyEp7BV8qtDa/VauepzQx4QIaQuAJ1YGBYGxc9259r3l0MPW9/jm4mytcH
3GNFA4Ekcon5dBbmJ0f4bl+glQPsjhsv7IenQmNYw8RGRmIKrFXpZojkQ1kzXBZvdCMPP8UMx3KK
3Il8btwK9GHzDYrtS1l5y+ZR90WoSFT9qdi4tyrWuo/g2WjshVEYmESvPkil3lr8Va2ggH4+T2gf
XT/rWxOvf7I8cSH5CjgWRBuZayi6Js7XgbGXKHK4uPLgIcbRE5k8jW1Et4e58IfsfJn+8tlzF5BU
wK2V9Xfv0WDoEeOQUc81PEC69FJ1u3DEVoMSnZIaNOVMgwobDt6PM3NIhlTdP5ceIDN1h0PCEkDY
8b7nwpafbCgdj8378gg0FPMxd+vwl7YGTUPm9eKWcnuPqPJGQ1YPgGX2OOwRnFbBRINcDTF4mun3
HGieVLe1jrJ5WiNIO3xppFYAS2WFWL5gJZZGXpKLdTjDkZdnov6JLlpE5b1nlpDqUEm1iePCC6n8
/ZT+irwzyA6EwBNeXHBfLvzpu8S6Y8cyXDr7Vj/lI4vSf9zZXSrsb9349ClgguN68kpGNXopiFYD
6yPTCkgqSgSjxVGsgwH6WAbdRWuO5VY9wvSER6t1O5T7teZaNHZTmc8TUDwLGL3F+jKsAvhjTO3e
ZBG7z7afArRXXsMi2EcW7kS48fMdI/1IFvgJURkKFxjU4H8J/jPtDNhy0QmWjfrsE7n7+irTrFcz
iPdqxr7cywOguvSjfBvYeuZ+PoPKH1Qx/buQzLY6/yMBrccQr6EKKt7GfdoGI802TfAc9YK3GY/X
CRDQ06mqysW+tgCRzt5s874s9KVxQY5zQxswLpXLN0mmDnAfdteRN8hC+o9FcSCko8M/u7FjRsUp
1cP3WCleokK4BRaGx0JjAh7om4QRDGW7+zLDdGy39PtmDy8odZdFY1+QgmEjfFXlUWRf/4CIghlc
u/LvRdu6fFGtomUghkrF4mYSe+n2ZQlpqihv+JtC3yrXPG3CdjqHbpV7Dl/oPSJmPC0SLaESG3Rd
i2ll+8nQcPJlGKoHtHAvI2D6lGvp4EL4vGOG6MRiyla13LIqgY49Jao24KhCvlghe2icjEF9j2l/
/MifH4+IR/afuPDUlKcwmQGHvUkVpIEdweMyBQsJ3KsdW43MQhgazwjRKvCvBcLVEowjrNXGNRKc
Z/mgPItLacRrxZWMHfUt+E6fwIr9RRAjOCk7tUPJxVhx8ZfU23ZQr1Ql9z6ZTQrnRmLxXuhnqhxT
fw6SFZJp6Eh4qvhToxTH/6e7Pkh7M8gjhrm/ZvNfIg+J/vEh6SOc4YubvNVS33W3HY2PYpC4oMcA
FDxblQzltE/9+VJ/sFJxNOJ5m4u7D4ElBUpJPzWEhK6mS8wcqyZ5u1p7GRC0XgTwo/7wW9EADzYs
UjSDHW+bU0iYkXsLK9Z3kY7IsVGQo4ol4m7PAzuUVH4UUQlufD72It+ib6gxVgWQL3Gz3zZi5n+D
r3daXZ2PQSP1lvdEmuxhyD860KNIAyggWnoM0c/c9bYM9jQ6bklld51xuuMhlNZVCk8ADAxZf/Bf
MAKpFPCd3tjP/d8GxWY8Zda2K1BbCv3AEepTRU2cvJD4rboCHYcmvv6daCVi/vUFAKnwkWWAxH2I
O03kyv7+WRkQyezr5DONFwmpdBweuig/dk5MwT8gYnXWnJbPDJ56FrE5W4jHQVWCOZ/P2coOYT2z
7bOFnbVvKRR/gxDkicn25b5CaFEbf8v+yOZfOHXZjdyMzuHsRXeMrrN6zAgG4J6LMwOHm4dFSeBm
hkS2EX0IkW7NeVWmwFg9oWTT5ozrZ0YLG4QU+WpCNBn/UD0TjAUyDqrOclR3bUKXr6PaSmz3ERhT
ZYP1sJ+cZfwBXUYS9HqKZGS+1FdJil4ICPF7GsXNa+2nvNRMMY+LjQgizrGFnoS4TcDOhLYDanz3
TsoY0qU4bUAFsHO1w5iwzM/oEz0nszH+sCxJOFX0F4LWDWsB+DR9aG7b3dwoLwUuVnCorJzhwF0c
IggaD2wsbxoHARhZnZNfclWYX7YsfZH6g6NuGjm9D7aWt2lEqcvI0XjnmpP2CMJFzfGPioIlOoFo
JFrMIJ9lNZQFyMCgkkaanhXaaNcpEuke6gdkYD+kn9Z0KpIuXN1VadAm9Mzqd7vKjd/jRaWEm2m2
gNtSOmnHgGCW2pOl9GDnlrlpSXNx8RHSzejBR4LG6vdm9N4jvU2oP62aa1D0gXX15y2TMuu5i4Yq
9C86VD8zfjb95uNJcv8qfTJPOmZfnBFpX8G+K2oEJy2DDP9aIIb+FOAOJWOxt8N/jb5qg/9hI5J1
yUoWaMlnMcsFCKxRxfcwscDPizckl+wMr4GjrO1TmvesdKxOmq27pQORweZZi0REOv8rd2OX0X6m
ZuDloOJKV2M+oZ/t/9G7dazW7DGIxaIw6khzvIvnCXcVdd5FeNSjTGHXKHvnHzY/6+nXdzbQeLMb
4ROYLHLM1HvF1vxRuDbaTv0DHSYgZ/ykLQ0sojRu5LlBnnpJhEdvvy+V/hhB0PxhLdohTlz1dSGQ
NT5lgh9fW0Ang9TXQht1II6bKT6SMHvUExfcCXVjDWTk7cKN6keCw1wq4RRY2a7jzMDIaEC+OhlK
a9k/N2ZLthriwwNCVFD7sfvLtc5LtD+3DObdeo6OvlniqgaGF4km15xQj5nI/fqu1Lmb8l3Ek4VU
vXS8n88qveNMSLlFxVdEpp1Eh5YfpchcnFIDf6R1s8l5eDiR3i2HE0j191EGZLTY1ZbWpPq5HAN7
UMrzeyUOYB7M5FeTsYWqbZaWxoQiB0WdSNhRgG32BL+gqxVA5XIURFgThySt5DOaYx0eBkJ8ulUi
KrRS9z/Bnkn5Yyk0X0IFf3/PUKaDAovjlRJX7Y+5XRlUiSltA4b9slp4W7TYu1oTQIEJs/qvXfNF
AkWAwsQU2hqI27dR0j7kg9ESjJ1lR7kPzsi/7RrrifJAF3pm01WGTkeVGYh4XHLzgMUN2Aeg/fzU
hXhgFVEQmupmMLR9LvTZQKQOo+VViGUK8ShneqPLLS/w++GVI5gp/J0XE8UtWp0MxSqC9hsGX3zu
roeHQG3itokAxHUs50iqjwbXtX/5QdP6eWbIWNhrL9E53VCoB6lKd0QofQGGEPaY1hX4H04LLyEl
bGROab9vsAngl2XYqotcv9XRr0zhAVX+ehCwJIBgsNPocJSlD+q6v15KTLHgkb1yC3S65GX/40X7
cXnJdqDEfOHPcxUODX5fLBySXhbK1vsUJGHwrgG1bvkR4IqUdBCAZ9KxSRmbVxpQQ3g6xExY0wZR
q2du9ooEdlno8JQv+bowb+jsVzNTPmqJdXDXTWoSLWXlwekWV8oW33QR5+9nFchZpTQxPMBOP1Jj
u+2DyaPA58c2vjRajTFKGYZWlRRjjg9O7N4B/bPeqgZ/oyGUDHaDKtjUUv9MD8hOUlSHPT3c4Xkc
XfeZz8Z8ElARK8xdDOOBfv0km5GB2H17rjKvoWRBglfMjElU0x/gOTiNhzg6mESv51Wy7Hqcx0i6
3vhMGmVHhnHFb/dXp3hbBXfRAhZqenv85Ot5eZkMKJK72pnwiQoSX0Duk20jZSZHDzw/ThVklFSj
A8w3B06EkVxVNmYBj6NK9YQwsfyfdnvxvVuiIPHpOorPBtyk66ojSDde1g37H8IOxZFTCPq+QmjK
UYu96qg1eJF4xPXFHo09Ty9KVoJYW5Ignqv1NGU3WESYO1kBu02XzYtBS4URKfNpzbVcP3TjHjlv
AvfrzPUItFRspXOn547jdclOIIZvUGebcqz4GKuA3E1DcHOV/B73CONq9uaiveebaPrrGNgLm63l
zMlvw5cxL3FCqkNzF0HxkMOIGob+8VKlutlJCYROftC4ytz+5Nxei5hC7pYFk6axv0ROdDoRqTUh
zPN1eLiUZrQGqzVvfqbA3XgFb+XgudSjQ9ikkhxiq+qtEWNcigg5dF5L6U54ieJAaiti+tIyGtnc
h1Js0dYjh/KWUPSm6alxHMnpurpoTSdUSgZpRLhQJ9U+bYSDz9tEOwSZdUV5H+WLm7piVnqJqmnt
hjgrq+wMs5CBP9OmsCov+qweghCuxaFtnWYo2gAUzIbCHnJ9pxk6dGxubwz6XGeRm+X9agoZvO5L
nHPRevdoUbBiDg5kwU0g0xHut4Y+e5iwyUWcGDQps85wqMTbkw/7+6F5XEbIBnOl+8PbPbjW9cMx
4RsztQLQFFEKLm5t/MEk+NCUZeaJ6m6WfYVkjCHmSGIQFsFpGb9BrP/aXDLEw/aqSC1ixVfA1NkK
xylawIGBW4RZVhOAYFX7xf4Dh67j9BhK/TUPxB6IwTYiOlDCN7zptYf91xMaOoNEnyIOlBQzROU1
9895Ras+N8oTMMcWIPE2+BWConNT34r1UImgZDhqWVoxRD94ygnkUDCHj2YD/wQUm/Fxuo4R5AUR
ytXfCUf8dyOGP0HCGJoPoxfc+fBJuxNWAOHk2NYpaTkCnyMQXiSlCEat+xk9ETiyW5O+euYHNAO5
trch47e/tbgWpL/QElmgefSRGmcZLzDPWFwAy2XhQnBMHi2lMYEF1wnfOBvQElw+JqdgYFeb/o5o
NeLrjP1Iyf6QnL3ag1C/bV5bSj7Qoq2JiOsEs5its7Gb+RCvNIlUyQE7QmwQ0ZQMaVbP792vnsnU
eKDU4SYrWcDz6ArwGTjA4h48IJRBuyKc3nFeC5VZLQMlwSZ7WJ75t57e+eP5LJqo426FOxGlHyWJ
1Zc1sInnRnTEu1Ta3T5U4DRrKl20yvfJQM5TQIrr7ycJrN2gZmM0IhG0PUBbkx8LhUs04tqvRZih
rHKNRxVHL05dCLXRV5QQQSAwfoCYmQkYatqjr+vxxVgQVCEacnWNByStW2bTAYUGJ/rigJwTlAae
Es0zC8Z6SWEEUqcMmRTQ29ltHarJRIbwiTx6ytcaGe5krDlTRgF7+hjv0rIo/wL+5GhsnW7RlowI
vR7pYglvV5pLvuWzCjTds+s5nCSbzjjOCQwfdRalAV527A3kjYrwqXL+1Vk+z45XhbZMLw4qXHOo
6zlSCUBZSkVZMR/cx9e7xdafqmUSORLrQr7oEG7Ov7wMaTOZjy+21joaZAuZaa07T5h6TiQL9K+j
3dAmLu2Ljfw3D+pv9lc741qTMmDheFuSbWAO/4SslVwh9/8LktF+xzD6lYLIFpsSMDtuph0I4VzK
ww6IUlQCYWS4dHxLG7uTsh+jdnltZiMkZtGJwSwcAzjtDLXWzcjioQsZtaSmy0+kNyvoF/M2xM3S
2ygFHyquIepCdTF1tk/7uJtKiPmtR46ulmzVC4ySDBTc92EEK2jS70U660MGb/sZoaPqJTOdo8GY
bWz27sdRLhRHbb+NaXZZ6T/WwvprjDEYbgPPDWy84+IY+br5SYmZs4bwKtkZWoMzzDdniFY4zlqZ
ZW3Qzus4UNtH0ycsdJVy+Zp3EE3FJytCoO3W9dDy8F4TIcdxChyYdpGyWiaPvuvyir48H+C1iB8G
k799h8hTVfnxPhrY3qbP3+M1Fuj7RMOGcObUE/7zlYcsHOBiMd07ULjkzFnh5n8GHmZ6hAuXA1cj
o6uQAb5apn0/i93mjmc0hSgtY01Mhk3CXS7Z2xZfjUUjpbf9GHjYLCN2Mnt+7bbRZUZ/cClZfEWp
uJ80UId5RufqFuGzPX+fYA4q6HepdQ61NJYaZWPh6eYiZcJv6cEOcw5lCC4GGOquknFrVydWv7Oi
BIxSy7j2iNJs45dUU/gnA+7E4ynL3Molz+1X0uH1TDhgzMrQJCk0+iMEz7Q0tFUW/isrdS3V+uKI
NLQhZonVs2Mk4e1179KxlElRZLqW/oL3pFLRwSdP0AdpuO9M9L7pDK6+yW92+iPzNVvnX3Tz3BiL
PigPB02YY4ZMP0+7fn+ItyveSux04/IL7ilv2C2yLmIcmNNe58zVb9diMVhZuSLojeI9T2w+H/mT
/EJPL15piMkRQ/1jB5446/wII3vrN/1RPQb+Wt1IBIOnxEYbzr9Kz0hRIgDQPD4H9EWNulRCiNmO
EApcsuyCKipIMSaDB54CfJ67gEf5o3Lx6NK9G++voIAQKR0XycFb0CNe3RUJFeN1u7Av+MSeGrLl
GlN3B3o9Apo2Wzg6CBlvSM221LmU+v+thlT2PLO+Z343hUwqYNnBai9Q0gfnmKoy4fayI+RYWm17
jRjD3nuhHBmj/6mojyEmwPQ0NrTkPerpj4Hyh/ntKLw+KGj5nt4MczeTWztrw3YULa0bn9O/39Hn
86kN8OAw/2V9Jcw2CZs3fh2IwkEDulo9L8tkOjMUwYbvsu2yjvllutJnLcA4aQZje0NmWvTQOaaf
3PZTLCZYuALmTf68lHYPYZZWhyr0WK1TVGMcV0/8S0F3fu9WjATDNQcDEuM0UdnCaaOAGw8Nrpve
dvkECt+25INFWUOckqUqpScA255ZeOO0ZnO9yk9Wty8QblWZcycVNDMhw7O13lyy+YinhU6tmC7h
vrSzp10dl4ZyOiyP+IIM1I5E+spSFxjPjYXRfOq5IN56fh99fQdjaiOhhQ2xHsAuRDdnwDzfghMw
OXHm9oa9EOVVwlgYmulIoymYi+QENAh4iZRS6ARTiDNgg//NhT6wKbOalMooJm6icLbh1Q+vSQmE
otVJbDiXTR2qIatZr68Zem5unuJnTfdnrHI1zSSXLUon/nTtusEhfYR65XHlTa1viyNnB/BYH8+f
JaRC7SMq7qrWBVTfgQKAwywNZVQhU9uIlXVA4E/OftmLS4HRcJDGJjNkHxPGHo4G3g7ebNuxLUto
fCorkDODLtOlxFUdc8JENV7nlB4/Q0UT4mOhVHuHQ3KUKLd8FAiocLkWRui17LjfTNTW7xiAnqyt
/I8illakDHMs1/cFyeQ7or9lwGayOy/lWkmjrvSHdMTBb2an5XRjaruxhdjXNswvhxKYIWTbBVtn
JHAe5TzGItiVfRjUGsWVmHvyj+YS6GcjzoEJ8hXKnSLItwMA/15SFg9AaOpyK4iKIzClmTzeO1z+
f+59uT1zHxe/OqvZi6+gOZsAItSD4ugp/6/heZ5JsHIXfIWnLpeZ8QO1ZJ/SkCZ5dZqof/jfj7kw
Eb4CKJb41SVPTEbEycSFwpF8YT4fhUlZ2MWwaPeU/7REWQfvXWVLjrnEW+xTI7FlDuZmhtvJ8Wj3
qWL9tv2sCAitTP21IvBUmY5h7lTbHg+cDB//6+tgTsIG9/zobA+6bZeF7vXwWyYckq5MZ+7toPPV
9QdNvr1R/d9JTKgMsRvkGu9HgZgzuSdkvPDhCxSO6xeg3IvvcqZDLk8UNZhGr/2JemXYfVqgPPTG
m1mDM1sO+cRc9E1uKZQsw0Nahmgiwn8PqTUVsBcw27sTnTOY1bu5FEGJ9nacyCoq8OGX3eoP9cED
b1oqBiW0+3ToJFBdmRtc8PnFmvU4ineqpguErinMZ91Ef3SzfXoY/nbQ12Z6C1zhvIO+aIB/8137
cVgrhpR5ot0M7ekiRosxN6JCr8Eb3VT+Z0e1eqb4Rl5Pg0C9pEvd1kUFf1Hg9mMW/xPzzxEDtfY3
Tv429Mfw5tuu7apfgF7Vq/2ygpOPPVxRgdkdcH5MtXL28jTgDepdXUvdrOLXII4R81hzKBiKvsAL
jONzBIA3u129lluTgcddKOjauG1Pk6/2AR0BjEhkUgUhB5PbE91XPX2htJY6hdhxNs/c7Lqa2JLQ
H6i73IffFTwU8Z5k6doHvXE/VmSe5LVnqsP/+JAx05sbzRHWknBBYW8Esyt53rBglOa8DVjKBrRQ
3FtehfHI9JYIb00E990osMZpNKIDLypHVgysp2qpeibeDTLwiTRSappJpQQK099l8ga6kLOFsHWY
+3QhAiTIdmFaOYS1Jh+6/vZkDwpGE1LQ55jqsoIB4ntLpeOUWsOGDCDZeT4fNqr7MFic4KtgDYM3
m6vqZCDrSawoInhHMAdYo1V4SPTZlv8pUB7qF6M3AcIOVcVq3fajiSbfdXGrbDUbwDCJYvW7tFVw
Kj8pAoABP+NOmmzAv3T5LzqxazUDXWQqGb2hGaaea4c7hEzD0r4ZsSbcUojpM5T2Dc6J04YG5voq
zURYAR1uCG23I6JJ0rMWYvkpKnMtix2ZpeGr05H0EGJq1865riWH4tH6Mpm2uldnphlZA5adbbNR
0MJSv+xy052tkJ9qEDL3GMAjz2za4xM7ORNohAc1OAeRzpLB57SHSvPjZG3n8u47Re48V5aYnGFS
BGMYtH0y0z9qBJqnq1w8MgVbaZEE213AjSuG8V9eE7op+8MWLWO7kbVKojR1rFKsWe4LJaFOcQRr
5I3MTssc0nQP6grO4WAeY3PW4UR8+Bhd50xxsZsWphl/J9Yq7WAWnxedhVvAk1dcjgQuO4LaTi4w
XsuA4X8hnI4N9TMdUze5ESN14kpiJ7KcgvTfvoBPcLxOzVx2TWtKU2iOBTjcK7vMjbTRZ4HcAi5w
bCqa/TgmJdTMAR3hyaU4cvHxH6tXnzkE8Haxz/Vei9dWPtLnTdrFxEpu9/ePDEFZ5SGRuQXvRKR0
liFjXAol0ZafnS0DOJvSZ+pdRWYCmpSnP7Xi9id9SIep2LoP1uFr0lF8+i00qe08P6xALulyQPE2
XtWQY7TBnOIGjQtYawtdKD0k5PGFn5E7uCMYZU/CsiTdGP2dzxir1cSxHTvpU0FEiiCTKZc7UPFT
IpYAfRsF5bi4jyvColoHcI+uTJU7OVEEurQOmXUJWRMo3Bk3ObBmP6EpbueCQl+Rr701iC/khBVS
X+JENlodnJNTaRv7VNe01lm4aDkAyc5DykWy/R4thq4P08u+tJf9FaieRAQ4BrAoYH1OaAOZXLaA
FfEu8513m7qRFcYsh7Uz403SvLao0rd7CZUuqFpLPICMJo8tatYX0ABCThr6AcaIFUPmQjsN3uhL
aWyBdxxJjVWxoY/uiPsCEGpTjE0UQeU9fvDHjhaaOM4gpY2CjhMEyWlpaubFlPwys1TtFm4xmGe5
TUgDVFbw4FfBBntoaquhFoBPtV6LLCN8zxnSXMTOnk0ca+KTUKWkTdxnSTvkAMD2aYK33myyPNpN
sERK0mwwhFM09hLZqYmpfPpSUcmq3KFFf68c1o2Dvmn5i2mfSe3XSn4tncCla6j30mMdA3UQxZ4C
zTlcE3vnMXg1xY43WsgmeHZto08MDnOVNFc+3wngCHsoCdexMou+B2aPtUMPASN6jcdt2EYGs2m/
Lsm7Dw6UIpkfLfZLBa2qhtiFA8OgwAZG1VWO9lgqYcWlV9XDsW0BDIpEJy4ynGXcttQ97P7pSz4o
6IRui0CjckmnCexE1F1WcyVo3M5JTHqOnvF1Ssv3i+U+g7DQxLSjJCTjpu6gQziAPUCz2h0kOGEL
deT/XILWEOPNZEK3KH75b9dJKzBCIPmp2irjV0/NgLZ6ZiK1uToHDMpo8jK71Fvs/3xEokTC1Y1D
iIaGT6Aoz7OKgphWyM3pXpCKrBuehlGhVHfTIyMp2NWh6h7bvuFe9teh8LSpsPFLvCq54tvBP3Ht
yYxraS4x8aRIlLANApfCrSQ1IMndGzn3FJBopcGg8EZByxIz6JSNbVQ5oFBvmiZSXZnr319bH0Ad
3SryuL9jGL1WBZ8SqLDZgOAFfNJP7xOqW/WVaoRCUQp6BeONa3NInQrOIrvnIFBBZKaba7/FZyix
yxTLohMriSXiXSeHsK7E0S528kFM4+wtocExPpLgxLaqqGywtFoZ7sYIC7U+pwGpGlkKEA8k2HNN
5PeQ3NDVX/Dh6G2RFTGv4zO9shDH4dNmYzM0SowMm9+LFrJ1+l4w0WE58VaaYN+gLDt5KYuT1/Hu
ldPRi1+hZOwIq2OmWQ4ITlKkkxaAPuzVnUmQ1toMiBm4BBF+7s43xFn0pBp2UBSayM53Ev9sz4Q1
q7dq5v3vlHELp4SI2NK25jNCybFLGtylBO3jUJqQC1JJwFc+mT9ecKTdiEWKsU9vLvZZb2YfHEn7
8trxbupbk7wgh12WaUcOWRujXLCsIrqGxkP90kpsJs6Hh0I2fFjNiHGKqS4KzYTnoHgk/Rm1xLaE
29AHD3o5ImKpir1cJqQhTSQ3yrd93UFrzu6kNeMxEBz7pz3Py3LoESzx+QI06a3ONeYdDmED5ZEh
uEo/Ksdku+0XQrClAjKiTemr2XGzA0AK3+ViXeE6bc1BPDRHTobcgGKtYrc1EbS470gNflKt45Xm
vWdFPZLl6NYTbHUbVP8Z4LSyzdMzji0rgFqCj/mCqr4wWv8LTKwy8QZsDOUxcPtNXXBgv72l7ixi
JKJ4jWk25hiTlbv647Zb0UmIPoXwd/noOwceHDtizNvATC1GLLNybZ64fVv5vaDbTNeLAe29Sj63
XTOULZkZyK8PtwFDkG/DOrn85sIshumXhMx26Js469tpKIVXPy7U1uHZ4rAcxbeiFN7UhVdmTtNr
L8ICWvHXodc2HJ/ZsVYPCSeM+GU/2nGAg3csE4WI75jMGa4UjqErOgrtQQ9YVz7s4OPMj1povhug
JwD5wV5lT1+LXp5XOVm9LS+U9grOHtHLcVrclN4Cdf1S4tJLOooNpqL2zI0MQksJXEBi5wwX/58K
gT7l2R8ogtcGmKcbpnO8aGoTmLLkgeKnbJU5FYgLV5bv9dp+fREQLGQvKWo2wBNxyKn6yL/GNYrE
jrN+6xyVL3yFgsXIEVlvxBoS01uxTY5oeqj8+hz6yUEiy+ilgSNfaEXfWITwZMo1B2aqPUAyqo5Y
XpNl+lSAIohvHKjRH3FsI6eMVoHxqeoi20gvni5yTcwrMLSWO7Qi3e8FgMC2I3t1i2ciJz4jUA7f
syUQQVuxa+MK8lOIyuH/Y90gJxulCPDhFDqmg7FNAP2JSnoMi5K5YLWXfijcPRG1gCNdq46483at
a61uFRXVdkoDuJcqRCLthTU7gbe/VH4aQ24CFXAJwzmmzfupTQsl+6S40JMEXdtlS2/jmxh+ubyf
MudGAmK8Vl0UEJXNxNvo5NM/iVzAhUbNqMPXFqpbvl3+sp2Hld540j2aeEVylpn7DXez48spCIJB
D7HK3qFelFyp3L5GPLgq2DeFXoY7KIf2W3BrJLkg91gKLX2Zqt1uslzdoQlDm86dcqT9RXbpd/Bs
NVsq3Ko5v/bcNip/jGOqly+Rgc8ZbaZ9Dc5qMeV4BzJ7YJpVuZUOI7YwxO0GqTnMm6tF7uvCOqj7
akoVgxGYStbGGzbCtpsMPxxkp0LrSv4f5xHJJ+QYrnC3bcS/W5AC+CLYcLtT5uB32/awr020kPoQ
VnqebQ2jv5y+ca6GGLjCsph4qQ35Y8kBMM+PkL1WbxzvlNt3TXuZ3/XM1uqy0BCsFkyIqx0lUW50
EtPUMBk6JnCKEI873kbcTIMIoo3fGdBJwPGtpy0qZLgcSobXPYqa22jFMyblgvAWlYo4oMEuCg5C
Pj8ORYm7XXBz8z0JuoEUJa4oT33XYuvNe9sh2cbo60ke4gj2xoyoCU8qLgY1EeZOd9qWE8ObFjbh
e8kjJxtrrG43po7dWtDZTVYebu3uA0higPDQt3NQ+Die/JTYzGxkRTA74a+P6qNqXMqPO4zUErTo
oUG82DsbROLvu01snUwGvIq7+2ZyMWxlnWgR73LCH2wW+/OwbFv9D5kyyThA3XqPdLU+/WNsPBUv
nGS1831pY21gSbMByzg6dsq5utt0ZLN+FvqqFYUYy0yuMnGBHvyeoNgpWo2oUFE1ugi8Z1/7TAzw
koC/VYUc3pQMuieO6XLLwrRWNJ7yWXRnvCrTlKW/RBRhryVzeDgxWSqta+g6ny0nqNOB6CAetWFh
Xzc2VegwDvQyF5cTEhhdIhHoVXNLAfaUj37cC3F6AsqqsqN7rmXRIlBXWYnJhXqHnYYakFQzGJSV
nSk1hcHiGI28j7ZHVmeV40L6P3We28j+ASMHUKjPlK2QPKr6jS13mGB2gp6ZJTJQDWm0omRnMc16
JG/mQFL/dbGuQyKeeccztuec0gu/m6E7Hhe7h272myvoPat2o9vrEFaSvQhBV8/YbmVtYp8By4bR
o2KTDp6IByBH+4Pl8alcFbV2WAoHhERZ4gBR5ihfPCUHVVC3SrsTBqRM3WaCeT58kA6jLg1L78M7
FcMxNNpQMwTKQRz8YhpfYvGD4Mk2m0PMK3h9LUEXjq0mwo+/UJS0HEa5Gw+3WMXT9gGABCW0rBAM
dnFqfaVCjbDDfmM82shmfGliERw4CTW5UXmpAJlyuIeg0y7Wf9f6pHRRGvr4ouxa/j0Q/if3eRnm
88HC8swnDb6J6Y2GaBIE4rGZh2g+92vFn8ATW/IQU4AzSNgre8QaHnjA2eM64WLiwnKxJjJoo6+P
F3UowWILe50NvV1PnH7XfRTCfpOmY1DgDPR3HVeNq3x/sYs/gVtkCRFXthgyvmreGwa3HslugGbR
FNjMy7UxwV9rgadTL5v98KJGXM5mKSnolLHJn5P9VHTs8wIy77m7yCRRPaJ2QqJVk1YIMIVrPMLo
XAJP6cLVoudR6q1qBduD3NznXpsy+fewLsRc0A+NlKNJl/h4O+i7Ua+2V9StrIliJCF7Dek875xG
4jqrJaad9+kCysKk7cp1Aig6M0vxBFgklGgJ1RqiI3byhv73YqUvZjXbAN/w/gOvqVaKnZaJYuGg
ikvv/pj/iAoXG+DPRYL6tu4iiT3DoltNTtY7fJym5ZCJ+G5ZSKBsIjIOsRUSJY4M5gn2irY5jZAz
eb0o2crJF28d/Z9YFMtoqZ1pamvuwA3yC6ogkmtw1AW2DUEwoNTFFXRDg6oqNUjsqZn6GeB+ZGiM
xip4QoG8fzzEnyoJ9FPUTQNHSZdo0foQXw+kmrF6xEPnwvghU34Cc3NVTkOvheC4vCqmB4h1twQp
q7ObTqnPsNfIVghijjNyFWzPUX3P0rkUHSrQzonRfWOb1oAD84NlstyVKg4ywmGF/AEErHHg+8v7
GWTfOGAKMzqPXcYCldZMi0/Lc4IK9+D3v56zajg7OLE6Ra74uefbcY2btVXMv3M7So4CdYZBv63j
OZgJNJZJR/XBBK7HZA4lyj/ZVgAyUNKJ/0a8hJBNGazpfBn8rgJVrP+IKHY786zOQ13WjymgzDLj
yZSWRGK8sdb6HeQySOAn09iIQnyWD+IT1t8Lo5zQD0iVtbWpfW9HBFn1WH1k7PRXg6637JIHergl
jpW3LZg2uPeNsnuz8hTJyRr0f9fC8+wbj96ub3vaLZjhkwDZDy0E4iF7pYNq0HffUSZptmAUUjb8
/xHkQCQPeiKX7pfud83bQ5bdVnEtLUOp9f5JIJu9+MWBl/6yMmV321wz9/eielL4fokhycPLCWqp
BfJkZelEDJnu9Tw41WyBzXEXwfSLMi5QL0ZPr+nbThvzbYNhRS0/q36k6inUerD1T72aBYuRFJfa
n7TeuMFTumKY6hudYeT/uATuhPJVVtEcdflLR0+EZwFKNplLauHYtfUBNebOliS3/fwwI6uThR2q
wvX8hm1In8h+LC5UhYMG64+49Pe53/xYScjehjzRKhVtowf5rdCIhCcELLVTKERXTesyxFodKiWX
mU1k05pUAemud8wDCWaWMlW06dWbSzcHBONwA0ODJeibnwBXqSnbpV0wyTwI7WO1B3QBd2KAr3Oi
MrSrWbDoRiAXsiXPiRHzaUXuPpY4QpFj8qv0PRD52UaFLQS9KXj+YUjro4Oh1+xpIrwqKh0TxZhr
34OV0tNepHsU2zLEXqZYoS7I/6C5hz0nFpG+Quyik78HhAmTe2iblDTkHx55GS2plFsJkWwjf8V3
Rg/ZU7ppSBIh5ACvgFS/o0IHhKqK2wW3CobHSbfgPU28USD8O95zKROy2ysjNyT15/rdiF3Cz0sH
1Rp6ICrdFYImnYxdRLtysgkfZzQtu9ReWqyCfpHktap7DWV1Kpz5T9lt/BVfY/E/Av/bzQG7axdp
1EkIQ6QEYBCM6NYcyznTnQ9hTGVSj2nguv4qzoS6Ljv/D7f+4zXJyewuuzH5hzupp5lGEGSRxa2H
BPovt8TiPmPPQDsNqO0sacJcsOtSfMi57KI2P03m1BRxCKlcEr8dwifIERcRSDhjz7g3FGrS+/CR
HaN4cBqXnpY/yDIpyvVRCULMgH/ATTM6YEGJ5iVSv03nlT8SWHydvKI+vgm98wvQLfd/Ha5BRKZw
fyMtRHEo7uO8XAL+hGft0+2cYuryNptGzn4A8IBmJxYekuX6J1nXkjwQNCfdiLK7/BgPZ+I94z33
HmGZibdAjQemnvgQRjWesFEfnl+szYjsOWyvbL77VT4jYyZrfEXCwUSMQGpvHcBSxK2B4fYR7ISe
cgXsUra44SlGTRpCxnBExpzPcFUmud00yuQZqg5wttN+FBi5XKiU13+ErqCFEFXEaRHXbSR9xuF9
M0Eo7Te7PkoplJ0PmPPizF//WjA7L71ribEYDNkFluePiJMTBZNKoZTNGm8E9VId9Rs8lZXd/Una
1Dy837TtSfKDZqwFQfVoeo7V8W2saIih4ITGPrd3E0sTqS+RlxF7kwgvEzZsUMdCWezKaZkvTR6J
LgHGZmoYvL8u5t6WBRVauYBGlaQerdJZyiQgKWBaChx+7Q+irqYYKjB9atLgA/vSIKXf8Ir0qsn+
hTUfRiS/BHwXybF8Zen983NOFN1u8r8NFkL6LEJ8W398eoerGdYronq6hAyGtuCPS7JPRciq5mVL
AV+MWFZirvgbL3abQhtVIVfz425Tl3nVmeEElPFuO058sY6ax+i1fxDOdP3mXtZNP6qUpgdhn+vU
xA6/pkV/emTkh9ZiGHEf7R0MEqsAMltCjCCDFuzZYLHHMUoAb1tyXD0dvMJkcCWK4AUDXA8vfGFB
t9ixlewnLwHJ2PJ0+wdr0XkPC2W1JXEpMe1qwDb4FaLoBMs8086yA39BSzn4QmOaZGdiIwRq9sIg
j4hyageneqB8klUFNDOSLvwV3qdxOanhKn54zl28DsZjZBIdftmAvUaVaeJJEjOGv/gSsH3bEujq
0zuc3cd0G38LCIJXB5k04q1VpW4XMzEnU/TJM0SxVzZmR8Vj9/frVdMw6jDII2pF9t0wsHY/3tl7
ZSxP26lGw9uNsCXDcMV0IC/ppJyWnhIxTPDBhQkzScjDAznMveaPKZ+9bgaQjwbkbi0l74FVznTR
Yd/C/b3H1BSGi0S7Z4yS0rZLcv0heIOyYccFd5YR3UkS97ZnzkXciRLk52SosnANC3M/m6aLeI1j
G7PulRTYWr2ucm0TLXrUw7IIbO+GDbLcQL2jv9qABx80M7OMjRw5LemlxhBnGk9sW8GJ2iQ7jL+e
DFctgrJK6V89VjU3rB7deABnfNGYGkGfQ16zfH50jGzBNjItJdkZPmTiWqD6kmHXm8cAC6iuRmI3
7tL56R42aqt56KV2MamalG6aMLeXLHfhb+fQM9wMjiMB9R5EO8+Kqfji+LhJuQmRI33E/7rmrqOC
fPkwX20DKPcNPubMh/nSFEqzpKvBDB4iRaUi48YMR/nyVoHZJRpr/3NqWw4zRQteW04WCDBpgZcG
zf/x968wcrWP5jQbbzEDMWfQd1Mn3ni9GjO8ExE+H4VdysiSSsIhwqPlPgy0OGdkrd+YvlALCh4D
8j9R8iQSdNuLFmk1xt9tCzebjH/kdrCVfaA3EFWcTiwqcXT+rIqNP+/0xr28+tLsktbEM0SKzVNU
jZxJddueePBMlR4vSsqLDoaOvfiTr6HkENLOMhwERLprEhomWbXzAk3OMfWLW++xQztKIVPjadAo
kkID695TqsxNI95SKeGASjO+1hEn8P2thXy/5/bTXUutXOJ2+0XXN5wCu31cqKECKF/t9hSpUQU8
rSvn3X0DURaI3jt/qstIpCTaNc5YLnmfzezGHzkaPryk33DQap2iVdmsmq8YvxmXw41TacU1EsR7
puYEx/WiUj4F4roF3MQRlmQl0c3eKzm/sXT0OYcmV2o6U1tx0+JrzJ+Jbe72KvnUybRJ4OT6mp7/
h3VneO1fBbbO2DGWLYnGLzCc8AieeJiD5co8SPjwWnxQ3+BH9d1NiBSrsZRoiv82GaUsCx0Ww8+Q
Txio86B6hIQPj4l1JdRHRs6GkMVPKDLu1+11AftWQFNfwtkRb82pWVm65yX3gt0sWA1xv6fVzfie
2W/FQ3vRobuRDT4SQiTPYNOL+RYoofIGY0JYOiIQ05sTf0TsaLvLaa7ki4keeTcHKhpSyWOHsNUt
35QnhZ6WAFamyEcG1tplYTyW52I7Z4heoDQgWxS37SKFim0XJ680HmziDmBu5vJJHPLRCPCwlX5M
SaHs0Zq9AoaF/3ePTfrJCZq5arl7GBGuEjFFwg2ubULJfNFV2ke7MsSsp3koD+34IYyLvjsX0GLr
13crHOihs1ziZyFcWHKsGRZCReFl1OyNKyys15RNothxiqyhgyREbHunCh6Um4hw678+0mPwj6jx
U5YDzT1aOrKuxh29npziI/fYA+Bu1YeFp3ShsMlr5zh8/Afohzi3JPn+mTWkDi6eCHNpajgBbD6W
NboeVBlQlzIgA/r6SqFPpfp/+SSpU45EXnxfNXloNvm+5KwdFigOAbpwb8t/Mvdf4s2aga/TlqPt
W3yY/mAk2WgQ9NAnFgd7bft5XZFgiZ3FW5GyBJG+QU30wdmyqZlhSAk/AZIKm47vgBp/Yn8JclIP
94zDj+f4+/m35fyjn0WR9nNWF5pzucdKg8/TrPIaO5wpNGFqcwmzCNODjyNWAFVhkVRs2iwTEDR9
84ZXP+ZHIzYs6owOuxUbRV//GdsOt69OIL2qajWDeZIDMVtiCk/3F/om/iYiwY/I5n49EiNegEuw
Hwd3SyJy4OAvYQRg+3o99XrtAvlOVMOLnfyZe9i49uRwegQw0YDT7Ff9RQvmn31CSZcEB2HQALmy
fB8gJbVNGgYqymCNUCkbUVxm6TB0N4SYCQnodWhFWbw+7mjaMD31SkIRpglfejXRVTARcbEQoohq
8PZbWLUhdbzTmglU+vGhQ7UKW9CZUQDNUR3wyP4+PYiGVhpjjXxXGVf0ZZ0sfex9HimcCvwlnUKM
c+47+fyLDZ552ehJuwXov+jybOz8Mc+4K5B62zDKbDuImsW7iN1ZK8k1K4JZOdNX+idUwiF3Q7YZ
Vq0h8UCviXZglg/7+8kdTvPtj343KsiNpOMTYiG2D7tUvDI4ezbZjH3v5VWJ9dCn069lWrkRHE0N
Q/lXY9PS1A3V/yYU9iNpNkLjzkHiHA1ZZdv55E0LxnKOQ9IpLwtIj1674m9NrlqMDy1BYAV/InRV
5bFBVuOlfKDYlCWxc4e3bIyftLY8AmK1neZ0WuW85rJEPydXyn7+yDVnPJKfAvOoNHcQxyk9GI0n
o29GmO83pLa3Eg3TUWe/tHBw7qR1t3ghhPxBGjhoZIS/TBJGa4pIX1Dg59pr1coQeZOWRFFWwof6
PBIuOxkhWvbjQfi3ZvhT5o2uRc9yHWXbbIurBF1In/rZ3CRS8kxB/x8bMSl717h7tbvZxW7lqvKs
jWbdzkxmpZtPW5xLLXKmNsY3isuX98Xe6lyO79CV7F97zsgJ2JXlwKgjIDAVBzZAJzB3inxy6CaL
20sLb6/gOo0fLEIYT1EtRS6umPQqU2MVHcFP3BziK+rv+Pq5F1mNwyFM00u3hsaOo6sFL8lAZCX5
SA37Ecxq2bWqePuHvBppsOAKKjmi8k7oiC/hM6uSKnt8WKZ6GIG/FV4l0GBpldHi6GJULLBOtzsO
0o8jerB79HNklIUOjPZ1hvv0cQIxoXO8tWSRS1V2JXTaX9U6vZ5JfNQ2QA6UqvaXpfBIaMMCzHWX
0Uiqm1mll184SH5PZRX/vwRxt2UF1ySx1gp8PoIrMLK9QFJX7TzTCcOoIX7G0xDQh3R5Rbbb6xWY
Vm8mzFuMO0kVyC18WBEk8V3WuazyBffVEZ8gt9sIGpG+hikGiL9wVqY2SC3Lbki2JUkVthfo5bxF
cy072jxW9oUhu5mGFohnxtASZOXFOZ4ENhEdhMHNIYPRTnd9lrSq9lj0BV4v38n8zmIMkhSnrTBe
TkUJ2L116dHBu3Y9J+KiNebRBvprPmZdJ1GHnX1qlYxLS4OM0D2tCVD3xDn4kyrCMQJNDaGJGjp9
Ee+LJgUpGHB8xtPkMBrymw2ZDZ1k9z1YSpjwymeCh0Wa7K866JBkMY0e+BjyZ2FJJr9RxGOwzN7v
f51a1LyMllTZVx8zGIE9aV6NH+gqLWxfwaLX+438M3kQC014MqU88V97fadv6P3BBTJEeiXojcvB
gWhMAuMIcorLN0gDcT1vXrWTBIurwEmxbqlMwxVEPj9L4ba/xujMEldgFVrlRBDGiBr1GrYGOrKz
qR4J+kRFNOJOIrQP2GwlaO2T73C71nkbXN6ELzohlnGOMT1wGK6gQr35J1z2D0vP+WUGJsfBZROR
DonR2BHiomvL9lr6vERo1Oex+xIFe44kEU00AQKc1eaHNJUqz7Un/okIF8QM8qGo8e+Sa4bN0zLQ
R5MzcfexVAx03LS22f1u/ebuVkN5zh9aIK4jo9Qzr34/bYgMnU+/oeU2J7yUCeIzqdAMkXfETqjO
2m/6WgtyM/vBnwL1qbjfy5Zr/VsqwPkftowZ4+l+Uk8nE0EfPL9hWE0HZP8GN533oLT1YW7KVIjg
ag1Vh47lSaJw9kYR/PTR8p8Nw682TWoxO4QGT/wD7T76AqIioLekzV54oI57OiVbHvYmJnyhhPSs
ItnSNeDvCJ9McdvAVL8oexYgPZthBADvy6HILYOGNb829vuQhbwmBtK9gpDQAq/8yDFQbsmizpST
pzTSrEkj5fFEHMR9+sOk1CmUDfKmnM5NJuPbxOPmUarRHgGU/qxVwqrwH4/w1Gd7uBjtJIeWDMc8
zg3RDt18JeGtksKxMPmnDXyFn7GzZl/RN09n02yBLpOunSbSsiuyOxHMM6SgFnYWlnkj1HW5Blyp
vl+eo847FUJOxv15Ktno5GchXeeat/ESLeaWvre2Sc4A1Pnt24aVm/zR50KhdaqqLDLE4zD2CeRq
xZZxTgYBMK5RCLcARJ4MeUPMbAuiJbnOw8PWfz6Tej3Sup+C/hBAKRWuigHhaJUCBN28e6TZic54
WasJUw3aOwRXLQCyBlcJEUvbIX3c2mAxTY/UurEgAaQ8Umof5c1GQHObG+sk4y59Tn9j5R4DfoCj
qG81RuLbjY1DQT381SmiS1ov1+OrMjPn4iEbDfxqybbell6OLmIH3hCUPW77u/oLYw82s4DZ70a8
S1U6QkX9hs7CzhNy6gsOv5Z5Q4LFtllLA7G0ckiZTcXdyiWjbz6T0bB1Y8nkbcrWnDPyEHjG5yvX
8Q4G/jPkbGHkjwUFxnd5hy/loOd2iKLnt0ZciSVXz0Ru7FvUYl0I4ZfRE/wn6DnAOz3+JgoN6oU2
z13L04+2Q6ss0mXvPs2TqSyfg1TNZiyqGExw4pHZQitOvlOkfMrZ6QHAFyDP4WFJeL3ITJs4lUSg
Vju/2+aiHNoA/gyfe9SdVvYmOVZf6bOizJBLe5Q5nvzvSRb4Hz4dUm+6aWGp4r0lQA3ykoYCj46o
11I03aLUnsVibS4jTGxyVWKC/wBwwWw6IiWtRZzKBNwYdwwDc/0LNaDeMky3a1l0NTfVtS23EimQ
DEwqZ+zMZuuRpHPVfutLdShTDLsINH19RPFmdCuD0PHT+fQWVhgO3scjj/FzkQNT07vuds7XEpCj
Tpuo5SthVUs3eQWkYKHTQ9ZXcWYdKcU5geYb1IFsczyuR3GJ3WF8arRKBF7pPUKX98IaZU6yV6fg
+NquoNR72fOEmXQVELvBxBDn5tPIEZyciwFJFl3cXUnxLIuXoaYrWq7Rq8/T/6axrpug1rDgAw2i
EyWqOkY3w2ou36nG2xcNm0ILE/p7bAhNF1L6gM5TIiq0r12mazQ6t21kywKiuVB10N0HkYXcI5GP
lpzZE7JQESGJy7KfK1gSj7udOkzSmwLYO0FyuGw+y5i9Ixv4nWNVyICKolsRmOGPvB+n9LZ3VhVp
EUiVQSCGv1D3AxfDBi5+wVVt0VG0cGQKP1WEChoD4Ufylf72+CVwK9aon4ca5AY3mgS4yfyLY9s9
4xr77WUo9eeHc6j0XBtZiDpaBje9hXj4TtoVxSawwgpx0E3rdP0is0WFwKNQ0BgG++nMcw+dq2WA
djVL7lS5/caXghRhR//Na6r5WWQHrZJ6O42RMeoF6IpHcvlSUE6+hsVjsZ5q2GFWQuTClH9n+IF8
WIVfrkcnq9M3159C5NkGLCz/o/bRrhgJBF86xpFEeowSgZK0we7JZtizlW2MlUuhh4hrtuwR+fSD
6QdQD3iq+lh1hLIfLFKCw1Of+qbUb7QSxRYaTEC0t0GG/5/DSIwiOhD4WsV9GMrCCHX8yFwWGrO8
fZu85uuk4m+EbUvNpV8RWwIvA8j8bjtJgZnJ/Ba54X6dPaQXZ1Lge9Qci1nbzy458vKnR119g9yT
sDEONvyD3rXZiQDkgMrxVQdllJF/cRqqU6o9O3+XdJR1vM3LWUkRAykbuAC2pqYhKQyKf/z3hF61
0rJQe/Bh771nzzcchJ9LxnUG50EbzZ/xFbkgLxljmn443Y4mHjnxwSFSIP4xbiRqLxVOnAOUJc+G
/QPEu3YfR7NbAgN7TIThPPntqWE2NMj9STcFHo10Zu27qggHWwaw8ubmn/wkk4HxJBfNp7l/mgkB
nqJBW2z0DL7DxKU84hLJCyKbavr02oIOB1d2Zzu6FD9fM0C9c5qNTH/PhMszGOg96tdcdzRHbKQk
bMqzm2I/tn2jr7g9QK7omDMX/Wo6SZD/4B8sjkzKmw+KsjfdgJt8wSmDe448JV8FaPvbwUaCNPJP
V+31FPnttDuwuy1TUFg9Ex34TiAIBNpmR5KpWjIDzol1ksOrEOICBepFAKAKpB919MkkW7gAp+sW
/dAoCjFyHQiRhus6OvYFaF5P362k2TnZ0Vxc2z/UP7+whszNBPvrqOxzmO0ZuMgdth1GmUudtsC5
5bsfVB/PiF5qpzZN6fr+J38FedszVLZDYMPiSy06dT+RFgjq0Tg+TeE4MNutGfG1QLyOAzlqPMxy
M1aZnlMEGBe2sGpfouOYIQoPtRBpmnNjqS4iyz+kXtpOV9PPurHdPGaJMiUGfPoRPfXKHKFCCeAX
IYTmCLPlNpH2csE1JJnS9v458PA2MNKCeVmZDstTTWERI24CR5MOfLwYjYZF/mU4ESXYKUZ3Hckx
1ElLVCxm1183f67U7WY5TXWMHHVi0TipeZLpsjSEx5lMho+X+r7AdkLRw85ARTKXg8rNJnkuPW0w
ZJz/aP9ycoPCgjaG6KE2fBXySsGj34iKqlPQmchRKk6eRhTEAWQtRMhx0tZZp1EDqm7I3haaPqDQ
Q7AgcUW3Cq52baQo3Fqh4e4VWIxZ5CnwTOUZgzZaXxrWdmK96KLignIKTvAhTpgpPpjAnMgITy6g
xyrR0CFtYGBn+48QV4fh4GsXClVW77oHUmp8Eg6oYKNDvfMv7nVlFQ1GM/kPBzMgWCoiRWLXdNey
iISQRtv/ZYaFkZyPndVmrAzTaQEwAfCBkYpXjpHO4qEgTHieRMHA5KQOGekarEk3PDgNGXkRwWQX
n4E2LLLwhrC3oN+hqjhoiEefmYQ3LhjSi9WCmS5IfD/pQo4KlCZ4WDyHJ89Kb47R7fcNX/Yzpk0j
96hHVHrspAJQGAU/MvviwMuqxb0eYgAYy7oiPUSI8NhtmnRBfNtm8xg22aFOfTYZw4HZUmq5bMcU
/moaczdq9DfZslxNwkedNuv2PG5CQNK7tk4+3E/VLYicEv3JDfFu2JW7YLbzbFF36vq6G9F1LVCO
4GSAtgKbdYWLFN0BJXfvRNpJLUwZ/V9jFw3zv23pKDnNOjHSzXHqk6rud4ttikZxEKD0sa2fZCHU
HgXoo+4b4CHbF3T6STzddmTP9fphj0jHgWvZVO53DVeaiB8cZICIaHluLZ3KZSPVqlIuBtfItOEn
2vogTA5M4b96k/VJ61ZkGnR6UiTkhsUNiiyHytOUxIlD8V1aXcIo7QN2XU9TeyuQcJPciCCwMsgd
P1G8CDzqp/KxZkRZRlgxiCaHt1GfSlG51/ss8u5IAOony60skD3P347W+fbi51KEgCSnmWqkKI1Q
Kvd9AICICkvuMbCdTwxAKHrIWOV1JrnvISt/Kp5UdSKM7M+4673svhgSt1iqM7rqjajy2yvUJfgb
MfoJVa+pS3o6hKzaqppxhLvYht6D6+xPES2xOgrvhiDIqjjEwLaWkoHSO8j3/8o9kWq2KrXm3uwS
/InVD0LfZj8UZKM1BoV8DZXzqXiCoghBCcFeGJ27hPNsQ4rEpKVJgpiX8H7g9RJvkPRMUmbLxPC4
1qHHvUwut8kwnY9AUvOlsNBmhUiKOkYQFyrW8JxhVdkDp1vcS7ItkyGUhUDdiGxZmqinVuJucHib
zSJeOMMfLNbwVRYH9b3gpnKGle+xPOv2mqSMOTj7D7CvoHxldm5bRuMS2+ljJFtDvfz+RYDK8qQd
K/7OshdcrtLufYh4a1Mkv7b3AuiAVZ38c52INc0JzJkihKFlFYBpaeB9jTuoY02hMLncDsFQEZNZ
pdPfLlQzujf2hU6E6HG5r6w7V9cbpGuzItmRkeAOVVPosmPfiHhDRKyzAfmgjT6Ms4MNaLmdhtlr
N9eiQLq5VanA408R7euKOhMzDlDaJYoqguzLhg/CLWc7DqmfKZtmUu1djCHumEh4YVATuogF+iek
q2JnXoi0El2qzu645bxQpGSZmor6EOBQvkDwvGZnBakp15P27C8kQmFEUtJcftj9SKS/UYN6iBHn
pgjF393j+Q6tbqTFLa4iTk6EjbfNHs3ORlnG0YEYS2DjTQZtCaq0h9SZimrOj2NJ6DyzNlokz5mT
o2nGBsUNSt4eYPbDL51pMcIm3nxL99B7ablIzDh3Zv/DlWtRRnhfUz22Q5L6iqECBRbU287m9HIX
6hgxQD0p5/yEswR9CHgwffIvGQyu4NsmzRf2NpseX+NvYTRKN5YomvekF6wPgzLfL8jL7DCnkbm7
xbPZf6k/5b20CooX7HZQZvzbnT7NPIb20sKo6v6V+tIxR9pzmk4SpaLKWsKJm3On53jZmFfyyn0L
t96DpXRi8boY/WWtTTL6/GZwxZFYe/WBLL5qQDm3ZzHHtBlS4E57hx68g0l214VdbzCJDwq/7oCw
n+CL4AlHtQP/DAbrTOUJ3hFJUpw3UBeGfslQ8YxNTWO8Eats0g2LXO7A+HWRRPRgwBsNpO/O4ZAG
ihbQsZC+nUFTE+JhF3X79onmHCcMkblaAYHjOqymLtiEbriUc2fkHyvSbLJ3fS/uFlVsU+ESCV6y
r5N7z/D2l5ooqWHXAp0vhMgfnESA8BTHzQI7HwtCfzP1gW47fjUuJJGaDk3o6eHg0m25SaHl4yMH
Xm09MpS8iBsnXXVZUFoyMksL9SnxSYJYFjQLm/E3UfCoS1B2YiemGGoXS5ftOEiurBiDwjhvHdRP
+8CiQe/+3g0tPA26NMOtw3J8VJPpcjyn/+EUp6BXwzI2MEY9K3SDEIUQkT3huvJfSsh8YW4jX4Wo
sPen19cBL4mtOfoWHgmlUrwjPNr3cxdEImsNwnNQ6eQGBpoJCB1Gdd3Wv491QHow8ziLzCnDRn4d
y78OQII5Z4PkpCjcQnBxZVyyHN1f5ieU03c+uuQF854uu0FieSzlHy0cVuU08GBZ2C82I2giG9mo
6fBbZC3WJFFxxCFS9KBTyp0MJ7p3Ui1EuAF50EeHezhhNwXAXhxg3ySW9xzjOmtW+SrUE25UfIgi
fU4scQPlFWWTPtRr/C6g4zLMSve7aDy3zAlu5hpl/oYRb3F6FzmnbZHW3Z4uUStkcinjrBPUbZs/
l1nSXgV9PIHPcsybpy0GYS8R7HGCxtUFVCdPSw6JnyuZpOdktApMZKIFc+fyfCARud4znStJmsMN
4/cvJ4TN9Q2yW7Oge7/inO1ugp7mHQMDazpoH87PX8ODw48Ay1CFmihohviXIYSUrMhMkskpyPjW
dUOY3QOyGwIdmhOZHDOPPRJ2BQYWtbwKbBoB9ORg3hy7DWR90w9dB4Am65PRPG/oQc7kdFleqvv9
5jfbIGiFYCViQYmhdzXNAcDVu96yprS+lcdgg9r8q/YygqhR/KUIiaC+pgaC7ivrlip2ygM+Kqju
NIlir+fOAoAYKgs+4xokp3hdNUBQeXdEjUCVJzjbtShfkAwy1xyH/DfXFkm/TDF0fgGOdnxmfpr/
t4f0cYYiupGr/HGI0bTkEzoqF/WZXi9iZ82F54wfyU6hEttCptGVxBJq10NOf8LE0OXzrFHesh1k
xjRF45KFBsROesUfk6X9Z8sq3sUYXTh3qOaFVR28piKDPsSmDupkSJZg4KK5v5uHlYF2Ipxa6ATB
MtM6qESlNf2W0gTsz4zmNF2h47oynsM6SRXbwqwKXeFQ71p/0LwGddSd4DSvvraYy6W5hXg+daSO
AqglAn/3B0+ED7w6Yyc5ug6LxrGB7ZscuiSeAfW+sVTUal/ib6rUAy2oE9Ts39yC7PNQuW2JxtEO
FMfvlvokNelHa9BB6oN0wUfkIAk+iM3q6vTfeCF3izrJnDXn7qqA1/3zz6GpiE9MEiZbdexjC+WK
DxOEdm1iT/y0npBxgYlkmM3bz9c3HZ55mbRz7ydjyQvRrZWhDC+7SQ+Z4qgTtpRzDYpygjAdlgli
KOv93eiODs+4nugmk+tgBpoOfRm2gnt6ughfMyO/EgA2gI2AtFfHY52o4ktQY2aiN8oSD2v6duyu
cnzdP9F3OXkUPwsmot+/d/uSHzIHoIegZ4t1N/NaI+mpOfNao6x6avAuOiXrNNHmC6ukj4y2PnjR
jPy68TQBWUxbzhDHur2GdWQ1FcnRVjlytcq0gDHzjqx32d/Ik5OPi4kWgUbIy+/K98Vo9op5AAAI
W2uW074SVCockcxhqWJmW+otfabMYFIIkC5WX0Lcg84iDJQyDRYnjpLDznP013dV32uFrrUZlFkR
TCCwOROGlgmZ3BHxAGb5tm6a4k5w35Uu5g5UMYWpKnY0otCJ3tORxVWwBDdyCj7mHzgDu+8244n8
9D5cA+trasAT1DyHswaHVM+oRDaDgVGdG5d86+vIqk67pYGifyqihGsEu7OpE0/CTODG0B7oQYDQ
JNv91ar7Pu3y7nVHTpqSN30xyhWPDih1gE214Cbc0hR0r7h4dn6dmle678YzAfyBDa05xGdJOW6C
sKSTVaMPkK71Drr8ZAIA51Br7KF4H21mMWybo5X8u+r7JJrwwaVFyVa49ktjsGG/gKxdGcqoa5yT
aQWCprFKzcXo/5cqId+iQXtNgcRgsZbjHk+63TlJoO6vJX3U/XgKv3blK7UWxc3+IqIzVH36GaUp
6mB4RbwAS7kjHUJHSCzbl2TO34VbvItKOJY5z9xZ63Lztut6bVqSfPkYKMAsujGlWfQSVmgoG2DF
qFpPu7fHnm/cW8MsSPqk/jaax6KUuOTuUcVySMaDn88mjLGmBOuUliEKsB1cx4bxU3PZjI2NfJSz
fGCsfPYG4MlRFVh2U3sEFp2FBEIWKXoLH/dHvMQVrBR+DaavMfHnqvBiu0F1v8VZyDxBh5zYlt1i
J5VXqsylnZUIbnef0yRFeOhElVF3zqNvb+NEN/04HfXgaJ4mZ5VMxacXs5hFwtI5tQPiR8khV8l0
jfppdPtu9A9mpPX8+cMGDfGdRSxGeHLQAzAKW+TPRzDx6qzAXL8gzBXlIfTJu3BRnJnpUA2LYqfw
KeNU91GMNK1bEamIas9OzEY+KkfeRhAvCGpynH+5od7Wtegx0+L6shefTIPs2BBth/2gpIluI+zK
KJjeMGK0VPxvlkQXfxjLIDa5EFp1jwZ33AgwSDzBf76YKoJubnAMy95UX8RTVoh4UBx8jwsCn8HY
z8bVsQrVMtrZbATjEvi/Ev+yAGYacCQYoqqHvToO23xjhCxJrKoOVn9dXEM7K9fwSGcvDRgpk+W8
84QT3F6VZA95QivxfiMfwbSLeOLwergxXZGHljtq+Q/iVmofShOZlKY6Gyckw5bvbX9tYdfjE+8G
PGU2S//8y32eDiv1bF+kY5sLfKr13ghFziE6IVVIgU+suKGQu6naZoBMkJl36QL7qlK8yqqApqEI
4OaUpmyeOZ8u4xbVACUyy5vUY6liHLR6AjRP9XVF5RwgcyQxAne6qwtQoIutidBQNWS2tEEpw+di
3IM8RoJbIVVX1l4iCM8Ls/BnJ1+IGO9WFe53hgPKa68Uujgg+okRN/i/QRL2jaAX6chUNBqlKmeK
4+1lCnDbxlWHbddDu8vo+VxQeK0xff/ZuC9nyAdqN6Bp0+FG/oDcEcb5420k64ARZkjmPCqryafG
XUS/n7WMVzDa4l2gQkmLAl2NEynwFAVyF65OYuyAx3/EdEEBRiaxQDAnHhrejla0rfca4Y8d8k4K
myY7Zudayzr+SkWAh6I8Ti1VJRHVGozUa+3Si6yXFjX+KXTR2UMFjw/sV68pGZ4JMGHr2oVXvg9S
kNU9SF0JJEOyZgnv1HWiilxmDzm4tGykhJp1i4Wiq7SJ48YJ+dhn+KpuxpHzTbcRFJWetu8d76BO
eHOm7ASdP6cU3KIGePUXZ4SsOofD/iyKNAJ9byH/UYfPUqdxBTdxmwpptEwwM/7mOuYFkCW2lsQM
PIlg5G++6TVf95NtABfzmZ+fXUYxuBfUVydMZzIkOq8bJVzEgvcbAURU1OopN68HCq7LZL28wjoN
BkGmfTuOcxUS9LiQg7G52F7fvGNEaUkSmLoFmeKJPeHcZ8bGt5Owu3GAVhYWkpW1JeK3GIQ7vG7e
EoN9P+HDPuy2xAT9jQG8Pq1IQZQeWxrSdHF17Imf8zyYOWSPKpxcm4eBO90BI3A0+iNAiKGVPMGN
fOTW7XNctU9bG6Owq6if+dF0MRnUfpt3Fr2bjeUGyRmUaR3FZ24zh82WIkSc7keVMa3MKU/3Wnkl
kv32mmaeqzWtplN2/kPs37CvgmjOITg5xa/jVRUtT2HXVGho9GETyktbuoCVoWqSCKwfA0jdvoM9
cQF5IEFaX5byVg9dWqKMe8UL+X2aB6jIpFjvwIfxkpx3Jp/6R9k6AKV/nVeTW+2JSG5rlYl0KB1i
v3uEFRzeuIBnbVcPxc9uazg6dFOwzPdyDz/7d7RGX+wF0+P5Nn/D0U5kiB8LaAiFZDxbHiLOjBr7
Qrmu9ByxGVwTuR04sU93my4mnlpvY7K2y4ImAuOrCuofiSpMh7W91J0Dul0gZdyA9YExoHbqvhVb
axZBjvQts/htmPGdP2dCRfYK36tgioutVNpEYXVJRDdrMbk15/aUKoj28hMPzwJ6pZwL5A5tLwqu
jY47P62v2zRfjSVfRL/SzVC+lgeWPbn59+vNJUyKcsqXSfrDKNWEVsgp6smf0CmoPNkPcgkNjscT
smtx49/gO3BBgIiXdb+NZSaRmcO0EH7Si1AWwnUJ5PPyWoW5q71gKzYcYL/iQ/vJT3Ov89QZ0V0S
n1Z676Hv6pfkAC7mUoZoQjyxcAnh16wLmeRXUnkRXAU16MjZZefpZwoi7JmKiCGMiqCyV8fhmIMV
3ZO89g8YFEsw+Ja0womMx4dfBW9r2yBTUuwkt+9ger+iWQRi1MRilLT3CCD28lmJ+KoA213ppmr+
FvfjjDIMrH6zNI9T45zAnaj2LrzOuHAZ1WSXk5F8W4njdF6x2vpT7E/Uskyovt9MMawy3ttaAh77
iHzy/VM1DT4DvAi0YAg9wxLdAycYXX4bxTvZ/uvi8OJ27cepABH3gvshok1KaPX35ExXmtyrA+Gi
MW0X350hZRAUbcEBLmEUKhZoTnIKuU1iM7O51LHo19zn8Fc0O0o3VM2H2vDJB/ZzwdWm/FAn9F3r
BIaa5j3utkOsKu4eXU2XdaiOfTePOfxOmXcaxPKyzIcF1RNrqR571zFxP9goRA1XhpdxfHXsPYsU
3DETgOsEXrE/d++LNIab+kS2bMm2ZJ3b9uSROtMyTj9VQB/9qDhjekhIR2eT3m5HdAVSVuxNyHx0
ffGEvc5hPzR2uPplR/A6Aqt6+VCQh1hVuCdHOEYkrhdJ2MGrTqtHYAQPv/EnAiwtnPAHO8OIRvyv
Zrb54j0wur4qeplqDvzeIqF1K8ad+Y4kVB+1U7XYG7J6OeQkcgFObRCPJ2/JyAmTMnbLcWhlNW+J
+5zO+h9sBMBRsLz71O/LIsBPhSmsA1dE9uJrngF/Vbc2KLF6ssWoHsiUcWaAO/PEduIon9Cd1SCC
34K4hf6L35FZ4HfiDSKWC/JbeVJFn58ln/woS/JVXkxvEX60Dx+RGh0dge1ux/QhzMP2bkat8RPW
sFuiPA5vdfyUhl0sdua+rhS+DrrKb9FCY25vb9thkrr3EniQC0c33CUOH1RnlCTD71AnOhBoUAG+
o7SvIHo82FccSdaaZFOOOHie4cHz1SM6iLAkJjI6Ax7u5hU0FXR3wsYxx34qeJooUdslGr9i/Tfb
0HKCb4swh+7QrQE6f61k5oCL34/IAA0anDbexYqFrCvyWfh52By5lljyAVpvcM3CE/qy6dNDwjky
9ZM2Ua56Va9YA6DPF9Fqad4tXJ1KCe81f1cqbihCGmuVF9yRNAgW/DsXtoL5EQJOTkj+Cf996SMz
zPAgW659U4IRJOF21+Jjg+S+j4Nv1nUNrgfN73vmZGbK0EK0Aez+CD3EdYqTLQkHuW2LmJ5PiTvT
BhMyhTd55DcR59b44nM6bPUOeen7xaJl6OKvDrEc6WNeFmuIA8g/xtSTweQxWewBOuxrmKO4jtlm
9//TIL1Z9i6O9zHV8D+N9qqSE+CVjYDMAAALgagspj6iTg0R7eeaDTg3y448BqWavpDQ88wfNisA
+xd3XWpFvEQz9c7fFZKhnBSWk9Mp241vRWDtTlO8QEhL89EgHcveGsjzSK0gWsOSj3RBb2qpaBv7
e6LCqsxBud97j3snq8VbelvsFfCyCeSOAYvFJzxhAfKEiGnlU/JMYJI1ROkyEvmknt+Zld/Ue+of
Gey2iQja3huDyPe5RTdx+1Rai9CEZcGAg5I0V6yA3u57Qgv/TueWT2C3HRO72Vj49Ucnq1mRMjwv
B48JFUBicjjlIuMn0FGIP6m4zibNW0k+BeXs9iEaRC9jDivaWGrx4ZHhKzBmyPGIv4d2WR0ne2N8
OB29ZPI3EJw071xDqKm3KTAKlkI87i9STDhUMUDNcO8WdT/dqHq9leSu9x8L8Uzd8Hoxct9hwgVe
I2Gh5srAk0XbWcnVFYTRd8J8QQiRkyFudVpNI+NuTmvQ1Ny7DxOGHnvdXyiXBNZ9VUnzYb4EMntV
Vv67Kq9rkdywHBvw0cdzb1exPiwHErd6evHGi3gwHgi7O9rLCWWt75kEnS4gwSjhr/rJooul6WLx
6i/7bm8Hf0fxQHZSOXZkY9wiaA4sFTyA7vlgOuWbisqxXOJh39C5GhhDu1Zg25VaUmKVEtkrw9AV
p9/sHGMvbgv8PccXduKk7Oo2F4SwBYZCpxzPZNWE9/xYTXbUlfE2gXgxzo94JJOjDcDvu94yM4AF
STMlEnBXma0Omj2K6D79ub7fPbDFPiiFX+ZeBlxKkszLwXUVhhzk9wOIrhJn+0zcVV+Hqg5YcH59
vg6bljHsuCELppQVIsijLndXjh8hKM/wwYW4vXgv/Bh1Xnk8DX/NNhzj4YJp1E9hWJIaa7V5RVDz
gqAVu7EgxLfRnd2UY0quMF9Ds7wnMIohBJ0m7SKcMo5S/vpn8cLSiSxtkR830asuwbFuNTBWqXxK
7BPI/SYFjAIfuPoTH9qIfcnd0hBZUqJ487iLQOCRgxKZ7RNFPNOcqZafBxMH5brAobIM34o3bEDk
l36ceE1GK9k11DEVDTtDMIo9HrQ06bhACi8kNFsdnqtW/iG1Wnan9SgtQb3ub+zNqTIaUdRuEXWV
P6BVqwWnnEZyhhoVWG7cIuyay4ghBul0cHBy8IIm/1ikYEqntx0qvp3iX/0u9HXArx1O2gikGn9c
+wkaYNIc2VOmYfXI6tnzrdXIevGQ6Isu8EYpletRPCwWVnfihJ9+2llXgkfLINIFCoUSZrtp941T
Cd20gZnO0da5VoQkCY7BAkrCw9Y1lZcK3sipHLD716C49S8gqgBanF854k3a2vk7NlgRMk4hb9+9
pWF+8mNoDd5VSiCU4pAn/konGGNqFrFWEWq/SGJGwYVmekVzG9iUfr7bsBsa0gz0bp1ORdzUmY04
P4xbL45lRYLvSkacOAzlHFnIBnJHH8GaoH9jUSyKdIaaSFRuSBosFmlNZyp/Djunrp9GvQdk8rPk
4T0Clf+n+4xBZeN2dG/1ax0c2Ql1QKNkx09DLSMmimmfk2ca+/wCwm/ATL7HwCN2tT2lxK9bW9H5
kwcVGAQyiyunfwwm0GrycNpNRaRFJ3eRljvrCg/Jl6h9Otu+y06iJcPCujpTD1l3D2YEsoOa87Df
PQCGNTrNwhVdWCzn1uixRG6PCSf9OWCuW1ZwDvvwCRV+rhoDB3yhFRhtgja5XZfr5Kz8fa8+YyST
wTTASUhBgvjhX6bhfyRtEt1PBgu/nq4qsF2aMvcm5U1PAdagWYyhjh05HT2HXtAB/6YmOmUEsFc0
XaWAmOkXmxwrdb+5hgglTpLBpGc5Scg0+JeiIwlJLwvtBV2yeUqUeDCUsEgKyga6qxpDOuCPo93H
4U9mqXRD3oAbeHSO4bqk2frbzeb/a21rG3hsMw2z0CeWH1TOCUpFu5faO43wfj5KCZtW8KqIgFa2
6AUtcJzjjPeMYrwuXvbs7rmQgyp8jnXKnw06Z21vb02ybrsOYFaLktXv8G06+yN8e8opsNHqkjUI
b5IZffNwg2nNf1wy8Jbvhq2Wl523dKZSpVDPWe9qdAZUoMJ6yq6tWYZXoR4nNbardUm/mN5gsGI2
t9rCnIdmUAOiq94H+dAYNhUOJyNz95d8ygbvo4WLCTIkyx6levMATkPlUdv9PZhTMDB+WyIyGLwE
3rbroWM2n3x1++kiLYWv28EY++dV9oXCps2FNvCGnDZBYLHkORiprj3FWHQQgvm267cRYXLdssHO
O7ZXx78TZA3FUBVx4qKHGf9ivaxn6t/04k4r+wKkFEbqfKFJm7/ltUfs3YkXFkyGWbzoGHJ4k/8a
MmGI5kP87HNYj5+QNRhPfNAMAzyiWlV7VaCd3KktIEKg09aVN2cEvCxr33x60i7hn67wrYcURpV+
HFcwG0O8t8+b4LO4eSkaKG7eqMamsi0F35yGiPgVsR/1/KNuAhyO/uPUSJVtrltgfB8JFNorC0rf
hxIwJShnEoeo3W5IZ2QunRwuskugOAYKyLet5aNyQ8qA4xr7Z3LjE3zLEwCfSly+DQr7kGhHrc73
IAQeg3w7OwyPy/YDJC+r0H9mYzEKKPJAtMV/O3YEp2xkUN4Zpbwkx6OdhueXfsF0BTQnNeP/v35s
l8bdLpRVyCueoGMgokuRQ16OEj52o/rkUWoqgnYoV/0QgsqOxDt2GQYfUBf+HM0EsheH01sdDvxp
L789H6LRitL2LnkRAlBk+hfLUGi5SBD07JHMJEP/p1eJsYQp4YSh18QvHe1Uy3K0tfdOkp5aHNKd
4ITTcgFks8BewWUNeDqEV/UZR38hU6eYTZfOkvVWJokWRGJxsfJkYwwetCgupHDEjUngjP0eV3XW
TUYofFQPx1Lcss3rHNK5HOvNtfQzHfxdC4SWyDGTWXdcCuUTRqyhPIDjrAif/gzaYbT8TdAolRxD
4w74VcTam6Oo/3A7Kq6xocd4tK6E+qG07UMNCyp9DE1LVjsPd4eS4dSzL8VmQP8BByi8BwPsTRQG
DAHNd+EJ+tILBI59jpd2I5izzKJjIGJlWmEGeRW6qTt7+CS8u4BjYOMaUccKd9VtoknxE2sd9oiZ
GuJ6CvmtU5AJHSeiCKRTZ+jMesjYBoN9h63pmlWry9vOcPcq0C7fhPKoDRqujzSBoSbBNnIlrToL
XQd1XTg8eqLdu/gdweiaUuB0eOJlvcrjiH5/qRwP7f2dhwfKi5KSwCTdC+olpLGcyROnWkULx+SU
YvCnJ4cGYvAMxpmCZOzguHn2nw8s66kVbKEicceLQBt0ms+z09bzfDroAFGAjBPIMxI6gAUS2gC3
LGoZX07+WZigacXNK8og20K9R3QPjeH1P5xwKDyjsGPhtLdn5zldOnLkQkj+JrMnDrg8lp0NFWow
g3WUgNJ+1Ua8lp6BxlzAgzg8XE3SaSNb2DrvhcIm7S/mQL162JCw3hp3zJ/G8P8FKEcLTDamALPk
CJMgIdYOYrcvNJsSmhNKtrvy9/4GudVvo7eVdzNEa1NJCBVVTRtViRZ1F2aOZV5a1gXN4CKpoUpN
D9H73tjC2BRkCt7BPbc+kaqwlcee01W/TGFJiSvQioZF6EEY/KcOqv7fsAWTu9TkOYZ1bmctcAe+
yb9VRISPbWczkgloJMtctcWwOcAWp6OmJXVU50Z9ifmiKRK8KMI8LE10VgE9zjs4LM42jpYM9V2j
E8qmOScxzlRjITeN2fpiit9hmXodvIMbbC/Z8V88fJv7GAjrLs/otIkPigtfbTFJgSrrZC9bpF9C
KhWUcXMDSjXC+Db+Y7aupp6W4ooa1Lj7hUdixWu4wFNehIpkbgLMqvJWMKGIKfZxbpiTGhq4Q+5O
ucJUykRXBZVFMGzCyurU2rc0xzL/LlnIp/InnKTZbrT73LnwCAIoC1pxdXijxFNAMkbTxOS/7KAj
fRO1DY8Jc5UxQnbQ9qQZwWoMlw5R2QSUyq4bZi7X4mhYXMT88HljDdg4NjYxQo9SfWwY/Jy08htw
JUDVmYQz1cOFLSPsoe0HzfN3VtyrAlhYtg7yBF5RdBDu+D7/lo57j+HLODKTy/YKOLv8EQW4RehP
BwMwD7xITWWr31gxxX1QyU43B6UapEmrdt+YO0ZEhAoBIO44xjSfLkY3zCrIHEW92oYqIRUyt8XH
vEQbsRanXrhaGHct8fCBGjL4zAq5e6TL9ZbFQ3THnRYh9bYQEv+uy9YvfdXQYV+9JP/Z/w+e2Mt5
zJVHD/3DwzCxmjheXY3/deQcy3lkBFNNBeHVjJinP1augdTWsUG9zdzjlFk+c9agzEgGey6yh1bK
EvVDEwxZkR4imbfghf9eo9MTxRdgGNOZ3nmsR867nbWWY7hMyOvmDlMdfWmutos8fbC7xPv7l/NM
dSKzMANYieRlm0L6zDJrDq9iElE+54tZpfGS8vceuw6rPY6gO3287L8fn9+aLXtlHcq+dvlYyuOt
fg232AmRsu2691AF3/dVrUfvMiiEjWhbChsFka6KzyblV69pEcgYLXXOJOD1NRoeTOisfVZYIVai
bLyuNQOndxotF2tc04bE4UYUczT7+9h8k/Lxqxqli6mC8W15gLm8ZgBcN4InSusl90PsZmD5PK+C
KBb86+7FAE1ggpu2hn/sadMtfLi1UczjYMkJ4bDrNNFzVIEhuodpTY4xKk0Aoibkyhw6H8E+6Qzk
Udg+3sp2BBtQ4Z1eMVP9TF8hwDnQf01jBMTpUQ5/zCx5E6mgb0cDtIwpG8XvCFUAGkKZH/pMcHqd
0zFKVfNYcgaYfvaDoGq2zZ+nonJcsmOkIEK6moselVYcFHtWcuTeMdyEtOspRGZCpRivahV6M4Pu
5TyPfU0s+viIPuMbBfYB4Pt92BpYWcK37ZeDEcYBvjy85KnOvX2gqfXT9DypELi16gP7AUasVlNp
E360/prEO1RGz/zfcK7gDUlZFwC/FEFx+QJzT/0RIXHUb+dT21AJ6ZFRruz1bsfwYx0Q51cAfddQ
Tha2Wtb8hnYWiH+qalVbUviFJgmHBAZuHR8FttghCn6umylArss56THqA+6bDVg9WDddCfWxiq8L
cx4AABIYcHe4trhEqqSvtkCp1XUnljHymP4OcPtnBsD7H+Kpxd7ExeQnM/yhalmwLq1TjPFvuCIj
BAa+ayhfnLbOQxf+N7L1VTp8SdigO40S4jjVUyNB+WFfp8QGcDmUW/fXbE9sXsyyf/7hDOEe7jv+
+lQ2Fcur+D/Mgsld8qoJt3plTweYuIBOwu+6raKdDO2T+i0Cnr2Kk7o22n/+hKwnS5ybhleI0H0u
xSzog6rnOobVtl4OxtlCQFwfTpcTAwyIzTvHfaoaI/9nH1gZ0gtsidjhfVcN/jhXvjhYjNwC05PQ
6y/ZOjRTM7r/0DlKi9Ws8aDVroqs35TbqyBi2IODhapR3K8OQcKXoEpU7RDKfCAO+bduPNqLMoZw
SVG87+6b2y3PNgmUWgSnIQ+muspzzcy/23hovQ2ZRkaufOgYffSCb/rKzwl8AvmhylOMjbACE5N9
RXiwmtf71+SU8Xndu9JZ0KrylB2F56MpdhOYqwKX+lnIXIgwrYSdMDB2i1BtyvEYcygT9tq5/d9z
FwlCTNSKsTawba/11G0NN4nxwymjc41shuXeY5pYn98ittgQnzjM71ZgoXh7POGuJJSeK0KFsLpZ
7h05HaCbm4urOZTlZqI/h9ddxnd0K867OBrcxK41J7oEu9hAvJoWST7Peg4HuPFXkViKdFTceq30
orifnVYDy2gyXmWZyGlpEa1QeoyRktxXittu7gVBIpK3BHG4wFOXtRpClm2CiQkGHZfrln1Y/cto
EaeY3i/8hsST4K7cFmVSYfSF2A02gukT/jyaYKjMEWsRddVWDDQEC8xU7TbwZVgTavLkGDZEqhgI
nRF7U8w+/+0t076hdPtokY8rg0ZSGAieI1U2sKf16iaCA4p3MKWZ3kAfukq8jEfrWaQZLS4rnl6D
SC8f2FtDaAQ91bgEaowlb4YwiwCSBWYar+1XCuOiYvapfXyYA6CMReBAwUl0qN5WZqUUUIXdmylH
pVnl433QcFziIlY0zn+5rFLu7scQ3ZiBrdVkcA+fIMqUst4A0HE/8jMTlsSLT0i4B6DtGyKXVId6
xzyODf3Ipw9Sj7P8PbbuZkR/JtgZw1Mq+z9TlWTX+YcovUcX0cKCMW86YFprrJpPaFwpvpBYcNvJ
YpfWMYsujdKoIqA/gyAzfe4dDZiKIUDsVWEXw5FWgt7RIMtDQTYxVvzWpczSeb1YZKqgC8ryinPW
P2CPhbNMTU2p6YpLivjmoQ6wdcaEPhZimCEJnvg0b3YoMNXoBtGXx6V7Zvso38AE/ndqMXhFHD9k
g7+B0h/WhRuZ4qRVcBi0YM19uJEvz0zCaebaypQIKQ1fCCduownZGjthZRRhedxcip7HzHgMhuWH
ThXYZrR/XxA65GW4QdYGIR/s7wHQSA3bVc3PsA6aEXkoEr9lku2s9HK34gj7L1VKrRfezu6qXgWJ
70UyC2p+7nbuhtVDhIpawZRySWoB9DxaWsKSktDaPLHn0bvqz6BvGlOkST7rSbDVXKqAT1x6DQix
eOTYgwOEYshBmFKs/7G4fK0hc7BkOImWGkcHZIPz5Di4SHl/k/qnBbJ9XUcqEi+E5Rx5tb+vwXEb
4te9QLVTbWw+zV95XQFIaw4nGKy8zGaYnjeiTWW0HPC4ngywg9p7CrVZ69pBUQEBAxVogxfcTSIB
G2GvgnULzBRxYGEvXRnV8VB0kzR2pcyHCTaneFVfVLCtvvayZ6E2z4PCObWEuJKnTDlt/DWUMbbH
WVnYLHdh0vS5UAA35Lc5gxY7JtYZTI6HBZahGX9cHFCun+wd8QTancfc+2X/Hc9QXSXns/sO31FB
BcWYiwwq0gGzSIiDuhWZyNVZus8l266QHGy/yjDcYRSf+1H4sMBZvIiCX59Cba1Vs+HD8zlMI9ty
W6qIxHvrp0YmObQnMJXX8TNn+bEYAHqgS64KIqvC/PYXQxuknahAdQ9Zz4R4scildUR/1a5uDo9+
Q+xohB6WnWhmGNNrKxhtSRGHXeNFw9IC6KGrNvOBkk45EW3v2VACzU8ixGaBrmTu9aFRwi5FH2Op
byFjOBBow77+FnM3KsxxXRmDeiN+/Xmt4bC8yVYsA1eqhSlXUjctY/8eDj2dq6GxYBeJziKFJwJG
0PgWpiehRBrl1A6SBpMiRBQkOkHQ2fd8w8QJeMBWzFnJAZHAYG6iWC899gcmuDQF7iMBOY2oz7CX
Czu6S6SWDjWCcP9xLu41PQ/Gs0DGJF2hPifrzXf4jDzxKeQtCICcvK3rHsZhzVs8Yaquew9CfvPH
TcVeJg7Kdbn85q8wUJcYMNo9M9OFH9oTA1BY+yDStWSa7Ou8uSXOseWxlqegghz2brswwgjSphDr
3NaTQdVtl1dluB3+9FSRe5uAggdN7ShS0wmYm2xOCv9yNnNKH4tYNiDgik3DedqJppSdfldKFoSW
SiOvyPzh1B6kYUhuSu/EDgduEutG4nGjab6xru7VQ/P+HKqfCr1wBca9Q8cTD6R1XHhG1tg+RdbI
9ntnvhDXUetGlTNL1s+4CJLFPJJXig/fZ1BC2vOK6YJd5zTIPXFUIXmAqmeAm/32tAHmCZoCS1uv
b3aXFhS1eyhU75TMtZHLPx3R6cZnd3rWXrIogZe7evHqQRb8iyPNgOyEjdHH2cwN/Z4cPR0Ribs3
wIftDWrwxasjdQLfCrbs8cYQsfsCHsyYLLmOTOqxK5t9jvPNAoD/83k1T3LeLXoe7nf1+lPGc5h0
zwA03fLzrBhzuJedw7PmkZwGE+O2AfcoW6L+eeAEVkr1yp7hbuuS8BVGLm3PfTKg6R7zEFB8FghZ
jjpxDEM5jw46KxjXHAJfgTHkxNK4aCRx1nBJdmzy9x1yVtW1ukWesSudC4F6PuZDj34ZwycbI6yC
uncaPNq6Z7Uz70CV+LGzr7ItNaddq8yI8Uc6xGO2THryfw94WW4qTUOFLH2V0wBYx5P90ieHGemq
dy7eB/wn6YAplGNUpXNelf9PdhEBnSg0mZ3j4Yg+3bKtW/tatLJKGrkcdlEZDw+V7Ug1EvP5XD2f
VwFylr+41E0cQiKERPIc/wjr/naHYxINYYe7acr9hJlGFG1ZQNuEXQ+CkukxTGMOMoPV64FejQZ0
Tt8a23el0TPb8keZ1hvhAgWMPmRsNefPE+Hm7ivMrE9n9C/kX0WVrDg3e4Kj3Bucmz+WkEE8MbRP
045bLSfrV1jk+8RygQ9x/s0sGVptmDCMDzUspjbAYKnGAjaWZUUXYf6oFcKX1K4qmFpbu/lAFkoO
4QxC4tjxyiIIn/qqA0sRtuP66V/NLustjBzuj2BYJo4irv+lAktvmmcyS3Ta655m85fRr72HOaFh
pDgaI3jhr396lRJGoyT3DLSMYJfaF7DDGd0qw5kCcFwDLS7XSV/6Us4y0hvYOInr6r1lW2v8PGbQ
DnqzgWimvOWznDlzxXBDP/n3DeBRW8Am75DKOfWzDpYhaaxuZB7p510I2Y7xOaAgSrj85GSuEL62
w2C6M9oIyFKBLCKt5/g0aUTw5iSNQwSj6RzztPsOb9/IYHvItvEJvKuSFWoaM8ooc652mcOa52eQ
T3XiMCn2BLtD3MQX36CjnAoLsRLUdjJtiwcraEMh3jdR85VoOBbnZisFVzN1WbLwlpl2WTHcUFph
cjWo/ptvnRcoa8wFXASwBlA3ePBftQ7TUZU3CaosYiJMvsqDYCWVUqO7De9cxEWCH2m6BtfUM6vQ
+4IC/QdVJN5LMWBrMn6KodKrN8n8NMGi7dwjIi/RL9D62DCZOMvJAhHlQ/0COAMctindSZHAinSa
mcaZuwc8evTpK9eqLk8zaq7wFcr8G/EtlKgGRKccB0kxSznqHKE1AJ+I0S0jucYx+AlQyK3S4gGc
OHGqA3u4z2gro2A5W7uEVjg2ZMcxJY1v3MkTq/1GrWal4z+Iob9WrOa9fXefURSwg2XszGma1FP2
wv8/WCjj0LJ96eooKXZU/aXsj/dFh7K2Q08B9+98HxQbQ5fz3Zyrm3FoHMHXL4a7rSUJuH35eFl3
LeRjdZioZqshv8XwRHSOShSzpXBnlYQF0RDyf3hUIpszd0hL71orRgrEWNn8j/W3bo1UrTYa3ROT
VAw73o2drACMHETkihnACT/SAcv6E7xM5xmzYEUlfK/MR7FvnQN+/9CJR/nOhUYuLbqY5UMxILUz
ZgBao4hXaZcCTlPEAb+IgKWeW/X5k2D49DPziIm5+qXdpPwDniJPjV8W5hXctV0SSJ0xZViBnSw8
lYIBP4wrzgCDw2f7mYESlmPI/MkM+EaFJUL5g57Ya9pYG54JIOPvKlmiyZ9vh1W9zGPoiP/JmIku
KzMsfFdLpfBgs6bK00LyNoTxBxJxxYM/p5htef3gu+uDHiyz8l0jPQVYZ19Q8rnAVcVODU3O3aJA
pC9+h4GbdygiMCo9rfd+/dePm5Aigc9pZBDIOsXkivNnLmoD+40LmLyCAjObRVxkFd3WB+gbU9E0
tNGo3DGctLfb4Wdpu7OJgz3I7h8lz1W8emwRaC20h3b4muNQqXvyClGgTNQWUvymNCtWKXyKmrTu
DeibrRMbOFlg+qnp6KAjCLdDfafHJVuw75893tkO6DccN0m6xU2FPxYl6YCWHnZgdfVpGf46mK+4
wMpdz23tF2jIrQv0Hs4mlbWh44c2Tr9snulqjdf3r7ISo+vnlvR0yB6ZkSZlS8XT3XZF7Fa3L2Na
wBEc5s8QOLM5+vSTn7Vl6Tsfi4y19wGDGyRYputcJoMgTiYav16qadDsTv/2Vf5XJ6Z3HdzfCBHc
jHUsSWHi4MfedrX7YiNbxAM52fxNKh8foURJXM+4rCmcSy5jTLeXYJ+PMcbwN/6j/zCPilkTubtn
jJujWJZ2W4uLG25qS8LJbD8fXpaSrBB++sTwxaSAGGc18CsLZoxoMEFYCDiUMXwUmCbklzvRa2N/
R+4nW1pCY57jjXqNq18xhFcpTf3GLNzRjnEbE1hkuYY5VmJHCC3+0JcGNN6fgUEjTFVuP7C6MTgH
BLfVh+s4/xSNdQCm8BjpSM6bzJPc+d5hnOIi2Z9ym7+FVvc5yCQB6s/lcj9goJVbHSjfjvpkxUDE
fbPS0vUJ+9mRLYwczSjjrTxExNjkjcA/K2FRUlsh5lji2VsyZstXjyjW+2mjGoDNkmgOrXQKUq7s
Eb1VTMaqa1rv79rE3j15nL/xULfduyYkkOW491N8RFyjRGOVCE2krvN0eGbk+2mleuaFIcjc7Aet
3x6hHV+Vxrrj1ZB2i/cZQWEq+yrGvFQ4Wsv6JfxeAXypv2hhq6wzVbqyxxn6XrEd3FDHrrFoQdbf
yDKBV2VAhyDEr5DhxyXVFMRIu1ma6vSD4Uw+0igCyukQzpkcbznc7AnhNZfXMXG20VQyblRy5AjF
f9jWk1cVo4fVjhcclXWYsFLINBYB7h4RSUy7GC7a0zJ2VqSTyppnshFN29baFJI23iMhIDMjL4WZ
gHoUQ/KSJAQtEjHis3uxOxiZ/lrfHJ7/Af6WDxeTzcjKsM7E1FaPKT4/ZhlgybKRmBkdfiT23aJB
Fdk3y+yXZEV/jYa76sMfZeQcxWKX+b4GJmFQk628zV6Bw4nu1Hxy/VbfWF2XNQev0QvnXurLDIyS
qw9EKsZdFsRjL7Abir8LnKds4DMP62HeRO8Sltu8diMb8R/0Dn8iKNBMhq0+09ayboqN7TItwp6V
RGiZ8ZbsC62owI0PoG36FOH3bk7oceYl6qUFTRdUEYeYrxHAnDtRYfgJi4gaHZDkZC6YpKxrRz19
vlsJZT6XgOXU1zzrRpa78SmuoO4f/tXbe4jluF0/iPqeE9FZpIsmD4hXQ1JXZnhUKzWn3R6fal99
gresxNKaocjsV2FNLasLrN/M1A3mISqbrFdWpODM1mlL6COgMo+EvTkU30x7CBzbV9QRFJbs917e
+TH3zTRxaeEeJF7HkFj4/f+8xUK13SW2sPZXrqlJT7T91oYKPEApkqEyoj5VbFRqLFZBVd/IRtwS
MFfRPUIwt5B3Q1sw20HBDAfbtktBi4i9W5mZ7IMmuvg0OvOEAWL0ytic0AtBrrTPWvhn0jP6lrnj
wfR/iND5RePhqmTkXFYv7dl1ir+qEXe8BRYYxhBnwOHJNKPFhwzKbynnL5w9ZK2ZxxwVVs2iaL1E
cDmoOdxP7DEkhuQp4mU+i91gH2Hnj3ZxN8npEbTvdd79UYcvICHqZwtllUf3+t8y1Q01a/UI/gRm
OwcjTIHBlD+WryEeiKIDoR3IAr6c8JD9t0HILRDp2tMTK9kmds3QNEYVBZ9izmgjdoqjmQsH78wp
e1FFOt8uOTcQj078JJ9vmu8Nxp8m3lHdQ5cWj7JURa8cAyILm9w6gxeaoOibJfTaKWqN9fyZz/wm
ZGqBd+adwUjYW7zZl2gCm/yzydnOEVb6bTvZWNNOz1gk7YSkjgvLWQAUufc4/hrnLFtuchzGrdal
i5jagwThgalOSrGJnZbJybs+joxF1iHc0G5G81uQzu9aN+fpAeu7PqEAJeNv4yxmfoE3JpjrBEnK
q6zqABh0JZRH6vBTPFPNyC7wbZqhg32fOp/7GmMjQHBL66rUtsm9QUS54DIlsPNBzsUwmpyB+dbe
pbnTpWEH9s2jnANjMbrx8VFjvcAAFjLpu7f+li2iNwFBkfm4KWKoDHG2R4iSSE6MFpmKfWDFoHM9
4OmPNe+swXkDp6i5gbwxbwKUEEM1s5uqyKEJT5vf8Hsd9xI1E9dOpWTyEsXVSG2g2PW0LVurM4td
7fR9tO6uj4//7gHl3glpq/ombWIyRYQu6IGKG7MIFQjZOV18W7g5MSD4H3JmbfvHdA/R5MOjDOkh
+LbIB1dgzSQbNL5dAxfT4n92o7zYWebozTOm4RzhzJQR4WUuHHJTm9VBch+DA73JZz6mgSV8CLuh
H+FZLWT3EvOMJ64njHPREhIo5tVYIcScYAz8ukfvPlhYrurN6BVk4NLboHJORUIQRPTKFUtm0Rbk
gkL/qIMH9VnxYVb1Y54c90+HrB9zjcH8Dvqge2Ji6V9k2QHmwnt5QyV0aBlZqzyrsFekp6NsswmH
M82+8GJzmzLER94/DqjQPHaBqIFHvCwHC4B6GpOKFhsDkOACLc+TiMy0sc1z9+iKKiCVyU9Oc8MJ
I3SUEvcbooXRpXOVn4yBX5RHBU/26do2nv2e4SzajSRqZKjaLOk3EyVm+C8Px8cqxoMXRR7FV3aU
SRe80zsivQRwASWcZjuZ1Qss2ORyWFggAoXgSPx8s7O+tF3mMU8rnj7O5O2ZktroBYX+2B5KlvLk
dccXiWciyB4dThcZvcFwhuQTsljEyfMjV6j6GelJPdtK2DvZwOJzBaC57AC2tEe0Q74FI61sSXj8
kuKqI3Ic8LoabAI5T76jyMFOURLQ1aOJKGym48MUH0Sd2f5P6JdpQ68dSRvXxYhrRDKPmuv8dPoM
aWnEJ0jRG1yW4MenxaZQCPmueiVyf7fpENWQmC9LlOH6Lk565QfzbC4T6XN5dbgSJNuU6bfEz1JU
Zlqayn2WKPeokY4rj3jDVAOZwIuKtpt6hIQnqNcqlLC6bp8yZEtSevQCx1CckOcnM3LXcJxXNfGD
1pAvZrfkJGVQmMmsAHYjFryqR7M31Edgsn7ZLx3JyVbct2yPWdeRY7fh1ncKLbxi1Vm6Mm/teU2D
QROYlJO3aUVc1xLppX5z/PTIBweReLYob6ESW6o4pwAEuy6dZWmWoazhUzwCa46pHnKEQo0UWlKZ
w55mA60/PVruOL9wV6qGfw1BYecrvMq5sfxW4/Sbeq2FikZ2bsHNP7U6GvK/nuyILxtwyeDOIcu8
xQKM8qNPkH5VJ560NPyhxByTEMWo3LEAIqsrsvVhJurhovURbeAPNT4qK96P852IUI18Ox3DE6/2
En+c61TqcrmYdzNvwfTNnf0cBfkVBqWje8BvazYHMFvtLW6WCDw/jb+0Sksp0cq/3Y5754ZuG/3N
0uq7XmKFoWZedtqeOupi8Rfn+GbQMK+Owzvv8xiNoqUcHCQCclPEQzzyxvx3PFbcs0XeMzqKu6lT
z33cQ6Lbf57fqUvyHOEe6jiYzN+acyF+AXRtrkqn4MCZYajnEka0ZZbzE7DyDTp7J9z2x1BB709g
uQgqrS3Yyn7BxgVoC4VncFEGkFCJZpLYu19ctGY6AdOeykh900NG8ZmtMv2NzMkViwkSt/3AxaLL
Tn0fN7uUXuUuu7rwZlaa3j72St6tHzGyZJ319PqbfyH+vP5Eg4KDQEnwEULQahxcO5BVa20eIDbh
KWcZm/wHeDa/q3MAlye5Q7fJnA6823xf5HWHcdau2dBMvwmqC0UqCwd04y3jfrzYmWbg08Iw3Upy
ppA8Br7bi8la/2ZLLPqZroQU9FqeDMBfJ5VNyBiY24G07ixdQNPK1GV4fRydj65/DOZ7ig0xCWJU
8kbdHc+pPKbhTCnQDOcXUIbomY8kksYK4Lv0SrV+eLf1soctpeG1B6rEj5L+S6m2RDAoAkvORgsY
Opb7pZXzFHiz02pVCF+HU49n6QuQWpia6xkprT09CAHiob2nT5mj9m/uMKiJa3ozqRk4/ABvYNaN
fJYmrVZcw272PPjFoHXI47svxvsAUvyQbf3+tVWZvoxSN5Xe2JF0Njtbq3kf3erpnjZWGeqKIfhb
/rBrBbu1TnZBFroWIPPu3zEmQBMVl5eTMb/Pjd9lo9KHiElOwgQ9T+RcuFWGpsxSLNGQH6p1GLax
GYCFdtksIRDhA4fn0n0btZ5cHpanWzLQ6hb27h6dJeMck6Qcgp7LolokJF+iMPgW5ZxOsXb55YKs
sVc6vLN1Ccj2p0rJClQUUj8vA/7yHzaKNow//F3nprii+fkFGzYWCX26llsA5A16j90cwP2UeIU5
r78Ivd7YElhG6svdjitGc0jeo5xpcAsBNSJIQei+ARYRDRYQI4ryGM0DNnu4OXtQsPMx8vkoiIY4
TQ99IW1GD5VjS2P/ueHwMCdpIPrw4HUmVTFyNMwO6y55SPaLvLttmb/+Ndhmk0nbWj4Zwwp1DD51
RLBOCX9rfgxyF6eBgtW/RzXQSO89Sm77OoVonHE3YUPJaj/sHe/j510SVoMW/+uZR6fb69XYLIHo
puU9hIORdvDn8AeWUHAeAz092FLTnqUcO/UwPqmrPCjZcGQRuwB0vNWl5ghDf6cXElfDi/dmTQ5A
5zALxbWgfKVKcDQx7Q25OCvSPtyvLFg5hiQMHAC8Muqn11SUIvmHm6Tg/Xqoy4cXKIig8bJyZdVg
lYpgcoDlV3Rm0M4/wUiNgMQyXVWCUvT5uIraFKUW18nw8y+6bguPOIPr1YTnmYx2Pf5wHj46pUtc
MRvvVhkgeqIoaruHw0ycue39ZWM37i9zqGIqxw4rJVkwM3aFYsTm6HG/X6MxODlszRChPOTIZnPS
nNWEe49gcbWdsapMH76ctng5m15Aulto2pVZ80M2eQCwBp7DGoD3JVclUStjdgF4eyWfulxYx1Q4
oP/ehECr8LqXqeMzcdPiBNSayPWET0dPy5lTjy23Yj2KRn5jmDu/+fgnrzaJIdPYVSaCiOxoSB6U
Wx8wcB9bP3Ts1BADlCVzWNq0gjgFNMkbq6Xf4qnPospkI/P45OPURzYCZryiTk19sZ00dhtQLPLB
WN+POavqtxWS6ZwO1Zy8b3G3EC2sSN3lsEI90Fw+OaoYEqYTF0HMGhEjltcbspKiE6zZpbohr/Rc
fcQEgSf3jXes+mMetOljgIT/JeaKrkraQrIPkEztruqjybvzBqXnBpfWb72i0+zAj2j9a21Ozc1L
PzGda3+lP/QYl0wNCMKsOQpFkfofaIzB/vxVXGox7ewHTs/CK7gzk1W/DTxZRWZWsNPprsBDwyCR
F2u+m87T1k4pkvKzZOjZh9MlhftgEsjtCGPNQqkWbamqz5SH01Mk4bBKVJA41rOtAgXUbvsL4wMD
o2jPPakyVcr6jUyv6PPew/70lirkjZ2HXwMLw6LbVjZLdzNyos5fGwP3MV3yw+q0QROoSJmVt6RL
Q42aabxnUwDDCqWJ8HUZQ11q6Ya+w0EEhQ2fPb+gJyEc9UG4voNGVzBYea47oAvJ8lRTb6xW0agx
KG0tcKUAzbv8bgHim/nadxNjY8HmdPTz293ROJijC1r3TVTi/jWxTBmSO0ch2nGq+L/2CkplkSPO
ldFvvNEi1gjmq9xLTwtjJobObcDobMEqewJ64oKcuZRAoa8qu4vnFm34ozm/CNuSoq+WDeIQkULq
V9DSYrOKN+zINZN/HybLyO7QIFm6ZnLGfhWxkZFHBzVEBxADc5fhQkuVMUBpSXFMPF0GEQ56TfpC
wxZo7pbnHyP4M9wmryiSeLn1xL8/gLh6eAYqPuPZnrN3CmaoD+NP1XjvzWX9yt3QTUUZ6rSBj28x
wUvvbBWer4OCWBK+j153/6dWny98Eng/U1qe1kZirOesuZRifwxF9a85Bz6+mjwwK+SXxstq3eZO
J0r8Y44fHqGTa/lAokxisubrAIEJJOFb1ILIWngzbmaWh/bbkTDN3h8t8jQyJ32EafLiDcvm44pC
AbKxmYj/u99K4/vwE2Ay1ZBwZ5ufRC0oG2HQBa/6qxpHKXr71dlluQhZd4/LwJ4efWXYY7VT1j29
3j+D8HVGhKinT3vunOyMteVKOEGQSl8IAgS/LYvdHB5XHG+8O0MJU5EZGk2/i6qS8sN6wV3+U7b6
jV8JZcaJlw1in3JInVgzI3DUleprDTqNBFHIxa7WolOVkjQ9Wj4p1tPaRtBCgDh/m1iIwbp7Cuaq
ACQZfUHx10xVFiz7D6xWJX5jEzu09oJCnecWcGyTpqHmWEORi2O3NRZpfQVwsJlTQSOiuSys6eQL
t6VUgYKAIjrjhQTn8tNFT5gte8hviQlMO7VFQ6uS5e7brgRj9imGnBH0vY6ZWQIbc2hprs3czIGx
WfoAHYH/+JK8rFP4bU9qNOY2J6hH+inWqWk65XHI0UKDeo+o39rWnl0F37FP3E7BdtO9sfKRCJ90
u4k/FT1qqiXfKqRP4CSy40IVjhQWb3mqQ3VamMhM6LmKpuZcqIKojM67k4VMyvkfmhTscNZlBN2b
B3QQTXrXTtPyTYChGh55UfDl4u/0pth1gfk3SId1DM+TouYQxVJWKjemFZs2GEYysSzsok+wGDeb
vDV3Hn86Kb2Nl2lys2PapdIdjEvsfh3ltyaDw4xnH86ai6ondxaakdFsu1LYOMZ0IwKrhF4ZmmCu
Ft2AokKthvMY5bZd1zY6S5dmZJT6YAEojRcYtO0I9OwC57eIb1XwuGrWfULMY60xNEKNfdZHsIjn
F1a6ypam7s8Gy/yN4LCOHuAK+3b12IUFZfQ5GXhRLWJBASeUwyv/R+7CRW8w7px6HNZDzrlzCu8p
njNBB8Mw5MIFbr8+e4r9JI0Rk/NPM9I8s+LHs1JT2+j+QEogYSH2vAx+X2XA40S0CV1S4JoTE4Eq
5MCK2OAw0Mc0kk+KIBfXqpeTxMZOFoZAqWB5f/0MyVDPbyVe294p9JADMXn0r7cvOJq53BlCGGcD
SSURHFpA1iNirRqV4wG4y3jtwrPWwxT9y/wvayg0CrnUsVuayHsM6WKvlZjQiIXwGIrgs50uOGb7
dadDEx6lladCqS/zI0qe9+7qBXiXz4lTi3PXrm5HQBOlEhoYE8GCUtn8PEd1niGgAszp5EeNRKbz
F3wbsAi9kYVm0RiYkaFuebZTnwfRz+wRLJF66oWzk2aKKvcw79UFF8gGAjJgk+O4jFJpHpDJoX3B
y9gmIqkophg+kv3mvtAcQwWX6NMP1jYVeGWnaPtsrTNpAigZJKWBOXg/bOTUktOKH4Z6AWXKjWIl
hLFsqXrQY6bNqTgg3M4yU0UJwDxdG6Ve0BGc0RbGfrF26cOHX3u+Gfi07RkIs8sPu2J/pyYNJWoJ
RzOrsBjX/YUk7CuykRe4ZXOHPR/MO/ib+I8Es1zo+FStBLSGU0T/4+3sMVHQs4EVHkc+4MbZ1Jlp
/tQNAnUhy5vlHPVYP7b95nS4fYmHGeo05Sh5cRnsyjvXCX/0IEojuMUx4A7CGTtCWlTudlaE8THu
9f4vwEDQBrQnxKh2uA4LOdVbnj0jMc85jrMRdLKvR9AG7hmR1yTNHItL/QBftdaDL+B0ILOPo3Ct
Ce764FCcLEP4UbsDbryrtZPVa3Xb3bnNoRuY302Vcu7BujiBLLDj0Jw25yeafkz9hvW1YtwMnsEe
WYS4yhLaTg8xZURVNflNNT0kqub4q/xMv4XTk+qZBgMvBjYPhhGUrbgxIKk8iYen5jPoN50VbSsQ
QttUkx5vn9kG256vLTcK+syn0WGj93klOgVq5Bg+SzEpX0W3Ns360LFHfipBEAZmSiQK2/MX3FGT
pAWJFkc0cubtxiSu2q7PO0Izvu84PZSRCQQwzNclW7hQnsEyciR1LtZpQaaGKPizvfzEj0hXXR1T
cjQywsP7osyg2qbtP0CZFZZN5F4qzB/k66d28LG/WjcIiOKrsiYOm4h0P2zLeqc2X0Lw9Nj4mhmq
PqgvZsb3msNvgfbmVaDo0haeBtCsm4lDVB3N9QOrujTp8gkZDs1JnYnT4dWl3Lpgzk/ctcMJvN2L
RDwgt63ggEXucB7fJBnZt7TCbsldH1Vkio25VywZRTdCltgjVMQenYEE0eniPreufvQt47kYHhpx
GI9dbN1b92Ge+WbXTPNqYPkHBeNChWZbjGt21Ctvf4l3cQJtdNfceiKGVhSLOMWPgXyE0rSfg6N8
7l0OsQbolsJlsekpp4AyXH29cwA0ohJEHo30mYMdq7WHl9NFLoVFJ4CNwq6J/5kVgfEkVZN2QRy2
LRAu7JUvgft5qgwwTspOwdcboDWIRvcuAWJcIjMtBnci+qVH4ScLkLPIGVSGGRxk1Spta4PsTzxw
ppV778um0gTTBYW0k+G0e3w8rmduUxngyDw4o9JgGY2Ly+pGzrdheBsooT9M8+uhdgv4gYlMDwz9
OKJPkxmY/EKgzDFjYUbxwysqERQeZTAGra1F3NfGAxtQ6zre2YsPi7CvVszJ8Pt8O6Ma5cadbiao
3BWMm7etMZ6h6sxy3D0y8IaG0rTULDVyDE8WULJS8RBi4RwgEdT/+dPSsLE8IpIHBHMgx6ZCMwOn
a0f/9AuH+wf+r/GFIogsxP2cXiInZ+7Th3miimAOTwEGPigc4rdQd4vLxl0LSnqf1+Ad03Nw+lyL
YUxMckswL/P/1XGVGex9c0qP2bNZo3wVXTtcwx8FsRiNucVT1+R8fOSH6BlGYq3dT/bIVISET8qn
j3wU0SaueNOa24P6f6z15EoZCmv7GmXsKtgKBC2bucYU9eX4uEhxc2jXTI9waY+V3rwMS+6vZzMa
/bRBte70woJjdYv2OzVBYutgW64HLMbYIZq5y6SepwoU1LMqwTy1bN8iIGp1AlxoV2wfmOBDv2ox
3d8WEcAxRu7jOpXUm2OMBhrlbVOkCbYd9jLWM7ERzWNLXmFOHYVEaMWH4VkPcB2sTbOH/HJi5MWO
POg5TIPcxCHEvXQANwN7XQs0UnaN91ULRRYJHOHoX75DhkWEHT7bIWEj1ddH0d9bFdoHn6S2eOz9
ZFIRbBSL4Rj/DiyeSfLdnrH46nfC7LnoOHFMv0JxD+2qEW7fkOGOq1mVV2GgiHw3JI4N+BGATY+s
tA7se3LFsfTNf9yKXSRR6Dkj2g5d8COv3yjSWK7pWJlF/vmEkVT5UnCXkkez9Yt+cyl/9M2cX/8F
Go21vDsVyqMKRMq/sE4uatHuHLL9//JXE+trxFP+CsPo7x6TlabJYZvdajHJKNY6XHrQuCFS4gxX
0FN14XtpxMv8NQYrYfCjE67VZYy5wiR2qGZCkYhVaoUN16fpfwax+EmETw+tv4J5nHMpkcXE8rgi
NjczlQuaMjPZ3Z4v/+b0EYCFP4QM2ENSiGPsg5UgTDQbQI+CVHC5YSVeeLD+/zeCiTQsl5JqfZlc
ZKbg+7ueVe0tfd+/VHicyWkCPLw/3amgLryyDq63j6U5rxorayxYu1qEXv4ZsGuZe11ygCeV30cP
vof81InRwavsArDWuXpGHhNkW6G5efRcae5rwv5tt6aL0OU/YwCs4MxqVegZkMRESM9sPo2jkcxR
T37upt2XBELBpXqw4wbCN1t7CHylZt0wgWbMkJ9eI3Rs+J5PX99CWY27OBVKEx3ov4htZ+CXVTUb
DfG4lgpjOygQ39G+4y/Jb1Vlu6+HRkEZIwF2xAM91f65/qf8a4VnOZANwx1nLdPgwbGOEFsmXPs0
h3Mqz7GhnnsEXg0RLhcuZuQxLVLXlGagjoWy2nYvbWklZCe9p2wJOksXRPnXXj/HEK4JGrD4Lh7x
dXe9zEwJ50LnCairzJc9J0L+8PxtVL9nPJUimssReCfQfM+FUFr9quUr7VEzxJ+VXSFh4quB6tij
wLNzOTuuyrYodzAIWlxEOYf/22qRSl2jRTLt2Pm7XN1qMSGcX/IRDKCd2R5wNZIB0yC9Tl9KePUS
CvTJv/aU2kzzHGpCiPhSL9SnKCgwbUn2m512WZwPyQHbfqqA+D7WLGcynhwkg5TlfFUVOQz+j+8v
agmxLIu5cOMD0pYtK5AqTXoAS0id3vniNCi7TI549WBW1jWmHvPDEXqna6dEzilbzbNZAxKzj5DJ
eLG8b24kz+5Z/ZltGenFxM/0BI6V+nttUsBVtXNy1q7oF/AFMOHe+r4nOLE+3Ig2FUbxne+/Dnj1
lm48JFfqpFJ+an1nXcw6+2JObqP8YDL8XQDd8PL/+jfbub9pwpWGfakrNgF5G0UzzRCYKaHPC/K/
cFzZCI9DLLt256XdtVUO6QVrAwcRLg65y5VME6CkK+nj4FTsnRGm3iROWNBE3n2u/ltjesnLW95J
fT/CKjUftfCYt6gitWatS9z1VdrFxXXlIgwtDKQr7ffys62aKl6OMrb1be0/H4SRo3NoZRvlhyhX
NCj1qiTCaDj2y/CHAqp+2Kiwwaj7mj1naG+3OGxUPZ1Y8W5NwEMY0q63eaQyNlkV/8jRKNGJDDrK
yFdcz9bQj9YdldXchYm66OSgpa5oN+/sy2pVyosCd7cPO9ZkrnF3LAYgndoyzfX3UHJbu5CAHN7/
ZkyGAhHPGYqnCN67TydKTKuCGs3wbLzhotvQeVVHVb+vWR5QfXM4rMXYJWfje1q4Dt5TWdmwA/a3
ePKMgxiBBbNGef8n2w5wYIetQDGKKtvUjliJ4Q625jApAEnQ4UJ8s+0u3dZktOOBNMft3uDKZ82J
k89SC3sdwGDGBEU4FPUsMsTigga/zwTpljC+yASmFobMIidJYL20nIEZteRLhuF0hVEjf74TyBUb
qS5qYiL9Cz+unRdO85wi22MLo1PdD3K9W7zoP3/RkP+eHz6mD90nwLnZaD/XenH4vnQfzEaqdRDJ
E7TWIDlQ6jOuP3mBJdNfSjx3BLqJFPMU/GCn5im6xkLfbsSMGeBCDQHyb6ldT1xjpcArLBPhKUc1
Z2hJmGqoxavBznbZJRZQ2zxCR8eCO5fAfbyhLZN5MReWlCIUW7lXyrQxR2YsJinzi8ERmAq/BHU5
oJXQh/F8qNKeStFrqaXaaufGXf3jcCl9H49g/YPzF3oEP1FwBhp4zcslMOxAbBNECNooA5sJaSGW
i+KOkHxUoAnBeh+/ofUSHWJRSH9xzJAj3LuaoOwNKFTpUSiWx9kJghDTjz5n1LIwUgmnU23plha9
aKCiQt5lz7bYvGOA5VF2wnrHAnQUY28M1tItm5JezPYEUiUgjzJoCTZF1LrrMi6LZGka6QNlYXbI
HRmya9XWHsKQ8QDZZqe190k1m/j53Ol1kIdusZh7WX05K9rl4FZslqjCgyPCs9NPuVKlv6jm5Vjr
v+4QaCQQ+PXgzOGud1Y6wmM76HQaw/3WL9xt6Ip2vs1L8oosx5OXerkm2l84KlAFlVVxMrvDu3Z8
TvFPPuOmcxcKmx6Dszgv3sAehn8Qs3S/l8WVIiLAJCYfILTZbUjziDsPmvWYQF5VGwlfN2d640Lh
YXYjLHcG2bawQexnmynWW1EnzrjVs4EvurNsQoThP0MDeRXr29qrzo8fAmAiDfV6nsW9wT4IiR+k
TQIwXNGFVAYp+85T1kpMVeJYGOjAb7iHDYtKnV0GgPViHzu8gcBMEYRPov7WR787KMaVuy9YuZ11
t6Z0+ec6T1/fvoign43ywygw1dG4L/XL8sn+WudG/R2+SB1gCpJzp24AapFN0AQXv21d1fGVu8xG
dbvJIWOBmPxe9jnbzlohZSWtnQQE8U5Z4rqJTo2nGuwYEUWuDEYRGx2UfDUQ3D61c/chBpuSbQYz
6FCS2ZQ+76sO2zeMip6ZvHSfQLo66GgrLJP3hldezDx7YmLnsSlo8+o0AkqxNaeiFaH+YS237hf3
4FwK+Vb5tSiw7CiDWZQ6Bv0eMUIWEHZwT1NOT693xbsUk4eEl9wBqTMRxAVb+4zp6FhTxei/8Dhy
O/47igQcBID4Wl8mUUSwVErg+KVb7C6BAUpdR+XQmMv9BbPUrzIeRInh6wZ9KXd/gd/dohpXoLXo
W4sRbxqBZ3r5RcCnIPNckKHJ58yoYeA1wX0ReMvT4qCBYa0C8jXcoeFucwce27W46hAm3Fxg/JnS
csQvr6/2xRMt7Rx2bJdUAA/YI2MTnikYq8EaT1qH1Afrn2Q0umk1xhqg5rIGSkKChbDWHJ3Flw0+
N5m8ol9Gs0w6ZiHcb7IdmtLQFNylnZpH3oWEnvZdU++eY7JKxq4b4P/8285ARlEC3Dm81v0+0YHe
BYJO7//YxRHoRDD7wLfjgMLvIiCk+1XE6w5B2qnSeSOM9vpiYtal94cXzN2zOazCz5jttw1yCsEg
jwtjX18B8BXwosifSsQXmgj3iUakzkXsj+FQgTw+E2mr9vVJG9D/O+tZm48znlrgV1qZ4yiCeFG2
3BOpl9rSaDfh7RHPOwS+iCPkHbPN5TwYJAc0OSXOs8zmFwNccIYVDpOQvhBX3yI+NjwUQpUkOebb
7MAEmYnhizffmC52W3fDvzW6EiHKTjw8D/4wHPAzDWI3DsWxI9MBb23q4MTD/YVNF9V1BPy6h2Ck
FzhyuZyfHQLzD55wt9PMPmwp+N98x3rXsp5WjEc/qy5dt4dLhd8p44ovxT4cygte5USlA3iJCD/W
vmWZ84iruKr/xcg5xFlFiqQFxkZpOeCCV9tF0drPnaTALVo/g4uGKwYr6q0O8jUn8a74kflrnEbS
WUF/FnkFlgyUcUCx9zDX4OXMFYwA/3x2BNN5g8jgv/3FWfqq83cp2mV83vBEcTVyi+AfZfo2Lvgl
fcSb/l+Wgzy3NDW/+5ZOAa0tv6CtLiUrmZXA47GwdjecqPzva1PGrGCnsRExi2pNdmX5SUFsPfna
YrCNP4ScTZuKr6FTzPrZCx0hnUx8hQBaRSDQiUN2+pchArVD0rNEWTo1Z+4idis7E1Vl/NH8L5Js
EgPaI2VShLjNg+X2T1DqlfiztfTD+WW+moCGwowPc5yRc0A/mxQbCNUH8NGU1x38Dwkba2+5IJp7
L2r8thfK3jdKwdG8RKUwLPM6YLVBFrd95eJPHI+F9Sj+VR9vLmom1ocX4EJIvCr4oDaHn2sT1eaf
dLTEPCyIzwg3vynKy1Uz3mt89/WA6dZHGZVu2JylEFcwG8/ifw2dLXnP1Xp3T84RTHoRetJZ0Awu
giBS9AwlKW1hdif0OGVNggo0JDq/RsyRjEqe28uxyR8tC6OXb4/3MxkaJ7LraHTSzDKm0/7mRGof
uknAikwOxsk8okysE6gzmKbLnNv7EKE1pMmyZF8YDU/NRaEpP5JE9uZhFIlogsXDq3bmUoQPjNjM
25ev5EDU1iROu0YElR8PUhHgQgv0q85UitALoiNU3eyqcy/xG5zjw0ubMnRjAZqTqsPr3mhgZQVR
o3mlvK/MfIvJIdhPwsCYSIDStsS8/bq54f9acu/OLavAAmuvff2syYyHvH5CRSfgo8u50SaLUVVO
j1pVNnzJ4Vqd5S6ZNDtRuZQQ9wY7oJIAmQDeSirZbg7Lxf3Tf28Y0R1WlCvyLLddp+hoX7XAlbpf
zGUhexz9bKp6N/Y5EUUnMkm3+2R8e1K01HKR879wpWxekAoDsUIdmYXWSe2nhbXJYAT8d3lkxFrT
AzTFfTUecGlJWJyuHnz//gWKqyz5QYlyJ4ujYE9s5CdiPc7s1HPqMbwNuy+gPNnxtY3blMJaj+6w
xwcqsWlDxFqN1gwBmEej5MEkOY8j4u5kio6eZ9MdbuXw8HbdxF9Rp2+soV+RAaLeNPQOSXYevK1Q
/lnzdQkGLIZd+cX73wTKPnna80+jyARfP+zxxUIXka8u5FitD6PIR6wKkcV4qb83Pf5BKrgK2wOe
0RA25Tmbaw4zRsANczhHhWJUrT/DzKnwMTXRvgNm8DVxTVjS7Bg+ctajYv5YIc54e5K0y3Lh0Vk+
0LFG7vV9dshCJS4JsrTfY6rz/0/xDP+XmiKsFUrT1VNImRq6UMucx2cl76mUI7sAuLe+R69tmGFJ
4BRvMA/MaOsQKOtT1JjbbisEpoLrYxA+kg/M0PZWjFgmOIvhnZLLD13vCUbtrZLOa040QB5RSeMy
GQaxgZm4ivterMcS3gNKR5VruCt53Pq57PjRXc9Au2zasmb9cpPOALpt2+CmucY1W0/njPoLuMg2
AvTpzkHJluGMo2MbK54nbq0clIP0Ss2hcx1P4ppilFx0A6ISfplwX0UV0Lwx0BM1PZUb2hL67xeb
SGr+mx9X5ikeFSnOk0wvBMAkDqLs8kWG1Brj18zrhvlW+ft4WY/VTwuojZERU3v1Fm2B7T/9yf9b
u+PMX9gzKFXtdhECD+yKCHM5fSPsoV2c6BIGzS9g5kAS/2ayy6XtsN0X6huHNdvkhRgzkZkA/dYQ
f0Mwrj9nGMnOeEGxUu1TE2OV4XzA09t4rW5kDXePwV9fUxJTEt8SKnAf2eJaveBUe/aKw54U2mO9
TIdYwEfvJcR60ObN1G01OgTvRtSCiVcL/I2+c380e6JFecOduB21bCx1XRfSkh1yJ/ae4uik3zp9
7i1FknUr3Wjynopxsr73FNBD6pwEBis4Sqwl/UK6d941NFj3VUZJYaJx0iFfSyrVftfnHLhCNH+o
VHUApIKGMEXawcft/EgVQF2Q6vl7llzBexSaKDVJlwtYYdCW1AkT1RPPnuUKuzLE0VZrsRi0gApB
KyaHOtulnkyDDii8fPg1d3UzllWrvZtyKAsCNIMGKWX/AnCV7keLDEmn604qxBx62rXnrj5WMTqc
m7DW8Rorwj8RnYQJRBXA9AiQG5F7mvkq6j8cjfTyTzyTrvHx8gcwGUD2EgDsxCv1I4BlJx8idB/M
HbXHm7eWsm12h0K+BYz5H8IWMi9Iqzjh60dYRPEwNrUBH1dmb1gETd+H5NuBm/wCFG0bnB/SFgcO
Vczak51NQZRKr+zuFwVYZ7UKtQEIt35jhFLDo2uILexj50cuvLStqV8aix4x99JWBPua5LvfS34M
eh94LoUYRxpt93hqbaj97OlUJS1Y5fPAD7YmqVI1e6WviXv1kJ6sD3QBpLGgdxhvJLPxW0yLwR9D
6YDv0e5b3LeOllAhkkJ6fDUSJ0/ZaKjc9pV+M5AwUYtw20ERYJeVfYEJLFR4UcPrGZPma1192gpd
xZmZ2hETTekGQjhsets0OEgiWeNqCjVxJ6aneq6b1qFMw316cMlDLCy+1VQT3kbuwIb5WNZKfDp6
UMFBRFWio1xzPtD8QrUoyO68EmV+tquDHahCztbLzWjmVE9YHy+gaIytng54pPZ5BHVF2DJNr2KD
lHPdie7Egl0gjPhpjitCwI88G965GsyqK/oE1B2o/x2aUxlud0IWr+MIcImDYVTI6IMn2khTwbbR
u2muzrSArlKQ2usjpp/EJ6SOZ33+R8UswtqVMrr19Z4J4w1r9Kx6xVNI1vKVzCwnbZ5Ie4RJrvck
6ACTAoa2IEDvNMlhF3N0RrCbUN/FLM5NAJ1YD39LNmzJtxu8mJ406JIUav0f2cLkkNR9RTXRz02o
h5bf/A2bcWjrUMsVpI/IN67uMpMjC7GVrQEtP3akVIwgZFcmeVeILg67Yt9LkQcCIT4iG05fRtPt
v46vqFT3gHFPKDyLuqmFQ4f/v/YiLqbc9oFyREbXqa+Yy5Q8A8AiIo2d7nBQ3rjvhnK1/kQDE57u
8pv7qd5sp1WekdcI0VFqlqbddUay/rt0Ryz5pqW06UDVSWQIOHxxdPcW8UcFAmZNfeEtQF2fwEsT
g5mjlExFR+Kq7IrE7oaa00sYJ4HN0OhP1d9bZmcF6MYtwg83VIYK29GXM9KLmd0pAx90tJLOWdSw
En1HoihPevafT+4VsV3kSzRveoygnFptjgeEzC685s5ny7Zby0CoT/Q0lqplmjMxtja2cdk5H6A6
mB4VZi//o3T8yXhsTJpbI8YXxUuxq4ur42LaRo4hCZAR5OnoyULyO0QLP684MnU4jgtGqJ/8eg6t
Gb2cQHSC5veGL1xt2UpF1eWg0W1iZbOZ9AIx7LPfh4y/6JWi2j9NxfISvVYnFcJyFl7YQ+PybFw7
a91wKlv/ENij16C1C1i1vcr2wAncDGIeuhedMi/KeSjyB7WxnOGwdjQmNSJ1I2j+9ajvNd/v40LV
aG1REIbLtd53lJproC6cBEEFrqDwgERBCc/vW2kUuaUR8ief8fTtUSbp3tA8bdAqe3Eae0eDP6OS
7jERg7spjTlkUp02GUnD/lzyj9O6ShY07nKZsYgYSzLKKN0E/cTISPSi8zTqWvhZ3d9ti/3Xtc1o
L8UfBLqfpjzXfkz6gfqvDhFGSL1BuC0rv3SAP/LJlxODRW2LvK4dnWzlpLhOCr0tsUhXCLFpk1yH
jzvY+rKXSw+HbJEtErGXj5CBmdQsPLXeBrWz2B/IF7rM+XWuLVlD+mCGev/F6OALBzVF8+quM1Yn
H1L5Z/TkezfCfX8UGGk0fkhkgmVtcauA8LIfWEKqnFgdk0Pu2D+eqKjaFcFBpYZRIs9jXwv/EKiX
GPLFZY2COuc4rd2i7MhpToC0nUouArWRGorhMzwzfKJ6zyjr63ZFJMAR9nXv6X1OoZQ41Sv5+nZJ
kkI0FxDOAm+osfSV7YMvO3v/y3Fn7dJ9uFX0FiEJDFw4OT+TuF/o0lkb0Irhx7Qq/LJhk/c/NgjN
ADzUh1WLWwlY43s7rPXw8XdpLEbho3q2F9dal7dUiAbQr3HnmlcPJqwdyc0vwaRZ7EVFZV2mg59A
TlelFMsvdd14njOyGlC6B2RCdS3vxVpRtFWzq8u5fk8fJYU7ni321xQDeOSqJOIohcHcFKOnYm+Z
v6v/LrgxK1xoRKq0faYF66+XNF45NeFdlHnFZuOaPg2AJ7uyflpmIoL4VTTxnrzySLYt10nZWDnp
H3sxMGaIXPFcDyb1aX+lEBij8nsjmxLh58iMrC8L0XpPNQF2IDrtCtTML87JUkCDlNmEEDHyi1Tw
K304RiR916F8NqzyzsYnAmgos/b8lBapwSt2nGp5Gcdr/jwOX+4Soxi48ymiKktMqz4FfkXQgVEd
65c19ydLajdrXKUS4CiqP0rWnILVkdL4u/lyor+wMNPNevH2KJuX/gSsPHiMDBA2+L4PQ/1UqGLN
UGAakFtASu6RSC/u2XLQ2G7uGdYIvigHT+fS56dAe19AcwZrdjeJybQ1bI0KfY/Y8ZN5iwgfU4Hq
gBvm6+u9vI9XL/kKg6R53NfmyLJvOi5I16yXknjpueGTvUJ7sgE48m8OKnKlyP25JZ3gmiJjVGw1
kkNF7ckBl9UIeYRu0ZF3bVOKBlkzCGnrLndyn5YiEo+uuRlESTzyi8/BtYddKrlSyU4bps3zFsoD
j3x0n6XFZRR0QfD4z30JlHDvidxYYdd6BvvtjpUHZUPM+XodxwpPUtaOfUnOpazDSaTcTQNyHxWV
dOdLFfD9i4MsScYRtYqGLJSQQwJjm+5AfU8RmeM4W2CeLAKwicGjvL/26ggfUZajFUVfHviQvg5s
TwQOkdNOYK4ECHThgZEpYA6rbmIVipvVo7IljVEZWcyCvYWrkN06XM2tdtoyjFgeeLTcbvAiPkxv
qK/xF0/tyWYJJbEyQ/io7zx8d17gWc0dX2saPf/rmRhDNQVqDHTZX8ZuA2IG/FgJnodBGiTV3QEd
rHEWlBv1RQDGO9RD7h59/rZlNzmQqqlMdMPG6bGmnxf9h6igZ7gobBuaP/geltll8fwVdPH784Bz
jjrFdwZVjlsV71vNoMl24H89zappCqVwwtdP1TK69i3GahQsUMXMkFru2V2pFuv7/EgWBP7rjsST
xByQNqdrezO6XI1mt8/fLykGNIwYGat//WvSBXSWfxdxkSQ9zfQ+G7PNHa+UaUtauXsa4ZPi6Nnv
t0ll1iBNvJOCP2vTv/4bU7JpQCJSWDTAXXqAf3w++s0WsLEpv54wVeka32SprNDTbiVY4xgQTpkz
GeX0EU0hv0yo3SzT8yZl+nfvT/8ooFJw3yMCkUWUFFXy1jTvp/kA50wBmL5IgwiX9Yu+qU4Gqgdw
NinpjscE5+HFzkGFwhkprkQq6P+9BsTac9A6c564xyi1EGg86Udh4dKWsbyEAelyHciG6xRKxfb3
xu7QGwsca6zgTKKxM7GUuM794iiGDmzm8weR2+R3wzdcYY64ErJ2s7GhKnRdWH7lLv0Oo+eCQ3U4
FqT0jefbLvylgRNEbKFWH+4ND0cTZrOWKsnyULaH8NEm1n1LAWWrXOvkCshQrYehA+AjEpVNBAT0
l2QWNdwzr0tpTflNoYezsePY09R2INqbSo8ANFZkYH0UueTQr0kpLESwlN74rGWw0y0UzsmEGPKz
fw6sggshRXzHC7luT5DLLQa3Peom6dDm0QyJv3u4yWVU2WpwI9sxG44JeerOa4R9X5GE1c1k1flS
GrjjQn/ZnvgNCpjg9K2cBnloUDP3AkAMO3lcZWHEhlI9yxDaErRfK5N5QSFHgWm6G5PCh/pF8VUQ
hvWBTWO8FORg0Lf9JSDNdLMcglUCZWUYblkX1OMQjXCwi/towc/NbQGgINv6fHRpUiMoPzkgRR60
qD89Q0HDL9ZCNyV7XtRw9dYQqDoyWgyH8R7EqNSK/Lk61oRddX6Vl5Nx1fZjVfZ9tdA9wNUoNIIZ
2pLeIn+xt98TrQOjjYYI+dzPoiXMkW0buXZdZejo/Jn/cyDwKQfoyUvxj8SGMw+yyhTXOSlBiN8i
8NPguHr6z4XkwsJhJzzO3uhc25PGogvBl8CGbOmOAnSK5EyDJ2/bBXcGOIFJ09M4iUiAmCgBQLt1
y8TNDhJm4VoagL21ngjxiwCI46NUBiB6yEsg2Yask+ZC2sjFSPvJTSW/NQsFrRKc77AggSOjlPnV
GiKJqd+mJuk8rkRJy5kU5uraCWC6/S1JHKwMz6ehc8fCVM2/p+5fqFlyjE08RNkodboyYblJxVjN
1yIWddffdi2VS7EYvAPgJQIxJkhTNpdJe737+HJv0pGCu+qo9HYHjDUTeFAa7tzk8Sk2jk8naADa
rzS4PE7AYLQKQh4uVPWS2+sW9j/8q5QBk1DTDt3+fv6p+qvvImCl2w/uh/takAKCRQ2Z+OZg/UQ+
FUigDVBOYOVM9giXhAS+IeDM4xGm+Zrk4WSNhKuTgG7C9HPOC5BgP4LVYrxeQS/J4cOSXJ834R++
XhrnGhkOpdNhzgbnlBNuTt6pwY8mmonAyGxciTeO60ljakSgSmh2m4yA3o0xtjM+SpkR6c4NGPa9
LRSnKbyzSj8KdNmRDrynhN2qnZyrG+cU5RsZ9VwUszqyglFta94g5ifw0QOD+LOq6zNhqEPyHWgj
WhBsdiVTzN18lUg1DuQdmjwdmtJTmqYZX8IA0hJ3dWqbhTEfXnNjaO5Ww/ImDx20DrqKx+LNR4D7
9tI3V55t4OJ9jP0y0SIYV5CO9ze+Ul0LgBfIphTFDSJptyA9MU8n7w7T1L6g0d30jTfeUFxRg2ty
upQzkYizQQCffm48gNiZzJS5PiNa12T7A/hQMJnKYauOusywEI7WapkRQfMm/g8XTe6WJD/49/IH
2i0MTNuJQ0/wQ8DxTysxtrW/sJiclmU/FbixKRgFmgCgG0jEl3OraEJ8blS2sIYdXRFtRb2HDIdu
VPV1qKgEBI9J2fjyu50StGF7tp534PgCxZMR2DPeFn6hod+XC+ob2UGB3RYsG4ZSOgME61612OqS
KOM2dsEMp5bhPNGB5CePofyDxK4vECe3ZNf9Ui5mWEnwBWpqRr+615a+XSbOgb9oKEwHTlqS5ynU
7kO+XvCagrd7UVvW294Ety5tgui/f4b6pFVxnGdLIVX4pXONe3gpnRfqfMJQPzNWmwnDOZ1R5Ihz
upMSIX3wT41HLViDj8XZhwCSq98Gk28ulqF2budcjW/hLRRbCVcLiFWT3c7/xDET1NhFHbGbfb0Q
RomnBHtOMMDda4wKtSkhcSKmSVBkBMuSYMDE4Oy9E6RZZw8dXQt1OTqY7Bcu3oULWgGgpXRenLtz
cn0wuFv/7UagOYe5XdHOibLXzpeLbzrnoB9WlKtoT31OZGsN3GiIatyojL3GSjzivQwYETt/4deP
IY/guRGBI8L4GVsL4XJCFLbCujGkB0kmMPMWujusSzbOYCyQGogPMc/THXt99GY4pocP3EyW5H3N
3n3kXYcKly8zfnuwt0eRhtr3SXqC3epZPDh4l+iIamlaPBH3nwWVvr7DMsWOWgJAMVdSwnRFaXP8
jDEogf30tPx1c28bF+7nnmvJfPyvH0bEma85yBfjZVQramAs8O5rvR4T7GGLPuvBqp12zN4natmk
m7tVGUK8VqX+gfMkICTBjnHE8g+0Kp2moZmSzsNx+fvb/NA8JApt1rwx7QYt3BKRpnvsb75/djAG
0dY9XiJtQYX0DT8V24Viz/aZgqb8q0JXSTtx7eaSUYJp6ewBGc+plk8ezp2I/IG+i9UvDtkPCcVc
8qwBtFMGWVrh3E48ac/om4AwmhYJccdugJ+u7c3U7/LhPrO+XBQ2KoO/Rek3tqUL76eE5ebCWEQP
8tWjpIxQ5rWDQ4Mb/YBnzMgetlkEMX9KTbWo0g1pyTkxIkmQ1VJlZrj4sw9oHs/D1TvY48GK+KR1
lSS5yxXmBT/cEW019N211NWTrERIgtDyc0DEd/23HwXyXhsEfpx2rqBT2zUDqJxtwkKIOmHhlsOe
A09zdAHLnHE0mjpwMX6PsOksXO/6i/BwxgfoBxCaNVo3JKwexnmroBrQ1YGgxwke+iuX5Mre5BwT
H6ngr8LdZnvbZJPspJeSPKpTIIRVr3hJQl3m4VfhcrtIkmtdVlB4c52R136G4IuuK5KydooqE3Uc
DPBkDz30QGKMr8xvPY1OJHgsPxwRDINCqiTYA53PqP351U+C6LYnBjISe7U5wuMRsyESFa8Lq6yQ
ZY9jcnBobDv0NbbDkLXOvG90JkIptZSF+Uz4LHVs5mFG++3bO5DXqHvBwtgEZ8viUaQgOi8C3AAy
VygfqBNHBs/LR/CzUHbXGyZXCpIPgl3802EIupRtUNSCOFb6FJCQRGb9TJoIF/5niZ0GCzQ3Rhus
vZ9NlheeAarkpRjzvXQLXvVi0IB6g9O0uyyoWziGn+cPSxqbae2xPWlwnXW5Xo5EMqR9knzSj/f3
O+zigz3qK6nCyVsOMZf9wYqrbPcl8OCpPfd23q+kAolyjsf7ivpMuvc0vKtfB0KUVrLmHbD3Op91
734awNM8wMAkmiSgQF1zhMvMee4Hy0XjEK8jDhWM81kofNsH8V0r7rBZOzlX37gSXI8XcrBdY7vT
LBM7aCsQljUiPksyVPoqBETeApzkO+id21/R4vGKcQxVBJnU7NZ3mZbSC5eBNG4U0tvIRhgw1OPE
pb5Yf1YO40hKgzAhwnLzvp/USLoUrpFbJMfopDUEqRlfNEkRRa6zQiQzoBS8EYbn83TCbfD7eCks
2Ffu6X4Cz1lgchc9CIwrZrwcNFqRovG66NG3XKAkK7HG6VkXCVTmi7XZh3tJ8svCEGGPOI78klKU
46fsYCiD0p4vV1rK4aP8SnxlDkYDmCxC1vxAfTbtBJYQcugSG6HQP7Z/KKnYlTPfWxmou+DA3gmJ
FAv2UrrJL12IKBtXZ5k1LwvXq+NxIO1OaGMKoVI+FdoO2QEVn69p5utxbW1Csho3sp0laBElgKxU
n8mHBGU9E6M4b5k7NOyE2N45PLEMnz6ZICrEIN/vhuK0+PfDOi8bzHSRC3x5y9jEQIMctaq469gH
OzclCo3aIGPJHSEf6/zTh4n8BOJqY1Mz6GSMe49xrDP4Lf03/FTpyoaxYYPlfsxmxA3wOVj4Q7fC
Myj0x6IpAvDy7wOi6lrqbD+vhez63qM8+8BUTLrFgh3Oj4e3DhgA38PWk/pb89dcMAbh4MwpHvg+
cpSz3/lojEJHAPcOVPksxfmAbOZ4Iy97rvKVa0uL2mn9FHaOp64AfbrvcWFqvI6WTrXaXPhUTFxO
Irqmzn1FP5VQLrxQtJr1J7wJ2CSz7/ftazu6AJ7+Pg15r1t7nwXeOn16Mm6SW3L+THyn6LmLyqkN
3jSLpCjivp+EkUppM+uqcFpnACKAupYbqMXw8eQeue2BUpTg9XoKFKHb/lJrSzIa0NX2lu6CDN+0
LieZbfXiH0i95v/wz6GN+aWU7IKqaPRQiVAb+qf4PMPWMLmSjp8WCniNa2eMmriZ53m8aq80Ikb3
0R+DdmQkM8jqHzDlrxLo7rwNAPBQS5y1PcoP861mr/z3pQFnuTDh7Atpka7MVljPQaqVwnDy+Uhb
UaOfyDHRWEl8f0BuknQ8S4wmzBXOVzxdNjQGp+qK0pqfT0PeS09Lq27ygMw7U3qRtSr2FKXWHQKA
zWO87av53hBT6RFw75pnEQpK6lZywx0wh3taI9JAagPasHvPuOPbhvshuaryPQCnh0YHoS+iqIsk
F6kSDqaH0Uwyg0LFzFkqn32OUM9pk6/8/Ua9xg3uvZ36DxeVzW5LbKH7Qkjea6r/J4pSJ9w7JMo0
qk/t99UnqOK8EkbeGFCsKC7gJIpzpAppieL2rmLDBbAbMloSTbyH/CcbdB5ANZXByxsIpzdMw+3A
DX/MdZDsd7uT1e96MSm0I/NHtLNIBfcj+RIXFBvzKUOPihgCD5rxpvnMTU1ikb2HbIBlxtiPBxWm
fXd9Y0Ih2d3dxWh3CtQ71rCfic3Hsls6WdjXF2VYnnb+/YQbYZH77up81TRvJxqGrWBZtjcRpAlP
1a9uKrjJ9Hye0tVstNbq5so9uRNJPqR6mBjTx0jJsq1gJ/UxaOp4YEyapEUK34SS5CnLeDJtw8ly
4sxa7RXMhby7Pp3iMTWnnNki3gDgoyFOujci/A2m+BkJF4yLwNsqSLOGAPDW5Yok70nd5ljslAq1
wwiNwcUVGeYrsnl4woFrIDPkl66khnDgHDMQp4TkhCVuVdlqfRZB67WZbjSfD03zqSH4VUMzqH8M
h6HK6We4n7ICndBlgj6ju80+GTTNfaRQgj3E4DL5Yy5AdxIX9OnK8yRUI8KYUcROJHhHB0Wcvfvn
fek1WmiAUog1tj6NydicH5qpXi7e+2gOTKDNDCfHMPBiVSYkEfF4baIVjkT9RuOSGbqXZ5/QY3xa
77rweKfOoYjQp8I8FqjHQ89TXwjzTywIkho7Z9lRVDs/8pojejqMpsixANBqvXalGvtyAvXxTN6l
ixJ2OQVUvpUOv9dwFpmU8XHJaW2Wea/v5sGHDx6HS+nV1PUQBEC4RTBwmGTukNDnktYuSqWw5JBD
+GWheutvtH0SAN3exbrU+ihL4cZtgnyvvLBZo8pDAsLJ1oejSvR3QxVANtlKLbHkVWS3blZ6Kju6
MjxuKrrdlz5OcZlj5rPudwKCjasNSOtZNFuBi/HehAuHLx0LMCK4ziu8BK9KXHQ1aFua2z8J8x1L
cZYnvXzt6yUPM6TQiyLde1NpGOY+UMB7QxcgdH6Az6OgH8kM/4Y9FJVO4u8o8Tj365kBW1zDGCue
ptITYcQW8+JbVTGHdM06qfuQQuQb5Jvgh7r0CrdH4Jx8C6MRjOw689rGt0n23ImcthpSajxdO711
BW+coEz82Gk9C2rW4gtyKwZgDq3IWo36RNo/Ry1fCdJ16fo7vOKFKL+r3/0gHtLcKeMnHfW1eJNO
sHEgZZnqIlk5sotJQ7GxZo/NervpExwMkM2Q42tV9DtkxlBa/prg/OtooEDrkJBzwrPTJ/mcZd2s
CxkKcvRSHqhwSAqOsKHJVZznU2zXSBsqWNLiyHhyHNx0VcV96Mt/Y4zwM/CogqU51HufrrTV78rZ
msUAiPPaRFYtbJFYk6KoBaACwpS+SoJIVHpujBOWDut9a0mR7yIb3mmrg5nbxrB7w+iWYv65Pt9J
avK3vElUCcutWMcoBLyijMk9hngu3AhOjPcfUBulTy5JXtYW+df3jwAyYliwl1nUgowKtGFmNHjH
x+DfmqJh1ZcDx0c6rca8if3pA32CcBmtPnBxiSMdqR1KKxWDjupGWXV4jIh/AoOYpo3DPZtU4dev
xhS1+NxUT3SvpOewrpKDbztaIuG1PU6M0KhE/RMguaObPY37KbqqGg1LxGhPP6bYEvNtWpDrfXjz
cVBDFw99QG1RIWiS0Q2OsLRF/4fQ2dQB1GTdZvNwZ+BuQCi4wo0fiB4aLi29u1sowE1RuelpDIFY
lny/ezJyG9OCoXgBFlmP9uSh9Y4IElI/r1zv6K6vVk9tY+rO6TGANsG1zV7zrA3lR0+wxPoRh8EC
0iCLIUilrrR5CD1qxMivGEDGJTUiS3HS/ARbYG902gMlTNDV3NXvI7451SF2CKpyxNUA7d0wuJBv
kYgO4NNJ9RjYKfrUG23y+uSMWW6z34PdCLVPVDZRRZFlnFdVdRYkZHQN9CVRTHogMGqxvuAEqvEv
zfhOoGd3ulfRVos82i6AVtsWtkQEQ4awv6YTiKjLCVAqa5mWtT3Nv8ILISSUBNS1SBxk4qkR+giH
qtwyZmJWOHhbtHp09A3scjuUg6N5Lqka05iaR0164BrNy0SUX40x23qWAjrYaw+uIpFNot0LwMXs
v8yCKqSwlijPQe4T7r0LaibqH8jMqWA+WgKwPEQQho/3oMLWMZ9w+cAYgCgEuXbjidNY8MNo6sH7
E1kMA7XsSRQJGyHq+yGGya+0DSAoffK2I8BHKMC7BZywX4smSqCnO7nq7A3O15BINxJjQ/UyPZ9j
flxgm74ORGY2VZojeXhX/4WcFt5xZDrV87vg+5VvirWU4lW9/RqLYqAxzS5/1Tptq59LTR/yMe3T
i+yMgKMWk7a2HEhcKpOu8DghgcA3Qcq3f9emrVdwP6IPuA+YR6PA1LOKl7XIhZ5+7nolpiHenIFy
TneJExLdtwe6PzJPu9o6XnyXe3TzNZKv50JemN/jOJXzB9DNivBHdW5Cb8Paonw6UJOJSGZU9x4+
LtlamKgjk9i++O3Q24BPT2X6g5BB9ro4oWYyJQolw0l5RCziL3qTdg9YUIIr3xSOH9a2dUNWUbyc
bpabdiRAIMy6enxPf6gQSYuSenexm+eVbpylgNRQFds+vT66PeoF+i0oHeMUPGYDNe6nz/0ji0g6
KrZEqaSjFpOo3GLM5H+OOhL/KeRRSh8XNZglGtl9FZ/es2sFeR4lnK4gylz8xvmXLfhqA2rkQFly
CRj6XCKaSE1v30OnSI1lyOTNlK6oUaCQoGU36HPczcEmQeo3zOPOB7YefjRRA8vfYQBb/aVXgqqi
mENx0y9M7m6X9P4xnI753ooPK2cPcCXRirEL1Xs4+B2X1jesArxfvfOtQiLZjqrlwpyfLSOdN0YL
vcaMwFKpVNfLlgkY1Be4KSkOEzOcm5mSJ+6IeaqwNuiqwoTHlWRfRhW+9+r3iOTqanTXYnElthKh
ADJMgvQG6JO1AwL3W1Jxndzpt2u8RtIKj1eAHzsc9sDy9/jXuOPtIp5uPhSMEGrnwGTGL2InnEgh
FyD02oHv61efI8c3Gl5qY55E2rRXtCYjOVcon42kiRVwsvBGdlzVl0Gw4/JkN0njyW0FbI4vXoQk
eYJ8EHDG9SsMBMdS5b3gk18qKBEir+etA+uWQwDub/QYCJaIVruCSGq8LfJMl2WAORve+BJgPV6E
99/qVNGk7YCZCHO1rvjMaRP3OGHtSSZFqiLqhspdV1yioHh9LUoVJpsnT+A3xBBh+tdtawLEl+TY
9+7jJAVEMJnuj5Xrhk91+gNo1HE/vZ+lvrl7tR+tEdylJoAzQApsPBXtxGZiUgO6pXcK3BQi4LrQ
yC+jB3Sd4dnPnOBBevt/4LZiWLzVNexP3QFWKnbUGCm/1GRwKX5X1to32GibabOmRUpaahS4Boy1
BADmVl4RcLChlBlt8DR969ZLpjnHajD5ehJKDPI9TGc5a8PrMJUte17bw04PDq9XyYHaqMa1fo/R
so88ukEEL2gOvh+JmD7KdBMHdyG4DEv003R8MKmC5k+Svd6KxeTYCm4iSBX5v7wsZ2d0wUhtgNgT
vGZYfeK+2VH5NxEXrXSd7aH7igI+nsJYJO0E+QZthwolYhUg+ut9nw+b7x6SucWyTcxmDn/sIbu4
aT989AZ1CZRXtGVEtgyKSUyjrC87pjXHdN5JXfLywcNyu/VahCDbO8J2qFpjEVRUngAYXlK7OoB0
aljoAV2KFsC3sk9DSFJEY+jxbY1hjOrbBu8dvz8I7P8MvPUFIkrNi6W+PnIfzeWRnlTeZPKA/Z9e
C8aG8hrYPtLZoQONvJ2KrVwwunoSjeOUuBUEHJhBhrhkz7s4PX78+zppeUFmjBJ9+qa3My9yc2ot
kCGMs6hILiA/mCQjZn6eJboPftsRTgVH6Nc4Bzwl2g5PBWLfNrL78q97nlwG49k0xPXWwRrvMKJY
yYD4ZoaHTR2ZkAQveRiBrcadV5hi+iZqI6BEr8Ge1dZ1bb2UA3WjoKw+qjWFVq8JMZgaOi3aPopm
NVa/a7cFerJeqxCh2JiqvZSeER1LDl2qXnNcOUgtbUhRR1CNp2DkHyVONFN3qxDeL52Tlh3ef6kc
l5fmR7Zl4O2OzawFv5ziD6tkuTzyOkWgk5h7lASLAZxoaZZNhmi+PkMSz+F8jSawUOAL1FmaLbCp
nWanIYY7Q56vSiMbc9XhDq1TkKd+fbvi/jX1IYVr55SKK/BGIcX/MQYi40RwYOHhEwSjBpleGkCl
Wghv34ct07Umk+NiUxfbX5IWV7x6SomVBGCqlOXkjOzVhQl7FuoXFrzEgHdLRRFht9vU+nL93LwZ
qzADQxul+qlwmo2SynobRusGi14+gD7iqYlIdxsOGXgXt6cEfLwlwziMFD4e6IXhI9ZGX3FWnfg+
DXecdWcshfvsoQ2g2I490x+JPif7ioMlrFRnKBjuFHtfCNUIAZwb3zYcrqywvys+Y0jAGlC1rbUJ
S05g67J7Qar/TyMaPQc15U5GejpNSVRjD2vmHEZRM312Upkm3wTYL0SRVkZ9u5veP8f+I5/6kqf3
udz8OGKhx+Z16iHCqGimKMZ0gVyPSjiJbGsQPYP/NjnekNqjrGlhmHOpAIpmIXPpErkEB7PbDCr+
dBg3CO8RH1T4H74YUlWRE2fE+YrwCHdYsD3LvcD5dL/YqTq/rJVez2WtPQCFSTQiPxA5olp5vjjP
OqM/1075FbFQ1snrs2VNv/FtqrksHgoqaoQCtf95DhoB9B2BmWEp6iIJP/mJUeV6G92hqpUEZ6d9
8Ml1exNdr8LDUi6ZGAjrqS5uFGQqEujkrm/PR/TWPQvFcWXkFr1Xipy+Es+EndiwA4vUGJa/qgY5
d74k75h8zQym5IfqcdwoSh7YmcSvrNK8V30Y0s9woQcSb6YvVshVIWERqFPKAimY+4f8oECVcKwy
ZSV/lo7UZv69JxuP9kB7I5KNa5Xtkk+RvuQBD6pep14NgVEN4dS21EOa7Mhlwmrq0rZ3n/g6vVKx
2rMFfRQRjCsxFdPubEgc3JJvEiebYOTyaYAUKtDQQr7vwV1+WG8EA/kSvxtGkX7WvEz7Z3Sr7c2h
8bI37UhVTuP+KazE7t2h2+fh0WGHWO1GmbZ/mN6sEjBYhANmGcbUwk396LWv/z/A/WLZ0DqZOQLX
x8ww3pP3zs80BoRFGHUcyeQWt7dkePSy5dd/Ydyhh6blvwnQtCG5qe+ibKlAYGvB2/lHOdQOy8Hq
lyZ+fVbXwODP04gdLXExqe3Qw14nND58xrMHCSEwt7jRUvitMW7a10cLgSrDmDjXFM+Vyl6r0ShA
RUXVXLidThLxy/jChnhloTtae8wGg6bTJ0GLIGOWVNBmSSQ6dpuJR1Qxmwek7miYjtwxXr3Gj2M0
YwVM0pwmDYc5FiIovYZiy20XPDH1Z24Th/Is0aT64mc5xaXVo3h6CjWBzzbwLBPbXUHOAoA0uBxy
arAiNvEpmwQ/rk+HK2hipsmD9picJfYK7xS4wqJe6f02FPw4oVKZyXubSdQeWbzVFaxZrijxccSy
TkeP5IyLL2bWUjzEQvI8KMcHueSZGkb3gmCXIq6miNOZTaH7oAeZR0VwtYw/673Dn65WrqvXwIt/
h2sK0/Fhmo5vrHnmWks7fQiRS+OSGepnsB5q3I17o6Z43mi4j76GYCYrGJZV8dn5xXqqooDPkNZL
MidpLzCjSVNh3yb85R8+0DEox0c3SIM06q1Q9H0av9gsiVtTSRRm9GXChHXe58ft3g1Q66ZFY/tq
Cxt04juqJfcAxzTPU2GTY/ZnutDINOFKNKMBa+/i8FUt+PkV7j2SzcMAPK6KqtUNyH1TmGdtbrXO
DdtMZbANcBT1EAP1f7O64zx5y5oIWEIJ0z7UMkoLwiFP8/nZbqx5bVsUUBzDqBv0/Apb8tMrajJk
OBT4NkUl/57YPcJkgjRefMY7BTjAo32vgYtsxC/AfvGVf27mi8ds6BgsCXobg6yxWCDBwel2Bsay
f961ZKT3LYsv+wsgfH5tuIRPOEomj3tMEPxcHAZmMuSBHncyV76uFjysY75PmyyxMgg8WmtmTsEa
zx10khBNTcuIy2K4UC6+I9Oxedso8g1nR4pvNjvmdNybP1BscCR5ZjJesdGNOEWOin8uhByLqpqk
67qhMv6505por9+GIv3SFi0hVSzys1hMgJqgASWSDHQCjVqt+G6XLZzblkH2dtlt6F1tG9a7gJks
sCz0jM7kiMtZT0rphSLcZCc4tdsX6aEAsAKnON0sk59I5jff+o60n4bFK+tc5l8JHaxBVDyj+flH
xrTSMHEEsopS9VkqCBdqpKkZR0mcGULoSPZ7G8M3j+YiriidfXc/M5rKlITCHqo04ZtVFJSN3/cK
yzUWfbfOogmq4BW0PQy/Zx+cD/qFVV/vU32BfovEQ0pi/gAwe2k7lDY1l+lwddPE6GoOBAaG/avf
NOK5f7rAfhuxtHhawrwWy8M/ixkhxfCKKtjr+B0VdPpCUu2oBlbnjsN7JvgrjsxxIx2cqu8RTbXD
QuSBJtsdNBdKSTnK8MfLjbrhP3QMLlFWrXXnT1avUqjogJtYmpbuXd2NknUH349T6bAvS0CfJv+R
Eu24iEazAhNYtP+xgNPgVs4p3WW0GeDjduUUiSwM6NmPjgqFKgq8TWZioQ2eQoUB7EjGAAbSeHRt
fyShCkgEh80Iih+TaksVgZ+o2xmrABzFZMb/3/zohQmQZSOdgmtefNjnqi+AXoWG15xgqnal/L3G
IaA6riCzcX7uUblzgfiPCUaakDSIz7B9lAixlmbh+xMRcTxW3J9lDLjG/XItYRrpNAq5MW3+xDw3
ZbVkw2XyU6OiHYK0mlAT2iS2IZDA1lC4Nu7b33fFQk8uyLA579EqbRuwBBzrFfQUbgoOkFCtioyt
yU3dPwISzW2DoG2Dcnv2sM8EApnEqyR2WcE76yyVsxVMUg71kg+O3Ekn9GKNDvKynavln+5IMFcE
yTOqhhinHmqeGPVVfs+EWXU/yC2fK2yC88I6tL232Nuns8sj9ffmp8EDjWyDFvTKmJFXUoVGyxhK
2JYiO6oOkkLpY4EQIRGAQ8tPf7SS7U8OoDcRu0KywEEc12wiBzHo/Xz4giZ2jqb8E3BO/4VBq+Gn
PDin+C3fOKqrOqyThSyVjkh6P9XyWb9mbE8M8Xdn4gy2LbTHLMwlV05hpEu+EWZvTG5HRhVDRdch
vPejbQG484GzN+lrIBCGIsiWaP0NswDG6IDvhmCIdxMMH0kH5bSzfPBtlTxPpReGHTDPF6DVDwph
5AgaJmZaeCZtrD8rnP/CbkIhVT5fPrmUwtpVq8QP15JobmH7QfxoEa3U+hXnLg98oleHfhxniljK
88ub8iUz9K3QSRwl6sQoJCERBIEe//k6JwQ9dVPmYGDr2BGUY9QermKKe6+e5kwW4fmxV5A9RFBA
JX4zE0XetGy7ncTusd3SElkdTkTezMH9OWHk57bdZSESruUpWBaP5CM96c+S2b0RCdZJaWqdZOmo
27D8NF7J4pjVkdebzUNhUnDi/YLXmP25xOgoFQXa/sgdM5Gnh9dj7ujN/bY4190a8vHg7IKoW/IF
I6g94nZWXmEbbLzWgpMY9juo8al8Q7Kp45HBraJZhmGmUfhN9ebOWTyvmVEkdRMd5Pgt4nT7w9xb
7LpULhVYyaKAGNB5SdjW8EEzMq3Yelmh4Q7R0B1jCWp64doYjJ1I6Tk81x44V2OzfGBoGHcFv/bU
mQnDEK4eC//tS3RwNS0edQV+ZdU+CMVVh72tPn8wGCHIZJ+8xG144r2L/UClwIXJ/PBQgtePgddY
ApPsHp3AYI9RY5b80uAbdY9yZNSYQP5/szLO22NRJ3afv0mPTL05nmQGwf/jWgKrM/RnMjGyJTi4
E81EMbcAfYwRh2EUox48Rl3G+TLS1Fjc8+YypDVYCdSZeuM4TDge+xfvR7fe7pIa5G1DMo8tZ9Ch
W5Bhtgxao7NBWDszZP+6THJ3eteeK0Eo6hZX+/T0yaUHozqgBMoGo30wZLszzEOVOQT7M8m8SPgy
ROuJ2qDYLqIZrYK4iPIlQXNF9ft+XG6/5cE07xt7+qcn03FraGJUZQI8hzfabdYgSGltfa4pFP85
mrmAIPmW4H3jr/avd+8SDJ7iR3cQU4QAZ/zl1fWri0MpelNvmfzgyAsFkHkj0sqXrC60mO+C/kgP
gNA639cl/tgcYRPbpaT24QksO8pPrkdFhz3wEvnJFWA1/u5VNCzAXFQehggc6M98BJC0EtCw1NcI
+t6uliiU0vrzyq2X8N+AlIv7IxgycfM5VUMxSYluXidP0YLKJ7wclzMpVVinXKGzk6VtVzSrGqss
4a8nhyOlGFJCKR+3+lzhHtT+bqlxzoSpTP1xvYC18plhAD0S3BIUw1LZl2ewzaKse0INDRNa+quf
Pt+hzzOthgzavKnLbdXPPvH3u7hJX+Swi2yxQskW8U09b61uwjoCQzf2MkNjGNinbgQeQyjjzSVo
MTkUIhniYSBPmaT/6kwcP6Sl8RAxB126ab5epIaJZXlZhiJKjBP+m63aKv9savvMnFXpzTo6N9Xy
2D/cx8cIpDHf6//kjqh6C+BFxXD4KyHp44XJqpsDKfhTE2hhx1XmM+3jMGqHqaBPJj1024hwMB0m
QFHcWc/esQBktlkywBUsNv7Il0n0solgpkJfCbn6B1MIL4qWUTmRNgbhleNF61Q/pYHNfBIWkxAx
a9wRClNPU0GtNUGyzbmLfpoj13HDOaKjEU+u6xTTo/1fTiDUGKDimsn1cY4bec43sWV/YVEdZcQW
hT7yLNFpCKFKpZ93ep3AjBCUBPj8u1Me5rl6aIz05/Iq8MPwcrsHVViXjBgzEUQwloEcxB/00rD0
ngjYWBm3wfGw0cBysTQaK5ic/YE9mpI3zSe46lIbXCsZgiHo/QATjmLX1fSsgqL0sv9PF0b0xVZF
qbC2BUXWyOPjl0//ut8RtBm5RLzBAWIyv4RYi4FGqhteCjyiSwRRaeX51Sxic0zswL4Emk3W4P4T
lYgITCxUtZqD5xvnn+yojmGjdSqG2CiKZJts1gknsOCk8DAW2pWEi27yGTEQU5k+l2bAeP0i5G90
GV519qai99sczq16ic1vMZK0XQoIRPGlL4OcSFOkbgY2INsa0978QeKEZFM2YaoATlB4E5spvfLk
OvIxLtAf7Zb4MnXQWmu18QDfw+7KVGK51n0YZw2Jj8XHOaNYZhNrwpsamjLdoltn2+s9Av7I8+DK
MZCiMxFlS60RninWPpFGwnQ5g2eKPrmV80S534N/4tcJAzYxjaL+ICvF3XHmHd+G3RpBdTE+OQ2Y
albjw5fajeHUx4lxx+EeIBmglB7Fuy/Zm0Vu6xGVGTnnahucYcdRcU+MfOC4KIc8XPSdIC8yNr+5
KFKpYVFK8qJ6VAWzM66UFIzhzaXaN62YrxWyKsntRALefeOAsUw4IqXPONzyoK9CzPOOm1Gl/qEp
Ax2cfmIisnChdVp3NVSJUyfSRxpPOYN96hQrRy/PjX04xL4zP600wFWzY098kokaHHDOoEVkcWPl
EvjhOzYSnAnrSNJe8zhoDIJ6wWM3mX+tkbqzZZJU0PFKBaoOf+MDLmZE0nAqJMhMDORi/YCAX9ZT
dGVSidebCUppkxkvrVByAE3kYt4lQoyOBd3vvlnCVdNMFT1wHtBygKzMmuNlmBfn9QwqZY4sc/yM
ZFr+ovLsWNvNQ3tjXyDzOBgxZs2srDRswxb0bSh0XlweXjediSuCdLofSUWUOsF6d6EaVdHqf9JC
elLWNzEiRVB6O0/HNlc6Y18VTzPZzwzajtetmwjoO/8he8Fanq9NV+ONVoHANyOguSsNh8ipNCKn
S9cC7ONJ4EXhVQ/B84kr1ElJWt8hWXzISk1PFywEHWUj2Bg6WKyl8/enIYJsrIzM2QrPloxrnZz1
iibSM57WvnWfzriH2fTDrsfXcja7mDq+ldf5+cuAjTthb2alEyKEoVy1Ol2nv1Uz79h8TLxvUmvc
g4g4PlbOim05ZVro/ZQAhBNT+fi4USFvlSNApfxz00aIlel6E6LWGrHEtwn0EkG6myKnda2+ncpK
uG25bCqrPEsGLf9EQzQwO0HZPerthsAp7/kebJfirTVdD/ZT0nZdVLtkZaYWl2UzMRINcwFamfZn
8VgBWsLPqjTOhKnrJsaZCLcEHOdhld04qbCBcqlPBKPSmNAfvxEX4eK4tqSyLwmxIZhlAH5zI/F4
G4kn3U1c24PwK2qmiojuXKy1yuNE2azb/nXiIAuFB1n+u7hfT6ph9sp/e91iWoMga+gR5Lz5XgrN
hiqx794DII2NByb98vpT2WZ8lb4xz845httYpDT66N6oJane3D/3MQLKc6pZCCccjQYFIcnqLzB1
sgXxB/7Kf8Sv6Rt8lfoVEL4rBBhchvYqwg9O+RmIQhn6u9fhk/9L8azOtFl9H927hFrYMxvja5yP
ydiSEQpNSCk+nI0mSWYAmRgu0CgBVhuJnVJ8thIccSsyM9C/ijUcYPZP2guUOdzrQXcNH20qWpF1
ERyIGUCt0RHVrwcxgu7IqzSIplOALXt2+z3TscmWIEVNfY8BIrcC0FI6rxLOgNZH3ntpLMdnmU0B
WP4jNycI1m/H9foN8tEKcBkRedvSu4YCR4rETTpJ9GzdtzlR7FS6IhyiNJ4SA4chmPqOfsJGg8Sd
EJbG9S8pvCZ5jK66YSJcE1X+R86XxqzVTOgNyy/Zv7r5UZPnGkbRpA4np3ytmY3vK8CGicTy3Kwk
j9MoEiq7yNBhZo3O2rFYWwn6t70rZT4zb2Fnu2wH7RAtA03i3SD67ujy26lGQb3n7aTi2J0EkOFI
4drtfhLZeXcHhx2mN6aLSYua7pJTztKnG73gJ00uZdxB+XkKkyMcSG2MYAXGbI/AozIhxVpy4iPu
nXUQEshNcKjVqR/amzS50RqCOF462dWhJHZM4FgZ9K20FNddckhUP4j0hfFq47HzgKa4ZyrWu8pY
hMUVOnLqvOqJd5IB88lGzUUarL4guG3UD+XYOU74++0QNGl/Pz2W5m4q08/qIqZUHsdUs8SNjgSJ
uUUBUE9zhWppyuk9xhVMlfNK2V168+j1Sbg5txvCi41a4gKServ6MtiUdZ8TU0VL1PY4vuHhzh36
t2CkqSVFnT5tura1iemUiae9yAw9IIO9svMZRHuZrRvMiQLqe68P2Ifr0z9fTfq3d9yRi7Qe5zUV
T2zB7pz9Ni3O6YI1eN/zvGUMVJzWNcpy3rA/AkaL4i+j5X927WQIDQiMxehr3C3e3osceITfz8IY
z1+OcuFdRs79q08hIupoGKKMXcf/mr8TS8fuJU+Qee3v06PmXjeZIxjLDx2IGnKXCueY3A/o4hxe
MQSLXhAQDI0+2Ar9SrBkdDxirmiHblkojWJCWnlGl8JJZdzPiPPrOz0SOO+Trp0mKm/jhsLOfGPY
x/FUIhPtD2R/d7itb7xWaJgpi3ukPsU97bc8RF783GwVByLf3KVe6IbEn35RRNZv+gwSjVLsYsrO
aFWoPWuvvI6VgyYEtnbnKOMsFSomZxZM+fjdusvHCsXuup9w6RR8xbDeYiKSbn8+hECvUV1EtueU
nQ06R0xi62jiTeMgWTzLkBu8muZD9T0rJu6zcvq2hIYBQolC8W7Hs2JlwB5gI/UAiKGyKspxOLmv
aq9YZJKT+bsarlJtShRnpkEigjHjz9+bUMQCgB61SzQm/mK5fEXAJFu27jbDEk0gnCIoF7ed/bqm
sPcj2uoP0aDlvnaiKWGWrH8mL/Yvzvg6yaR4EigIcD21gqAD0KKyuMD/+wu2sGAdbB9vfXuaIW/Z
v0eGEJcHlYPH0qklmxw1SKfiN4KjkiYiLkpZG222fmlrPNk8PKOPpWmia2d6vblIOdH/eEzTDmGD
WMuPdQETdDuGoZARl1bkx6BvHtH6ua13tcsqxdzKnGoRQKiDBeFyq3peqnbPM66hiDEgW0cGdbmj
r2tFx+RUlebJ65KGe4UH71ecvN4HN0+7JknjZ+uB05AuIukCXDshirCy4m3tGz7DaRdOqRZpm7u4
d+JedX7HIVjpxu1+T6UhjVcRDkkriM5cMQOqCIHS0y6wO9W6SdXgyw75mHibr+9b7cWYN+kIiCti
tu9dYzgxJALWt8hp23rqT7EKeOrzuhZA6FHU9q2iBRuc4LIxfg7ryHLDVgaktW0vCaGz4jPejYM5
HzMkvKCF6/P1ZjIvJvfEIOEt9Pz+5yp0P1X3OkTSOxCZ2hMNJ49XcZ+3Gywkfh+bO8h96nXhiGaw
HMHl3Er0NqMZvphxwoSZo/6EJmU+rIGXKwK/gcSLf0NFTw+lJgo150ulz332y+iQUAt5gBxtm+q0
ciopr7P1EuuxNkcurk7rUNlHFU8zFdvEfqLAjc9Wg3wUN1HYW2HCVitln6DQZrc2BYL7Iu3FqJf/
nOuppwcUlEPCwYFdyTsH4o2rPR+uPdxFceeffN82i40N0O5LaG08TOvrWNUWp5AG5uVAfmpwJLK4
McxX1WsxCFvMxo585vEhQJyQ9r9w3n9ulHrHvIrw8bjFB07mZ7KFFchTM9xpO9Pck/1l6ZkN9rMn
4LX/PZrmxQTW4SPYHyxtrDjW/lm4PejrQowB0gBziWt1dTLQQu/XUqRQrT7v8EnzYceAnoJibkZA
FtIKIiWWrbDZRSP08w3468jeG/Gd6opo/anj2Rey8nP5CL2a/cB3mUTHJBsVYX1xNmrq2f7fW37C
z3AmLU7r+FqQSakEiEys6NdZvUPPDy7cYqaJV1RwE3v/6rhTRo5i7NdxLbouRsfk9oi88pLzS119
DcizVq4TflPMKe9pzQv8LqRqhsVR3aB+41zzpyt4dnRAULDEYrQPU0/KQlfc93ZKcuzDwBOJbfc0
riEsWrQnQ68srtuL5nqgwzbSl5Zfv7ep+SOiTHQ+EVu+Zuq1OVYAa22a/LGYmoQSiY9Kpwm3/JVX
nrgUi6ji55ULTYRLMxrCZPcOa78m8Lv1I9WioB32yFbEQ4SpKp2qoBAQ40FQzTcF3roLH5iraEFQ
KD7x+6FOr8spmNOpj4NX8zzFDIpSXUacoYIdqLb+wpnxhUqcG4mOG8Hzfv+Pf5wgMCCoZxk57me5
LMpfCnwwhV19xoJQDW+CmTFIYMIaL+ji29nJtQ6nqx0Dc8OURW54Jf1dYtmqV0CzuUM5p2uujaSn
YRn6gwduv4NCscErcPCbJDh9BvfB2abhy9cDTErF+hyTTWeNJNFnV4kCL1xCec0l/2p5g3LJiJ6+
/a1tNWP1x50vXJpVQYJq7dtMIZKX9Qs195U9ttYZtN+XEQYe7evzzt7ybjr+UB2OSrVO9+QLqQ1k
IkcwWB44i7Hg/ufOVSd34hSztB30GrCH3Ihi4auzU7T6ty8/R6uoY+MO/+gXjZz7CsmfuEFpmSuw
KyhvMlDDxV6fUwba4HYh4WmmtOAmHL/H0m+dHTJC8TfqtVNgH8+JPEaO3ECvz0csZY3JirWtOxRW
QPq1omL6zQbRjjf18jLzOomSP2cbMUKy/ChQolmA7wP4ljipxLmf7mea8nFP/Z9LMzHkYlTtQpdE
7avGBYN5eag0iD4/ZQz1c4CUV1vmr8ic43udyMNr10xwZzLznaIiXACmZDGkSpPpKGEHDlIm6t9s
urm0R+5idSaMGdJ/Qnj/tDWSRNAswqKa17fNLNJ15DW+92GtDFljwIUHWNTXYpIgrb2y12xNTWhz
zTHk6ammvBGXU0vATfODBB/qQSQAUGA5yvlGeSoeUfwZZZd7cV4pnKYPwJFfTBOK7RLYTSJ5dyf5
zCMl5pxSnxMCsYW0SrVep+7A9hBDcrJdqJ1sVZHFXeIiqjg+MZ1gVO8JQziCdN25YIb/jzt/y4uh
ijrx+E1kmbGzdPaZ+DqfoHeuncyjsvQi+grUa1DrEjQd9nQ7avkhavcdICp/VjODRKrXqwgo/A2j
MYznJ9bMadMQj70O9yit7BV2BJaiFwpQiCJqCKk/qO9tPoTdNWsJmupt+zxoMHenTvJHVL9y5a8c
lcExyDHi1q+KvjhYglFInAkhyP0yhC8y5VW14bnlv4QQid8u4l+o8r1yFlgGQOjIO9ionGVkNiI+
AoTUhP95O93uK0QVSoFIJFhVMrw/AE6pWXWuNiUuhgPs1nK0RE01M41yHgJh3f+qaU8GbwDzmMZ+
dK96nzowWuMIDLCx7WguRecfOLQqJPMtgQHoR3b1jDlbgitxHUKSJ2QpcK6Apj+Uln1zmfjh8vEG
WKod/ChmXlZO7tc8R4O9G45MyIz1oWW68FjCd7kpO1/GWe33eK5pzZU4ZwVYGmKln2oOoMHBhpLA
fGey/77zno/xS15xjnCHmiXyU7Bcth+h5yZPy05ULvzpleXKfIgf05/tERim8ZvbpZ1CYaVENUwu
0L+ztoH2cII+zn1aGX99yqWSS5+iPk7EGBHor4w8y2n4qwo3LKrCR9i36hRqv0TdTpHgWHO3O3Ne
zB6B+N4mTCTkbMNROFG1K7MdaatLFTUwZijporh39Gbzy3y5FWWYwbRCzGdFta7rraSo5RvwdyaQ
KWkztGrVUCS4o3858xz7wtLlTNIfoH2tPtOa6T9UGFQg2BlLvIpCwi/hz55WGfC43lyMP8cL6ygr
sJb6DsXlSzgR4HxAtLSHaOelO7sKJqJw0943cBQ8X7wXuoREvjUEMBW1NieKUWjUhU2yJX4EyuWx
WARaNFeAtCUgHD5MQlSu5+CJMMVkK8uAOFttLvwL+TsMii155x3jWzQTRFe2hn5fLkHZcS2mGH/C
v/ocHycIS93TjL5I9Q4gLPFpbYHbMp08CQ8wGMmeXWC/0ohy/cWmhjZVQ7e6p0c/rFJAlXBhWYdW
6bFhVltC/9TmK/PyUKK0ENtIGZTMvulRSzN2haCGusU/MslqvV+TmJEp/qhSfs//WJ3LhVyBvdIq
atSpnA9gucQoKXq1kk0ilX6JGiUX6IoFaROAnT/gEq1FFX+dterw4m0fktuXlB0UaTL1GTokWHoR
siQ8HF1aidgMvpSIGy9+F0P7Swpfpvw8fHUYA4WTThZqGk4MmUxutoBI1cnZ0ZQBL0EgFGlfsBRx
Fs/fkHV6PFpvmAnQX4vBMykwKoQHHTIpxWBxyvHHRVx4kkuzT9Z7IVgYjV7mVMRmlYM/xoXUBA7x
zh03p9PB4yOwrKGEwalTloIXmDP1lk4P6VmEidj+eGdN6XKVJxHRqeI9tc5ZAqia9dreCM6UgRLA
YRubmkyssXVIUKsTs+vw8rkohoVcG3IXuO64PFwc20/5KB8LBN/XFIUcZYzrS8BjFOA8jXg82cjS
tGVfW1SBH76zZynnEnzaq8RyvhIuI3HZuGOIFkVQb5GfH3Dw67n8Twq/25S3xpBJ3YNr1VUcgnFQ
F5+hXolv0uCapCXWXBwbXSxIr0M2H/KieosOZklS5sZ80uiYgnfTmrW8JvWySGjsnhI/Yp9+RitN
4iKQKsRYWThLlEIh3xaMrAv0Vl0dHGkwwwFVmwOQWzLACazE00QDnd7OcluDq4Xi0/GxnSTF6I+H
TsbHOTvVfIsSoOV9GZBn/x0SANwWwWIAvId9IttE63dTQaJrmjbXVmRUy6R0nwGyEVuU9Z141LnK
ZlxXqTVwLJSUX0JiXngA4bGBwPl4KEzZLqAAWNWf8iDt33snI8tmUuJcjKt3jM+Kv7zlktUoVjvJ
9zZ9uN/WYISFQEGo600nTZKDenjzlQuysgApFDdED1FiSIitbdksnXhRt/0011wpYThxUAAhCYtW
PQ7Zs82Qo9F+qt6elY2eI5DPBF231f1RKntB2UYs4ZkZu4wA6Yjpw9tspJ/SyPs2924/G/vTxh2y
mHZZTRYDABcml5nc5XbZkHh4lLnNZIVJvhWF9puIqslBqay6pzdO3hBOnW8LtjC0xQlbi+jc2UgA
4Yu2Uwv/tN2qax37081Z4spfxqwqFgqaf5Tk5Cj95ERfl60fEJioIw7UeBMfQD9M1JYPDaOD6l47
jl/pyVEriEn5+IuUE5cF2wC88Y0veqagM33jX2OTvhy43g73PFlsWKwfCBHCAtCPoR7CfzjHWByL
dqMv72+bMezYiLIXkCZ1J4leEzVteSBYYkLlYeR4Lg35zocmAqzmbbJKKnDDx85YND6Lu4dgxRKe
WcUrniKVeeV+JixIP24xJCfPYeJw5TovqRLu2OUMzxso9NGdrqOZiZZPevoNIWBWLNHoxV4MNJJG
d3UYL2FN6w8wPxepn+qNwuiOU1m7h62dcypEWwRjoOZnr3rISU3LlniVzq/TPnndVNExyaU4vytZ
mIhQ/V/Hb2VMcUR9dob1yymZ/zMyrZXXWsC2u/6pWVhQ2Ugxm5DGcjstF3+vqBxrA3tMCiZZSWq/
bRapREQKxAE1B38MBgfq/+VL0K7GMK7EWwIIe9RJ7W30DxsAuQsXIbonIMEFf/6bsJfVS87wi7SW
w0NtG2QJwbyjh8jxRcdaGIz8a9neGttcpIwZfCnv9rVjkJwUEoPXIvQLVFk4LW8Siuo2GgNGMUhY
+0nghXNqrVTYQ4yj/w+O9j+l3PF82uAaSZBMtZrt0MWgY/YUmqRXETAKz4bSvvkii/LhXxC0VKw4
sbwOAm0KLiKx+0LnvYdykIP4G+cNm7bOftzBDnR9g+g56xlrpEWSv2XdNEkTupzbs7vcg7EAiCPN
GWuRH+MgyDSEHLDJrJ+JHVdy0hmHehhHGVqtY/TAP9CgRD1igzTIJidb6rWt8eRQMfWeClhi8rt2
x8TVpr1DHMes/Xkfx2NcI9ckoDbWNVowWVvDiuJvC5Uu00lzhJct5Zqx9W/pxlaGNeCQHksJCBr/
hSajf6yYDOyPbWxLKVzqrgvnZvDQhhTKcoCiBqsUgqvyhmRlMcVtr+kwAaFFZF/I3OnebGyuWhxJ
ArzdI7K6Dn/vpkqRJzFUamP1K/zvuhOI0z1ZJVSj+C7yA8xJ0JVqrEbq71kP4O7QKSRzwqh5D3+V
p2r87t8OQSkYEGJcAPLdm5WWjRA5nU3au1sdU3hqQZKOBqIGBBPIBUc8eVkfnVjHwEG8WNMFVHzO
nQMFY0pX4ITBXi1r2RjMNqxfbTv4xb16e9abiJihORF/3VlIa7vU3kMop/haVwd5ZP3puKGrkYfE
+KdYKBGcH5Fuv4sTBsQuhulniz91WFPLTOp5I1HXHZFPAJIi947hyxh5tFZhE1i2MBhxAWiF693h
zdTpp47dS8oV7dhTLneg2TctlAlMUTEosYcegzlGxoW9reX6VvOizTmvGQLnQ6Lr3l9ZxS0/uoO3
HZTJBnFojudHVax23CYrlyLpMUzvm+1NpR8zbhjJpc6sQYpI8seCfdeKCP4f/oyGb4+v69kozyrS
q9bVcCpLy4y0UsnsvvJKHbAyOIXy5mgcrsV85B8AxLbnxmQ0vtOFQVE8ZU4bQwRqQBsVnVwFsVcJ
GGLxX6yCKFavu6173sELpvcHwRNjoTRLoRcesPRH91ad1H/tI/H5NDJ3AlnRyLKggQnHWhy6veDC
q96pYI5zn7Uj3CUpVXP1VgD27p3ptz3wZtJTDy7MPUwJ6lUPky/+g+eZrmkDh1mW9hqDeHOEhN1V
QPK8xt/5rwJSprx+w+3g4toGGS1ZPFVMZtCCNBjCYdKLwJ8teSk1viGjO1quHg8etbhpVH+ojMyj
Sa3qk8tjp5cAEon7bPBp12BwY4CTFmpGDF/pMithZ8nfWl2fTZVYATHBQHoiGl3QpXXJWSDws1a2
5eItbxVPtd5NpMvfzubwDs382D5y06BbyKu0NCRrZKYGesoOdhpM8/imuxiTBh4VtVIhjvG+/iqY
3H/EzijG/Ja57sMwPFEYyatjXnsHGXf03tUfPSFOu8Rw3aDk1XoErZOz/9felGaX7NUZpf8h3lgP
hGMd1E5aWg2yWAY1NlwqevR5upxonA0XZ0almxGQbwL4DSuLBLgSSD94YupeivVK5PYiKG18SaSo
XOPDODUKoJ69Ny7SwFwcRg3dmXPsvkxGjH9vmtyADCrhk0yvDuu8JcjOgkR13n8KZNw6cXKvAGhg
BGeUBc6Qb73YKM5RFTtAc5OpstnadQwhQYrT6P+yGqgsO7P/qxE32Hssn3jyOc2JGgIO6palP+UQ
C3Lr+R1gvv5G0w2uE4naw7VwZc+HJIXEBwQk809Rcxq461EHUDros36JTDqI/vNn7SVcNqXZsM4c
MSZLTzcffOpy2B8Nb1rQOVW8JGzIgPoFVpLERXCY+Ba+MHZihQZWUN07bzW0iFIc2a2VkDeqj8Gq
+AAiQPL6ynmnBKZWNSP1xy14WwuQVV8KRkop7H2jZNf8Yhx/7SFH2v5HNjGviKxJ5y0nxpik50Bk
jMgX5yyk5rPV6JmP0ZRzB8PX4E2bePvqHRGUF43qDseigU0OErAYXt1yQRf+nBz1r9fjPW48tf4i
x1eLyI4IrQr9+HZz8pwM4GE07zea6qMr990WZ6tMsCvkX3BGHVlV7Qto1XQ8BK8dqYAe32IgLpNV
rPyYWvadLIMjc22sbH3yfCWtE8QcJfJ+2Hln+Dj4vW0A6mmMmmPPmMQ0WuMHUeDcdx//UhktlAXN
QT9XQ+2OBFHeYOcQeCh3SabJv9+V2QbFeSNA/2mSNgUT+IcHHC67quH2ABzgKiciCTr9OrTbvijG
t/CL0WcRlwKRQpLJhkuOgc1vlykrF1xR+YIpHaCCqkF56Op6o6+9yLFzgpBsm8sZIqR42yyuub+e
J7GIGJVGO8mcr+51Q7uJtTgZE1S9pI7P4rI3O75dVT7icrVozrgFJMquGD/QLV9c6lr/U2cOQr1f
77Qg5tPfYVuaPMFyWTatL1PDeX84w2GniJd+bzeUEJx8v2xl2ZbARGHB9+cO1v5XXMUo/b3e19fj
ZvfiFJO9vUIWz6iUv5tlpPHVMaT1Azqa/zteYrTZ/tVsoChP/owmnEPHuS4hzNZ2u6A9qJsBc105
l/VK3XSOnkv+GjM8FcNNonHVKLBZ8Qz1uvoAdHAXG/Nqkqu67f4zesL+1Qgfcdzu7Fswo35NvtQJ
PPuEp5b2+rqMmJrAINzuc/G+yLlg5PE9n/XBpljaJGb9bMPh+CvBra8maF4bqor9p2+ILJOcALEL
GU1CjvhTPMzFhZm6bD/zz5X6ScvxPEbCKDjlsi5we47xwcdZQhIXClGYo8TQC21Me1jbLWSqQIwv
Yds4czrlUfeNmV/kkavTfn+j7gpgDIn+AWjCws0btudXvJ+CsPBwD6L8M9CkFz0ElB5lZ3K0g7/7
pP+C2RNJYjU//keFuJBPTyuqGN+Z7/rF9JB3u2LR7qf9O8KdvKPlTMOXL7ZIqVvVlzN3a9Yjf+w3
eu2Hk96cOqP7vNWY3vFPt+7QefSKFg0kA+rHQc47WksW0DPpn7LcB4LG0FQ/1isjSvPo2APZASb3
XbiM0xcKRmuRZypc74lZFSOtdEWoyN+ld4ChpgkcIcGPlMxuwcdXy1gbcbi+DTbs17YjS8zlniDN
byt77NkyJ8QNCd1bjwiGND/hly8NA/6IUBD9Ux2wJZDx11VW/OmU4haSWxakrWDVOmwX6tDlriNa
oFKiwug2XNh4iIR86AU5yiB9U50UJLv+YsjOfTx6FIvQdDjFijZzKZWaIyuW6VDOOD0lNYYIbenZ
JOWyVclEpLmu/6IojoAijs49TMKCdGhgwj9IGZaXZEye7HpuCRSQmmyk4EEGZDNdkgZD//E9rqLV
hh1Vc6rfhxHNVh6fp1/Dznc/KsFVVHo+I3YI/B6tn5Mgy5A1EqkBFFK+Fr/MJdjMOmwMUzxBir9h
MrCX42sxqRbA9Xb/XSMNx+F6yoPyml1aj8VS+1l3Xr4vZagg12tgENVT2/x6j2f+f/IrafIbMMrX
HDlnCO7u/FGIH+x1kRszce1jP7mqo6F2nYsfAeyP6xoi7Z9CDevBx7Y3h7Fp/ymwiFe0P0oi64m3
xL4BM235nwVwFdwFqNqJxbBsWf1Un6rZGzBeA3e01Tpg7btQ8XT5+G1rfXx1lzdPJyRIr34gq7BW
KxmMvds/IIClzXy9XhdUsXBCPYUy84IBkf3fi5NEFldGih+bzg94SlzR8sCMV4NFPBBejDancn4L
yNLyI/9DNPSoRPoBhWpNV/G+5MS75zZwhmIa+CvEMfg1kn1uLkhtfICTcgV6Gx1wyQYefTGoJ3HR
C93RcitJDgJf6Uxu3u6FNJoCL5uRdBFDdZN1sTZLLPARJoNzZI1v/h8KHdjD9ugwiwBaNdbMA0+y
4CMdU3HvNZOF/yMLbvzxgZDTeU0okCHe6CVfnw7k9t3AaerPGmJAfhjDAXp2QCSReNwe+9gRwK0L
pbafDSJPzKXGEdlb2u5qJpSm5S0NeYZrpy4jWoeM/TOL6JSht440J/u0XKm4r3QWvRKBhj7lbSAO
f6KWK1CxTRXAVMPZ9UPVc8R9rtIarwaIZ4k7uru7JsPcb2TW2VlJtREwN9zxw5Af1vD97o/ztI7f
KyQjpCymbl3PeZzDuW9uwp9KUY0ITVDxbmFxB33qSvBmTZ5So2r9aiVzpbHbHn1RuMSrcnSFg06c
yRTfzsQQTazUKwWW5yYOux3Nx+Fu1RO9tty+sYzcaRJNy3PQdpSNKK7SUSIg2zFKNoMZbXj97yv4
TZeXENBlAtW0apdWR5y3GBYkpMXuz17daaHEAXdzhhLOC2SsLAVLLlZEqtaRmgwwiLDoP0fACpeK
ZP8+PARLqXtSWMIQjcVVQEe6uTdITuYGd/SGnOe+h4pT94/Q1ZLtU5ToJn6mwGRrlIlHab+LWuHg
/0gwzt+a4yr8svwh2uUNXldCaIYGwcqZ5Hzx+anE6lG35btcJaoysgc2PI1iMQn4QN1w080wsapk
d1LGNmCObraK3qNRDGT13Q36BWVq4BXVsL032mhQwGblsQRk+Cm5vANBGMu9fh6VUlJoxDLEwpqG
aVS53CSzGwaPJDK1JnDa1wFI10T2R1EH64KCL5M7ZWrtMFzdkkzPFDpvJcOOhaivQARuikSeOvo6
uAKl7VcRi2Jxno84A7kJVooxRa+WW/jMtsZ8zUuBUEHxPxHkSpw7fw2Kr+Qedm19O9D3NTUlyijJ
CjzgKss+uvVske8/Qp6rv8fX5PGm2Bm4TWpB3HRRf+4vbZQHYyGZh5+kmZc4CWZhM2526rY0m7dU
mswXgvVggXYtoSiO4VRjQEuZWsTuh6aADrZhw4sjc74Jd7dWMjnv8xe4r/MDKPf7ojheLfxWkJ4v
Zdg3sz1w8eAftJpIsW5JPkFjRCqmr+ZqlUgnlZQFb7acR2fdKxKN3I7i/yf3X116gvk3QiCy3zKm
fSt99vtKpyj97eOoqrFBj7H6OmMfyKiEN3llBRi+tLYWk0nCEZLg2UFNtrn9Tao32jjRXI9Kxer8
V2qQxhnm1QE60a6hCaZjHsL7Qoe+xco80O9fKfJP+X0XGyBgwgcfeQvib9wgb8QO55fHaFgsbKck
vcPXHkbA37GnU3h6edkHprwbApTPkv4/nK747aagkeA+NkY2350XgVrRCtpKsnwEL+Tw7PBw5fp1
An91IiZcPSUEm0ts12UCS4aM4kc0cStwZVRM0zfI+qI6Gf6jY6Jdc3A8Bk2IFyJXh+yO4it2R0oS
snlz5nPNOQb+iY2IsW3yhTMrogqZytagkwAoKM+kA3msEb2Y7eYj/GpD3qoFVqJwweKeoJEsqXkE
N+0BOtLc8hO2COuO9VuKk0B6HyPPQOin6eqHE3JtVWioHySL3Kn27/mjI3hZYgofvgexi03pgfNt
jf1p2rJac1Gl3WQv9yeFeqLMiETV2ZeRlhlClgHM7Bj/xmQFKgz8INQLButRwz7QeGd5lMBGN9Ef
QUrpKb+QeedsCZIl1BSce2cX0ARFdhnGIIo/1tX4+EaLchImqWFajKFqXBionD7R5ss8QxIr0J2A
9wXpvN5XsrCb3SMBtuS5nLLlk5BwMxJ/+9P2zVqVDxoEgACFzFyvXXHYiOHkmEotgizLEugrHRWh
+zDTQWa4ghEU5lSMeDYi40i7VhLFeE3l9pGIb38pKABv2Qy7IJRfyzADjRWEo2r7OvxrXWcu0IXq
iNlt8i6ym0jpb3/p8G9ndeNwwKtaIpygJRpZPgVQe/uwBQ2s9MpyGIlpi38EVUpKVxo9I/vz57WP
KJLvplflFCY4KvPp5BF2HPExdEgfpR+nIxaRDk6rM4k0vvo2uQR/gHun4KAneMbXjV0McTdrX5Lb
8/wsuhBCuqgdUDyKluk1bdJKKF8fpOypN05VV3IvFZFh3c9H4lHvY9sLkCfTVRoFlHrir0sVWEiJ
E+jpAOdZ6pU0CyAXQtKBtvdO4/qJhEOxlrv/nDFVaGD1UDyerTPpR7ejHQLbMLXYIBzuroSjkUtq
cR1uC5xxTtxXEpt+aaPtRW3wfimuA9tauKcDAjYw6CbNuxYdKjusK8GT7jOEiOb6Pqa/2OGC2T9r
zp8aHn6UXZhyTwhFnKbhLu59qZF1znXGO+yLHZw7NGzpOaWx8M1RynEn7AbPDzcCyt1W6RAREP+X
i/E4Ul0oYwvC7ofhLytjyp9miSo2KwYGk2Cf72+nmfqoxtgaw9H66QC0AaenPA0PvewhY1rB4/GL
Xf1jpGung2dFE3lf+HST1GD2epWTBp46wr9PwzUFj2flwFl2xpbvTm46VhSbVLVkc1F5gv0UpKnf
1CqSmcI0Gdc1umTnLvBUtAJbyT8zWAeti1SQVg2A15aKUb4irSeO5NeG0i9xXN2zEs/9vhx5bw1f
jJhWUdrCMZAyCphOLouUT2VgVBTWQSNOhu/uJSZN9j9Pz5+Ce+288iOoxynfwtDBFWTdZJCLFL09
nTU2Xj/L2n5HjwfXjV6IHwCmKgc0Buj6PYTIf6kabXGtDunj+aY1x0ZklBasHOEGidYl58EeA7ft
Yh69IPhtIx44WToTgvrRQPLv80d5kVDDllexb6lmY3h9D3UadHQKyY7YUEoOYk3KxLlXbD7eXkS8
r/VTz73/iMaxKqq5XR1PFJ5N+CIu9X5EZfZqO8PBEyuKMxajb4vgCUMzNnLMcI3Xodoxx2y19zOw
KTg2JC3xfSlpIRsZTHNHVUtdyQ+H4e2tJpZVTMLg9OD7iNul0eQp4XoooVVvVoDXfKcZLafzxK0u
G/+m126t0/5rDEoO2TCP18bE/X7ihDglmojuod5yPTNeMdrMx0TKzIswTFNlNFzkS6TcXaJwaptL
IIpc5Wwyrgf63x9p/FpdfNUp4XXF8MgtZhChuz3d65ctUMvg6U8VZkfWYBswXhKoFkqJaDGqqGBX
IeVK1OBmvpnNWy+sJY3R5Bv0U+9DY7HxQH1YfbjYnAinMsIBRjvyGTYVlLsf0bq1+uK2frQnsXgs
qTR4ZdYcyYChdI/MCfzYW2DVUHZm4+h1Zex7bZvT0C2hG7vOj2foo/RiX53zsxNvy62QK8hNTLcT
6WvVl3omQ2oCZmZyutfV3cNOb5RgopwhJBd4j09jKmm6YVoejaZIb2V9c91n9cbpn9gVr8ZXO4mR
ZTlJLH95Q71q075aExTMh8t3T0uYtdy4xl0mzZkzsAN/ruhUwu9Dhht/6nyho+tL9Ae5DMXNaShy
yjgl4zVtrwFi52IevIqMAJZeHRnvdzhBxNfnIULtyjZJHT8jkbOe7bZUL3gVyXak3i0JRzQ0NMrd
vaHPHCjeUqA1bxt9hJeL29wANBoXnMsTVn0yCGAJjOGPD5Im42MpZU2RAKvEv6gPy4G27MA0faUi
WBMKkk1Ws3VMgyvIGsETRX8q0Armfp2gMAqkfKQEcNSz1djqKJwMoCgkofSqfQH2UXtf/tWG1cKm
UnxXO45VzIFhyXFkq25rUzQ5FbR5HtCiHbG3Pn+USlPJen01lUczY/hM8CVmA0o+r1kGvS7luSBz
fqY7jFXBFfvTxk9icZn8/rg11Zjib0cCaIMu/XLn7d82K6S6YleXNz05DH4LyvZuEBB3FaIeFhkl
mVrNV6wsyzJQ1kYgSryeYrzkeXQGE4NZvTJ3bBFZ3CWLe4SSxngvcialUKy+kZdWZYRWZOaHVFvH
azNImbI0oH30BjjFaIHZNA2Vd9/2zNQY3b0/lNmh+ZBMUBjHx7WuHu5Z0qQF5/Gg29kxG766gvHv
INEGOiID/KB5Jo2fseGGFJbepw/3YrtupAKuZdZpN5sUvDH5U0xa9Z95AUiMxtTSEq+RNVJKeYNl
DIs0aF9lBBKNr0JWa+3YyGYc/cTmdFHP21wJW5/+m5bnbVVmicGD8d7R6QjbHR9sYM3yAMeV9QKK
XFRxE7evaxJfWiUhYofxsVTbi/uFf1qmuC1sv/7+alkgsABw0nEa/uPOtYdDLY2A5m7J/FZSFJpM
AevonCPkM4I7nH6V3l6n+qNM4ksSb/nKr5Yg/em88pm8IAkuFJ9urLRXV/bpAJ8j+xa/BIyvoDr6
kD97tTrXK2Lq2G/lJZqNhh+P915+ZsJC+tOFbKusINWjQeDnI0dAp2a6TjgiwBZPVJmzPE2cflu2
z591pjNQe0U/VgUAy2uJfWfRuacISmI+gVrnZJdHbqtWEGEaHAQ1StSIQHVDKJcPrk8Na1K5VTQu
JKp+U7ylhDX/Sj/TjV+Yxkzt2n9sgNPXHXoZs221uWamY2NPkJ+S/xJ6JErtER6+EEzJ884+EAln
jANM2Yk7KsCwkdF4N7i4leEmrpRsqcRCCh/496sbGpw5QYJ05nmw7ETB11VV4Jseij/3DzWennij
t39oB390HOyWnX0G3Br5+TUivEd1a68fzwWJiLVDPUHquuV59TZcYRjbq7OB78glsppm6RqW67n2
UCtD71w4nbQYDVL1Y9ZFBqVy2cgHG9u62cGIsoPRvhuBNyMqsSsPluInLOygwq7bWhh0ZaPK2ELC
dMSsLpJHq4BwvV+iq9XGrcl4XByOgxco/GaM1YAQHfDoHgWbq4ufPKYFKzNd7LsbAvo98L/KW9NN
fw6ZPC5sWYNptSX/D8KIik4FO1Yc8QXzmT75U0wqgIttCAvpun9CB9D2UN7OTUyy09JTkJlit50E
JCaTINWg86BovYSo4kC5YZMn9jYhahBkcf/Xe3jUjINJOw6a25imidvMW+Zh14xqjUcQSA+IjdsT
h1q6xK/klVS59AzcCzmVge2ZbwrS7RUPSvdI5mG2BFzDxVMHjQ2MJN6GbuMFYfBPkSCm1kYcddi9
ilLwhVlwVIGFOrjuSjAOMru+UBjZB8keTTwLorVBMOz7uRzvrKksRjL7maOom8zXlgL/cvM/L+Mi
S2zelxbymmgtkXBZnSYN4DySMUExUFzyiEILr/yE1mvHG69m9Ka3+U7hvQp7ewcI3XcVNjqDExbI
8vFj6EMHkXii7MXuxW88zfHhQOVqWwd/WAy8jHU3NzN0Yngl14T/P6b/iSyT9b+Q+a6A7Ms3Jmnt
9jvhoVf1zRgVQ6Iyd7v7amz0806HsEY2N95ulJHFbywNjbGWXCP7vaFqQIIofbHbqAtJmInV8OEA
M33MQexEgLMc1M802w9huclCdZvB53s8BSIksBClM8hjV4c9iTlG9tXG0cZd+t+ma9smtZm2/yLf
DySpU9iepT8Ds6mnudyt0TVDi0rXFyMYiGyNr4OUcS4BRSwuxExXKDwj6sLh7mMQM0hkUHEbKJeQ
AfMutxWCsZOFwcATx2lZfopn0dAyLprAIqKNU0da86CoJhXuYMWYtu9i02UdzCG8gJi6/ERrq9TL
caSQvr0du9fTmjVMd1JTKpo6Bn5ef1dA2CxXjgfuwD81u6bmqqRZm6rgzAgeeeE6a2Xs7+O/3ziv
AaETYphZ+7wGNtER9fPMJdCZZQQxifXAn2lQTsvddg9ZkCeyW1l4KqEbF2mgvxDJZ6PCIa/Ke7yS
pAMcWLMoLr1UHJRw634KK5qtQRP2ah+P1HDNWMUnReFS2WEWANn0MaMeTjPYyzbmhkagDuH/zUpN
yh4y1qzGBye/U8zf2rhG9j+RoMKbOis7ZGVSt7DjPr3uPeELbGmEujCKEZoJYCr5AIsYmAg8ClGs
dywE+J/QO4EG9vrLQg+0tqp48wxkryzWfTN/zvs1YvfV0HjubxhDgI+Qx99JY55umR3iFccNGTtE
Us8WY2zeE8muffwqxN4pLM6OsW3gRMyvAMcx71owmBiqb54+evuQSo7NNFb3K74zKnfeZGVnVgSS
TgqE6+wsiRn42KD3k0IHhgPVUXUu3bK/qBIaHfNBM9hNWPiVFmtOkXlWCXPLaPKrYqDQa5CWUPUu
I7017nsSbbYBFVXkyoIE4IxAYvTrh7UIDnnndpZD6wRt8NfWr5s1Ip3aiFkW/5dsBg/qFW48+dIi
/eAIkRN767ISCnTjXCtCb/oRZ4p8zdkabu0VQAQD/Un0YthBxZPZ+rep0vuL/ZK23QzmB9FY673B
Zq66d4bjJkfZ7JhYJuS19QgFNzNdZFs0wm99f8kgZw96i4ylKC9ZCu6MLVewBMA4HmFLDsDVYjQG
jbVDBqe9hyWOKQYwhUlsjqDMhqHMbx+mfMCdkWskJkShwIkntS8hMjd4mN8cW61e+GDFdAJY6oym
HcSURIxmWgskfBwdhfdarIjfTiRhfVvBZdPS+um0j+YhKrvuKzRX2VBHpxfcCGVIXZAIwX9OlRdT
y9RAdgwvifa3s/YdRgpQDHOXg/9EbcriYLKgRY/CZQVLmRzRn1U5KK9ZqXo4onF5/lPRfZcgWBmk
YNPdlngdsRA72kBv/E8wKvs4An/XxXTWPcpKr4xQEZ1Q8rhEcxidO/aGwfFg1eecQaKmj3bYfonV
h5NhoTATMp22fD7Bbr7Skz8f2Y0edMYvHAjSieuLZJPzqoD+X1VJ9ElaBNGYbFDcAxlDMSxuaau6
HD4yNS9Ew/3pKzmJ/eQcLxd+YYb4eEzxST0Rgs9DeeeIy3recNV9g/oHsUfNbXZxcuT5s+kPP8cI
8IwXgSvyP/IkvFrIS4uyRPeYvOYiQDoYM3vD4WX9c3T/d0Si2uq9gJqDDnDQNviqBu65dSm1Qa8h
MLj6wBoyjfu1vJ5ex9HP3e9iCmK0Q1eQQwhMzGNeBhA8oo/V3pTm6NmloYHPOkY1pTDxYetFexmg
vCeDavDGVCsOLTQNWUStfypiGLrxu7qLjAwCdvFsSLlDXHKG1Vw7GSprQU5qwfbzwIn/VqTOHExL
oN6zTTFxt+tkYqIkiws2GiCbJzdCC2H6ffdiJZxUP80c6s8RC3GNFmCct7+J83BaPtYuL56w3FX9
vBbZDlmp0cxOJp5n/+TSrDm60EZETi2EszwaMTuCwJ0lIbHWbAkVQ8xChZeATFvp7iAL/Jo7/ZgI
m3lK9UlqqjHEEesEKZpkao0Z13pAdTSiT96WQvBioP6SeVPTv02lYFXr7F9aQw1TqptCh79rV3zd
mxFQup7gPmu9jlxEDKW98iICzm/6UliCGAcJjR1oj/BxjD+cl5vbURBRHSUCKzSZ63MKtx/VHXor
rVIQpr2jScZXkrBKJTQpCkjNVrTZxd9R4b1mAtBYkpK6pXJWXZREb4/FMK15ng31OntNGOyRtbbW
jXeINXByqeldtjhbxp2PKsUf+SNQELF2XiRKDPs8oy3SmkQlnZ/+SPGXEqXaPwOnF0QUDm2vM9tY
HTk1Pxoz1hBEO4FpdjlKDCejHvWy2QG58bdHV8Ufgx7+9/8B/3LxogX3VvXm8VY9ccIbC9SZ4Mzt
Hih/vd4Om7VO6C8iONZRGNKbZIagmGEyfkmx3IcqqoaddjOrnLLTgg6h821EJFmLwCBg8cN14KZQ
O8lOBjrc6cJKkEhuFos65vZ8IjOb0YRo2uVA4oH7Jo9BVo0XZReUoLK5/R+kuxGZhq0oI3uejBEJ
UBX8DLtDXwidMTh9SsZ4uqG3c3G1FBaE2RNaADpDfInxFGbd91n0/0GJJCmY0Fsx2YeUYIP46dLE
zbQTWHS9NzOM9mEztvtJQDYNr+p4lj7S/IbmusgQzdhHEArdB8GvSODewkdYXNQLMe80zvtq01db
F7UMuIO/hSlrTjE77wW2spoNlAz8tRpEDDswJBj4DZSyquvTmCYegGoZ8P+NKPaXGJ6g38jpqfUX
x0hHCemqbRGZnJkcUYa/FRxSg9YJX+w1VyK/MoQFqLP3hxjMY1IwP+iMDl1KIbRrg44dbs8HYsyN
DLOAtwAT3zG2UVGGvCcaNtYlcQRVpVeo/JelMjt21D4hXp6qkS0znJJ+YyFblrZo7O9W87bTT4Zr
I9pLCJtcuTyWIBU1hjhvQ6Hhu6AxI84qTBwm/5ZkwWMIcOxLDqcrAR9ViqbZR/LpBACregabHVVy
VIEz6jxyyK8fRukCfsPp2np9hPsgoz0/8QlNDHvGYBSCSuYwHgcJPYNMDPuCEyTa7u9Dvjl5Le+2
EHgx2ev0cf441OlYlPnv7dCPvMe7/aQFQDeoF/eUE8yYNe7xVZlWFJqNpdb8A1MUoyMdEJdghBnL
/OooV9ZHudXXnIUUlEhqpIiR5yQ1DopnXonMbHH7sxvRDkIlq1C6N7IP2guvq2STiLSkT9pj93LP
5dIjdUJF7ijfPbGcqLKjqHqQ25JGE1JICOe3Jb6ov7I1zOn1topZht25MeSSPxJEfIQ5AmvDO0G0
AXUqzr9UtfTlq6OqZaRFZ/dfSOqx+vFQD6H5NRSq1IGLRbgGjvsmlSuSWLBPYihS/5ab3TQmRuxX
04E1Cy9ymfflWoR4CJlIMbi9kCKU+226fEkDx+l5TAmSrmHqKlW83efCdfAXsmzF1/70wQ1OaALm
I+HTYsCK0JCNWTnfplNuObdj5yVrQ2dwdsbKsLJfz5wJACNuvQuZmPBP5OFlZgnk8vcVCE//f944
+s+GyXJHs1A96gj6t7e6EhaBejgKqcWUp7WSn7oJKYs+ENj5P6sfw5T9FbXXo9u7QAgqeM4FA8Ik
7kMALZPwflvIEBaCRs1GPtFIivpwG0xOWBhYkvk94g+ff2yV+vq8vv0rD+wLaegsqTLVsToPzRgN
mnPWNEbrg6YXJyBc5eNXqU9I+hYzRxYU999QKO9UG0854C9r5mbCxLxk5qS1nl68jf9hcnWiTtKX
4VkZa0XXckShail6EeVDjvXJ4FpOlQnyBHT9vgIcee6BhHiz0j66CoH9DDwPDXwkpWfL1Sm2bxPQ
eG3sWXMnQaIcNk/Z3UaXpLx+ZPXOhYIjrdnTgT5uerZzAplieJB4MDB49l6Wgyer4zimOMDQ9QQp
+fn1nmQuqlys5FsSzneGTL3/5DpFlnt9F6la28CTTRu71H9LMXyuZwj36xk5fOocKdJ8uGvqcjJF
phv5TbjoJF3CKPW7i8Skw8MGCXB7MWC0R4Lh0ovVSmSJQfbKjft1BhGxUw3wFcVePW2yTVOM8alL
bzKh1OGJilL+TA+fGzvtC2S3NoEJ41bHo+72ksoIsebFxdEh+915GPFgOhgM9WItsG/7rthWWFpG
mBnhMf3gQVEE9HcYKa2sY3IZEL86MDRlh3QcmVdelaingltkA+7eGoXQ7VxTKp138SkKl1GHEsoi
LKcETAlbkm2Ruc3+rqZwcRKPqTViDCtJPgr0oTwKY2je+3+nE3AQX1g35utD4r9g1ZqpaKTAdAjE
ir+aIN+tY4ORRiIr4nAtbs4+m1yD/XPeStBj14TC/I+fJCAyH7I20YXukkZ3uutw8+YOI1PLHsuT
GGFfMoz2RyhrOV9wNxIi5zzfFkUTTTCfPB+sVK6zg4uOlJH7zvpe6GQZrth00TmmOk1iSssSfKZI
UcGFHMuSVvPqA+kZCujCvDBVa0yO7PbeEhEORKCDoC6//xXHqvtGswxP+/obdNVxPo4U8zFmg46d
cqh0do1Ja35fzNW2SJlFkohowVqCEsgCOW7XpytXGyfLfAuf5VEFlFGJ8IheEpNiksirJXymbMfT
ttT+9SNXReiLvGnz8tsdxNQhkZ/Xn5PNMFrDRBg8ixlSCNlmkJ9XgffoY7orQXhYbvzC7vO1Lv9C
+48RJ5GFFzBwU7zqzjEGvs01SJhEnoqzP5M8WqvJmkCHTlzuW1lxaQUNGVobOHVkPfQMam8N7F4H
iLxfb6oBS7aQBpNet5PFkbrbMlbEmadD/FujmPm8ydrVbtmRAgODf6wv/g4n/6kSTcvKTkKjldCb
lOw2Hi0sw9KWOMfE1674W/wRLFO/+owqifB5boNUVf8GtyAUWfOmWIIrpIZ2T3qQki7wFmaAa6Kq
2bCVA+15Ir56f4dANzBRMboD6oUsdij6Pcn+8l2B902eOyTsfiycGDtgoS0JLQT6uub5Sgj7592E
O+R6+CwR91jNNz6uLrb+wkdwfVQAoy2mxCZhY3gQVaQVnDQt/YGW4ZJKatTeG5KRLAlUV0DFJKKB
RS71iHf4/hNQUBdOHzkYy6xY3gwQlPSdK1Jod/GMJgK0hTYf1BOE90euaXmcsY91Ix6qb01AoNA9
RbFCvnbd0zpcwFazX1tMvim3HURYLuEE9Qiw1eq+c6nGayK8Ca0NRVyefyUW3U3gFHM0ouSCtdKn
6wGHLhGK+K9vCItqAOCDbjvmw9dlA64IFnwUJBqhnRfD4F+6DKrRxUwwl79LnqGReVczNGpcFeXq
nUKUg4eTU3D4XpicxcQjSMCBEcwdhA8+U3p0NgSaisP/w3TNiuDNrtP5m33PZNtw+bKrgQ3WPKMW
gxz7G1q5+QVIN/RYHvjdfCTWM0BrY7ssMy961dvsnSOnH8AUJGyMQb1RTGco6yMQBlPFr1lhV/Bv
GevqgQwB9vdbB/0shTvQyKa1lvZ2VwD79qibZXXBltXXonz/4AWeyEvcBPGhXndLJaE9WLptA0y8
dP4JteZ9v8XIRyeeYIon1IKdX4ToA2w/eBlzXXmGkpEJu9/zfb8eUWhx0eADfCgNDnJpbGthnTr/
pjC8PjTv0xvPXt18v0B1SMd9k36NkBTmj+CugWyyOJk4j6W8OgUaqWflPLcN1rhYY4hbkOhNOIAo
C1aungtOCzsUEMipvz9uBWr5LpEeuzrkz5xhhNCWjJInUB59/w2FUCSPAEm6ct1wjSUr+bsBlNES
BPKvZbY39y0724N115nJSCrhgcq1y6KK/lCknpmDEmuSXd8XvaId8PjVF5QCXSSsd4FfFa6/MblJ
6phQxOQF5nOiHgqpUuRogLKnDi4UB8BYJlPRVhG8gwkslpak55ZvnioBdZUZyr1AnZ5ME2eySpSb
1Mptp5Olw2x5RRBO3fqLXyOc5wfkVBE2Fg0lhRjWDOcDOUTpxMfio45cBYaQwf8UnBblNvz03sp1
3KBPLQ0MJctvAyd4tNHiZ3QgR9EyiNqKxpX1SO5zCni5taSA8jkdhqwrtKSsWoJrD2adCGr91Hyv
Twh6f7LiTD7iBS0M7z0bCj8TUwFUtJ54Sw81E9J+xI4HmhK/ffXWU8n2ghXQiyLoLW1jr9T2jHWg
1YPJ/e/k/u+aHVTwOobOabiB2cJhqNoKqlFNiY2ZVnKZyILIs+i1fx9Ku8jXrawSoA1K/OIc0JmG
xZ2Kw69jgjiHBUaYlGRRUw5t4zDkftHPR/Q6fgIkgtMkQKnDW4Le+Z6549qexm3x9lq/npi3vwnP
lloMGvn569KB2JuHq3s6coIotTBWdHi+/cEKtJX+uPzfPgIjZadrNF2wxE0oU6DI9ODVctWOaPkK
KnncT1Xtr4iyfU29Wf2hDSOKmySDNoy1pKL4Wxm19FeXUi0ZGVwu5pUGA41+3nB9i+/4j1H6v9p4
GcgrXEa4o0643qpwMPcqF16D/FNBnoCZ8Yu54aLMYc9YHOokVRrt04kYAVzo5v4/1kuVy9uyCU1A
4wtcAlfqZDUbUfH7SITbiq5XaRofV7YtoPGKplPp5MknlzINRMXNUvei48940g/Utr/g6TA7pHvc
+V4JW+mUR0JB13d5x9qaylVzSy7BbQG5YvSFAmGHG4m5OtXcZtd04AIIV/BvBMSxJN2H5X+yKwMU
f7OZsCRMH5SUkVzZEV9/RFX+3dv5GGPdVDEvdmIekh1P+cXdzX/uAzGybAwNZY8TvKBoF+B6qCh3
76qnvF7HDFMXN6ue2eNFai4VQ4p9IjDKKfSxRNkPzozjRQC0LHZWH7sKiJzBeIVhWFQdTJ35wCSd
UNIszEp/UBY59a3lcH5+mDVbwtLgwZadIVpQKzuh4dLAaRODbQoQnnhU8zLyCDnRIODgstl3rrjM
QmNcwIrf9H9L96PPwoVnXDGj0sS7pj8abzV9M+PGobcoAmUqG9ia0RIYhfok7rqnLolY6TQOewt0
kTVHjgccfyzj4Ma+ZbOYARBn8vIo7/CyWi5IUJo+pu2CuMqKA03Zh+z17Eo15Yfvt6viHbmhkY4b
Fb5Xn0Rs8wisteEzoEY9LPl3DUhxw1tCHHnJnNHCQX+cgTryEKvrJlkhxFF/PiPmfZMUa0qAz5FE
HSnL/HPBBu3M897qKcN/XmN5QeeFgUfHm9YpDS8EAPnoT0ZmqS4nmTehAfgGUttRWOrkapVQr11i
FkwiickdMcaj4p3NPn+R5HtRov++mdGE8RZRVqxSgPSIf1GcoYkrAcwTVPrID+o7wfTlJbipWOKd
SylAq6U809C5GCeMvdCwQ1H92l7Ik6GzaqGAujfpi36u3Qc9PzlnP4Hs/15DH8Js7hnP3wl3F4Qn
Q1zV/Lj/aJMYxivNRZ6zluXXvL0AeupGPnREkjenNLf0qfa8vgkIi2+AY63B3nrEX3tSowxGM5QG
tjN1/avCEYOJq21IeuYWqmMNa/YcUs7QMTmzapEwl+slybi90PH9wXLeYJMu57KgxgHwIJf1NlCk
cohi4ofZJDEngk/TA6OVA/MEIRlxCoXKilANiqnmmJdgJcA8l4loF0fRhwDlKvQg5ts34RkjkbWf
jDWRj3R6pgwFfFziS/LFYYVoPiIE1Q/btwVyQopcw5ZVNbgqAS0fbhzylhtfWk62z+4VEqRFPGod
na9t1TwybNUM2/Fh+5/Ej8FkjJQLh2HPJqdTPe9SQB/e62Hzt7D3a5SJlEgoumgJXK5dIQeTCv6i
/P5GKm/rHLkH1Rqzh7jKUla+vTxRlXggr3HUNDAEc8y5jaGZ8AVNUxfmvgW61S56h2yybZ+7KoSW
rMLmNdfBEob2AghqeOAEIK4klQGXc3ZBciKP3GbRVU+W3PdPJm9lzqUpsLyHQQ+BjP0PRSd8fJoQ
3C13frgILjYrYpiib/iVqzWWBc3rwdXPfHrDnsfQwcqAx/xLGSEVH5PqJtI+Rm8CBFrepy+Nz4fW
PysaG9wS2prl+5mtKzdAYTV8EVjtU3mfEJmXe9qdDkcbApC87kbnYlwF7zmuwpPQ4//inhp0gnj5
AOaRUF/8eOFZaJ9Yy0X4RQr/1HIRRJfTq60U832RUYRg+hd86VGQzPaxkX+LFjVCqzNS9K/BqjCw
DFDiD6VRrIvCyI5yjf3E6KnCqrI6odi2+ECtC21faCzidVpiY9UE1Je74qoHV+A5Tow09gA3elHj
7nMmPjOYWKsdvj63xmpCPBovcI+vXK/cgbr7AB3UkhFnBWSMJ26heOeuW8F5bWWLEJJ759MYc+Ub
2Mo7s1klo0tUYLoeZKbE5IYl0uV/HUPHAcZl4S1K/v6I0mQ+E3sM2yWBqzK5zXcD+pj68LLutBI6
ARn0OJ9+EYcY3vKHztaI6nuPF9kQoUlLDGU4gwmzCNVMFvK4607g61Ng90gM6Vn/WPHiUwtp0RVF
KTOFXRGs3GUuZ9WGK9meJ/ivjo32RxK6yKf8w+IF7jFYHEyjfFLGdJ6xSq/2X3tdOP8JRkjzZHSK
aZseh4QWRDOZpiafeETYJe/jTsujD1IlVA/Z9UwRs/m5zPP0LIIf0wetDsimHbe1jHK4qOxJnJ7Y
xG1MabCJiVWFC3Z1gN6SicheDveN58Y+XbRjBxrJ1vBXfJhu8Wg8mQGlbzLEyshIZQVEzSiBt1uH
LbNX500wJWsjehfxuStZG3Qh8/NgfvRvbfuUZUOSJl7xfvOIXkUoZkXyu7zVifsu85HmMdbyvdrs
n7DyYk1WTbF9VanLEioBQfunqzqhO/Djg6V+nHrG4ZgBlgbjT9k8qkcAWnucr3DgDfWRzSBdtFdA
CD/eV9AmRCeiRqTClufm0fs0TPoJ5PeZMk2fS0PcUFHfV7R3AnszV7917seadtK9rPoYghG1Crjy
YPbCPoE7ZRQejNkSxi2i8DJLdbV3+OHnL/22is5KCthhpGUaQ5YAgkAnZJThbAfgIW5457E4hAW3
7X0gQvyQThBo1j2u1fy05NL3PYh46xK7qOhKGBcQHEbIxLnS3QARurD0JPgz8TAnZLKEsG0fuREt
2edh8/Lb4+PkmMy+CMxVzO4yQbPNJYmHlAR7iRuKB5boxMAoriAvIYlNXnMQDTU7eQFr/XtUFr3Z
PyAvXW8JKlBQYzuIj+7OTHgfftsGZMOK/971wXuVdxh09gWRZY1JIqL0UQBtS10y3MQnAJhRjXnt
lGjXkpdWU5hTAH7jefOG2rfkvA4oMXBdRvblXwOiRLVLXLcvZ96w5NfLQD3uFYg2wpUevVuKUI/v
xPsxq26l1WdBGJkQ9iwm2kZ7DNj+M00mUTqlUj34jGWlRyjJWHlvp3EBy/DoEWfluQO5EjFgnQ37
jAdbNyDv9Pf13EOTwKZ1B61djawEbqQCe7+gSGCDghIjh/YyHKviNLPCEFCmWgn7uqpdmjh3aUux
AOVlAp7UsEzWfM8U5F/dIMGCue+f5huIrHfsJVNuM/Iphvlkxvs4hurEnQi7QQxBbMdCFLaCNL7J
Hy+ErwmG3EqU7njcUXbCcJM8oVd6dWBgPgDHg4c9TQdvjlEIAnj3omq0K5PVGGg8r9qq1joQxy9w
5XL7fLO4CNbktFg8vRLp3qVGbLQ0+HiPv0qPuWUZjamexxEavHM/lJ2V9/ZD/n6YId08XNKCDy/b
sGaopTl1PKFgYKvRAHhG0/deRTKTjNlv7BCIgdg9NOPfLglz+xiyFAARWxPe88oQc28YosYfpqTC
1H4eKZUTmDA3dNB3AoAre5nMsdyOzsQ0CInruktQUi97WHXhYu2fbhs+wd1YRXEE+wvgsst8y8NO
jpPduPkGYfDKt0PgTkW2QurFQkvlJua0ZnSIlHWBKL2KVfz5CUJveCUrg6D1zPb6NmemX4f75z5/
xVqC6PxiZORHkqyiYf8Gb5Sm4mdfYTjbFXUxUcDcEPS8dBBZqEZ1LY5yR54woiMM6ojGPVmZw7nC
o5BFmNt2bUZ8FUByv2Pk1VLxERPNVzC0QWIIuKVf1QitI2BPp/xmgf+gNFJbfjgTOEHIZbqV4/MQ
isWQWdhT5yHjLcata3gne6VKDX/LdPlrRff9hYkVZVTnYb/PRm57dwT8T2UgfmjX6k7hLv2RTdSO
iQ3Ezxe3g5myiNik5dyKojw79dZWsytZ9Q0g+bUroULsMAfHYzK4mHgVW6YnB3MjH4Znpp1aoJ3R
63fLvF0m0yaMD38th9YzR/V5RoOBMa32unlKsz904r30xPf/08s2NcRFP2VtqFkppmcYMIWPkx7R
run0lDgjsjgHY7NO2lapc4ohcTHr7q1e6YBgJeVBnmuFC0wk4vjUeeN2YtFB9pFFQOMItLP1BNJV
grKnYfF2FCLoA+nsIlH+qmizwJHzi7W/wPWeTFpB1bcvouUqaeUs8Fli8RsJlZTYma9szeieBB96
KC1KKOyfYH6vOnTRkIUF022L9UiUcYP5b4B82XXyngEFV243DkeBWw1PBHpsYvTMxBMJ0K6tVAzl
Nto3gghq0WavkJiQ04+CpOBpPpXDsORkJYPWIcM4TkcpiGszTJwtUciNMLFGdKJMTkcPr3OjAGVp
ndM4heRBYBwSTNHg2F7rnqaFyoCO7UbpCT9m60a4h6O7IDJUrVPJVxDMafsZMNw85j9xCSdkL+f2
W45RGaJOTBcZdEHu5cqLjZeCAtiskzYOaxyzSpQs9khnVYkFLgsSKnOqUWdefymAHyeRAF/ibIA0
RJCHt2BSlRLUO7sQT8sZ0vQhSYH2L+GgESds3F2KRfVNT/CahKoFlwNRf010Tk8zhFjrZj/rx9nt
ZW7AFWro/+CX9J0EOdJfUSb64FYsYp4s7qD7D1C++ospf4FxmcsGr3TRazJkXL5osrUJysushly/
OIulWhdFht2bGlTPqj78yEdvz+tN7Tzl9p89s6N8beKOQG5gB6CY1uYbMii9Y7fLihuh1BjFi8Gt
D2vYxx+Y/RnNHDctf+6tFC2XtmDt1gkqJmYqVTVHzUp+lenbNCk1ibZPOXM1QwM2ab09bDr8Is/6
uIm8j47bao1+hACqR1yOElA8760WBN4+JhSCaR6IHoOvHA/rJyKf9wt3r11kksz5POLFBuyvmQUr
XnDEaA33dFnel+MBMdRgJafcJ2W2c+VcG5M6NDiRsJFeke9gwLNgPwH83WCNVXW9hDMCwx33Jbdm
7CZ/DkHt1bB9v3Ii93wyhQchE1X2pJVp4NGmDQqr7PtmO/3uF7QsQhOFvBq2wRcoaWUhSKXNUeVx
MYHTqH09yLeT0cHd6BJy4Yt1sVX3PHk/emEye50Kh3tl9hV8OyEbT+tHZLx5SQufxlk85oQWrvbc
bd4zRMRI35/H5vJoJrxCIcgTJYAGUNziYVt12u/xmFOscUcbDK4thFzB05nPre3AATZclBASr8ch
Zad0dEJZwXbC6EkrxSCA+Tjo1GS6liGG8lv32vBkGaC+g5tZEaTwQ8lSdvtI9whY0tf43gbyulfv
igjyRpvx8/M3K0F/CBPrsgtKpyqIlkTFCy7XhB99SAf3ERtVOEl/ikNOPec9y7zjYFn7bda1DvyB
zmOKhuVUdxqiQc7alDfS38nvqL2m902JsCOLxIdcCSd+hvx1IwORTjSPVB/l+/lMh+GnWVJdAhGB
8TnlxvTImuOFgbpbqX3PRsSShZke7eOjyDkDxIeljHpfx0RI5FWK2Uswx3cK/Lp4TExB+/EL/3ul
kEgE3oTg8B6LzRAUInD0XCTjVyiZtss6e5hajHTvNvQUAn5Mrebdsr9Obyv3MQMXMF1XakKvo0HG
pd2dhyuNb2gf9uBG1SY8HFSH4O+KTtAIr1wjg64YjEnghiOQTe1wTywHtPqvcGCpR+oSemtI8uIP
TmIalAV+HBrSTOp07kG56+iMQ37tHmmVublmuVefJvOdGPpzefbNL3/pjgv8suJ6BEdZ8lc4gMCY
6TGRovEEkQRpiI7oyqCXFlqQqZEQ8GbaMtranQyo2a/YX4WjTHTjryzVcsSTGjecWgaQApfOr1aa
+CCfx1pumdVrA0QPLiZryAh2jbGJZ86yvmdRnmFkrGN1r0LHe3vfkupMV5rOpncga2Aj8u6L8+Th
cnQ72LflZlGltCnYwUE9yxyGzvcTCu84w4MNcQp/ReTvinVnCxEwaNDR1ZU463rWOxHXFD89WHl9
dtIKy8sLQlxg94ukemoZfkIVO5am5Xg0bz1u8M9vQguhbPhYeRWXkTMQ3an23Q272pNnsLjJ+Nnq
3K5fUijQyHorWbsy7JeERCDt8GQlKxZpQwfd5aaK9x3a0BJYu6CUp2WnW3U4+gy2+dPI0rQpqb2z
RO/oaj6MoUucPJktr+6EkUy7UO56llvVLtUY8S1Tjrn19rbQmx1VyPYrXQQ5/9DN9j1OenuCmkNk
oQZhMeO40epusCgXVNDcMVOnZ+s/7WF/FHNLTWc3uVSpYgfBn9MWpyoo77uBwwIRjtNuS0U0IemY
ETuQS/1vpsRRQLFxx4B2i7aAZt1FfcNCavWayMjTJMoWQA717/cTeKw9wvRCMgumEIyI8UeBAYBB
SlBj3J8hXcWV0ShY72tVFplzjyz4N7D90AcARRTVW6077YTmlQVwA50r2byPok2+xdxBLWVyyBsb
VVdT+Xh/aXKFAnBf7D56SHN0orTw2J3fGLTsV3hG4B5QxzvcMJltsAGg9DQXIlQPXAgXvTwsOZYe
ZCNQGHUa4vAi3HMh+Eq3HyG5ajG0GcPtjbok3pUxwmuazdLy+ZEKwjeEhIWexdC95/kMKWA30xFK
llzx978n+Hu70a1ud/WPCGVIxM7d9zjE1Wm0aQmbbLeqZUZ87VKkjghh+HwEGSbKZ5Ri08lrp0m8
bUZZjSphkp8hyS6s1vOKkh+e2JpQBQbqw2PmF0MUUzZj5hZGdYPU1if5YsShLwJtqDAlZzimlKNE
ER7I6MMjOgOwBO2yTsEQ2GAqFn+0D1bEHPvrQHAQZlCTkVZq6oPAI1L5KK8/r5SNiEdEynBmpPxz
uCPgj+moiZEbi+NdfwGz626Ym7XIVuBVQQ42ouy0M6KCwnsjGa7UjRzy7z4cv2t8TbDPK1wL6DJL
a1rQYSKrSuyKF0NdasF6pdAGujJ5RQSTEhYHlv0Y9qkbqxYTAA1QcSfqKqzycUTdWnMaKOonAO77
hqNoc3L/nJkR0urI32uOqqb079jZGsY3u3qbylUbFwBrpQqyLKf45YApZ+NbPQos15NutyeDWtFd
OHLkGIxYgcMVc/64ZUnPnlwxxGyxCI6J/MpvI4AbX4an7EEp4vRyZYDnqPKtPAat4kCFLYTnt6bV
zPTkxXlNNjhSnxxFn58bhayL579tcwDWvFkRWxoh5uPJyB0iP+IhkwDJrY9s/cdCxgA8eCoY5CuN
EeM7zeK6wT4V9gRcoFksy4LskEFkSS62YYE4DxPxLmInnnsVxaXGQ6xxT/vhIHPLvZhEOjb+FcVo
G8jKwyvvIhIIAMEmBublcL5maW1/zMDWrMwb7PFLVQijzLXeLnfuKFWWAuE3PiorqRIY3fB715GZ
0ZTHb5Gg+bvk+IjwGoodf6OELkbwyKFVtRQgiQ2eFC0al2965vaHMEUWVu94pjmbyI06TlFAozVi
9BYdnFFldgLo0XXoiDtICYSQwamkgxz6wo9Ol4U/yw8ppf3cLtdGKE2cLB6L0RAMPnWXc8FTcMP+
KTFpxCDAwbvXl4AIn4QM+Nu8XUuzo47i1eRqkqHxtEZtrNynKI/R15JaIqxJMvnGi9ALiOJkhiG+
i0IwycfaXW07xxUnh03WvzHetfZx61eLbRvM3kliWmWEnveyYfFpaiQtmBj3M613mh6sGDShwAdq
WvMJgx2wce9vtlhDlIOmNuOWPu7ThULOY4sY8X01+DkMdRgPS8pgwtlbtVnSxCeO2/c0SqlWO9Wy
9QStFGTyvrx9+seHEVq5n38jkvrfdS+E+7tJ30ctPOCyaR/eE39eMK8TaQSur8xsoiwfXA+qkPSv
hrXYc13NlaoqhFHC4WhpcMwMgd8ewEzBMHOwpdw/GOPG8hS33p1Un6RUdYvrbUVyUT+uCR4VjWG0
WbrAQOVYAO0YGTA8Thm/NwDkZCnJevRMVz8U3WL9u3u98Bf5oQg4y8trtU3faH0QX2E8H0eGy/C7
tZMbhGDyV9oEbmbwIbGTwE6FaEyYQzeAkAmSj/6MCuJs5lD7KQ/mhGYDm20xpJa1RGmJUyZWsQlX
oNuZWw17u/aUd5xczlj/51Zr8wE3NUj769h/VzUcLjyK7AwX6WZtCoGzoTG25QOo/MCi3VFEoFqE
wkfossyaq1uVP923YpbtrK2Zw90uYpYpHvAQKAnyGU4YihgJFWBBosS3eWguCTPT5dIS6O3PDK5F
UaE6A9j8mUBCJnbZx1sx5mebQkSz8xDaaEEcZxU1NIRZgVgMMljTvdepqQ1SaobFa/lYU90GmAu3
mO9Gtd93OdySMwzNokzwYktjMm0g7279C/XeZvf/BcoDWbItTDS/X2ObOF+v1ShyHos6EQzqmj93
Ac1rSHJ5msuF0jk5j0t42JigQQAihhv17TDSBRU3rFEJ4Wt7UlDJ/3N9m3YChZRyWYoK76ne6msr
nl3nXsiFdKYx0WqNen7ihhj15sAycDE+VLwfv4JJY7b7j3F05UpiLeCO8WKDyEi2qYB4ku6LR+Du
JJ9jwOlOIpNtdtGeOQBJJ6rXuMgHwc9kGrxhMXUCnr5NDx1h0fbd6VxYiXsB+KjoLo9ULQkjo2xL
ZKhqfBw3+dL01FHTXZ6AVSgHpllViX1A6lv/xQ8/0ZWNJdnAsrQPI9Nv7C7oOnA9jGabMrKNN65l
MEido6bAbFvf8KCdpIhNrXj5kuosTWCgVY8eXBJqIpax26+YVMRH2WybBiAHq9OJ68fU5slJRBPD
1WVqutxQFwUqtzlU/jwOvbi0uOkwjTtWV5FMdynqjcSz1FLW9c85auyHcz71JwxF1oAH60XyLU8y
455e08gdeXQTrsbEKfVvg8Y1MO9H/3RHN5FGDsK8e2yaZUZ+R6X5RTa0JZUEOXTiCvYfM+nutwTt
W4Zymfda7yr1AcMHGqVJ8q+AlwUX0XNS59qT8OSdqlwe1r3rRlMwkwSJLU59qjaW87ROMYvL3FMb
r+2N7hrxrALxedzB0FzAVEK/sAsgbeCAT4BV0B7v6TES29d4bOh5rFZyDsp/idf0/eXGNim6kLXW
LWY8YVOpMspmcDskRqk17XNOh11P9HOGYWWWqxEqf0uPAUGCFyVR/unzeY5/oCLt15LbP8MnZTxL
JdGcsnXWtNww2lV7ptVLHRE3FouNgIQQQVYv446Rh/o900ubXrwp1Kycqti28SXRNE7N3DmERpBk
RKP8cKFCU3PTwOOyb1JapTNQbJpaEyzpcCAPjjSOlaznnS4XzXTbSqVNabPci1K7tu4+ZazNQ9pQ
DczPAyC9w+Q0xPJtcfAzby/5bLjKvRjdIe0FkHxGi5bn/LrYZaXD7+Fh+f0+lYyftWhOwSUpoPOE
JHQsFpZ/kabONz37QBtjsyrg+IZHFrNeAYPbBUv6rQYRiIra99KeiyF1mas31DR+GoFp6Z1kkqrV
1ePidX8HC0dT/TLn/xOUVxool15R2rkJ6wTVSG75aVSTUVJi9L9JaK9dL9VUa+TUXVhx3IF33Jwq
8mRf47C7dbgRJ2ALKgVU3FK21R8fZwHCwloFdfUC+sCZpTdsRA/40eZfcxmQp/mu1OKXY7mvJahc
swZfwILUP3obA/PGu0/dPoB465M5XmO3jKDxwj4aILg7DKBe/PMCmqChfEftjcvclth9iPIFgGIm
hKJ0ZEVGOegIyr9VK4RuHv0cb4CfqvsjMC9vL78O6F7IVRQXICaqImVcnvNJc9J1fLKuCwqDPDCp
u+iwVj6WOX8LqBWuadlg8GI1C/XbVcpfYSS+MrXjMjS/Ag9RPm5SK3+/+evDAPwa9RTyZVsSeeWq
8Huui5IJu+4ZyySOhPr8Zmsu0Z5z7z/o+FE7qY8rg+MPV1nJsCElxwXGdsh8V2/q6nW1PJkV6Ij0
SnfKy2st0GCfkDzUNjjoEsLcATA0HHvsmktqG2LHBW9cLLzTeTDl+UmCOROUCixkyd+3ZZ8XLVuR
0zHk9ncrRAPpiclQ1c1Zapm/tA1LGi+Pv4lVr0dPOG9lOMK3UBwo17X8sbVbsn+HXhPFWclZD0MR
NAd8AjM2aWyt0j0i/b5AHBtQ/IPCpq6bVOZEuo/r2R9Tp/aAEeRNzYf+jNzW75Ll2fYjuV1+fwNg
4z3C6vs2p7R3Mq+kXBeC2p1cpfxviu/xZnqw+2EDKcAfFlraxqDvXgD7v5aHYpsN7KyLUQZu/tJ6
mR7X5JROES7ZuC6Uk6tfFHzk3F2TEB5WQJMkaFCt/6u6IuU3DnaGTRWYodMJY+0K4MF5oL9vs8ZC
QYjEIjJF7NqWHDpMIOU+SSnwhN8pHBJJfzAyR4VOzUDIR343WSjDPzRN7OWnHFGDLtVLr/cPJIjZ
ZTqQ3duXt8t97uq5kXr+6gZBBDA05ZW0CiKUrfcXAKmp1d7zqq1i5jVDN55BmOoHthYZKNLcN4dn
/vOBGORtpy1VyTtQhn19n+49i6uV0/cUVcBGfl+rEJc+dkBpwpthynbsTIPEB85eO2H3k3Uwyduf
Qvq3LPEJjWeYnkFKxS/gO1vahZP/xs8+tKz1+viKqX3pe4pDZeoI6mdevA48aNvccr1TnzaTG1Y5
ZAGWii6NKjicDgtZAv5/jlAgprmvBL9qQ57oPzy+KnFnpNf9SSiNR99m/e6lEQUMy1jFW37z2yiP
CxDBMysi2ZXco1fIOMYaauLoihGj7s7QTmpXr8p3I9Oi8iWrdtXCFPutL38QWBz/aud+q/3pS0zY
CZGXkcM2xYke1yXXhYnu+oJ0aLmBB9BwJgMO1bH6KwTWx/66qzXF9FeEJ/9Hs+5VmXXUB45HmLY1
k4dEhRn11cSOIr+mvkSBfUCJYrW38xA3FoX8GosItA1kc4+vjo7k7uEUgfAngyxJHFY/WaLUatZw
LPaEFH8ifbP7FRmPZPHEzzBwACoF45Q/3HALfOFE/OWs/UrvE07sp/PxW/Ia6N2UxJtzmxcQYalG
B06glrN+BT1epfZTzpkXhL9Fn2miD0x7L1/8eeEQ1PMC5C293ZncR0QTURcOtlR6vnPyKeq5i6eh
Kz0Ze8pEgul233jUx+7BtDhvP+vA8Vjkqn+Zq0mUyLNWaf7CUeahAZcfTYjyHjEubkArLKDdXniD
VRaQQDW9LVryZSGHjVyJNxKhrUQoFac0jp2x2k6eYTcgaI6GhAMYSgVs3kwzuePqcSIPLiHYCiZl
rECIwK8a5JxnvPbRj/C37X8VcZqhtru4CbKM3de+y7r63Aa0JFUlSPyd/MbEd5/1enUZQaruSgMH
k3ZhWMg9iDMkGd+LZ37q/+aPgBgK3n66jpyhhxSY59FspFZ8qocNZHIdd1CPtE4lhvw54gVm+++y
+4RrqpLYD/yUMXnC3pUVbQKinRXteYxdiezdtta4/947KMWqWPTxPXcxBMsPk6SU+3hTCpoM46ES
sH49dYmTJi1/NOtwz5F7a/XLvNigXTm1HyMavSdXscIQUd+L2tDMucswaLhsPm49tWv0qFv4CHCj
HX8/rpgKzy1LcN5oxQIxwqOpVV+5T7yH0VdJUyB4GizDyRDBnWoAgSz1HHPfPX9oesDOnDtUFUqT
4p36OQ7yyAiIwqcs4WR/MDSqu+3KesRgagcV1Gv/eKK1ygNUaa3m/uAhlBUmuRkTb3+1dTZWApAF
MHGLsMi7NeUMZpEAHD5Y9N9HiZUytZsGl8k8BcsYmdDVbXQYn3fymBOBlpcGuu+QCfPEaW5gUdWt
hiqJHQLrQRkZhjITCGAC7qTxFOPvMnsB9uSJ9EKZl5fTvNNWcLZJLtMXogNcn2VkvlZf4EB6MFpo
L+itaZld1iGQubjgU2XETkY125DqnU+XiMpZIu01g++0eKcWHbuzWTHisuQ2wWL5UcLmZcf24VJS
Bb36kww88Q7Tx1GDNHiAPoGTnPe96qXUqvqxKosuMcImUTCVH5QTrWH3lbJOU5QsuFycjozYts7E
FcYSUvJy5IFE8ZyNE/sn1UBu0UcybpFDTiWe+TLl94oqHifWSDzTYS6j1KF1moCpI+oFv1wPBIPc
74/lNHk4biqTF+US3vry2I1Jtocy7JlwmkJjpX/AYv4KiZ3mk2vwJD9e88O/7edKdnMQdbPbQkva
vdNgLXoIWOh8L11bZp5G4gYVPfwztMuFP3Sa6zotZCvVGlNTqUQiyCbZ6JlR4MzSeCRsfym8TLsO
V5Xfc3YnQ9p9gohhIuBZ9dKnPPc7t3HW5FHb11JuyPTTyHLd6G5T/IwDm82pPfgCj1QUGTNwi5Q8
rGvHtdOWTBXCnX13d9U23TOxl2yFw1lPCbZbobSdGERrWMK9tAJCxjrU2mj1RjpNaMNN7GoyDwO+
8f6ZNpgWBejiMJBkpLfrvCiTkqquMSVcXxEOTZOvxmVNHL1M1s+8G95f+ZmpJHxNzE4tVQ4uFg3z
LSgNeJCsCK4hwMDVoFh/GSXOoJgfYUJahyhEg9kQZQHHhDyJbP+WY9Tlj2MZ+cZ/ehAJ67OV9ouM
Il60EpGgvyQf0NwcpmJt8TqvQ7+IYHqY1yvodH5APZ9oBDNvw0mWcptu7myxehp6OirGU7UgVMJ4
IYvjje8EJuNmkXhzgipJCOTh/cJYGqh0goEs/fTEKLED6RA2PZUgGr2nrjobDQjZfQIYibPHhGFp
w9BBl4BL3goWuO2MdsnzFuZb5dpf5pKRCyTIUA5edOT/OKi/Z+DerpvIFPO0d56aoAPDQIpl4fO0
g1zpYhoxEr+I4+4dyVZpiMbGpDlTshzV9UI1xa8s/tuIXLYdW1stR0ibreJxkjW0EGCgN+rME/3T
P73/S24jWKADzjEw2/5chpVPGHP1dsewyDNF0csWsK1TCElOMlbgz2avvh6QDZufb749oH3n20Dt
XN1maKVSf4oa8tE5AB7yCS/1gIzxWZD2OdIZMHP3ogCf659AR6Yf4ck7z7d3vjsRjt9YYMF1WB/p
7SPjXYdcGpgLtULxmoADSZou+9gv3DYVxviSm3GsvOTZ+LVX/RwVk4pvx4IDe/j7jgl61tTAFosd
2Ja2lDHjXOk2MgnK0fogkEnPyYOnWgTw5NSc51+8s5c6wWXbUtz7vJTTPFQ3gDX6Dc5bMoCDysZL
lss6SD0F2DQ3S3Xe73hOTIkRC2r2pgPqYjaBENrq/vLdJ14uBXAQl4bhLfqvI0GpK5Lig08C3Y/Z
eKSPQe3SM+GvFZPKlWe9u2/7YWfKJ97IxISPhQmqg2QP+ubr5KxfQFl5QtM31cYEmPfytxt5Le1W
elZ75ZykYNHnwnVsLtUNivCWGRWKgfWyMQtbynD0LcRNqxT+GOLHxq7M3eaqY7znMhRZBifEwxig
VhpKcX9cAlQOxW8r6PPXRE7zOgEkHks4R/V25uC4j6WJ3xBYaR2/ere4bCOEp40ZMiaCx5RD6/yt
iBAN7qJfVb0oY57gxUW0bjcbm2aPAdez4gLyGOdOPddl1XFmyYFDvaKryqKdnO4qXYUX5CfgvZkY
UFTLgbR7HAUh9YGfN8+AiTtjyhnyEiQ+Q4u9dObycJ7oTh24kJBOQyglor/nj82pT6FeHFHNCkuJ
tyIqpPEhcj+GEbmoqukEnpboKXnfi8hLoDAZpAeQb2OJrElmqDTs03TSw0R5o3gT+RMkCM8eoTvO
bY2BBnc0FlGBjImtSpJMbV56oBw2etePlBXJiLAyvzXflNcAsp8uzhfNhn2T0k/x0iBCoCtNfbzM
p3YUoRl0oDfdRx9GKN7fypp71Su+83MQK5VzloUD9YQazCFV7cp55yCqcJks6APhjwbvAMMZntwS
JiZf5F6RXDwVv7juhz1f2BnuRbB4QC2Cxxt/reAmO+I5tOeZKH27EOH7p0Y7zmWTM/soIOw/JJWD
NRbkv/7egVH1UJGW/j1Oo9YzFvGv3GtVsRwzdgTeY/KdIsoGnUv6PPzf+TrHIyKfvn9hui7w5o/Q
+kZnCfzNELfo8Ax9wqhqcIlMxuMyHUptGVj0cg1yXWDR08JS0mc/x5mDoSz+CiZxHbM+I6cdZlp2
WNvZ98TDDgVtuM1fgp0E+voHTI7ntqbrbOlmQV8Gaub2cQVKwrt+HJbaOxwKdj9gOng/QOhUMYFs
I53s9Zz1DQRdxvo9eI2nP9bW0QgxH0yBa/MKiBBMJIAVwk+cYP5z+cOf1GHDJYJ75gHHLpAUb+jJ
pJDBk3LCXwIac8n26mL060D2fnH8FRr7FZZE+lgMAeiIbdeoAqvPG0TE6uqyFVFACW59ODphWuD2
JgNfO9EYSKF2tI0XVIn+2VNpEWSzW626QrC8MvhlckyocK3/DDRaSEU7msNmk4CX7+BHo49I4phi
dKRGhMETrRU5PZPeb+ishNHGkYNAjyq+M3RO018nd4Kwl1226KXmeyaXndjmTs/wGdlEYR3AS5D5
R/HLCuBaV0FSc7dJqwgQiIKPDIDj3tGzQLrfsW6ZbpmRnBCW1P3shOcCHwMy8hv+zA1POQP985WI
fTldw935CY1uLD4oOyik/BU6P5foUY0ryIZoNC3Msqh/9HjvuQcKxWZ6SDEVDC/WV2JN4cA0qsu+
sJDekT3dniRwmzRg/SPZVgpB4lMSVtHXKRnwmdTKXTHGMQw6nJoNH+GS3/Zv207Q/KYflXR2ZcqQ
UzN8Vd2kW3W1xKk07/mz4gy73uYw+pHCv24MQkv2n1d/MEPiQOZpb2qyGLTDyRdn8kgZrPcr+Sdm
tbf429w4cRnKjoBuLiXHjgCmbdtBLJSu5gVHn1P83O+cKCP0lRavb+qnTbtGxcTe9mHjYfjPbqhH
92YFw3y9nNYWl9Mb5t3k5RZ8fzsR5SF4sZwV2wHYtSuVq2g8+TtW1b8ODPtPFVnWeQs6J/OHprlM
5bAs0fXyP5GXpiOxdoxUBqS6Prnf9g8EhHcxqAXTTKEbWrA9OrBT3R2xCCn13tNoVMgpkJm7W/lC
l2XfnpQ4LDpjVdbMhfMHyzLXqyOu9m0JVYP15dbDNOk7RSkvSdDFw6NiuN3T5IyTwliB4JGLTR1G
Ba++/pDYSYWKFUEUn6JUAxR3li+fZDNomqVKRTmACr+tnqlaWTHYrYI/sYQ6CFro44DN5gkrvO4B
uyx3po0AEE8fUFdac5wAGI1ZRN2e7jsKmsmmh4H6RjPrfB/ZpDECmYLjUEcuPvQv1AlX6E2W8Sv2
2a1uaIkr/8YXk78a+jsuC/5lVqCnO5WA1OEXE3zy7hr1EC2X0CWMtSes+4tfW0UkvucRSFbqIZHt
8PboVBbEtm+RCvTCaELGBoRTJOLoj6+6Wum7AOrzKMCDZcqd2+n3OPxPRAeACuPpCdH86sbiI0YI
4koHP7arW2EjaxRcafdM2Fs44vW//nHZN7UOFqcwdgb8hS7p3l8mbS16Ob8a5BieUaO+qwiK/+nz
Hdr+7HLCVBNWr6zaR4a1O2B6faAEhWuhKjc0PcAgnt4nVR/Uy7eVpDLtfTbyqipmnCEFHlC8ytNv
0ebLOcemGUxHmzt3FnSQqtmiJnGtxBU+XvUpoZoqWmW7q72uQnPo+B9cNTea04bB1Ou5nR4PiZhk
55yO0ChFZjIk3mgiiKtW5eHl2exGYA3kKgU3VNSae33nFnlwAbp9q8p9Pn9QHpua2tepBA5uM8KX
2uAP1XduuQs+eQa0SZQiyVtRIR6X9Jt79aKmR8p3N7Ce57WdRy0qke/188B75qx/+Y4mFsMY3ayl
aloPj1w1cubcwY2T6mRlB7kA93xYPRn2SMvCMYrC1F3CShWTd9IUqixST/FRFj8EsGTGdDABX1Qi
m3PPrHTc0sllf8Z3dHZqBcG0C5huWK6AVBsHkmZt3mULPMXDGuW3MPNJPrUs7tI8PgcZQ1kn0FuS
TLCyiDvyTVAugUlP5W5iL41NBEEAlRN/rbMnD+Ax9o51TwZzzxRCMEPDoG1ZOPHkiYV/k3FOIBG2
/NfAryFHFzis1rmf7WHzDOmumH4B/+I/QVrXliVI/7cj0GsKZNEIe7sxVm8cQ2iOmP3CKb/ZkLzO
rct2zzJyuAa/ray3ImWyXUPlXp4cR6yoeGUofGIlATwj2cZB64uXU8Mf/EN47vubAYrxCuX9d7F8
1kPv56YhPh3EMOSbdn4I9KGI7sYLwGHYihM53YX3jPwSzT+1nCBhA+W/qhQLFC6TU+gTv2hheDiF
n+YJWvQ5n/lduf1cwXXSrfuZMy9DSAlFOjFK4dJNjZ4ivCasbyRhu5KrKur7Q6w7O4pQ5mcV4XqO
I+hSipTkujg1iYesn4XMztDo5Ng0fjxy/vUKS/hdxDSy51zQv+TGxFTkAFs+7i0ijKfhy8nhnzEb
rmudE1E3b5qPI8KX+W+FmPcTb1QZNzdlX+QVBuJow7DINVfL6FaNhXRG+X0JOcdDlWljHP+st/sc
yK0O1nqUZSK34b+W+i4DgQBOiUX94tPHLVDD+wVRkgg78M00gfWaTrQIf9JRdtfB4LlTPG3U8XsU
DOWhI/iWTVYX/aJ6Ji+EqUkWXvkFxwcBRKQXGoEmNW5SvKx3xRoDTlQYzaWji8VtvPYAk8DMaANY
oivAKaqdmqAq71yQWsPX4giYx0SWngfP4LEKaOBfTVwgyADIs3T+8pto5I4utMgVXfPaPeCy1InJ
LRt/dsXGYCsUp3+JYjYaduoKkAiShA8wffKnDd7+euc6pCiczuYc2w6DOidThA1mUx+4GFPhIJU0
ueoHLchlWH4oACvDsaLd1n/o8IdFvhFevI8DrM9ZnU+r75S4ZEp/Dxf/I/7umeg2zGEaJP8BesaG
mavEVX8F+K+rQe3dGf0vnnyC+9PcXsWj9lxdwGHrj2lQ6DaE1770iD9eT6vkdW8P5SU3Fb3bJiZY
RS4iz+eo63vSk/QdMDwh5o/hVfqdJYQYORRjtml8LV6Kq1jqOp8PRDryTCWA9j8KRm2dZYlEfyYu
/jHzM0ygvwkbFHh5K76qPT9jyfjgk+qLJtCmgd3wgr2+QgRF2Y7dQQQ0lmh/Z8VwWzkZ7118PLoM
KBV2VT2d8rZ0QcHr+BoYRoX+Lb6SmY0SYvlIzGf2pZ8bx11E+U/Efc1TQcZVzIkzxSIZEohQEr6x
Zb7ZR/tkkXlIMc4kJKNogNrcSRROlO6je/mLqzJXFThQAcTXlI4EWcJHfoSCQ0Ea7HJQDuZNaiJS
+Mjr/t+EthsFujOO4fL+0DQcitcrisJtR8BxEnWgQ+tOZ+CAgWWfZ/w5MT5CbQLQ/+KWNOlTTAk0
Xss4YrHTdcKRaD/KeLsY++4N+5p21AKkgZ1DfOxnKhRkIqFX1AYwI7P/f+qOYkfouizyfA4R2wi/
tL8xnizb53Fl6wOlfIHq184ogYPCjK5PlbuZ6MKS9b4vhysAeURHzttdI9C+zLvn12+xKO4grBmo
7IJxQVbvR6+BzEadRAoKCSuFxjXc5v9lQ7pr7NCVOeBovdb7iR3xE3g9MmBMMCu9hiJkE2I1JcOy
DzyuM2+ma9cJpNvqgGNDK6MvckyE1FPCWqI/gjTSIbhqCpb9WQJMhAtqqJGuSJ22F8LRRSo5i+WP
5BkhWiGFbwp6DiJl9Dxxk4mx1NSBBKmMKa6G4vlfdgK0K7GC7x7CNbXssaIjW9Kw7eNnIWUgu+MB
zTqHOvnUn542cfC3PFiTgirBYMGtt2EEXHuC93Eg+ZKNqdM4bl49vod5QXOIA5ks4hcayX9MTKoB
QKFfp7ZM0J+X7gvBsqeO5pwtXMYXEvg0x2zvhcqkVPYbbbTXAuefBQwKcDgBpYkuG2L81HvMLfSW
2UcJy7jNv5lDgkUIdsJ4IknKM2AhN5zIUZeLATrelrSxwW+S++f87WvU+0mQFbYseCh302ccfj+j
/bii/3PQdD2eKs6gbsNCllJmnYvDiq8hlDq6UwPXPE5o2K/wgw2ba0kJz2BdtBTv3p4GpXTORZN+
9gj/bg9KAsLoHckernKIrVkrsrATQUh6kIsIdJvLW+2OwgXQpcVR06Kc+rJvb+6crUIZqS2PhEAj
7WtrAuHbU301+IYuHa/JjliWzXCcwr/DHa8z5Ec+FXxIiBhAdIFhZJX+3h5WYfid8ph+tmpDDq4X
O0dIQx8xrnBxwubuT7cSXwMOCZS3h8tHl82esUhaO7Zk3JApkPOKmnOvBcV4lWRiIExPkbYyq7C7
hL4MOIVJ2wvWH0SAI3jcS4iyKAROjz+cwKJCnYr3oZQcCEDT5FII5ZtB5Q58VK315+aoT5wKX0ia
gxfZx0rMeaO5QuvMc/3P1c2J6Xc5nYWeQO59gWnhOtOCFdNqfa1TAe+yhXDrp+0t95x7NZ+FIBoC
9vgqXUC1tzGcII6f9qIoNyXiIVs+lOiWT/gLylsOI/8n//vLZDY8a5sPmJRvT9sPUTP0qR5X77Fb
BuU070MAiQJADP23rxut/1cqbZnaSsKPpGL8b+bplQ3EfdfRNUKlstr5/5/Irdqw4grm82As2RfC
6909LAEKqaHelp/BvU75jJsxEknKoi0/aL/He64I+onnL77QjCLZxaWnmwSD3w/yszzVkbA0X4Kk
YyWT6OjMkxKTT2mT0q1YyuZ8ThtVTm1firi96InBFHOQTJg1mS6Gx79x2HQ/PJEXztVgVhDPo3q9
DOby8MIi9+8SFat3m0vF0s5KP/B0MHbN8iroex+Sd8QiBHIOdOMbSudT/ukWANYaUpUObZH1t6mi
uVqfSyOjxHNbyG7WevQJj0Wp/f+rjCIZ1//63WRt/Ilkc1epD1t0fqW/VWPPFp0E3RvzzCYfMaRk
CTr3l7414abdFpBjhdfs/fNCYtu4WC6ZCLPZ5s4bov13fpVDs50BQLpmMyx/9d+BryJi7CJU1gvU
lAE4nIprBHLnijy9P4gMg+5fAatRAAxxiBLB0eiiTAY4KR3n/QRFTUT1xS7s3D5N4wrqJtU66Zln
suIz4fF6XlHiMKbKDzUtXa0n2/l0GVkNUWOF5rKk6AOBmFN0AugGOFl76L4RZaklk2xOL+ye0yPx
UCJQPUyyp8y4cCY/eaI5iX+oExKs8kINIdXnj7CReVYnE0obtgwSUmJvW0JpohBDnjWtcIS+PN9Y
4t47awx2Ph2i6Xm+J/3i2uxRQKHgTlib0FS4Kain4yJfBnSWekEQHOhavYUdH5WUUd8KwhiTpvtX
0yVYRUgcxojbHfem6+jWxKQLMvJRZaA0X/qKMi/J57ub1MMCzwCApLbhQH2anUjNEbKgkGAm6N2g
D4RsDtrtpm/a7LkmxvZQW5b03zAunJHmQyIEx6dVFSeQrqtqaLS1Lqxo8geisnEdHJZKEyaN46bw
IZgnlFIolHmAASuxaVIfqCfOIlUQyy2orHuYDyMfHPMSgXf0v3nEKn92hG6zEI2R+58GcP2zA+uq
y5eAK+20REVNWgngsFTgX2296PXeMLvVd866s51eKTZHz7lb5pvK585xjZKLIjRTXg0/7+FAeqOt
kx0z+ggEIdJN79oR2ymtTM8tHDxa5MsoOHDMCYwpSVGp9MejMCM07xo4n/baSoIIMZF+B7mEfFEa
IyDg775kqgfBsBz7Ye6XYAI8GJfUjG8/yAURcRIT+Rnb4+w7Ejtv24GVnHlGcGJgrp+Hx7dMgAaj
SS9aMN64zsCg0A0zacmI9RfU90kaUygZaRyTq5LCb6g7CH810T9vORWD+bS3qFRvi3VdLU4Lie99
/464fnSP2yS67n5mWcmPKLCSH1aeaim4gFTnc6MNKOqe78jEaTL5fn30tnWt7GtqkQzTzLx2+ofP
KLbz2XBmn/4UNlqCa9VnwoIV292QjTnEln+cIkMriCa/nzWuVdMwq80zekvQ6NAuG2Mno54vflTt
6K7yEJuUaP1icCQ1j0fMJcG9uesrS+QVAId+EsgSY33TGpqXHkhOw4xXKmAbQZJAIerGT6LFbqoc
akAAVOBh5Ws50wQ7FRiJNgDRNIr3nw6fkK9F+YYMHql/XONkxrfkVyNBUmv5RHGMr4vuG2dwIa3+
mfDO8G8UUPLPrehPn6SWJJAvJkNT+P3rNat50O7srCloL6OL+P+0SEbetC1J5Wcn9tbEDp3HigpB
2YmM3B+aWVVxZAN0ynNRbIUpbXVUd2bmd6hye9oGYB2YR8A4iC8CTFUJTMvgfK7Ob/jz6iLVdrpr
t6p3eZYbdCvyvYMRxgMJxTSkIXOYj9K53amXBHKwEGMtvqqxteoBOvrgCRPxT5FeYDTj0VR6e055
DUB5ev2ZrBcCdQ7WaxllfmlyG5ikZXT5101UqD2ap++6ID0U9GRF/w4cjsPzZLHQzdTAbYyvp8ip
rKtEA22pFuyQWa1Z+hVqvHaafaP1DHPvc55XricZu46pm/w55WSCGkpu8TzuK8mOQlnw8qlBUjQ8
PWQYNiDtCxEnBJ+/T3wgnGk4f1zfnnIt7kCW1Cu+ExtrChwkRcGOKmTirIR1Y5D8wcy6kk3zhuye
/Lc31gYWvf4YdA7DF4kcCmFdUOhk8LOmz0BWN3x0CM+qZyRozmfyiYewg+RAJLWhNtHxuANAADkr
4mDql2RDgfbFnNeNOFVz+tY74dsBPF4K/KhbF/AzxqeOpzYqrPTXeCSCzw6PJVU4xXQ8JC1TlCG6
ku5RC5V5ZqLY9iQvLo8uNPdriz62LZB46XNiUt+s36ptr2LMQKrFCTl5dZ+pXKVOVTgp3Q0IbAsV
2s+urkTS75Z+SPnELkMh95BejeisB075JGP4mVv2Fq+l63G3ZrgqTZ4xbREz9cdjkhcKDqUJzODX
9Ozn02ozFS3ZGrHzbEJ5wZtiWnXJC0sxtXKXmJxOarJoTOU7WQM/Ixnj30WnfvR8L3HmwG9aJ3Ya
LJqANVMe0moZ/DFES4U0e4PY+eeZ4gY7k7A61i7MkYCFTiKorsUnF2vs3vT4b8XXimNTvLRJVoCu
d7ONJcbTaE4CskJ6mX0d6Dtr2y51DjNZVC4EA80D6kas2M1RR4Qx3P7XFkYS+Ot8Ti56FtEePyzh
jDfMS2R7ldE6UWyzQ2acufY+jpufCnrL9xoxdlRe1LCywFbJgG0HIhq8r4Hbl2q/cH5wXtYgchrj
frIG7nffJMSnNErUvacGKtsYtLhwIYwzG+odAZItVO14lRKkuzbFYXE0TVpCSfQd5o1kplShnnKK
x0EatRvxFdYGsZ1kMHtXdeQY2hSBmNrNAODifpmxxjSDvu0llb7+cpBj2VDqFwge/IRkUCh0ncaL
MQZOm9JvknR4MhAW7dH+lszTFejN681pBjtSpFnEGQabyrg3TCxlI1g2yv3Pq3RYZ8KjIUxwopkE
ez5Zuw+9H9Bppxt0zIthiflp9V6Y6/pB66DifQsoaLOv0LgxPLnlpyozpGiXN90S9gz1J/1ALzBN
W/75iEHNhD2GBXBn8G0cCWYCmNi6ZiDXM9o43pawUwc6DQa+zzLmgx8wZPdjnWGzshec8s3/jdAd
+Kg4RnJqHVa46pqch+toXQL5FeRGiLUGxkeOF/vDVQwRLT6Q/DH3bwZmpHfaDbpZPIXt98yt+BBF
ncQFHowYHf4P+/w/1dx9+7XWjP6NyfrWX56UdsvJrHEW3z22GcY3gCoQGOeybZX7YfAu2RBKU6JS
CjIQ86WXvi1miicWjm/mzkrHtJoqRoVY9aTQrc/xwieMhLztTPsYxzgxhTP1PyQYSTLRONTGgaQ2
gwC+dGFjn4j8jPhiZF3VshyQ/gI87tmZq4OkYd69u8DO0fvrqT9r5ry7eZ0BTh676zBSZodhYvHj
/6LW1Dg627RX1O84+h3+k11uPtxh323Hy0hoz2JgXHXTYEwRxvJOk/Gw9o8lv1yAUiyB5ZZEbNS9
PN6MaIco6AztQX1XUV9fuzeLYqzfD72G8tZrU840MRzb2+SaGo4Gm+DweO1gjClwV5AbiNO9yJuT
QXQufXmxoqZv01LwhgBgBE8FzEJBHc22jL4KLDp+G6u5/oCUgkcGIbkqtu0uGUfQ4rIghiZxZLfB
4m25vgCCNOQ0XzWWi1Q1IuBwlc66enmgwZJF8odjli6ytVLdgxlco1vpT2hSffFmtJjcHO+qSc6v
3jekPzYZ6GWpH2aPhQ5Sz7rJ1XoVTgTh4DNSBReymhD9xYkDo+jQUIIDcJ8OZqg6Agw+v7C9tV0G
h33Y6pHCKpyJJMg3SeBvwHmb1x/zt5iT0d9zS/jBkY8FKQ4qlv5/VRYgDTWW/kOEZsTtEiO65pmR
27vJNabkmpRrCDcjfYIFTcbWQ7V6kfGjwpwHVnVhVn6svK4KqAW+aiM2C0nBDFfiK6mQg1zLvb0o
szfzGHjvWwGVWZxvZZHssxg/wrUOZnfoAyd50tVC3oZnNRTtVhT7iXLOvJNgxyBNu0gRb7vjMW17
AepVJLQyZn/Q34tAlhOewjSOCUiug4sHccMuqX3ElSlXgjSSVIQg9p39em363OXLsx3xRBTAl4aG
yySFIn+OhckPGgRPEEDdN48F8eksH8L3NW294jAWZI5Iom5T+W4GNQDp2JZkAHxS7/8n49nzgTFM
24lzyCl+OxNFNgIOsxw5ONjEsJPclAjtzpo/NpzoQgYuJnyTunVaDQfEQqYEJiPFZEkJV/eHEoO+
HyuKiObm74odG/yMXJcMBtNZXb9cMqiQ6emGP2LGyEA4Re3OdSgWVHvUNNwKDi/yE2IX4nVhT/H1
ZTYlWQWfqkBh56oiwfslIgu/jo8xrHSDP88VHMptN6486OD8K3fIs72K9OYh1wamAVLDS35wXYtG
i4YJgk6DqffxkH6Xy6HsZ+WVKEVlkcrTnEAnimfwnW8MHn5aWTtKtzurBZy21bxnE+uEmMXsIL9p
j1aoOS2o89+uL2KgrXVJif0Obxfm4UCut9Wi74eWkXwsaS60YVEwvjC82Teinc108hCq4YALAfN/
BhcyX5bD8THXf9dULFWVN/bO81NsTTEmGSoxVEW8JAx5xEbLfUQ+TKwNgG1hGel7uvk1iaPimr8x
KnkuaXlgPF5/tsYZMiSwxCQBlDs2Yolj/UJ+/x7/HoL9S5Cwj+Lc/XiUBp1WsDVn3bNoanztimHV
KBRgUbtjJzsKm5vqiaINwB3gijNwZQ7Ts1w+63zcnYDtXINcCfZYAOwJtEyDta+lGLZ0U6Nsn9jr
PwsNWFKyVBioHQuigU15ogJSpBzp350y5qZry2xp4reqErfryCZlTg5asY2wAhXPIHAsmHEf+gmQ
r5rk79Ue0BqwVT4BUR4kV6fBvaNzWX4pXPSTPwmFklapbf7nq+2nshqNaONdfPkB7gklHNOalN6c
7gp6mce/ONdcqo/N6nGsuHsvutqx37/TDowgZzmbJHkh7rO4/nCTnA8yoILWB1cEE1lKqBUGo2KG
XvJF9rWVyZ6ISbt636gv0+AavSVz5Rs4rx7/66cwmEIOFrgvbNxDlzoRLfNf9yNVTrTnx5wQuasT
xrzkMBYRNxkTFyOIMvaBRohgC9t9/0YBVp8AV4myiuiKeSMMMGMDVURorVifHjwz6IApg9GxP30/
mH33dX2GUV00iKyZo+84WIjlDNhe1XHX6fM6hCIwjjw06NwPCPQJzIQEa5MC/df4goe3rC4L3ek0
wzjWb92CFwAv+MnEdo+uWlXo3B8TcKOjk922uYbadKzKY4ZU616/d2IyRRlLlunuCkeJRdMQqx5r
EgJ5ylH33s9jZwc7UakzWmoMoMqZT6ghXKsmzFgTooI8u6LmazVot/GKLadTzVdwRCOg0rRFNcqK
uQH45tdNfucSMOEcjvGty1+mzBWePjkJS7N0q8WlBnqAfcnQz3mpfopsd1QKMSQGoPojHEJOHton
MoMY3APWCS5JEoGsyxFpWJYbDZsO4EnaEX7+5IbgQjDFf0jJMYXw7p4HYdFzLlBJa0TdjVsg3pg3
ZX5fGqUtyIwe+ZStqG4xuu9HKpSrHlNYNtTaUqqueyG9ItsU376EPUrgR8HWBm3AUSjNDkbvvkbY
vaIxyYHuOGNWefuSjoiEdp86vArLW3xdYCEYiJacCskVqzwnDC/HkHdiL1pr0Q4IpPaNFzkJfI88
ZpwYAISrB7sI+okJclw3OYezOQ6a2WoOYFuf2Jtr3wDY1pPqaVGsd6bCOdC+fRU94L2pRfAy6Bcr
j7EtZVdzgcIYsjuOmKlMS/8L0pGHUOXqNH2gXxmyCBnzRQgghaymUo6RY/3/1A/mgzFT3JLYRoI/
aM9c41UsDg2NXC20jOT5mMlrwSApfUZJwWy7jF/FcPEwPOuIhHBE+RaPKALVd6MwpMDTfHoFYntp
bZzf8f8AVvKUs+O6DtoH/NE1KdAhwqX1Pn/sNtBJ22n9pZwcWpCr5C8JFOVgvHdCx8enIrLvLdJ2
+wIzUPU0pu6Jtq7qiQHLu6nDhiN/3euEYJC29O3OtBrvUq6hPY0rNZomd+nL0cX+cV8zezmDX8Tr
G2VL6TQ0yrL7MG8kS5nZATBLK6SjfPyDeBWxwxvoxV+zDpMt790/XfNJOewhYXBISE2Ww06Tv/nW
QPm9mEZyqLCHUoV3OiPTg9OInATgRIAlk6625J0+dqxrtzN9nqGg1epXsD7zwn+xRPeA07X+UcPz
nD7++NlDxxuNw1fXv2qVXtOV2wZOxsT5b/byOM4lqnet+x5FE9/usy7I8TuaMtNJyQ9fEJ9BJ6nL
owGMp6EcNa6inkpVOXuHDHIBybIqdwEmIsqj3l/tEJuzAeQ3XsSfleRF0burpzV80hjTasOSkyXr
S1Oq4I8SHnkrAlWYtoey7Vb7jUqLvzGrfAonJMmh7sas2NWD+MbaVM/njnTMuJ1LfsiD3SkImIA/
cv1FnXETbS+wQwPktQ+TyGhD5dSyBWZ0H97yhY1lJoGRQzG1gmWfu7wPjhFpv4j6Ia0jme1/Rt+G
N/LvhIOpea/Pcovxs7467SJrFFJ6ROMe//ztl8amsM1IInFbhOLLCWbI0yuutClBdvOMcIAY4NBz
2K9MD9+4+QyhwiokY3u87BZOvSlix6H5ACFq5G551MZDfsEEGElFpdHCS3qJUlCb8DV08eSYU888
y4rGzppdzhnBBU776pkr9dd6EGhegoZvh0g9hZmZFIilUIR+GgmQni3iOD5sNLYYepYnYoDuF/e2
BGKv0s2CrOFBj3ZOQoHo4sMuoSXfhFhikGO/9Br6IzMBmHjUpx6M+660m7hNfRUL2Zj+HXTrsk/8
sDY7/TwOeCNTw8jsFYAPMXiDPzMHIqAK/EafGSBjhPk9061ogR2dIkpER8gDk+WGezGRq2X4UYyv
j4HfWMtJn4IIris9rYj6HtQLZnIqV93QAN3JxuCIHC8o0mG4eINUrRYqfX5EexMRGzsK0+Vms6ez
IOgEcW+cQhgbe9OHwqrS46OchmBSNCrL6z+wrDllt0Yj98lUKxrl8CaET1KtkilUC2AcWS0/6Atx
h+0VucYn3uwCcexMB70GM7bgb8wfNKafLMdoD0QVZv3qgwmaHyOnk+z0kOi0i9YyIvDoXckz60ub
DC83OPmQ97MhJDkUB2Pw6Pvk64fyAudJR1kpOKT4OaIBprinAFaNhCxVTO07Lv+JIEbc9FIbE/OY
OBus0GMvYjmRWu20rQIY8N9I/Mr2vKn7hnXDhuMRyKKzwiQXp5G7cGKNzB5ep7jw7jlUl6oBmgUL
3wkSEMiqBLssnF2kvJXOt2HNH2+6HnvpPBKGeIThT6Cpk/pItRHeF1VCqjXBocsWPEVOErNvVZS2
GAJ5L7MdNPR4vlE4HFyremdL9/Xdulzk5IAxsf1fVYYaywui3b9udKHS9MfDzQlnbt6RoE+hYs4D
aPjSqK4S4il9g23IkdPnN4uVSuSelF0hNzh7krcopi0TS8OSNpxeci1WWXCzJCmJWYmtVbGEsPV1
KH/2UCUX3zd+x/A9VFvdbUw/rVB/xJfxF1wfgCzRYEf/NkSDGlKB+a//SxuK3YI6vSGjebEJmTvT
S59q0PDsECD2blD63hNPkAkOaEsI3VkSAIMCYouUTMVMqjJAlzQg3mcVAdxoQDUKSnqR74QqI6KC
0welL21YXTAjklJHFnP9KOAw+YFDx5QdQI+4cbEQbCLlO4wB38WI/phIYFTI7FOzx5Bd5X2mfERM
regfvozj8nsjaoFZc0EQUjG4JPAg0GFKZjNtnVixRTPaNcYv7musbzocf1tM6ffa0C7mGEfKQG3i
ECL79Pcrv2PMD88sXk9KqUDz/c4SEA/41u/2AWhKcwze/ENSG466Pb8oK0zyK43Ec+mK2qpTI1vB
mrdFj/anEPaGJ8QC4+ykcpM3tWuGL8SJn1oKjHW1PMNyq/M3r2Ca06fBiaJ8+Mnt3cjkk1ANmwT7
59kXSRdNZMhKiaHnm7ZxEMW9IPfa74AbYS2MwwkeD6m4dNmAbMFdowRuDGZ6pJfh3BALvUt38VxF
ggc8V0HVeMLnmBEA1FLpJnHmD5ZPSJC3BLfrNa6Kl9puCutNhvNX3YMaf4G6Na8QW+WAsdw12lws
Pd23dGQc6Ia0oFSzdH1axMMKoOTKnRPkIXh/pN1ZyN8T1yQDAFFmJKRp/8sTfOUeoEHO4KWs8iBD
k5RZBkKk2HfLxi2cnhwl1GCKIGakNqeYqlL1zqIcV+nJaD7AsD3+vmb7+QCjZ26YBtITimHM3xfl
Tl9ChOPHp9V0qmt44faizoFEg48yaew/b4xAG9k4fa+jjCsREB8uzLUTBQHRA3F39XBYvgp0v6ix
rk38VKaTggEFe4LXuZ5assV30Gvx4wP81xiWAzKKTVqsR5rT6eRrhwustRC1Q2qQ9q3wrWXt/Gk1
3Iw+LSqaZ4kHWmB7qhS63+Oe7qRJodpe0ZusTaMwPQhzjxXN5dcC2EspBjp6wFqYcFgo8BQkeCJh
0Rm95I+YCKsiMX5r59RX1Xc9SXgSoL7kV/RMC9oWO/DYoThPF+xuqiMqM//J41yFM4sq2TtoZE4g
0nytKBSYlMvMbvPQdNe7rtJhbssGgqwuOttoss5mIKLDXFVnz/i2b/BGgQcQ4XBD+5zxPWmbIqwZ
CAp754Ph0IHiBRRC2xjpUpN8G+vX+esGyQNTuplbLly3RsL0+RQhnYSYJQs2dsZ21oXIQCwV7L++
9RJS/NNm+W3hvzawO6nbjVFK7dQgsP0dMsBTnGwZxYYM230mPDfhhqDWa/QYQIsoqQOC5hXLe1hr
Zwnz5s2/ZjpWZ73Dgilhw9fMp1Bmi+tVu1UMnpu8UNkcUkbR8Rw5+VW54AtPyB5crnPMKKe53Ldp
NZ3Q0lJUQlAT+HChEKQoUHEyJigX3J6HFTQ2XYxw+0GVeXv2rSRN0iFbBz0ZLUZIaljxe9iXNgwO
qKNTa8p/t/8E08JVeO9UbREOpPOTebXCqjq75XmG5fz9IDkuUy+k1sk0+ntBsTCLrG4H/ZEQlY2m
FSIbcAKONh34XL7NyGTrATPleCSuPABfe0t0M3MGlgeuplolfZoVX6KimPwdCrXMl1Z4fobPnbJE
G6B40ir/3f4CWSykLKYwZEZK0r9KCMuYN12gKD/PXg6YhiQTAJ9Ph3PNfD5+eCdUnvBeFMC3ffl1
TuLGGW8m+KhzbrGJLVO1ztprHMIQxmLNk2jxVFlEHpjmmZ8WtCXhrxe8K46u0G3cc4yBbGNbmnUd
3mYL3VUU46vgcuqZU7noAYtOadEYFf/PyfVARKn4blUuTec5zp5ZT10gVCq1QBa7GjFPq0TwdvJH
gTjuCE9h9508KnMZV6xxueQxbiv3SB2mBs/GAtd80V75KEXK7WxJlR8FEMvIrdSXe0jopb/YreHW
UBx+BEMZfYZ/4r+2InzD72qHJFuOdtCu4SJw15mVNPIAR7ycoZD69bMWtz/davyw6MBOzNP7bIGD
BdZHPwh94b/HaCoqA4jSu84ik6lw5FJyrXlGzl/pLk5GdbEt6D8QztKgvbMTU9Ph3kQ/HLH0wBWZ
DSRwVqoEMG2CXA+zu0fyfiiMmWg0GAiubz6xvVCWm6AjYppTRaHSiqNdD+JPJWXgi3CzYIXF2Uvx
ZR2W6BFN00ERSrN+Jr5uXbhGUdaho4cwPUY6L02hV3wbiF6pmnUYXF6MUA8VmhdgJWYGcfi/87Mi
u9eQIgwb++gwku1s2vLhXqpHohRXnqdZzPIS2ECmbLhtcyfif34HSbcg0w/6zdDA7hV4ZuKfk1k8
bygww/gzCPv4Zl5Bvf45tbs2tpBwH2BppleZNNifF0TlyTmBTU+sNRuQHQ5TTOTjConfMThtuNfl
lGtXfO7hbwiIX1rGH6eKj40eQVgXaKj6WBJ3RAUeDEp93++RvW3zrXlm5yjRM3SxggIA24aizl0V
FPENTadu8gFUp755iciyZ8kZQnUxv/1U5uKJDsvogi1m9mbq0M+PgtpMCxtI1TuukeZPA35yyeUV
XUQ/jk3e/19/+oSxSMd0TKvM9q3k4XqpfLYrAaGGdRDg1yrJWeXzCH583glrL/+HRKzLDLjBKSbP
ldXq+mZkn3lO+a72NMY8SElNcVCYiXUndiVFW3lw8+2d4B7g3FXyF2kav7saGPL0Hr8cGVT7bIPL
9GnhWW5D6v+OA9y1XyqMWS+0XGUrdJrucz9bNzHcVrdhSqjD17j0ixQlaeD0XaMKETMs8FHS+ukO
GvOYKYiwDcu/ntCmLg+Lh1XjXZpk90lmKBOibBya6ycjUODqbNQiBb47iQ1RaC897jJALwbblRn9
96NIEnuBdPvp4vUXqergZlTmqkIjLTicHxgMt4XeXIxg1duEPss4Uck/iH1wxt8Jgadw0ACE25U5
S4Jix6qJYx5BuicQSsuFrwrwBZVZvi4hi+f0py3IrfGYI/XwiWeFvnF8xsC3YyJXVtHB17oCb6qS
G8Jt/8vaZrovGrb2t508XpN1C1SBDsyjPbnQ8+3GxZJqToNTeBFlssukAzs1061xZd4B/QvVBzAu
QIBX/y2oaIdEB+Wb03j9fAnG/AT0kSYAFVn8+ppSBmHG6Ji2lPdGOndIdBxccuOdWZ2WH/Vb5Eey
iYVLAh6+UsAghYLqX/HIJEHvp0tLD11WFPpHIz2lCkHUoX9ZPOrSkpQKQT0kKaK9O/AydETOPxNE
xB59xFCV5tP1Fluc+gjKvDhq0eyl9HhZT4dlB/SAhsZoV01stwX5CxxvS4yv+IM00ozHykJaxDI0
1fMDTjTuIQcmfVPcSgQyH+oNV8z0epKIfbPvWSDBqodRWx/jHYX3853UCn4wfFNIhMm8eoHv3bf1
PFjaca+vYV/DLO1zW3P0UiK+rRzISQNlp8YP3p01RGvOGCqeZ4wXQ5xPMwJvfrdpKssk1oLIm4D5
KnsEbL4HIPHmMbdaisvJsIAxOxh5PqRHPXBWW8wsIqJ/xpDe4+kGbfgbr3hWsGdR/68LZNzzfNIb
cSQRZtu3eJQIogd0aagJhRKJ1cbVjgoiTzAK1UHDd3FqbM7R4GFCEhwBDLEt2sxW3ZR/wEhRhwUG
iT91awEjJ8FtHlsZjy9+ijZwxWV3lwNOUe3V4Fg3vhh6s5PzDzxYdo/jB4MAv7YHSOXFgUkFM+Km
9XviAlfn8Ae9i5znjv0HvSAyRrP4NSff/edOP2ofd208wuoFnzW4hYAhLH9D7CenvQFD9bXfbnoV
0DxpgSz6VwPyT0khZblZUcOLI0m5ok772FNQWAlILkDZjR4lDk+EhqvpdZppQbqKOx+fa/PAe//J
57mcEnbUFwd4Xb0s/TiGaEhIxJUxzu908khZOT/gIqUk969HJ5oqHsCG4AFMW6QMoATWqy7uN0jm
ibxPPXY+tcQZLmW3FqSjTvwPNX0YjgbT77lYAZj4UWHt+CgkQeyRKFIbht4uxEb7dxAnzkOiyznj
fU592oLF9ts4gJ5zYndYQNkskE/pB+lXFT6ke0LQa3jRsUyZ7JBap6NqpyN4FKT98n2Xv27F4osr
WRKs2T6JEzdC8nSdS8c3Mkjq8J/yZpFNBVJtqf8J/swr8d2t/eTgRxnRId2Q9A7VZFvhVCta5vKV
sKELCoeor4fjU3VcGO0Ug3266aDRduDU3DimLOnCa8E9IUvQbgjAtrqO13dd8eBY/LVRnuF1wnbY
EQq5LzHgVyjJ7rJQEG7sXbvbYrbxlduVUoJeVOG0bm7no9GHPZBdIugbezVnOEgfNLjjNlPVKcgj
ar+EbLHjZ+tMcBOe6NX5pj7gKy1zuD/4BPO1ITiuXUwAJc33CQ2D7ZZyl6Ppphn33Iw8P0Sz/O9X
fXqj8Od9hZ6WmeNGItUN3vepzsDvBjUx8lgZZ+1xphp79CyiOgqCuhJtw+M4+aSVyL5Sp8uvT5Zv
Y+fPV9kDafT8HQscefoenL2zOL6+OmmaWY5DlYlX4ClKehuLCdQiZs3x8NIGPg1tMu5UHPkrsAhr
3Gfck8mBp5Uh4oFMdm7tCi2L4sAE7/+nH+Xq/Iip41Q/+jxqT8c9cExehT11SqlMn+fZ5fPiQ8X1
Ops7cBUGhfZ66+IVxeQZb6YV3k8U+vjYLBBTRldSvf9X8VerhBDH7xPkdm7ky96kazZazu9R328s
/NlVTjDAJs8J3OAd12BHaaogNrjTWbWeJX2jtcTQYE6Wr06PN7ThQRBBRoVQwNa7xuClo6ntXoiY
q/JDyYXe2qMVRpEr58yUsZm6T3oFoc2L//7inNlzPaFO2PpY58dcNabU/v2h3TiZPBwnLdLFuE2P
8aAVNn0usm3mI1UrUEhn23NBT2ndxaR7M6G7ltzkLZlcUUosQMZHAvyOKaFYAoEk+41aCMFZurBw
XsIxH+SzMJZG4SsNmgkWprFpJHw/ZDE8L2TzbwDw7LKo1Rzyc6KOMu2+kPi+e4aJ33rT1TDcA9vy
o5oqZs7o2SpfjilXFuN7ukgA5b6Px5Dja6Ctg7OQ1xbZ/HFfJ5PtoQvzmuVFJLBRJjjwXjct6cCF
PSWvKfgdm7wLbKLI1FoAaJHXvloaec1/23uotv9vqgR5qETdXvH7LR9izoQpS77mByYeGRQZKQf+
YLXy/NgpeMebN5MJKTe4hYYFPD9NeuvOl39EWMBdzXvL0LTdK7OqTdKCEVVqZbtzYd3Mp0s/7TEh
0ywTi0w3K1CTeu7cp+dFuDy+47D+eBxXZE4zo/eo8xSg/xE0hm7L1AUafE3CXvJcMTpBBbcxzHEb
3Ucn4Vi7CfdzTL1EkV0xUFNJAja+dzD1NTdz6YdaD92R0cSDUmd5pSacFQxAsvjcMaPqeSHPJxNQ
yAKTOQgHSDpTKa9blgGuh9gYMENA5Pe2AkUl8XFz4r+9EiqFisJFmX73vnfl9KOinW+uxxNxJOaV
0VzRH/j1AjiB/H5Z40/xBOwN470QGT6he0MagKyhtHqbEv8GVWvQ36AHA0E3e2RQo9MlYHizuWHg
k40azAOnApLD+CqH0Nq3EbxDXLeAy6fl3p+d0xzpeLSTXIuMpmZ+ZAWMVa46Rxzs0+IVgsW8UMdu
A2XYfYkOPXgO8jcjnQYc/XT26Gr7CrnBEaLLXXachpP/xSBDBNmpNGGgbKKLKRyNb9QCgxVyqYjC
SI4/jit6SMO5paVTlbjwjgGfY+DU1bTLZXWFf4RwiJ0OuDxik02UU22GCMbtpaGoWvs70mjQP8TZ
hL66qhdMchfcPCJvZpJs2UKZyM0lJstHL9ODuXqFFnRo1gpu65P1cFSPT990/MvdUcAwvw0b15Ik
IynKvDhbJHg2cYWR8zzj8GafuongK/9JgMy++AyfQ0uXFFZ+DWW4pKV0OcDcEMose/D2yimlgKt/
cryDsaptL+PcoiowQlPvKywr3b2JkvTDvw3i3HRfT0GJgHLRIq2C4ibTeB5q6Rvwv6dgZwOE80ei
7cZl3qm/B6rxSqmaiWKzdYk5IkuvKl8SHha5FCO4DNlH04FtxewI2aPS3WBWBVXEhlRXH2qaljV8
wNEmXXYqIk8bpEslzdMmkKL7Bw/b8oUeES7Yi7wxuw4nGhyFkwH8C23okYixy6XrGk6PqP5S6dfP
sKSB20T+6cjh1C4mdASwV8hIjDhcNSxGIILxOijSgRNAZI8P+ltmFjMUKeXDdwXilaNKrxBtZYek
bCaAE4f3kzMQ+3O9QAho399aqFD9y2WEjMthYOsJMZSekWdoKtDl666Ha6xN6N4pn7UmrrwsA3/5
gRV0uVCQ1xdkAnxlO7oxCGwRRVh9l2o7SklL6Tj+V9k6Yv9upZ03Ufn+vTyvtluw1gGYEd3Me8AO
CpiNVhnGT5l0aZRVr0FHBhuIpn/Us9KgFReknL1u7l3l5z8v+CBG/BmzCIkk/QkaAfwsa+PHwail
4FLNXpKB5pNR+NFu+TeLWs+6kWoMR1ydRM6yf9Qwb1eipsw5dJetoeeGhrxI8TbmmYf4ch2boC1W
PB/wGdlI0ac7JPWFNnImBOBnZgl/xEAYTlF8/ocW0qDqsuxTbDWlUVePFHtA0AKW4u+7P4PSo3H9
l0wR9fhsv+GGyR6tIQpImpjPjiUuvx1U2rMfM6W4Xd1lM1yz/rxIO1PmXsog/2gtctY7WGSBOum2
PRgwgq4MUkAOoaD4vougOFqG94RmeVbVY8I4yDBkzpZPSGpfb2aYKbUhVa7NiCxkNgDzxibbwzDZ
4Hp/9MDIJFDduB4HEgQo0W2dNdTO/AyhL8awlj+KdD97sNw2RF51DJoo3iUI06Tpg1MiUBRTzesN
go2a7DBUSC1FpP4Do4LBIeuvhflN0kbykatoQhKSYh/YEefZneGU40HO8vsQrAu/BTD2dIIKBImN
ya2E0iTuOrYZ0IZYP2wDHHGLUYwwCd9nOOhPOvF5Amxfvazo7FHQodpQmCdNV8T+wYCAqn0DIBsj
tPn+4T5ThT4CGAW7MCpXZF/EsnDbzbVGkLn6J83AOYkqt34KxiQAZ741cwKVziGc+jiXH+iv01iC
HjiOpMHuy85VEIPoBgDztFi71bd4cDIDFuMsaX4WuzihyWPEuDTO5hzNznRqmYX/pqwWmQFXlmkh
dEkG1Tffsyg8z032602O1/rEL44wdDXADUDyt19410ahGNfE8pci67p8e+D7U7k1k78fsxwH9f7C
qr+clOHqbYMMV85yZie3XrXFDckHQ4eaxkRA1wpv+C5nm7JaA8Ob1+u/c0g2S7bZwM8jK8A/sxzE
OvbTyhNv7TT5RjSBt1PPgzFrs3jHRyn4yR6TLrd1qKT7emTEynXGDjQkMBuasZ1GAgM+NmJoNgAv
gmkM3AqGc4sBL1Q3qRB2zgru+6typIxp5g9nouVQPq2WpZmBWzSj0mdnMSk+AF0SwcmmpbW1NxTm
2ZJFVcdFoQirCxI+Wx27CWTRnVSLGNuDQ3UwLNnP/cgfKlOjwsr8wUTpVwISVVoDrAT7Q0sclDlw
GfXo5Vxq6rRpr6yjx+pY4st5dbK5/fjfi9bjC5qfoC9bUyHHYlREgomFQwN6g1mFHQT/5QSb/bU3
DY63oW7IMDJitn6kzIy+bGvWA67GCxUhNpPaiD6plFXygCVU9K2uvgW3L94VGzg40Zm+k0yMrZmD
yhwlKTMshrP1b1ekA2yePBlNSfTtZNkFCjgIg9WbnzxMHRPRzV8FVYp2PFW/afIloPW7y+sU6ZjX
ioz9bfZhoPCcrbkBxGPTymNP084k4EbT2hp60Z4QwP0rXi9ByeNFNtCTUcRMixlCnSx0GDyXa9+4
B7xkmOPrUUhPjCWIVBMba3cBqI+JceGejz6Om+pPIhv+YsFI90ojavc0NbWjEg8czNzaMuMFnr2H
MTlHBA12HBrUm6BxP8zXgRQ5yfz3GnpSle8pSpOdnyvUbB4U5nHsH7oeqJqkp3BKpAwo0fevMLhI
nUWpg+SFik0dEofA8ad+9OCKgQSlqYGc0doA/MeqUNjv+3Emef5LwVXIMKtZ+hTMXCt6TxWs4Qys
cqSB+aIybY8kq0PP87gpp33IkttA0/kYvwWZWsTyRjB3dlENRcmgELGiMPXxPSwFl9qRSU7r5T/O
eDUVGo8V5/X0wUDhOZFl9bmcMVjKDxU71fgw+f6JzZ/FvNxsiGWRDPloawdpIsJHQNmD342KtpB0
IvSR86Llis8qkxNYpa79zcu1Tayu1MMID49PqLZ0Fej9ayGsYAv0GcRnfWuG117NHrr84/3ox51j
agythWVvpWyEfo+0BOdy7kWTg36vSyEuCmPgU1X8DCVGxKQbo7P3RIvy1GJpjAZlUX6zjzWb9hOf
C6vg5SzmWzBbx4foD45e64vLeAsbnDaEOciEUp95EbEc953akI/TM2PL/CofQdIihVOLcN5Uxw0c
DurPkTGGUgLGnh/nzbd6M9TfEEG90RZX5yzsgBzEy2nS0VZDEdSXPSBIz7xKylR67woBMvn+cfwp
TTLqp37xmsAAo8toGQB8jxT1l1wylJNtPJ2h6V65MVY0RWo9C5LcnjvzYLU8chs0BMQ36trTxnfP
UOA8Mcrqa8BA3wQajdYV/fE1eazgs5MDdf7d4CztoEmw8DgxjMxxqvuKie6HeCWtHt10/YLNdcFN
0gEI3gClVCA+vckqOxCE78E7grTuab8eTVxPHkbkYgcAfiVB9qk7zIaooU2yZsuLvh7eb0VXf6+3
r0ikIFRgXuf+IiaF3JOmWT6SveS+RDB6hUNi1S9kWpAv37btdTGTeJIiMrKWzBO/9Vq0Uw7M/g0Q
boXEbXVz7EXeBIwRWiNNR1ZDu4aMukW25bcZmwu+PHxBg6F5ZDq50ejkzB9TZ14eC8GM+cerMmDj
P2gmSCgWqvqBuZuWbZ2ImP0mBj6UvuKpxahbB78OGAF8EZyfqiq813+5LRQ5n6JOG5mWqWLgIUsF
HrYObPFN7eYGuDFIg98di2k7bTHbYCK0yFWyZrr0foHVRIn0gWA9Ow8Eyl9VektiNACZ64a0ME8p
7YKY/GNvIgwJwni19fiZA3lmMZ+s4C/Zx63hH4TTvsMkk/+S7l4jfbeBKly0S2tmyF/yIhFFGoZy
RtC9TXgVX29lBrIOzyUkYdjpHDvYEh2HIeuOfp/6k+GCT2P93SRMBdFOzyQBZXvFmn9JYk39OFZe
ArKhh+46Op0WmNKk1NAfgIpvqqIxu89HMVwDsbIzMzG6q6pwEqkQA6WSsxPsuW2toNnVkirkzNfY
KVjysv8fXa7POKTxdAHhveDhsG08Vok4Zjnj8zBNv1OUr8hsqCqCbZUjjuzjEPANLX+oIbIlACKm
BsHfEkBvn2/QN504I0Yi8OhVPGontDxnT3rG/icSbbIF2aswPCbcsCHame/j70/R2iVOUzCKB/0y
yKEH7mTl3TsmbmTuJ10J0g10Zc26CSlkA9br6Rcfj5fMjsMebRi/k7B27VqFyIbEfkgFVbgEGx4z
RBwGbHqnp5pXrU3PKorRzD5hKSA90+5FXrjYB6tOgcAqPB/RA0WQ4GP3U9xQvr0bQAKZj75TEYg3
6vjet5D26DWREp8oeDFw5vrfd40S172OMkGiEvENGNaKJ08MrDyOyYgaFY7BCf/94W0UuXfU8DMn
/o5rfCwhh02kmzlLQ1hwVcw7M/OFb9cyw0SNAegtV1GK8qg5691Gskyz5UGzz+L64b6NXh+myQhG
POOxyK6aiE47gTDAc9fh205Z4UXc8L3yLQggKaln0Ck3H5NuZHCks7E7LnrJn8Fmyk+ESFyCfE57
Q+9SGSPNSvqPb/bKf3ALy0mLaBdGrExujMIhr2xl7pTJZFszJuZJKIT/cOh9+09eMOLgjk8ehvHo
lecI+8ZaA9K/guDrgH8aAaOEfw/xBR3YzDldtrfGrJVdKfz3uT1hsO9I0nVy1hrex204eR5qjvz0
a+59IvoaxZOL8HZSTvDF3zrTUnvYxucHRNrNbPoK+qmHzOXlY3WY62XUoIFNO1aOsmcgd9QVgHFL
4xicRL7hH2pciQ7QmXN9KCHHCnz358Cd+7EpTourNLqKtcDljCHtbQrL/XNDr9C0mZvsw1F6Ck4R
pYPZ8orCaey1Garn6WQS7m8cjoZp0QSMAhwEePw3RgoGDX0CPgsHAEjl5w/ofZo7GXMR2OvTXAQy
fSIrEhVPIrTFoYOjZqWhXh7RJRSK8hTo39yY+LUN5bOy474LjYLv4xLoQ66iLQ4GSZNDP3nAxBxq
ZE8lqZ85p2WymplWfbYyvcwKV4U/Us8II8Uj18c2a/2a7f2aQnoRvdPjN8NzGZojI+WEkvxzY+d3
gIz+cAZ5QnGDeduuyB84I0fiMRjnsXiDxOXDn5paEpV51l0v6kvFgHL02ERL7yF1Eif/e2aBotAr
jnFQiWKlDFvqTawknwXgOahaOQDoV76QYu8WNDp64G+/9f1ISNzbbyY7TVJ/+LmOLkSkcPyREKFc
IY6OQ7RFNL5+PkTYMiG4t/Z0WI1aIDSm/nKfD6pXaOykoTjhGUNo/oNDt+yU4xkbPnOzj42J32AM
WsCohzGZrXN0BMhgAIfeGHaDxuAf3iRsw6yEyhvs7lm3Kawt0rSueFUvRRjDDGuv7fKuqejG/8Jp
q5VCEQj56W/YbbPpeNuVaoe1HkqelEu+tZaj5Pc+tlK81YYzZF2XQlRFP9H4RK6E9gBGk67fS2bj
PqlizfKTaYY2Pn4wOOSlB629nqSO04Dfws9n+wwSm2zGE/lhrmnqH8Z0Hbm/T1gUhy7/mIQlWs5v
jA/6XIU/vg6DRHdNDO2JUKabrnr50vYrZDNVnyR5RnOE3CYfTa96kp3l9w6iRPSMFeSnh7lJD4vC
ZdMjBvi+oMqBNf65WKsZtZ+wqFnDGnzujMbfvXlHsG/GzMHm7nBHBpE4ld0GU28K0x2LIiq+c+js
JH5QufronsQLNTFxvO/ZAYF3p5Rf4ZB+cwpnCK67XlFGmtjitejrvyp/IuhV5sltsc1sW09bui0N
IJ/6AcoCA8hARWPYU54Ew/7Qor7pZhUVdbfyk/8Xv/LDwnQfrr31i/xmPCuXejI9rBprUVAlnRFF
/TaC3gjmBj2qHHDqLuAdUHrfJBEtEeOnq61KujHrkyGlfWYn9rNJxTv19MEUVvPp/mn1DYaEhNCD
Zb1UIXkKbc8j5GQAfoAc9J+N+6Kxo2vWmFiIKFk0+wts0G0IxYyqoDkxG9Uw4wssJmSPX4bvdrdD
KwFkt7huoBE3XhSGLperm67UfMiVJ9sYOnMvBQiV7OOF3ZCM6ybKpMPDmIDLEKaCIP1+taF1Gvsg
4NNzt2GbMkS6gb62MdMRGDffFbjk+BNXFpfXR48TPvHRONEaqBolKWMeR12BKB0Cwd55PihBQRIS
nto7pFeM0KN8FVSVvYqYAEfNXSyD3hO97XoP9d1DyhUmscrp50iMsaiKIYjY4nbQ67vU6xDSst1y
VixCS+LWIaxFuCC74pfRAPdFW+GOe94nRCY09z16GFZTFixRLG3djGxhfpBS6EoQt5/m7z8bBQR8
eNWX+xG+9sK1uFo+YRu8VL/qNgzFiltKG0uOhj7hxM07LwRx8/jqhgLRJW68hY3XwQ3pTUE3RUXW
/drTsQNRpPTGwADoPH3yIbUsTyRg+tHBjb0+VM5viPQFNVDDweyWz+3nz1qHC3WUNWc8MfawmNNY
jNitw/9Q/5AnKqKr5PvPSv1mXM0GRN86W/XrWhYZiimmeZcms011NavPGYO7izfy9pVLkdMEUnV5
n0BsKylncDnMz7HsW9sOPmlZYOewxnlS0DuQEuxJS/YMXl253XFAbvWvVl0FoJNbiOT3lcRioTwo
Lt6LPF21EMzBZp9PwyKvqfEG7JEvEiIbBHJmVx/okYGix09X4RbR1tSbH1XhM58mEm327t6YIqS1
HF6z/4K04t4gVuSzTvYIf2DwiYGw03SweaNs+FTNZFd/qm+djgFmVDgr+KzmjWKr6nbynk1vw0Uh
XBBMJjuVjo3Uv0UauGCEHhmPmClgW47El/We+fSi1P9a4Sz1Kh7+rRQ7qR8FCh4/7wM/oIYlwvjn
+fHCtxUVgLexGif+2NGLyGscnBsAdfF2cJij71lJJkpU6xLyfb6hzGWT91VDmKCBqix5ucgIUxRe
EmqjvM9Q7C4eCD8tUHCDP3y3fnRvyTxIxfOm0n7o6jHJTb0zN4o0jAcFYHcO7rLcbNJhonESCLzU
hR6YjG2S3RK1RG66HsDx2jTxe3+styEKdRw7F0K1peNS9ZekpFG9jpB9K7ML/rRPO5xTFezg+tJQ
rvtKkYI/taJ9nTBou0CfAgUqiuu/SXJgOmBnOLQViplXPWifVw1yOCJcv9fCiLqWEPO38mXFK9DO
RVBUJdP8gojBvKAJFoSdT8bpUNXtkRVhzX97l//gbb7W4013d81debuq8M+eUSanxGuTVmUVqM8M
slD8Vb/rIF+gapnNqlAQ0/y9/Ctf8tFVVl+rzZl8JRVExvp0mtUnOfX7BFvNZv8Nx7ZOnyiGGVfk
c3U5FGxLKotR5L4w3lVXvclvKgvnP/A8U2tw08Tdnl8OfagSGZJt4EN7e9eMkwBvGTce3spGJhD7
TeEHIudci+BBoNVynh0p1yqiFNIjWTzE/lDgyHdJpg2GOMJLoYVVwaYk2sFd5e77r/GGrylSa4Qu
3gBt3Sq2VvUefgS4k/BWILvM2XQc/tr3ZAan1/Wr2JWi2ZA7NAc2RasUSzbsBTLcxyDNPNocrg42
QDbuO7ULRFjFsBRIpqIW84WctVfe4nSY4t20hLju0O0uc+z5GcdwyaiZTvLBXEtEHvHWRXlJQVkv
supQrMeWtekZnsDb2Px+KUyhJZiVyKKUzDi+S37WNuCPZ0CWfK1owCJMY78WIwj/7bhNi6401kZF
ow8/KWE7Ys69udmi12Zwfj2AniU+gwsWzJyjcBrtxdjMv3zhonrPooRhIM2vTK8rmXQoIzr8udgH
7APzm52yOzXrHsbko2zej4kWQDZimiVwycjCXk30Kii6GfMBfTQ1ni7nMEk+Jxk1u+2qIS4jQt0z
EQL4Z1MIAtJEzWpG57fUl9OeZqPOR0KFUo4oSe6+aZWm6JIhMF51KycMCYpVWkKMvyUu31ymZwkp
nE0pXuPkBsIWUgJfJIHXJJk6akqYbT94yXfiIv1DlILKasifkyDCbQ/I0rVpGmTWocdwrIJ2iExR
6e2Rq0w56LYP8iAn6xwOQAE7s58qAHzZaKjm20IGRK3bf1uy6h8RSAQZJ0zhq5kYKbv1AXYDoQaK
qhHUoOkMbOyOPZgM/PFy43jKWUviSB5C0Th5B8Q+81zKWhlx9HIy5G/4XvbwhSXRddON/FelcNIS
uSKmQVxWFRFr2bbWIuEL6Upf35iiGt+sQBgg2r/2GKAAuBPcTHXbevC9I/kVZqqWoNpXasVjcAzu
poEa9j9nUb1G+//KRobVfLMBnrk07krrt9FH1uyB/kkE60BCSw+umPzSqJ6jowHaSYrH9FftOBAP
sn13JQuEkAKYM+TPrv6Q9dHmGMIhoSOB1KAE668cpGswg9iN6odiGmsoJYuqytf84EApq9W+O0Kj
C62z9aYEeLi9W1b5QU5+DSzO8+QUSa7ySNfz8bj2RhSaeIlgNtdKnLXSPALOfuFdtq2R5060WeYg
qYylUnQ+UyXJibxDrsATRfRfOhaxnvlQg4ps45pNnEwbeTOBUdkbnCaVvVAyQeBivteGaVbXVFuX
j8cNH9dOTl8wZuUR+fGYeImTbFoBc/FJdLXdrN52w9bic0RBOiqChDrHTujjetJbqT8XjptjQzgN
He1sxq7Ds22xGR9wf3OJSk0zl7DBn2zufPgFCzHjxIi52vEo9UibVaDy2zxJPJOgYUdYGo+jziuV
hPcxXrAkiiKGEITkkhzf2waaOIxs/FtJzQZj/KiPkbu/AbLPgxwIc9XVvplWai9ANPjnn7uNAWNe
xuypcz1Lq5DuZiGeNhB5zwPbieIAvkpDz+5mcVIA3cOHApjlDT4zxbkcuOYS9SJ94RLP0CuKyGEg
MXsBqiqneNDfpgQgvudAHh6xsuebLhe9Xci77E89ojk32kiZw80Zw80dd4g1GqKTN/X4dci7KsjX
J/kMT1krjuIWsJ/uYh7RvMO481Q49yajlpc0qzWfYpRI+MLGB+s7L1r4oeF7wdb6DoQ2lP2STq5J
0BaFrg3qrC2E1cAqotrZoFiBV/kO2FebmbUz2wAj6yZVZIXgziphrpyu9WYu2n/76pjI0k+CeXfV
i3lYLgmPBcRhQw8Cm6K4hlp7f2f0lj1X9ftL9X34/FS8VpXAS3RKHivxYhg4RMiBYCD+jVsb6VEv
sIquZDbJrtfoxzaT9+4DVSXb8MpaWma7N+II1Iuz8T0ro3vmu4QQOhK7ir6Ce8EljLalZ4895p9d
odobJDKOYX4PO4Rrn7VxMKn+0HyH9VbQB1wMsdOdylOj7V6CI3Bi51wnlm+Nmt4OWSOENaSpwBVu
vfVwcaNNYv4/DdyP8fH5piO3e3oZlEakmWB7aAOOy4zovw5pHW8RhVXs3jMcAvtVh0CG9mxTCC32
qA6K8zKrPFO8RuxFqEXcjQVpjsHRD+8PVNtOTPTUMBkL68sSd4UF2GXJ5XwVcbf8UN6CWE3NWMZI
Zvhrj1b3tWBdvzQzeq6QBs9OebkUkQXjh1Ct8IttO1Z/qkcPgmgQkkUvEEw4Q9GXq+ASPgS43d9x
cs4xn7WdQKRHw7PMsRLxoQYt7GzSxM2u/mt+zV/bCZoA8ZMBNlOxwhVo8LVgP6Y0F6JtwQZHHEM1
x+2q+PMgFzTD3KckuVc1w6+TqXjx5uUF5zkCXY+55Ip6HmB6N+CKtEuVj+NSQlBspF77kpXIUs/y
rLcFwnkBJojt/Wbov5rF+Olq5oM4iwik/1Z0CjCiqgTtqMbBurT9zn0+3Dv/JcKtY9UH2NU+YFKm
Be4rAOwRKdOYQ7gD7gAbu5HuFWfzdnBWVaqm6PtiByI8Z5pgou9YFaNImLWd68M9mXfL0YVgvAan
RTqLNRSH2TCggifcSyVsZwqrw+qySIV7x2lSXUderkavIOFeGPbwOhRkPZ1jTRkOnjw8fz6tYcWO
NZm7Wmh//ESgUi8kFxr/luXJK7GEJ9gDWhl9BWMq+/WFB48vCN68D4fUoVjAeadjMUEBungzPs/k
rP8LGfKvMKjJSAjc9sf4JA4ybXI6CiizQTZbYKC03z39Cci8AKySMArk9/SB24ECkPYXwjkWhdk5
JBbxEfTqYj183hEXjreMIPqqhCVEBYC7JC3Gkv1XqY8OGMOylrqJiMw1S/4KV1uvu3H/YNhRYDbY
MYkGkuFo7ve4nSOqtvJ7xoFTecfIULLvRPF5DucaWddpMcALNe2d0+/rcI9NgMpzhhvqodfhnIy2
ocI03RMPGh24FJwnQ39UNKx3GJEG1Tz/y+cqchQlDZJfyk7pE0RAwKoBFprgYCsqSwS5K7PcU1WP
vhvxsk07Mu2dukoC0IK5vV0NttwLTAs9VWIUPscLYYZOfSyFKfTSa4Mjs6BpBZljLqKLLkbxuXqS
qtFGgFJpQWmwGYCALZ9XeWUCPODY5pDI4Nj/LRGI47aQlOZR1PgNy6cHEUJQjb7Vv6wgQLtXwsM3
tqzGN8eFsmG12S2Dd8X/GyiYC4i4y7QXK+YlAU5xuWbRsVOlCyrUNvc/VJY3roA9jsy1Tp1Ytord
2KLs0i4/LQ0/vQuZfTHR259VnSM/W0diUu5rpey9+0KxDPzJ8vP2VILtJk9IlH9ow9ZxX62Ih8Ad
hjP5SXoyFKfUFSTcY4kLU/W3r5eXvoKbJdETFRC1q1mJbnGfQ+j8QAOS8GqI2O7zwE3vsaOaxcS0
DsQWckqmtdvIbmYKIGgosaI94hDor4UYc0Q6U9qsrW1urNn2KOWjjDNXBL7CPF3aVgKek02rJaWa
izrDiIsCj+XUr4JkppKNfigOtD0PRfA/JqqL6Y6eYWFbLqO8APvrT5B1QAKBYPQYQrIKb3yTbiyF
bhUZTXMtcXFUIPOUXkWZYnneRQ/r++jUwHxqgeGuu2QbfL/VE3lyznrr/2CDu847zAbRw4H4hII4
BsJQKk15FKfbrvodNRWQBFpvjMHX7l3WvIOdnO5bSaU4y4lK5OQTQAMfwuvtcEksW6w1iTpb4WeW
vmKD2jwktGrtp+rIlGQBjJpN1jp9ULqx2imrheLtoAMZqgQzdvAej5rbBOw1iPryz3Xy2T7iBlcU
1ET1syLo+qask4SdCPI58Mfi5dDjH00ZmF+bOfvr/VpYYS7We8NPHyJt7LjLFVTrC9Uanwv8H2tZ
y5FOT4GLlvD4WwPCFbmH5aTs/fGSMlKPbd1ao71YEUgESgV4Xm4PQm5FGCrdY8Eqf+uN8RLgNgiB
V8kmDei2A9Si7y8vLVGjn9nCDDnZhVOEyo48JkxRkTMUHCFndp/iGdPCWGcfTrIbEfj4DrHyWa6X
/i+DkMW3laByjDuvNJooAY2jUJPwRCUGs9FJwv1vxzHUoe2XtlKqCZQ0sFjapMe8X/t7Ob7y45iC
gK5Gf0qfqmyLJ3x96of26HrpEnw2NcA4x3Z9YGAVFhtYwTTicZ6tEb3HbTCj3v030bUsX5mQQ3/y
fpaJxnkWlAfg17SZ7oLbt8BPDMKPVbX3GB0sSKgdmwrfih/qDx3bH0cKYM23uqAJbVPw1R4V4iBl
ygmPk2Jw3TmdVzcoRGh2GR8yWkHODJjzSmbpOvOZyrEQmbLs8QL18JYOYeuWkeC7zta1GX23AbzV
jndjnjAUbzIPPGFfp0MzlGNBxxMCx7SJfJlGA7ttvv6j86S9aogNuPLi16Q0HJ9qE5ddWJcwrREE
4LVK3CpLs+7fbOG6OloO+uMWr1QU+ID7gmYcw0JxTap0567aAN8LVDeoPKUfolTrboNp1CkV6WRR
d0IZF/TWe3UQk/Z56Yv95a8tYsJdYH8dP/cTs/KNHvQ895ysE6AKQRnJXRtYm4E3XM2DywBJ4OEY
kamDVmUBg/T/s0mq4+PifQYwcnc4u519lz7F5zxb+SG7UjvMcVFAwhG/oVBWvPwA/kPr6nDmWRot
8Ry8PZd0Jjl8OzB24WoGXmjp7dBi/qZX3bV+Dw7gvfn/IDS1TgkYDWzV1HR9zElF/3VKOorDaKks
KpzGFQXIapGRFzpkz7Pdn+tNTHOLFG06oMZej0KG3ynevBetSj+wgS1qLJnlY4HhM1ijAUuO/+rp
V8HVtMMGTjlCOwhwwn9gX1WHVjCK3zq5OYAwG7Xqo6vRsjttkVRSFg8wCIMcLyygo0RXOouQJGEO
fDGarWb7mo1ep8Xe35BT/HmBz/u+BcMHwHqrbuzN3ykRFMTmt78WxKSHQQv6IQmfRJQS4I1fkAwS
iLPb2XUMfc9L+KqU/+a3R5+xB/oUPqF4ubT3tYLClIVrmEmnHWTi8lIzRqJfgMgGmrJdjd3+1jdf
KHpHNXE+OnhSsFIfUSPHz4HNo5/F7su+TAlSdRpNOS5L93EV5NI0it3BANpWjFfXw/kswYCkuHdo
DoMqwtoyyhwEUD1QaFQDZHusUfJnikI1u6rbHG5qC3TRjDimOWwD/Eo8mwD+WiuzDoLTs44yh4Kn
lVvmbyElN1w0Z34v9+LX4Kb+EXXxX83IFczFc6bzMgxVhEMUWA99/WrVnJcVOdENn5AhxX3+zFBP
/pLfq3iP5S+S3LjyJeMXKzwFO3lYTQfV9zci5EnQw1RbNcgzTfp53jWLw6Fa4EYhmUjeayqmYVkV
GO2wOWgWf8V/mCnMqJtRjoxzoBOvqTpppNkQbM2QCbdHF5nIDj54MJRmq2mRrL4EX7IkMnNe9b1J
ZUiiVeatbIdC36TUuVcQ43iYndb8woF7YZQAsC17ubcKw8JwKPJ1JZqdzjt7Tup7043S++kKaLnY
cVDUyJABdIpp3Mu5FVwMOw2WmTKFc+5NgIh3ONge4l7SvOhr+8UjVZU1Hsy2fT0GMst8p39ldhaU
2/UpQCXpVT3pf6648sJp/m3MIIa5FjWfZa7sMbL2KtGAGFFRqtN3HNf17TcivsV0rZ7lc7Rb+E7z
9+d3zVBnqeVqjvlsPZVlKN3u7IKiUf6Err35XAa1njhRHZnCq4DEcZg+vJk5e39QfoJbgI955ylV
8gdNPkTcX7YpQftwbTzPuxacRn1h5xo+tM4vW1IdJ7mHBeFxRwGhuhf8lwqJTtDZ1B7Fvv3eGf68
+1DRxflADmR3gbBfFjCG9TXheUHA0CYJHKXUHucy6AJbj6Q7os/BWHB+xzrWwb7vj1iXoAXhjBts
8SaTODRNfnx3MBChCn4ZnCJOUZ55gMNteDBNQofqHbeWzQUMoFr8ovfmKGqxTAQroSfQ3En1apKf
N1OPgRTmP3FRsxJi28YuOAK4qglgT0DZCD8kCtVUU9s+F4tFFWF7frUZMOQaiZ/vpXzTZ7GJJ+wp
rTiH5GXPt9MSrtE+UWzCLfx5GklL4gE45Ej9prrPQdS/Knk2b/kQC8b/SDdTVSJsIqJI+TmVKOis
WliSGFeWQ6Bak6/D1qlV3GZmjHq1gh1fgqLh3UZlAs/5CfcBFqoHky3Ym7NSyYVeqvHhmeoqbZyL
DZGT68PHBAlB42da2zU7TL5nEVCe/iu4kQWW5X+yr1/dylKYO4gHseSPYA9p4bG1DerOJRKnWf7q
OUK6Tno6iJv33wMqINsLgJfK4rSOSRWiHdS1yP/KOQDpBxlg+lL+VHyXgnlyJNdNq1iWehi5moyO
vq8Ue0Me/a58Vq18ErCvQwXIlyO8983geA2dzRH/aXvoZWz8qVKLMd6TSnIQhOpoEM0e1DUAR4HK
20O7KYLG93GAwRdGjjHzg+3XXoBrA8B1coMHNKyvWBB4HA/W8o5Q1RXBNf8v9EK8WEt8DKWElGrV
hk4VsYBFXJ1Ljk4i5Z5KcyT1vRwjweP+MebbXyigkcKI/64ZEXKqm3w0C8moqFuxwDSmOvGwCsaj
pxSay63rcN4xKuBIrtDQ96jRoZXuJvFHfnXIJiOVpMp7rKu/nRU26ukdv6U4Gq0PF+mduVxKaiOZ
lUcjtFyr8iqruZbkSQOWzlp6WnXyd43pHAkF0ONkbuZzuRSLgwqQSfwpc8KpGh4k3VXmN0W6B9Me
ygXYfRe7SpWS+W1KeBo1BbO8EMVRtfNmSHCy1Z6Ujp4GlMs/Lsu7buN/49r7IDY0KyzzRQGgfdxK
/qMrkGHuqfs6iruBjSDpBDf5JMoRTPgv4iNCdPCeZYqGGOgxMwjP5FIoyXnqpS6I9QL5QKt2vu49
6vMEpC/PIMg3gtU/A6wFpQ6OX+IAX3dA9VpJQqPtH//RqZEF8X1wfVQAw5BIDtXp40JKDkIoRXdH
KA0pGM4HQeja1gBVkaRa6Vgpbi5G9IMDolU4/78jWaac8nxSWa7tVrv684M+R+UrT0tCtck4lOFY
O9SAhe372WhD+daOTDVLc10CuPQ24YjH50bZNmEYWp8FoO7cR0ks5zDRDeMDWM38SWFYvhlcakpn
yAEvf9eeHSNoSYe4gXSyLekUiYW2eaLJu9y+YtArE4az+ucjpImvHJ5EjHMvkIQXDF54QznXkql9
Te3KdgXhh9M05sD5jqyoPtN9PgHCZQANndbkhRoiLaOZRvoneHRqG7nl9R+OZx997ng/snejCbpc
UnbnGw3GShNoxsLLx8Zd8OZq8tjG9VeKhXMHsO591htbykr9JSvE2agTJA5hNXNhTA6tKIeOq6/i
yl/jizbCc0xZ0s92EUyhR+BD8iHeu5JNjWo3/SA5PeaMpiBqbsTAE/eJHAicvUPRWeQyV/hWBjsd
f6MUSCoAWGD2EfiL/9mANiBDExOsRCm1rhDS9ZvjA+58U/z/Vhvco+WzP7hv0POsH9DffeV2wJt4
/foQkN9tRtNwD9Z/gCGYqWy5G9SDTPWAVkVzIh+XKsUQsKhyl7qEasIRBkAE6DIsJT35yHKdf0F3
arAZmp7fuNCshvBaOE/WS4/21Ri/hINd5V3X4Qz//6s+sXPbW0wlephwTZvjD5oujRnCoXUDeEg7
aSjZCyKEVeyzU6sYBtkHjAIXQE4yod18oKizgoN9moxLXMNY6blJzT45cerbCy2sUZNZ7F+sImA8
fJzEynNt/myI3Rfvw4B/VWXuepjyGXgawtsvHeFDuyJco7w2VAK7pa1+5T8pAsA78lnxI3lfM4CE
JhpAxbRC9iBD4myZhbeV7Xu40cuQESDFYpFikv+q0Vmo4bmN00wmTnErlFkizF1pIdxntyTqOocq
Wnh6eIxF1ev9pHua2v1sxT77Ky5+q8EhUEakfhJ8EwROAr8kAJoBMHL72nhxEWsjOs3FDXlr3Lcz
SEWTlhCed7XT+fDLIjjKFjPcrmIPp6NAL1vve936HY6KTUaf6vPzv1rxDWF6uzl946CEdhuUpoTj
hAm4FRPumZJ+HVgzzgZNQYwC1KHe4Uj+NQEe/SYUCkm/3cr5UXeJaa6VABa5H8EyrZ/S/RYN67Az
Xanh4/u3xpSHOTO5tjm3sLf+Ou807Wlccc27MgHINOElGhWB3VnLuhu2JBxn1JBANzDGlC0sYYf5
c2Vbx3tBcDDXPX/F1S72RheZAvSk2AgGnD9Al8Sjc523YoBUb2WdHqaAf2hTUfjYv6K29+dinF1h
7SXq+gA0f5jRcqS7UhGNskj6gb0k/6kp79Q4TJL6YUtI6onnrl8Gzo/U/iZviy6Oln0w0KwLyQKS
RqYDtO96OxaiZrWrPWzGZYjJljCZT9Q31BBRX7UnzlDlqkDTzvHJzDLTRd4dcwJx3luu2wbQnFi/
+OArMZAW67EgrLq+Hl4CYf1l4I54iSsBSKYSADFNEgznyyamw1vKsgAz6pAh+sL4z2rE7+l8k8SG
KZDGVEGe0QVFATm2r9Bx9yu2DuNc9Fd8qkeC+xomK6TbQj8NaXHVPbwC//R3OwO+3sUZLH70puRw
dQjWQa+/HaOdYSqNfKgVXnU4YBFvPql8B9skAHvYw8jk1cJkcTfW8cMmoRlhCghSfUy7+36BExc0
/8sWZFH8lhtOioISvmvOI/GtVGJnVVjK8dkMQwEVTgTk63eVJYKgDCfNwEO2OYgv0F3lZZGeibA8
QW54cOZ+5Y+IYfUiECLHAiS2MdRnwoGQ4Om4x8+lB/CDx5cvJdttNcuVXWIq0/YDf+haYxlypfD/
6RAkMZzo87Hg96YFc49N3aPwbcamkBHNvioh2e2bBD1bLYaQM1821qL1W0PuVfMxADqtL0IF+9sd
/f0PeP9SXcmzRAJhEut5xJ7klHZtjKriG7b4TiHz/Hts5aDqnGhLCDikwzs36oMD4oMAE2L3LBp7
Ghl58GCr/2MsThcSPq8PXnrGSsYyVgHvY/+6jQYvIy7qVkGdu+ugLTumkMjVNlKZMliW25Nxbayq
ZCe6fRxdCc+Um81Osggq96WGYBMyZrG43jWhamHlGQkNSAGlKfCR8vba9cnLptevBhs2cxZf2XzO
P+cMTn/+An8a0RrSSZrywi8g08099r/FMKp1NkdNXjqmmf7ws4r6/oY4c/3MAg3C63w2Yupa8maB
dsBgKMKbn+s8sAG2Sf4GzFurKGGWZ4ZWc8GNgCiLHIJ+JciC9JgU24KmJ39MRoVOAHTeqAeJDWEy
BrS8n3ddFgjM1tN5YamYcY0D1ELMZWKkmWx6itzCv2BsEeJtECOGalg5zyPS4SVy3eDFutJ4q+AA
heylvxQ0Xjf0TDRyrV3JcYzlqHLMEP/w4HlvQhyI5dHaXohWLo4EGmtLXacJYkrdOek3Z+8Hg5Qn
hJDllTc19g4igMSc+K8L/EQs9g3e4Bhq2yU9qJ4kb92EzGudTNzvDRQfRT+0AzS5qZOXk4E2u3sc
aiHohqpjLJjna2ZxF3nWpKW/xxhYSBNnQ7xiGFhJLEu+K6YjaoKaFThrB3/NLxB1tWHsWvYdrgC+
TFdxQ20N0z6RMaKlI60LTP55XtoHU+Qq0F7uY7AehPQhi7mAe7RiJU6f90pEq6FYP8XucEcn8l0w
/pQY20l1rkQfJwWXeMxVi0Jhv1zWHsWP6f4Ynj+wFFWKUpxsi6g2UFgetlprlEbr1z8I1cLX53EY
Bb8CPpnVkNFlnKach4CgfZkc1BIpVhivLRuuvjwD1ztaXlEF6fqUB5wd2geJx5tDGdMq7RyL0dtD
nj/FE9cj62MQAKot0TcQLv4h36OqWHQ+yESNV6Ea8tGU3Go+4kh6hDX9BTfaPFZmsxshwST4neYA
+K6UBie0cNPILn95ZuZlkfxulbahK3WKFoRb5TXXN2SYDy9wJsm4KSqRvNLD+1pbvMovRE/HALsm
+PWAyJiFeVHNilIguABwYIGhrQRVoF5A10G0BcOHMhESmNfxTdbxEozZhZwJtnCn0sQA7dFV45X8
b4mtrWTGmY8YIkV4DRmiFNh5jmIY2/i99VPqPUh0zo3a2aT3bhwvCK1NnlFhGxBnT3wMqtl4I/2Z
3Xqdnisu27Hi6pf3C/celKZ4XGJBJIdPlIfODqvhReQD/tZHUKtkLSEyomglIQPsgH6HlZfgukwb
q1VV0O1WhJcdj541ENx4QBfSN+RkFtg+kzcxH1ZwWt5SH30Z5vwmLhAOxcxRz304gNI8O2DkcsPa
mRqcXej0vxcZ+sJleTp8LDLhiPZZaWX+iGsmB2puzGiAxDT2z7eaL47P6iRXiarXCRXTY7YaDa7g
1R6bYy9NhmV7QuAmonmfhObyrsnrIBS6nmvA8VpMoCcTwAqERY2IReznenCfBrdHMnxVPWcm/sOc
nH2AbbbuEyFZhaFGiRc1lNAxWs70ihSt7+xnnQmPLaB9W4qJ0L0ltxIHbzMNFExcvHIPCNIKQGa0
+/dvxBDtW2pIZMHpRFe+5Cc5EtyUSyTsCq43cr1QN7Tko2lNrbEwZEBezKNeOYwlz9J+higpUj3t
exC7InnLZ+S1M42TdLjTeIeVVWHsmDthw/ys7LfU1hLkTxoPzr8s/agVC97ydpBM2bVz/nk8fEHN
khsfuEiVh9KZpmAsBGjm6k6GjeKEzUqoR3cA9IL9+80uiMF3gHDqF+uqkZQcq0Wma+XMoBBHSbnV
2KBJCzQFUEar8CfqrGyue4ah3qm2v7VtvfpKZzvrL0VXhPg9X6GWcqEPyf3Y0qnQyH09lG16UnV3
Amlv3DqlsmFODjFCxiCqws/zAfhwW5gYL406CAZnXizOy/scJxp7zcBFAzztanGpmv9BhS2xGp6D
JOTvcSNIDD7OcGPnEMApiOjsuwMVXnvg1WmBz0lt7cTPBY661KAwZ1ryTAT1KFKWGU3JbF6FVOMD
jU8tcEj6PIkGpClyTSy22H/Wp1eyoVEc01TF9W3Uqn9cgRJGazEL/+IK69S9bEYDaO1En7zKNt+v
LmRTnZGLCOXhM/7XIktOdzlDCrVKdlkk7xjId6SUfu3qSTxwQOhxljOqXY5A21Y+oIDD3FoB0NjA
CK58B4UplFvaiW89dlyKDQXAL90gq/0dIlPHtUmqZK5n25JHywB7cIkI1zVvsL6Q8SKCBs8qaRQC
oPyKVvqzZpxpAv0NNJ2+4pYHi0hHJO3C/qTtcE2i6NuLflsxhcpd0zgt8leqAVJ5TXkKU4x3iCuu
uxSml8SaEt7FHDRvcO+UulJxpKF7fDX/7bL2L72HRxfaEjTCOyGbxu9wBNNYwBEmjD+Y8T25Hvrk
W5w+Kws7R40m9bhgbghJ+yRZUpXA/guNHBiurXFLYWs4VpHWf9pg4VDZT/kZmqD5FTC/1R0A2mii
1Ds6ZWBNzCLn3VxEA6peyia3Hq6UhF7EEQf/zO1jMyhlwjEuO3I2QHVh4gLxJ7zGxohP885HkeTn
1zxPKHaUYxdTtdyaz53GLWVW97Ck7hbou6XMT+bvqSP38jDhFNdv7o/F4qR6asv6JFaq7hNSc6hE
hcBm+NxrDcXLFtdKCakEgXW4eUZtMrIHL1VpzAOnrVh/T927GrILE5ekEhu5JFVWQ33oB9cLhTxo
Z+3h/2+fwR689UD4VjI/v7a20VBK+rMDLRDiUlGMQW2gJOLVzb5vMIb7sbjODCw+J7teLCV+rhUH
WEQ4ig6TVHP9EEJyyZVoNOuuKbXTHi+XiH7m/Opp+YiTKDkEZU9uas5pqwbufaZwEel8lRIvKOMR
+KDEpPzb2DPWd7i0ry3/39J9XijrC4E6xF35Ukb1vGWIIG+5rjPBmJ+5orowl2OeB/LJqp3NVC6c
axpsQKgHSMT0AHL5u52+t2a1yS4qEOna7O+00KklgqiVtcwcjyMoXBaOqdwj4/UMicrFOkTF2+TE
WrI20CnqPFlSbx7xQjbD+rfq8Y0+SP031hkYWsxZNOaxA9KAlMiadjJV1aJc3RCvgFEq/kayzZ00
M7edwzE5DvuAVHNwQXYyLhQ+w2SiVoxsseSjS26+RkZ3AYrtj+z5S0foeKCiMTw9UK6KpD36Fy+e
nMG6KFUepdXU52+JIWsMoDmjLqL/aIGD4yOmos9kEI0GASHIWowewWAERhfl5byIlbtu0BXEML9d
BEuiDF36uCYhWyp2tHnoLAeliSbsuTyP1FQ9B14pKcmh5M9tJKqW5OkvdxHjFuVy5/b0pVtzLWIm
SmBiztASkp7ctuRjZYQB+1QktHCAVGazYw0G+Lg7Z4kgsTFXRtlUV1V2bqJYAwAyX6M64ldrVsWB
5t9eHLAo71uhIxiDZBCnVjC51KoBUSyLIBpYJu/7iIGPUrxaU8PZBS4/T8L+MSeIbUn1FgX99spw
gLVG2Sr/CYIuxe3y8unKOduHm7odfN5S9SwwLOuXp3iemysbLajXQcjkvC9CKnpZyDeG/685aoD9
0B1Jdhh4f8Qfk5PE9TJTkW6MsS7COTiqvWLrrwGmQMPK8kqigxbfq4lOclFtCcjyHhbROmbT+gFw
6uS/MmGHNJ2UDFxhEbNnwe1mYXT9sEOM+ihTdk7CvUO1wqguuWOUSNuYy2aEeDByAX4M2seF1jZh
yVVi5+DBAg22WHMdYxz4+2bW6QbU0ZIgClIjPg6jeG8VN/9YZytvWtCcDqoNt4Py0VZfguMvbL4L
b0EjeVMQSZfM2pmpMLmk/7QeOYi1pLycay81QLoieIWKaC5/KTJRVekxbdXO2fhJuVkN5AwHW2fU
2/300O5H2S47Act68e2cusim+V5W42Fkng2rVAAf0ji/g3KwiuOEZS6BIgULWCo957dbVjoYq1va
UW0Wz9E44XhMTy9VIEcU8D76H3SCM2Zh3/+tEhR8y3l7BoIqpePP00Hoh2zIbXj3nfP/ymRsZvLE
JbDAuoVzyp3IWtLbvVR/rsNU6X+RkHOfwz6gtFKT7EIKfBgommAeoRiqYxYMRRagZ8ipj3m/fwrA
ViTlUIz3r+8FfvJjKLL0vkb9CI6ImtMlUr+Qb8tZt4Necls2sKaWbkdwjuc/TevZIkNZ5AdEDCQe
ScOet5mm3BOwcmwO8aSwjLZ38vtIXMu4OBR12RPIWoQBu0aZUmsA08LtkYSpOz8ZVVjbbXMQEaK7
RAYyxexgfdD59Rz24NX9grM7fAh71Bg7SGBc0Yie7+ArmsJ+GKojWLCLGW9QvBV2En7uDEBFwKwR
GKZsqrEjP9MD3Va6fLMpEy9h3gtjp4IZqMvBURYRpK6q7jgFl60NaBtiVW+daFc6a0knX+nyLRGI
RinBcsjbBTPA50Xmn10T6bvJ5pD18RUufmBZ4IhgD5WGGMjDcFEAr6qtX3bdx7Vg0zPVnpGqykVb
EK/YSsuvik1J0qBunuT+jfLYFHjb73w2SvxSk9NEv+6RJZGvIio4K4+mYUBUTS18MjZ/+8p67rjf
A30hfjT/7+ffuTN52KZRS5ACJPpf775rN+Us9cZdlyF44Ek/XJkUYY9ljxtbOj8K4gjw/1rQ1NMF
kQCfNDOiLwazLwx2b4J+zxQbqu5leqdRNjo9R7quJ5M68Yjw6ma7yXFUkwnSVereaXQxDumipU7v
HOEKBIkZPqfAM8mvt3InYo/6m+VUfbqSHQAUNujSIZNLMLucQh6et6WHqm7HOikKkqHvUdYJgzfw
w7l9ExO3bBwkMz3G+eaHvd7X/48iAz7cJMJ/k4GScwoCpfF803gXHfeYlUAli7HZZggMugR8+pZ4
n2CqhkjalskEE6bz1NWFkAhRfnkIx2xY4l7mxTExEXhGVbF3EfWER/wERm3RM7wFr5LDUKwbOsV/
p1WECnd6JkZSJA46T2nrwMVKOGTPOls1xFUpB4Snovbm5aLcqRw9ESCi6o9HZij1Jil8wNjU9xyP
jYws+nXWHe8s0ZE/69Wl/Fxe6o3GNSbbsm+nHvgyt8ZX4wQE0aaH6hmCKTNTK1ZLxZ8W6nKSAd+C
lfF+pvfFWb9f5eIsEhZeGUB6A8Rg0g4dRKVtNnjQJj3hQJD6xwDfM//U5zuqnPYHXB8bETQO0Wa0
bZ4SnrDlqfFyRKFLEh5Jahp+4jCSB886mbCVSvGff2jMEV7yGtOtmKzKJ/8pTj7eltTpEVNAtBhu
dCS67Ttk9xSvPbjsxKU5PPEWRKPXERFerGxA50iRVL73j203yFptZYPrlGigQqz3k2v53xDjMQFo
BD4AP6sgTOTmqXuITRlQEEyoDeocEb0hXA9ps4fNPvhdxLLg6HOsBLCT7elIVj4gZ6nWWVePdAin
Yd6HR6h45X8MbWnlPSQ1s1ciehb5pPF6/7NuBnsTCOCzBFy0b8ydF/lhw+IqW84HS/3c0B/TimyX
wfS7vJSmYNURrR39nB+HwsEAjc3NQDu1dP7JXDdKRRKYwxSnjOj++fpSmrtTowmLtrLgAMYQvJkg
LV/oVUsPp35DdmMXMnMumOXq7y7LpPO66OuqSkMjmH6SKNesCYfmLekuKTG0si95AQaz72ATsztU
ooEa4ZnFQE+AL+ebmKbMt4dsM5xUJufK3v1Bu/maqDHGGS8hJTo5InbM2AArRcxHo4y4mMP6fPfA
7neVFFWErqGkoBE03v06vv2ONlkt9DlaeXu/COulTPRmArqCDRQ8Pp1S3zdaNPxB+GzxE/31XhgM
0qZX9sYjctxh5819IxgBjmPg2OLDFvju9i5j7qAP4or9vFazJj0cYdx3cECV0kRUD8jsJC/W0Srn
i8JKtVAMJquL4Kv4DY6pSupUpt4WB5rvjEjiRdG4ORHueyIjTHkm3UZgaVcsK9lH3cOFEgsPScNO
bcbOpjOiVWDuV6M/ntWJJRM5aD8cEXXnqUPwoxr6XBvzdl6hVVGvOMWHHn21C6HsMvD7VaUjoT3X
eM3vO+YjJnRb6GSW8KOyN57S68Gyfqo/lpiL9w08DmHpKzEyoPd1c7R32BS2aNHU1bGcqboGkyCm
o+cVWPovMWpvHQG8c320A4dcfcK8zdM6njMVwxvXtvjnGazihFpQgKMMbeyi64jKKFrcANshvSbM
L9oGPUMmBwndRIqxSbuc4xl1rLtJhJd6OjNJuM3KpV/2S2e/9/uA29YBe7EiLtFTVmIBTHJj4PCG
J14T3uj02VpbqkUanDVxs/x2lUJC7N4aGrz7p2df/IBq0/j9FjZD4p7RLphIUfhlczpwGlFEqf+c
ho/d0VQAqYO55J9jox7c6gQmtM/zcSEuj25Z9U6Lw21XRw704cNA2oLmdwN5ZiG5FUoneJ1871RK
AqNcPGv1dxfctcwKxThgGty0/UJjChvO6s8fm0AB1xgMm+zIAqkYdEqTH0j0txN+FZMw3giaWXli
az7th/FZKLmaefieOzGw2rvfJmxCeMsxHd7lcuiXqR8KYzuR1cocBeqg1OWAGXEUpWBcUXjkFsZo
NcvC1bgeyQILrD3KzBmHofVZR4mLc9TbbSiCFagn0Nn2MIhmE8zIEIv4mLcQvIuKP50EJk6wq85s
vzNhuUpnctwDUoMb4jfvfulk4UCUyj3ruaVJx36XW/78510RweNILNnLbsLow0yWEo58CIUJYFxh
T1YtJK7ZlWNTk6KP8YXF9/a2guP49Nqz9N7zC6ehmwNIzVEKCB0bn5GQc6Q6j0ADDkI23/N/OW8c
KW3+v0b3i4haRr5D/rdj+JUhw29+OxDTYKUtFKvXqQelYJbk5TJcwbLBq/V87FwFFjrDHPGu4qxL
4YnBNlxSsoCmiLVzgYjfgeoGOxgzgaNkZZI2/rnx8P7CtaWPTTDv6Ue6DuRSL0zzMsMB20C0EEXw
FNiMCzVkHhnwwHF1wAVqjKZJ4qPyV+/b1ouP9rlfohy6EWs3BJQB+MKACx6d86F08vu/48XmLn0y
Wa3ljeg74Vq/m7obM3cFx7pzQb9XaSH888I7wQ7XEcHpmtE2hCl0LeRJnsxwjWJUBMabR+IkWfQN
hp2iKRz3lNxHFQ1DwrCegi2ABintJKartR937752FoEgAi5OBxIAS29aa1fUwEdJopoVHQmMSoAC
UIBcOR/Y4JG0mk0rzI0ey2tXCjQxEXRQYCe72qn3DSreCMDZLe5QqLQWNo+Rxdl+g8AxrSEAI1Pk
lVPUDzvxEZvTqAqg0sbpQRsHDx6+zE5Smc7UDMt2DVw8ANxhbi0d+CX6+bV7jvxPS9+8Hr1MLC1i
VJhzx0MQiqezITOSablIjFuRuK4BU34warK8P7qqC95qH5VMxc6CzwlxTUL28MQyHI/ouiB2EWfX
EgqfHDu96LKzFe5V5mNp2C9W9lVnUD4Z9ctNK+tC2eS0iJCsyOgDtuMFZtbh/D7SgudF0Al/jmTx
UD9U7rC146S/IBh+A1Z3FWfxQkVEtzMJUMVX31ejKS9VMLTgQ8Wt3QWbpf3Bcr5tJykrnAN7tExO
QamAmKid45T1+y5KpxIagQAwNjZhO0TrmCAzFoFMOKlPYz2FfcBXw/EfDpGS/O/jBBCUY/YU2wGy
Y3exK7+thZfxCVpVEeMTo5FuCNa1irfSsfUEVqGpQBWr503YBvxwAPbYDO3k4qfgXoLhyu+BH6wB
SyrsOWxmRe4Hpa5BCMgGJOw0BLW632RflWKJvQtili2Zn4MjE/Xu6LghirE8H6BPonI5+R0zKnM9
F3p+/dj6ag5NpWQi2Aw908gAbH9C+YWFuhOFn/MaIdhiCwZjbHS02kITlesTv/+o4AFKxAQ4dc3d
DMRO6CiNqXaUlKm1E0r4Ow1utVXNTsHGyHRgiCnPHueTkvO6O3z06T0vjitC2i7jPidQmMLZwrk1
cYfMOTREWc2Z7lk9ux3PlnPFuXKoYIqEcMBhW/MgVYtB7xOhELGO1mMw1Qd+fZKurFPVy9d8y3zO
F+XLJ6PdmGI9pBFnbleX3zZ6GyRIaShQaBWU+fG7pt9q2AJGXiu0+Fp7eWb+OA4PnTtkDzvp5dng
atf8QC+1bTO/ry7yoU1PGQwGrf+zpSenm/CKw2XpN2gW5znXUrpmoOyUpfbUjrFtGOCPRU4lb6jL
bPaWsWdiA5ZSVRE0nQKICCPrlMLcKFu2gHF34goGxzG2RQo70NuOaxH2hIAtt0Mjsg5Dj4ws9gpv
dBI4NloKcWrmPBGBa7TEppeT8BdtnpWxNUlG4ZYMdYm6BJUMuez1SADprwZ0jGI47RY89E0bPJVr
3xATkj/oSdYU8H9qgfOd8rY6AEd9rjHTwZaa8Te0kyf8wnkfKRpkIUEAg31mpXTIWhawL/oFJUll
s228RMlWmwdNOgrHdfPK2mmZS/WWJ0CaAbHSiWrAY/8SaPJPTJqB94pkt61vfa2ZAlruheuCFNEp
PpMOxm09miqnzqfbinaDN+keXaOuJbfPBaSvrtLH0D+AWCaIphQJnBi3yUXF5SzbPFpaiYGq+/Ym
5W7cyH3vGsxtpoWqfNs4SOz5mzR6jPU/tart1YE4AkkmEP7M2A0/VZ1qzTytB48QX/FpLH3Vz5Tt
iSlG/fDqC+LAhls79lDT/PZOQpChYB2IbPdsL4Vle5np3aaSZTjAwCQ38fSMYmff947w/N2KiVgb
s3luIB2px5FbbKuVhYOxlEEJw0DsvdfbpuN5u+tLfVVm/OZmw9bzQMikNB9kwF6hYSH7wwtKyZuB
pf9gPtPvlE3Nxs5ynJbdfqyEuVklgsXI74hc72Iu1Qpmi9uYXjySleGIUSF8m1XyER0dCa02KAnt
UIwNGB5GZ71aD67Rw7qVP30ka8yy3AAKnSjahye1DPCjjlKiBRLiwrFaUg8RNr9FRvRDf1nMgY0K
derag/gr+L2BXpHzdJqRcdIO4u/aXs7eTLr58njLYulo1IF4nDHSnCAVZtI6v2+0g1JcOuiLtIyx
d1PVoZDza7iY88iP0tvPJkBkbI2W1SQ/3gttKlayu8N1K+QEMKV328RUFaq7cYx0h5PWeK+93rzW
iAJyL8gfgvu86g2gPemMDUMGualUfAle+tY8z66u6zKBQkvrEGFISes4MzCVnbHV75rjgF9GPpk+
3TLpeHbAo2eVLTGpIfU+sxSNWasDfgTf1Mb6WUi6VcRR/hzFy1gfVsaodHV+DonBzWxVCOXZ9tFb
pLR6nxpGM9rgMj5o46S+i173hlKQ82/C6YZFrlp+iFTNIP34P0BxodtTDwuEJs3EE5difNKT7Qpf
UXstd/+PD9Bn1FkXnZ0L+HTbuERZ4TL+ar1ngLjMGVCzGphWXlZGeHBkX5mP/KiI2ISvXqm1heek
2fzcGo+HOr0FguKLr9S2XjVSt0jL31EZ5iwyNBImPuJnQqDgCteGbWMjoD6PeCqZjuPlZWPmKOVv
UKHDSeQPfD0pKKgiccTT0Cl5WtJ9QznGO+PXwyj5PHZo/88a50jxSiCUNNaGmI6JNd9VWN2NjqTO
th/on8N4914WaxcXNKNzBSvzejFkBzLpMFkCuXFouIF0ESdjWZPK1ST3zJWwot6/13mfSv5tGtuQ
NZFfpn6ogOLpxX3nMGL3mg9MGAdoQLC4czQiWyl9bCb9tfJbM1snMGoRyf8JJX0lr2+UUnnT53yv
LX4woEWMMhN4UbOB5dzvJYQr9XhuwzM+8qTSnLT/GAZwtg2FDnrjDdwHbXsEHeku8XSgPogQcYH0
b8aW1bD+LulzQV1U36Pj+w/HL2zkcQUOACk0iF89S//qiheuo8LaEWKPr+Y/YjvUuXi9zel+nZX/
XrUpRxFeaeCrSAEpC4FiAyVRyj2RyW3E/xHlpiqHWG8l+2bDcstO7pkVg3rOk1JRZQ6dskI8Ttsi
2oxiOhDzT1QSoZ4Pve3+2N1JVFCMeGgm18h4rYkDo9saQ//4vbmItzOIGtt6ORo20s/IL3xFNCcJ
E8+L7PGwgumnlUs/YN7CCvx9GTmKgAPm5+8oEPWxMiMfNaHbqSeRMVb++iMqkfa+LRjz47jVXuAl
N/tVgMhk6iOXorMF2C/hCs5wCajPc/kOGDQJL4Rb/tw/m1OuXPEMAUR2UIqq9p+oSmVTIQOZJ58f
ZOG5C4XioEByk/PdgGgzhjwT0cv5aKpkcwF9YqegXoVcIDzgxm9Cim+ex9XPqxx8nkVIXu/s21VB
fTrrLVNZfAyq+V/Oyxv2U36qiITIThUoPYD36A5d1IKIAvbAKE2M2KmzEOabUuAqfZKIJJyS8IMd
7vxvaaRX8W+l8FYpoFLGswfEq4wKcxcTphIumc9qSLXFCmKsb2PA+oDO0rdz0t1PkpM2fWQU5k0c
qTUxVyQr9p7fUpxID/SjDCr+/J+wfZUD62ubC0FiD0fFfQlZURA4MD4uXurCnnqwjY3JBRzu9nG9
kGMJjVfA/OhXrHc6WJ1zc0RDuKEWHqpeTMqnfpgUmdqBCksBi+Y6dNnanTB/slCBd71+MIyoxRlE
5h9755xpli7oEFQ0grFLywgjwSVkidwMTulcvjaGZTuYTv9tSLuu+8PtvJigZUjHaetmOQSPduDr
JSYWvMx9qC8cIjNBpYmO0E5pqB5E9ugOEjw/JGLVvLbKsMYjHieV+5pTS/FGYy0rgmftWLKGLt1x
7H1ii/GEm4ddn+H9auJsdQe0nN3eMK57ViJsAMMQnAYoOYjoySrPSRrceJ0K0F5pERewlqI97OTe
Kdkm/vIAF7GcJsJhOFR5B7R7JWjn3QlYocnvg+XEK63qkLxbUwen5ynMjEwtCoqX8Ow1Xi5290dp
NW/Sq6CSCyOLr4zOJXaTHGNFLC0wWZc3FvUC6F3vYC6rcxfTFA8YLqu9yHoUnlfpKGIVaX6H8oRr
U1hJdso9zFGGtspB/N/jfvABn8xGPS/IDLWOYCKVxj/Qj2MQSsOcyM2H2PCS0aym1LIvlRCVp6ik
zxlCDPL26ABsMlg9iVV9QllhITBZ+yE3HLLYYHJNVCCOrzBS6DDFv+C1qqfkj01y5K3yE26evTSR
QaI2ueagN90OHo0tvihnDEzJpRO14Lk0i9z3NkAloVXZLuwoG6l0bdAHGUkEh8ut3pN7N21HSSHe
nwrX0OfDDxkHxiAQp957lqspoAAASlCBDmZGjrAi1TgdU60wxaSKWNnOZv8Q+gsaiVz5hP8oM9lq
hLmQs8H2al3V1xfpM65+xKhWN7rCMG4JDix+3IU1g0E/qu9jT/5+HP74mcUa8BocebQl0oqIZZg3
JpH1R/T0WbDIUdk4RlF4Vg+PDX2WiTCg3g5gKVHrSEmmYkSrfYa8sd8xBnJiMAMxYvXH3AKOQEW2
ewLDmyNeXBrD/Ak8S7+Lxs316VHnLbyzFzSmasJsq6ccWsbrvqbhxMBZcdsWpejkDVqbhzw4ysSR
ySH50frA/drC9PVvzoKyg5a8sn9KeHQ0B0Dc0VLJB9Hb7UWA9Akas6hRyBtIwDOH71G872o0x5mJ
UV+h7Uc/WEswj4wQbMc9NmtZXsoFkfD50Vswb6Onb/r4G4zHukyENlGND0Upau4dny2SyuZ4EaGv
UIWD1DF4Q62dzXjUB+WGJ38ZRqsSQrPK0VPUaAdtRCZYTFFjn1S7HRTtwC82gYUongWxl08b4kIB
m3jqbPyyfm7NxPeTsT1QQILwttjzWlcCwADpVZ6yd0WvXp9R1/I2N0VA9/TjVDvHrgmD2TJ445Am
v6TXZoLhjkv8yXKQFNdyYXQlFbrznOA8X+FmgtJHfwKydTsCwmX99Y8BFgjXFO4vg1zabD3reOCs
wQlGy/2QeU8arHPWuNcMB3dGfGicvJC8Q4IGm38TY+s61L1c+3L9KPbfX5KqIMwDTanyesDvrwVL
cmBeFQOcPI10yQXrlM8Nfbbj4yWHtma2cHz58qvUm7YlwispYiPVdHfo9N5quwfo5Xwh82meikdZ
cerKM9VaNZA+7d1q5GyHEqtQNb8AORitHFr8X+WlMmt4hiexGUQY65MxlrkHcuGgQoJG1FkH0p/5
hCEjjDVK5ez08M15NXKA0Uqe42LTlDp5D3OoPb3R5QbgJY62odP4UKSP/zKSWz95VvhEc5YOwr3O
TnjziZD3nXdjIuitIppelzcgnwhI+Cmdw0uSh7wORi2nhzPFUWoQMbQOp4g6IBy0Psew3iCfs/aq
A/SUGvYFZ/jBwAbtk1Umhe1HEsoJjapqRnTimboHA9k3HTgvBtFEfFWZAOvRtA8AxwmkvFxao5dQ
DsE88DQ4ogLBi5e7MuLCZnGfS3i/mI3we+A//XqlJQ+aqCHK8pTKRmAkabvShjDM+87aOp9IW2/V
2ZEnZvzbmm6MspAFaR5ke8pMIweNMtUAIXlc48ipFvklFKULuxapwql3LzOYK8J47jCg2lO7qoxp
YWUGAAiuAoZIpECX78bFQaLW6CbcLDehlVx95CshEyMX26+81jdopDYe7jcPPjzuyC34VV5RMpRk
3nLM7hsMvTFgbR2pS6Z+NLXaBOeeXlatDdp43aLRyXcU6eaw31A7DPlTooTmkwDLvXcSs3UxG3vr
BrLeTSFUQc2+fqMGRAphmewvlEiWG/CoenSKWjKBDWUaF3mcwh+A/rdME5r8tbaWpuRGNYpozo09
lVSZGR1cltbVUtpYmWevEdHfBRVlzjdqEXTW67a3rEO4hI0n8vBhrU3aKz/A5+Q/T5WNGaCIuVbB
JYV8nyR4G9uaxTPlNSy5zAApGnkWGVlAzw4dbT8owuU0ku0yr12fzaAA6QFaLRkO9L9+rMMMRLPC
oimCZHmkNaSJaW2dU7qce4266f9ffkMTnhJENJLDm9P97R5Vk/eeJXcqIGxrMK2lFQ92gGZuI4og
wnDC7dESF88cWibp8EW1LLT025ZuFD74xTJcf+vTQaGcTeEtEOYdTZL2aIpyDiffGik6IF7lUeOs
0BwJ8FNuDbL45l8eY0w95zVU2KFIO7zmIZqvdXl1Ln/A5WxyQUIJAM9puAaSZnWVe+oxnrKe2zbB
vsR2xQ5BfpAZvX5Z0/8fJw2rjf4BIkuUCmqQW7K14TqEkoMsRScLnncBK3H4SekNLJV7pfQFF1Gj
MnLNNhTHhU86cCGknAn7wfqKgjjcpuAnYDclJz5LLUxEAap12J8XevxudZCFkg7focgiBAbTOPPD
pwvfXFiJ0FjINxV749uwjkZ/5LuLIUKYddHowul1PHpV49m3ag78l2mAN5JbWdML2U7fZdalmn/8
Z8bl6q+WNwemVXpF6fCw6Bb2istMxueqjDz1lGdEQnzuUwd0D4HROF/MQ2y3YQ4oCm9EylPzZYHr
EFK8SUs9ONG32XcZnD9MJk1lCdw8DKxGcu5+gIH1Zj8W7La8kbBe85bNKlUHrGl8tynb4uG2HTSY
a7sg35HQJN1j9H7A0S62jGVqVDUzSatXiWB78/DAjwEqm4EjESnlxjtDq1cwqgwsH8qSQgxskPvX
sMM03MZjpEY5DiCFYlnjP+3JhRzrT/jbfGFWddWHuYAbqyPo21ydQc1JsfAG80i9xw2UeXclHCAE
kse7NGO/c2IjfjiH3eA5LGxIcBx2CdVz549p66K9Zw3j4FdoPCSix5jQd0Fzz6IMqZ0/9yJoKT3M
QYQaui3fs1PMC1ud1IgoxW3CFQDiDhCpvtkQvjzYqhL1KudGZD3GmHFs/VKV4X57ccZq9kaHQjeX
k3oOf8mApGTvzx3Nop5pyYF2LVrrEv62hb1sZakA5Sd+ktfdtHEld6SIZEEQU/IrOgn3zvjlEwSr
GGj6YSGzbpuWxECuJHt4+rkFkY0jo2ROSjqSyZMUHeLNkLZJyKQ7qWQk0FvHlDAWtJANVX+jnVJ1
+YkVZ1QXVffq4FBUIA0ruWd8Df9wePH1dZjai6twt0vk/cfgRPtILrhcO7PJmgxG2aTmaUnHm7RA
lrjdkCxnHpktXb7kiWFKrk6j3nLqVsDXkZ30+KEeykEU2Vxe4vnDdfBmeMU8mbL+w+201lrbSPAw
T6MfZPG7U0aNgL9Pc9s9UWnLEZ19B605uXB6JyjYVpHj/ZRe/6KNgbi5D3mK+dg9UNfjKQsteis0
qtNCGDyz261woTls4nIbJLjLN/0UZv/qVktfLlzpVpRyB+LPCGFmBE3I0uDTeWLqmCj0t9xVA19D
DqHDkle6h+GfLpvcWDebL6AcMIKe82d04HmZN82S3xmekaFIhzveqX2+dGIQ8CEQhGn+F5mDhThO
/4DIYaDAWfwclJh3PO8TOjBRQM2iYstZQPgF/esQ49RFqJ44LDFhGNKiz7QnEIRDMaSFgvctzK2n
y9dUhfYyXjKwuDpUVB7F5gkoLgVTt60Lc5aLzaqSAp+oMDVL7yWiv5sqtP6x6etOA2/WQolEbABB
DSvbPbuCERUWISjIaQbSa4Tco4esrv60Qq1b2RaRPrrXwzqLxSJeUZyekBQhayl9hYWy9vZp+LJD
b3y1YK1YWxf2qN4BtyxRWGburf08CE85/LbjlOr7rK81kz10Mlx9eSSRV/JQ/kzJkbh/1Wx9c3QW
hlrOavzdbHt+0BPKHHRXFaIiRrNsIs0og4qgvfL/Qz5omtAZKRsevWeNHpuJDz6s6K9g6aMy/uEh
Ll6sO2RKs2QIZSX/M7HDGnm31ZPr5/wMM+1mCpNk9bEGaUz6jWqYbwn/fjRK92Dyd/UFMoPg6ld3
jE65TZr6A5G+Rt78fk/2titVX6x6Y82avr56AuWYAPDGbP89aPiz147xsLnykRnIBNFoBlLqRcg7
m166RtDudJlNeBELwQtJY9F+YAeyuqGS3fMOG9Txn1c4BIivQJV6xyXexI81HX0saAO973VAR9vo
giCxu8IJTSnPhZs28CdqylyF+yjZFNLdcMKqQyDYfKJnjRsmKmi8BjWjvorY+gn8TbVkfmqjGUua
PDWXkHrdaPMz3ORY67GerVlKbViwvEkmwWUcTFwFvccrKMcvkokaa1oxzoYNMFouO2v3pgtbyqhj
NLZE+Vhb/fXag2uzMMGQvuxMWVby5cobUiNVD51MDKfZz8DMSyJcFtjhjLSsNwlOgMEBNEUIrPmj
rP+8BTdtPeTY/yyQRr2YeeBiLPvVKML0bKReysIqrk3MogFQMsjtUFjjmPHdk+GcCea1SwRUlrIE
tYXuDxWAo71emdBgNu3f20FtCmbx1L+muz5K6Up7D4KwhYv+0C4xsvybSTmZsMtuXWyff06uC+E/
F47SOWLMWrQ/mw+Nx4W+cwCVHumTDdMgdnNyhhxL1v4oDW+Y2mnZ5AkipJ8CJLdf34djeR72LEtO
4PgEuGHBHJpTpSQGTK0ZYyx4EHkq32XuXaLgRC6oOBDSDHjS8mxHqRL+PdfHyY/Wq2YFJi8FG6SW
5zAAldjgSxjfiKwudAu7HRf8U69G2zTW+LZCRKaXFmB0k8nUZkGL9B+xooBLDCrJ988vWMA/DVal
wRZZuzB02F/hMApBrcKw7ZhxlULVQuCcWlYBmTMKQ6Ztob35hgFEnyWWZ6RgcbM03BYDnoQgM5zu
OhVSTYOh4O4n2TwNnezoXWuigZ9MRYf0mngwkvdWLRl6Y2/035dWHQqJRXx9F3j4EYwJRtny609Y
pqlX3Z0y95fDuHxCYgkmPYF0vBVi9k0YMUia9pJH7BLEnhp7OgDsoqqS+oZVJZtozLqf2D1xbrHy
R8uym2UBIDSrSbMh1nVko60zVyTB3XhHhF/HXir1+aJYJMtSRjtyxlF2xjHQJ9mpRGlRRWlThhn7
FLgiAis7qG5OUhN/3jdXKltbweF0PpzDwgTGGV9Sdug8y6T1lra/ebLm+GNq0T21kkYBMK5N3Gvy
22MT6fOzgxYprDftiXmKG5ouCXa+0JvuFwJ4PImt1WhvSG7G9yIffQHw3WyLahxSz5g7QxQVI4nH
KDDb0RsBEP6oK/mdO/Ny3CVGBmGXbmSQE2NVrCBj6nna1ASV2XVsyxwagJn/a7+Wbgu1N3JxUj2P
eLK3nAoixsjqqf04iGVlcDHS/TzJuH1OMLUoZA5brBW5apIC9ZIlkrLr1W7/pa4a6wMn5ClixhNh
t1oy0FZh8EP0bFx+11yBkQ4kC5h2S6Ov3UwcFyQ6y6rEoW9TfETJLYDTIIrKEjriDZ+G2CK+1Evn
MBW+zujzTDv2OkmIK9SGzaPelpmaDVvYHQ5q4Geo9x0HcPJjH92bbS5nTRyW/tfKlz2SIQkakT44
Zzv1b2n0oHb55bSZvyOVFqkFm9zdtV/mKOSHZBqRqsdSa3WMHD29Z2Nia8phZ3KHrtX3JqBvjW7C
/cV66eRBet6hD2uBC5TrvaAS33xgFIYr1TggdcLLLuuUnXMbHS88bqgK0DVwZrDTjtKaA38L7IL4
E2gzFwrXEV8ZlyMHgvD+/wRz67R0gkhoa12V0PjqgXIoW4mXSgrr6la4czoytPKDj3tpnYc620h6
cXBLoEM3ifZFUDkKesBykkTJ9RDhbca3ZaGFknQLCyXlmhdVH4IS7Pgtpb4aR7hIeCCLVrhMkntW
INAKjuUfZBRHK0mVneFjoFUUsdRMOw8kYzj7ueOil8izZB5vDsKLtZ43Hvbra5CYu2mfwD0WEqL/
ubjnOVmZ/mkXzuMAwQpKCO0Syx4Eup7kjMuWeUdbRJvKZm3l9xwye9+ZkEwj69+PRyktetjYQ8jM
aPv0OSPLZBtDmRX416VNmPpzTTyKOL+pOTkcvAru/6BrfAYcbXFmVTsVPrdF9mcBrwW1BIok4xFN
cMmfim3dVjBYb4AWT1La1oyuK7dOp25Pw/t+b9OvHw+WYn8kmBCTy2usp5DMBfFRm6i8+yv/U5XM
+P3PaOR0yF9bVpkza6XX9hqGg62JNVqkIDwcIMaW6pnlxLXYCxl5QAMtprf4Np8p+VXj1L+RN1eH
D6Lhh1h4s+mXLDTuY4yjJQW1/S+/lH4OChiXoBCdbewAvBZcwk4kwl/b1DmHr4ACSANa2X1ufDQw
5Z5+6xM/XNUwq4QZdwmK7yiiRCZUC2eK3W8yws5AuYw938c5tKCbrWWpBboPOXzX9CFjuCO2zeNR
HCXzkGs3mnvfdzF4dmZM3ug5+CrAJBC01/n88do663WKKUndnQMWOjftXVnexpd71rPUbfnLPGex
GcIYHXqpkIal5HMcMbvCcFDooqTzrLIJE1rN3QTsfK/anhU+7dec3E8FMHeGinuUOlboXkhUDCgX
sxcVKo+hKh7NkuZNKGlIKsAjZ/WLt2pOSf57DQ89bJSeleUaeENIsaP1CkOabj803YDjtHsghv0+
rIit2jBf/8eQd6QmYZhU+byzvxwonR1vtGknPX+NTukFz2YbxvY5S7CBYuIbdcUhuGBLVHpmW1/A
xO/4HxGDD4h5gT1cjJc/A7VKB1I6ih4Wyq6rpVdwkEyWgiszJR1Qprhfz0/m/cjpKTxl/OfHzayU
hR1NI/TnPHkxv62cdyFRkvKK2Mh48F2Mmxe7CYIYgYZkOKQhJvgkHINFEArsU4xGU712DNLpKURL
7qqrUF9qC9Bfv+cD/RxytyOiADbu6xywbXxJpDDjqpQ9M+6j8R0UOAcj2ayMSpO9eV+XqRmuKSnI
95dbtbNxyp9wGDNokRo5rgvEig3kYpjX3hO5np56mo+mVlIBXMDDcShDAF4//4PaqrCPfubgheuA
womEEuF6kwCsSOumgtnAokgu9FHSTe/9aF2R/rzIioDq1pcZYfkfFBQ7LPZD1J5GE2++xe8miSob
UYv80Zemgy8Y53aEMgvHPWs1iSd2DsIeuBa1YNew4ZJD68zC/Qrcy33aXFT64VsuqkQOqvx2Rnoo
3t/ydMKUjsb92CAEHR6GyYDl1COtYWqhlJBfus9bkm0TnbCjDITR1oE/KeXLhwj7h26QLDMTrgWp
pCKBmwhDanIkKYibnazvyb4Svtu2naHUBdHSCxzuxcbzU9Ko4vXboRXZy8D+yzgHGAxQxgmChBhF
z0j/AgsJBig7s42rkLNr/c2zUr/Lvcw7qeZmLllw1LvX1LsGgdGnE85616k36Mpp/n9wMR7BQOLy
BKx/usCgGk6xTupQ134Q4QGHcuHTiH9T1KwW3aU2aBvGgov/+8/vt/6gY+FN/Wv1jhSTgX0wVUrI
8fFEHTfr/cPduokcs4CXbRMGFTXjfLWIGRd4j7Y00MqO16GY9eTB3MqOStOjre2kfUKZh2a9zqYv
Vo+can3bD/wAyzC8zVjzaYvUa2H3WUVQt94mqJ9y9HQHubflYRsEZrFbsoBouuJS5TLxvnS86DQY
4MxpFGRxYUnUAV+WAP1fbPzld4lIh/h2Fv3RmRGFMlQ81vWdrSaiOVAUAqUd3nkTrDxQtIb1KO/a
/lYeDVtivvLN6GbhFvE/ySGbot+jaus97odWdiFUeq0N+vzzBUNwd7JlpGokmrtXvMfGW0I2uvLX
lA88USNRKzCl8ShX+cReAgzjjDoK4tXa9Dy/iLMGWBXT4YyV/uzmrKF+7Tz7H3HgXKWUPHEo0SIp
DzMbzRWSOVUL9g3XLt038ZVRfypJbVC0MLHXwkS3+8QFfDJXsmn4isp25yJeOecx9LkEBsi21m7v
HfVAAQUJiK9Jxxpxd7jj4oR2nWE1gfZRKYnYlSRqqUJP+XILPrEk0RUFyIttc7SZFCFmZIz1X6B0
010s9BdP3FIcz8EwQuqJEt+BBfK1/NnE9LS8Roi1HYu1eifeigFpGG3jjZVha4nbxrQ5GmN0SUF2
4Zb/jfDIqvv4jd5mxSPNJPVwh0fq9xSnP3GBcRRytBnr1sTGFGurQ45/NycQ1f6y25dY1Dwwcw1v
kh+TXckDJ/Q+SI6hUlWrHgajbJgiNwb/EYGwAcLB3V7nIhPuIzSKxyF2PUtKYsovdZwCE3dA9hqG
sDntqpD9O7K5zbsn3eExJum/TJ+FS4B/ei4yVV9wjFBmLeVYj4C1dIu9TCtnYxdwAsZRpaBkCfVp
7H0MG136PGQaqCd6z7vJI+fmFBdtRWTbTMXZcTvtDd5WjVlWTCU3JqN8eidfSJMqDDLN93/UrJB3
37/FJ8WPuGUNqfO0SuUcUFvFbDcwoz9B0WKiurFbLymvTp4zomo/vrhMchjY1N2SC7ReipbWAYQb
SmIPjeZEl8SpqBwlomLFae+RXg2Beyd2i0Ut4bZmXSFbd5ndOGli/3O7ntAuOzG6zztTXB7b76Ji
4oRXHEqLcs39dBzxi6xr3lSjzK+8mkH7Qn6KgiPIaX/lSQfTv+J/hOXRRV9dfaWqqx/qbojt3nWc
iq0uN/ff6zmh0him+wRZSrrlnTTdQ+uUhG2Onf4/KD57KJtFjEusMLI8+gcNMQo2aA2o5Gz3NVpw
vJO9jHsLSR72rHQOwRrf0OT4JL6eWjuwEDFwFQK1S1veTyo1IQ8vaYTrzPGCqR1NANCn3SuVg0bh
j+7/olMNyD9Of9sQaQyWkwo6ftiZY+NSwRY4gcdcQKQzpeUnFpJiZXPLMnd/kQQ+TMTLC/qWWcRb
2nRJM7pu11YtWIhB/7oExANLiHdzesj2lb3qn/5JKPK9FO7sWTAlZ4HRAvaRndVRkiR1VccwcLeG
M/IdEEzobqbXeF9iXLpLhuOA8KiYrmP7NWWF+bl9SLRtVNpB0hAP3IHJ7GGOGnJNDH3iygKEFZ+3
OJaZD8x5ct1cupci/oF6PYBY3aXCVu+ptZTBokYuo/db5c7X1p10mcFoiuh2kEYIG/LAiG0/sW22
vwG50VsbE1XrTyR8Ah5jlfKh3NaOFgJwpij4w4iIInJ1g7Sct/AP3/gO29Oc3bdG+4uf/UTOVzf1
RxUhDYOOATTHB8jcWL29SjqPa7L9ya+EsVcB8Ygd6w+upY15byIPYSM1nIHvKgpNKd+0O/W59358
lXwCiB/Sr0ZWMLM3Zm7hmLWlatTo94Pills8pG73Zkp2e+QcExEqmpuLHlxhx82McI7wP5C3ojLg
9AMxRuQ/Gni/yyQlsh85gAMUhqzTWYObdNHbxINFQL1ofEDfw0yEfnKIu+SXSB5e6T5XC5s+Pq+c
LE5SuW9JTannu1TkQ252Ncvcl4CxhHVxE0N46pKINrmgJXAHIzKzNxmByYjugGnRQgnH/sCS2hKH
6lWWSrVkuLKyQ0NFRGvRa2ifOgpIRABMxCvZRL/G5pxDkp/FA6Nx00hBIIgDjagkdpzSeYJSdwpE
wVZFsbfgzmydjfFPLaK0za+nYEGaDFuiovbwBj/D+Dkdw/yXBslT5bgXQwEmQjxFW117E4cjaYu1
rLWZQSvnK6LLa6n8ZsuOT/O9MhcZ8ltgINxi/31KYBWlqT3jI5s/v9PnmdD4hwQucocQ5LD+S1Lk
ApicmXHK4ZTG8r12uvsNFD1HQRWkenXEWMlyqNtSP6PJoLcuZHosRPtYwi2olcPkzZKQTL4UYmzU
UbzXUv+50rKtzIxaAcxHjU7gQu6DlJ5iULhMEs1MNQ5UWQhYh8JGQalu+jWFS2HZ0qpiIeMbex6M
LMpP9fip4MOUvEp1sg7TTnDaue9qCA9K9R9z3lMy3N5GYAZE+ecDK3m7VN6AGz1fb+wEg1vTYod1
z/MhsPbDIEXMHgrBtF8Ne8vTBohwFEYZWwqJSZRadIWPfF2COLKE6KZn1qH/icpnY2PQ1LYz6Vlv
VWfpyaDZ353DO/5fFnilsB6AixSc77OHUbw0UgoejXA2VFkbkZ8Ln7rllkQI6duW6KxC8U+ffkgS
vBRPFT42o84gMGFXh5Y3HRM/3FS9E+3fWhlfbQumv8llEPUHw6eNIRjNJpqZ8bjqNTPlg12NOjlW
ixkCgrp0+2mtfeOvCk9x6BzV20Zxw5bRP29mBN+TeSe8SAlZsHjOO9Kq2pQd1Ix6tEcO67PkNMLM
0S2G1fwPH1BCzlbDHl69xaSlGlpUCUOKsIJk0sWszYnJLlQM4O8XXWe2RimIWlVGpPyxvWWjRxTm
VE1RYnsi0tVwptJn/WHjOWus758XdsY3XU61dGmcYWm2WzEW2A7bV9PP+yF81YI1h4VMPZNyZr/P
XAq64F2e9etwMudeZeR/gYqI9WsQY9sc0nVyYw3U24H18QOlCzUC4QKbsB/YxLzQVreRmYGGRgRV
YU5UXotPsZTZCfOktAxVOVlci11vtSyhiWzXxV5qcJglPW3kpuJ0mtCAjLkUhswVeZeKAG1TTWWE
MAli58cINtddb1fepEJw96NhG/EaMTVTxncj3s7Q1tTN29KAncelpqW/36AOcQVBfvwH0zsXawZX
8sjttXK8T++8V4Srwz0rFTxeghAQFePQFo8hAedqXH/38Wxko0tv8LbilqSIGrNGD8aRulAQDfXZ
MwAw/1BgSjVCLV7vx79ZCOwINKKeaJEZU7qWjpeVjT/O3US1RojS4VquH5PGYT/avBOcwp/9xaN+
RyA0+oGOcpL1bJXw0k5VidLLVjrNT3BY31ZdoQG9ZwuhebSLdx+dwJicWdMK4QxQLIIFAB7G0x39
qXGEplMzKZedrlKqD/Y01FzZI6bY47jZGylTaq2d5Sw6ye1j3u79v5x8zffTN9rT4Yi3/E8rZ9Wh
j47QnJVQqkAtswcCHsVAi5PQswwLVwUUIBFcmaFiVtFOPntvxM1lkNaRf7hwkkN9ld0MIWSebUPK
QGQbgghZAMydDVY1QFjEHB0dzjvkNgXRWJe1bHbFYbgirBBQCs9pmFlPLBL5VbP2s088cmE6KURi
yXd0/JRg6pMb5nJ9aCDv4BPWVJO0YmYw3/rnxLbwMfqg4uNyLJm0S422FcSKoCkkVKRn6cpPCWe7
0Hh+5AatkJnt2EVH+4bzpfca/TYYT7otvVtHFQPyWIbiRJciEKBpwP7Wtmae/ZIFx7fDbMicL1gq
ELQzpgFuegPwefTZM8wbtfEAe6yDYsDAlqfiyntDskVuvjKLl4u1pBoBbmGCRSEXjI7amqUb3LFn
PHUomYR+AFCCTkrY8UsafTJeG6DNImZKGLeg4ni8mAsF53JLR/IBy5xqmtjygLfCFralaiViVVK9
xTIot7kNdrdSUiEfYRYOAgXdPP/hX4Te94HXuazajNxp6Q5T3a0CDa0Bnwvc67Cn83+223KllCu1
MGx0gDQwnIctEbtZ4xwRUUKvSLqExqTxry1RoQ3ve4G/eHYzA2TbBwKZEeLZr56KiTVd86U0EgfU
5H/IMkEKONrnoAhjm2f2rCLWvXjskynX5CW38ATjed5Ps/cGUuxs2Pil5R3tOrVaTzlsV7iXWKwk
I4Gms1ITw1hTFKoLIhQMedGFoi+cyggVXqGuDvvleLt3rR3wroGwYaUh+RFkMIHoHuyBvjoxaEUb
yfvOAN9LDtCZLmHBYzfDTXVIoF3dBnFnpIZ/vb1qbE/CD2FvV+2RUIE3xTgBgH4vpBq9AAHvR8Qx
Nhj9n2ddcS+AFdccpr6QgGwLYeePvortrix0ApCBqs4eEX/pSkcGUldli3Vb3QBtf3vVsCR8I61S
2i067gkNOUcTLlvP5clpYObvoAIO6FYotzWlyRNcuoAxARdo0jGuI/40m3qYSOMd2YJFCf1QH/fe
NuirxS9ECgqaLQbHxrbfU1AG+w0sQMiaGG3ta1CD3JBLHCKvU1KTRiKoGzLKAYeGz/1Ax/mGjOnD
RLY9FrPLgN6tYqgfXz7pL50gD86rPllwwF2HhTTkz73KXWoUd55FilA+GoZn33W8x3DaVQ1f1CkL
IQloKPf9XLWwPx6mDYDo30Gn/RpSDPx0UWleAahlQNiRrPgbe/dHC7Ar9BwfvPP/szQ08YiS0Jpp
N8NPw5X9Xi68hZbtNsazPyB4VvprJUtLLsP+4c9Djc0LRN9V+BXpDIF6SRHlG04kGJKl99iZ2jpF
+iBMRrHFYXeWZGwuy8ZlAV/mz46BLDjjczH1uUV9ia2V6ffGxXdH3QtknKdyCJD/okT/PF9/PbUd
p1fq7IlLALB1DSj9hdWTo7P+wXxRAhtseHhkStD2nBTEsm4MTyjE6apqm0IN8REWgSxf5d14rtI1
r3UmENU6iv2+Sh4ZE4RtmRDp+Ut8yD1ZDtEs1xFhdZvUi1jmr/r647+iAKHlCGWxvYo8I1eERnNl
Cg1C4BWoQpEDkDc40ubuaa5ObtAvdqY0gLUgvMmtqtITnuqhLA6QHk/gqMjSNg397WZfd5AF+oEH
bAGV4dKY2+kRZHlkqx1yydg6CaAuN6yNv6UQyTUcu0BsxoTCNOwRRNkwkoacpobNdjye5HMBWPSl
pkgyk3ur8qPD7qM8JXc/TmGHm4a5PT9F3Mvxk0jRlYN4SbMeeEsP48cg/uHWCMj0EeCgX99LIrfv
odehQPIoq58WcTKZPxLJFpa0c+ubTUl/FtFXi9Mq3qDTFDmtfU4VQF1bqzjPY8QSF+e5Nx6nHm2u
KfrYRBmjyT6WJ0hfw/UTfEl5wGQqGsItuXrOUpimdpaHQb/RtFX+3mV9+NiF3MpZ1L+fuVQ2X5gw
h4FK9r1KCRO9Hh9C9HFVTYq5dS+R+iltIvsIKPK/9IKJjoWiO14lB1LUG2ED3kL464UN2ZkiaZxO
EXyxXuazXsPUzD+AScdF9E2o6xSzxjwtnITW8FTdpUKqCvxXgMkRN7I7YLXOZrRYMuRZpph+SmNM
hbp7neGdlha8QF9ieZs4ahvuanmS8m3KlUzC2XjWNE7afJ/PkPGRng0l8YCvDBdAK13XqYz/tsVr
LZP2AlE/SiSANXcq/m8zzGWnsugW4I4nOXACHvVIf0Axvw6t+f9X8VSgtTaxnXFmcE9YgN8YG0Ds
juaeg7gmo5RnlshQc7JRGpEaGEopzxpN1qzCM1duZx1hakMXibOrVBOS8EgCI99T7kUPYYtNqWyU
LChQZQBIxRMcb7XHF14U7vXlr1Jt0Cb3er/wReofL3GnC8QK0bpx88F5lZK7qCWJ13kJKXBA4bs2
zFvzaFkvVRzd5yij8QDvauBG9PEPbTAAyVj2MeOjhj5MvPEA5U5PsJz9AVfX/Ix+wBcXcZS0AL6t
48WJh/5QmAE+03kEdtnsDem13ndz2bGUs1iqfRcO9+nY+dv8WJtth3FG/A52X3B5JNitZ+LUr1nL
+oeYNy4OqAGAbENtwg1KGuxT01+2upsQhwRrV7X6BbeI5JLRXDMPbD/zVL3HthdznKx6MfBd1Qyc
WfEtA3sjI99IvQbKgTWxE/7JLK6m/GTst/6He98XZX9g48vzOfDxLH9PZTWpULS1JQvnHcqZBf34
p/cxnibUO1fiVDLULlot5+ng/PUdDAnRvcS3PCGbRABnexQlVgu78/fWBWXru0bjCrEnVwDnTzTh
sh8usInAFvOV+GMlUVCtRsqvTeID3l6skDT+Cz4dh/p4ORl/mFkze4QMLXsBYcVVD5/DfrhRvvSk
OiXehioZlWV1JAbBGaFwF9RgGdSyl/1pVadeQ1qZKS+KAD6d+aa7IaZd0A2h1A8pTyCDDbSU/sHk
PCgQb23ts14nJEHtyAXYboiA9SD7JTMVeueCDXRwIs1gS/hVrLNkxPQ3iITs3gtlFvL9MUjPniCN
FF3gsoi9sqd5t84N7jKoCde/wBjbW9HbD3elcDfVw+LaH+cR3jCP7MUFrjtr9q4YHv5KwAyJdfL2
OlK0rEo/G0jkX/BruY+Mqqtg5l0UL+WleuabfFomJF/iBY/upL8iX6uenG8E21pM8jpjVvBZI2lB
jADooTuYUr2bDG65hDqs96G26wYGTB62VwBJhb57LwgY5XZpSPtLkpzRDBi4bZnpDcYPxxw0fhED
LhEVMtQwAv0H9/98YpgUrUrQubXU6zmbE10Q28vK6ZS9JqkqURE+TtnzWwX9WtwNV/Jof5NDSnDJ
Aq2mACvwHQjfM0/aSDEL3ZqM3rjGci5V/byJ/ZB+9Hbe1CYaSv8mZlRSouKOthW/VyP9u38JwQwb
a1pLPxkDOcGBjDgyvbDf8tpT1TVPSNn04m88QhHTbcm91uc1ywA9CPGdUFEL0G0W4lJQnys56ktd
PkrEO8L2j+QOyizo4wow1TRLgJ7WH6pmg3sq8xGe/vFxW+SIA/F/07v/hxeq0HsZ5ah00twEgFMn
Wge6KZafwQXY9p3q1NoSrbLVugFhq5+2t2jRbmhOufSDr7QUTpEgfUE+0V0zTOn8dKqEdyfewSsY
dXKessQR6uD10/TBwW7dBh9wMGnSOvbkISTO6fZiNkC+2WT2HPRfJz+1d/Ru0U3ysC2xVm28Yjg9
7y9YVse6dkllxqVlLCHQF0Xg9HhyPj8MTRdjrbbNUFyTF2i2Vk9d7u4zOV0HcToJVm687q1ULouF
yyA1hlI6jGLOKjMka/vqb8wZOuGE/ZnWNtJYIMOmH/1D5xK/eIDTNX6HWemgtklg+730JjYHFgVS
MyJSkqQpeTX2ufM+VJyVkcbR0gOO6CB4Sm0pYZnac8/B/TWOfXJFdqDS0jS4EStlnsErJW0rWhBR
VNtPatxgEcn62+gr6w3gso9BnB28885u5wSjuCskpAJ4c4i+ZZYs4K2C2a/LVoZ//s1kL4GhHYJ0
XMqtIGAObXEdLLb1dQsXIqrymiOtgkYYHemtX4dwrPfCwCHyd34bwtDy/1mHjR+yH8c10WaxtFys
e3HCeDtUUjUBP2YypFSNMCtT7LodVOvec/ebq40SvksE4t9ogubE1Kd+/EvdfkWv7VDA7jCzXUq0
dDDDTU4BV5pZ6Ar2YMbmcq009HAHX32639mjsbFT78Atg3nqPVTq6K7tIcOgam79bvi3zOLpNyuR
5I5cdV5XSi7MHgX3LCVHRcuQjh7jr9qSejRrpLZ7wHv0WRgtugEdw4sv0tzvIBhIcRO91S8M6Uy1
hLGUOfDLXUgrLmcpPI4/WY03V/xsKwWHR7I0JQFRBH+D86uRNlckBG9HGpSS9K4FqtoNlHi6K/ou
5kJ8KzfgrpBCanlidF2Zk2V1S0mmRZz5B1MLh0vXasRwQiAVKrILcBv+wR27Vq+YzxkbNZ2anUuN
1ay82ECcnfmj71X2XPn8bFt5gZmhgWbsdjdR1VjRn69uRl2EQ1Vzt14+oeIO7H5AwL0hzKe4AucT
HfA1rgmHf3W1N9DiRt1aMXeq8cNBcvx833r4eLeDMwbDEGXxsXfovk5/lLpbkCJrT7SieBpx7UzQ
gys5u+rOfpplKld2INQCDeb8lxz3zCSRLUxHnnNB1s/JlK9rMnYqs5VRLg0+S0KLpii0yGw1+UQE
Tsg6UYxCqRieLNAbGu5OVFs64l+S4TzZ9aMEXs0iO59NzWy15dugeBoJNyc5mthSmcvc1lhDLKzi
sTqdmBWN9v0AlxziOPRLWwTlu0enIVA9fPxhoFY+NPbMuyEG16eGJOvPmZzuXKAcD5u4uWX3Pe3H
uNqdQ0B/f56t9toIhvr6eUfd6qMG2OnldnZWqKdS9AxxLix/NmAUBWpl9xj9Bfpsc1hYeeghPCKP
3jT03ivmpwHFYVL+niL1w1n4yb4Ltql03RRWnerOeS5brukCD+0sbQbtqhFGJjX4tkSw5HRwhA4C
HBKcG4j8nIAtmRU/+z6kd9qnC37+Y2kCgLRQtQrgWtCpqmS8l+Hb0yK1nHGwoQgLOun6qVznBO65
3cc6/fQiG2M3rK3zwUbw0MDenvXNWal2U0XrutlvLSuQ6O6zc/b12oQGtzgsc5dHAUzX7DbFIY2v
fb4pwwxummdQAc4GsoPumOzQlSIHCqkHGqBM+Wpgq2CSVz+eQN2gj3FinFHsPa5gYTmdmE9z15Af
J5UKtCKxfaeIJdA8cYjKm2KpeKO4/I44kvvFbVTW2Zuh0xX8MC/Oh/IvWQcth5X+HiDkfYpnp4hi
xI7/RnWinzWQ/MhoRbttiy8aQErte+xLxMp/VLBt4dfQUlLcL3al059l7bK9Pr0JXB/hqlU1f1zF
je5Xx/KLquwNOUgW25WJBmI2nGViApoBJ8NnoBV+AYs+w27zTlMGdiU1wXUYswtopT9RkXynoX2a
eKgLenHKGT47eE94xToSV9vnGxsKRyTDeSV7p2BIbQEqNfYd86rZj1lGZ5XmqZ7xH/fXnIYbdqHa
L6MSOg0kDF5Oj8w4narWMoXLYQ1og2+OLlONde9zQiKR6Zy3DlPnd1rgsgTVi3IXrXsBJgGc0r6T
2yATqLjod4vcLaps0mVk2SkaQUV6Ge35wdWx9/CTj1CsOS6QcMObcC9L9My7RokXM/fyYwB5r7Xn
DBD/awNXSItvlNINoZl9P7ycICuuDq0TNlsxLva6fgicazKnBz8x2Z8dWzED4Qq5FDBiT+PqjUeZ
Uz23Kx5rkuUYj/vXHnZiVN9LEfJ2mlt/3yKHd/Y5Y4343tuz5wYf93OX4D7uaClxoqwXmLyBSBT0
v8g3fp8kFlhLI5eOdLB2x/2j0BESL1KDQEE+jFugzKXiniG4URsxfo+E23UvH8l+k0Wkp1r8KTYA
bBL84Gb/USiuva68wSlTZdRSroiIRwrGFvpxlVSTCjQnP5F/HGZgqUpRitkd3pvNO7BNuWvDVbBb
UOHkCVwWSACNzqm0GoY8Qxt/xXXxTpXB2J7NisNG8roItFdD8FuZVMybq7ot9z/ADB0cvWNGli3k
qrYFpU+TQcDI/Xsl94U0ZAdE9J4xlznHlQUgAN9ac8nePXjUy5u+LHOi9yMFZsp5o7GF0mjFyuVH
MtSHUjAKvjTTdDF6DMFDzbnyPffdkqOyjLPlXtj1oiJTi3GTqBJpHbFIM/BfulpkFNw1Gy7uYQHd
EITzJujFUVrwDcpcR10V5rsavYc4cMSIakvDfKPKrIqQUg8KOzw5PaoY+cFf2Sk/nbeYStVv6a1A
7CV+HCyoI8DPcbF6DL9Sy20Jeuk9z/gR5511nb54ym0+470ZDwoaLLTtU2xAHgTHnfMamt9geyOA
LPrYxYL5hbjUw2hx8TayhY7P7st7wgRyS/+CZx81omgYqmvAjt8v2P8Olkay6UkMSCBVxFhJzTcq
/UfUhvEgpiXWjNO9MDGrkhL/YUxZXaN0IMNGLrdMDheRBVbDjQ9zR3nDIHs7i5QOy6RI6p5D8bzL
TLtFs/scNxcDaKejtN8qU0jsijXrfNqlqxgQVMubZiwYF0AtAVFS7ykrtjG6pZFeZxI8z/y18rLj
9WWshhuEfUDiffwwfy1z9n3lDOCYraOTIgcpU6LVuWyOAagm4+pdViNz1XWy52SBwTElLR1V9o0l
GHgTXWBEiz4IyJNyssp6KCPLJizpb6ncZtiAaHOx5EZkK9dRhLOPdPTbkvUo/sSMp26xkzw9kmrU
gsWxgZtdVuwAomHXRUfM3jLG4BoGWCFyvAR/5RppuhRCWZLSrzuNoHcpYkOqdgScS1JNB7qPvBu/
LyYKUEojIwLVcYq+X7rJneqd+kyLUq4lSg987kE8ikLLDD79j/9Ur1bo+EmTBd0CMv6O0AoKDWAf
3GVddkvbtKGS7vp/8XxSbK98Gc3UuMsmXFk/xyJIJu9xUz5tHCsIzUjv56OeVEMdvrHwwywBMRZD
6bKz3wCLlMRVwdxzi+gyo9PbMF9x4+It/kjlonGqD/8m5ICR2Jv+vMQw7+FJoFxPhEnW2FAdOesQ
jYfQdAXMPNUaNFTb3uJrHNwGBz/IInFo6yHlyWm5pZqXH4iLhHgjAYspe37NhN5iB+oIwIYiowbc
NZ2NMDyDRSOEFPqoy2v5g65YNxtJuz6jm3j8CSM3Fbd0Kbr/EqGRESwJYIf9VI3RH++jxNPd7649
afHYp4m4cr6ExtKtjIcXLXkc/yAV85tUVkqWDzRMfLrHVwSWyhZ2G3c5D2xFMoVZXAgPOFKq6rDg
GURQ251wfylW4eTFTgVmuU2F0cRSoJChkCQxqwwYjSubZZtGWIFDLXpdQANd3XEUVqp+dSqocUQA
zmIghGFLwpwFFgUpsq/x0pxCzrZBa/2YAITESQ1CyDDOyCIFHhKzuA/sm2snHopbiOZLeH8Pjn1o
Yn1mXocGhldGZwrL4IAYhZdUExr1NoJK61uk7ubjxL3VrdK1L9M8p2WL/gqMvNnPr7VNwT1gTiVd
wtzV/8OCjFihzc9WF8YbD3nveJagbKpVIPJupdi/ydFkaHfjC/rVeW7K0MqWy6M4uYxpXsCxdOi4
uEC9tj6qtEZLmSsKn/RLCbeYkqB0HgUqy2Vf2CuRwtTNMbBa8uoa1ED1dCm5elSQml//9/xG0mjt
6Uxpnb7/E18oKCyOO+akuAfChwa4swD6zJvenHrmPbfGaYIr5ksZis7dQOTbrrFXz02L8rXkMBYp
LYNcumllSJbOPaRijkw8mW9rdk8VNo6qI7PDn3JV90Xj4lJjFZbDALQ392Wwkf575h9IGUFn1VI4
D41Szh9pMrSF00godYaILsBTF7Xsyuc8HOMZwM15NbAO678kNgccmaTyRzzXPpYiLGzVkA9hNa41
fBnLosTu7zM7qa77rNwuOV5+Oti6fA/n5ch4KS4f/Gh68OA3KTghyTr9ndrQvE06szJ8VQ6cr1zU
AWJwrfyNfLiCmwgnx98DHJUGPxCYKifu0CrNleFXhCSGYUXRcRV0Wca7VXO2n/NM+gmN72y58Lnk
frhaoh1XvD6VqGqx7U8m8blb6p4Ot7toCtC9thcB/Adnum9mSKjRDrwk/6yyEda5aAIDuB8Z7O5f
yicaOGJuQsFrJF3v4AitwANqZ1S5r/OUlmkkUWqG+IZKtdbh3HhzTqNM8N7jiVyqf8Rbd9ZWmdPt
SbLFt7vpOKyymqFLM6PHwip9OWAeYTa76vbnQmjg0C1Hvwq5/45lIIhqUEVIhN7NhVzfG+rD6trR
VeOgH1ENUgydd3+n5FUoVZue8yitnsQeYP9CPN65NptYl97TAPM+tB5CvXCeM9zNkeqdVO89m1g5
2mt3ayAQzVgkSAH4ZhvexaPYCszohUdir2JCFgJUl7briCOZ0jUFdaV9vkDDKHTHEhTfHCu1Zsla
jMflAfATnNeOc17VXACAeCrWrXhA2b82pJba9sCa8xVmw6FjWztLsgZNU4mwXw+Yk2Ug+AaSxW4y
7woUaXyP6btzbkW7MUPbTQWsPIAy2XtamN790tG/Q00H50TQDAVXh9Hj07BhFcqXrvq73x4K2T8q
vJ7qBiSaDcmfEExlp7wO5KeP0R+phziihZIYWriQXdM1wMKlhKGiHoSKUyb6VJyuUr4fGv4ToVjP
xEmmJFEAI0W2ocqMH3ZTHo1ePGtnh5Vvo5YQI0kIMsONveCLrPDXwfyn4eV6nxLH24CJON4NadEa
y1jjVECe/VAkPPdZyP4+ZcySSZThs7gcWGbGw8XxLHDbj3wKJemeUPtT1F1pqkokhAPsHkJspmcd
AJZycqI9BCEgT9E/x02wBV9ttXMQcl7ZXy7VUtXhNXyPHA4eyj2zosR3j1N90SaRWGf0hfNJyvBd
GXLccle/Slz+8iTRd5S41M/+uDlBUQE8kcjloAAA1J0TeqVsKZaZVIR/VpEPihU1PlUvPfhWwbP9
L6ameiCMSI8kXfucZomn8c1iwVeJqc980wQvxPAK3LwWjkPtQFmrftGNaCsYiiF2OiNbDErVm6Vk
jNHfjx0md8THQ8XVymJ22d5G7ZSIrwOsqlUsW37mSn0kty0hByu9fOw2CPoYF2SRrsEtfcSxjQqg
V+xSh0bYQNzoCRdhXD1lR75SYdSQsUzp5eskOlw9Za/JKKB5M9giAWWiBNNLH3M62Mx/sWddht8P
JcEilSNSe177+rAos21PuIg7ZLAKrNkMYB75ur8A1u3OFIjPT0DSQXV2gKfsqeUDVkCRjQMpNjvj
FEzPI3CGVqxHjtQuiauG2wB00g21mI/f+D/xZhLZA36CI5WGS709JMi0c43R1kcTAfTdYTs8fDQb
ImaIvB0UxWD4dbuzaznTz7OKU2zx+ijf0kjtz4+WBtyM03A9ZRJLrT0ZmcprmRsCFm4Dd/VOif67
VagTK9i+v/5ELlL1QJe/tDpbIWRx3QeKp++ENXrbC6VDNEaplUdCO5f3GJxYhed02MshriVeem5u
zSnn7Bp+zljEOo9mzu5u4M3Ec3aQti0QbhugpIVre5DMs4sDBt8tcOSvI7tMrQCwVUG+aXEjfwQ5
p23uK9ILcZ/z7RvHkSOJ18LpaRoBL5wIUY1M/c/bBwr0y/YDXqHIyOltjyZLwjt1VcSu57mbcxEg
GB6vW2e2JEjFSoRS4JHL0TQoRUos0hWgnYLfhrcpzIPtOqI15FJfzynxTmzOwieb51cKwELXAfHe
08jwDIOJQyOM+tdPY1T0lvsTcCWsdXMIe4SjRgnnMCe5amKVvTK3+w8oE6YA6stYbipWw5dnNTun
aZxyr/PPcD+66tmoNNRXRWNRaax+Wzx66QK7xIyF2WrmYcAsWVJVl9Ki8eNiUYbQxAgs3fCc1BFt
2mGw548fqjCHKEvyfDzLWzvSpRm/LCEN0LDXPPgmHhVSwigKg6YYz8zQtv/bzuLBoHFbm6eC/xp6
yjyE6xWlDQRSUTbdtiwL4K6z9zF4bXPSBZtwondNoulFojTO4dzuW/ziuAK23cUtzKJ8xVdQQoT2
9ehTuxdURCah4xULmswcDwvkhVcn04rZdWzBqVAHu4YmBt+Hgt4Fk4oI9x77WeI7vlxhGQwR/cP0
hT4Y7elBgXB7UEcKSqVGx/NGt9R8jwibSQIEWpx20606nTID572CsTZ/ui3o/+8+sxQrI7JWsExn
G/TdRXLQMmnFgJcsiUyLAnGgb8kYuNuVROhXVBhbzefca8G2H2FDNAoBDFCn6yqtN4mW1hzohUn4
nTxQoVejhFJBd2PcgT07J3Z6Q3BF0Fb88t4QWhNN1g2XDz64kkoTXmcZU/1ZwECfJ3amYqWambEg
ef8g8cgmsKImr+IIfLT7Y3+3K1dbISgAicnxEouCn2OtoSjLS816dUEJK4DbBTfBOeT+NAA21HTT
XMDEQiFwa+9kop9El921pceEPDIYtKnzN2W0lt2eEB8SY8rnoIIWhxZ3sniwclZW2DjfNenEdsTj
3RPu7vQOdRmVFeJgC2rNphuzPyp4dGT8y1CK7F58se4gxyxJoezgwHRShs4a240p5qiwIqUnugot
qP8j5g0nesQhhAoSIrKAa0gfqz8qcVM4ul97FfOhB/o7ksUQmOcZ8UoUbE4jnpeTePclnRYcv5lj
kX9pDJ6F72H7viD2BJNLIq9PGniDIJdI1dC9c0pbPfZL7A5+snY5CXqCirPO3XaEomcax1r2IGYY
2jS/omXFNsBPoqp2zXEiUNBXLqXWg3O3wcPxjsIEZZfx6yNw9nZOMwOio7bW3qwmqHnJB9c0RT1A
JT0UzBZpdPli+bdPpKr1q0YcRcgLUl72tjPchhpxHcbFcuNa9Nja+WLKaDqms/ZVsKd8A1hnS4mq
ZURr0DMVghz8AgHpaeXkTtz0H9UFcvIZu2Nw72C2wlj9031ecNuhFtVIjt3HRka5z9Bl9s0iqiOX
gbdRTi14uZIFO5khn52h6e2jjRRtRSdQW1CsjxrR009vFNOigyuJMBA9TTAgqKFHZnx09+Zef/wq
TFbJ7yHFdJ4hITJbWBvtmLR02ubpuDGtYlOvgfPMufi5XHY5LhEpsEXYqBVMa0f4ZvK2gSZVUwf2
enYordHYZ0oVZ6KjlUDXPEexNvleuSeMMFDRH23u92vmCYX2mbQnysnj2eTJIQ4oLiMVK7F/MQT9
ZiSUP0c75I9fIoa20Gg021IPb097cXP/XgfPNOfwrAR289dnrNCHGN6nFvJfwCQlwUoN3n4HAm7a
MFWnkoU9VryX9xDcuuA8dkW8ieNHRmUfUTBzl4QgqL/wMqkD1i3fVByZEOrjmsCKgcPovfoNSIRq
N7wN4QWx3VqOwBTwvHEy17ZkX6PKK1sMikPpuIcDZFSoVnTannKOM9QQ2fJqnvfeEsf2UhO3J1Ik
nYgs2vxyysy7tZDUf9BJ+sMdYvj3b+9ZkIiPLKq2OTaCVB76W3IQMOjSTunGe6Wc/avgLXaVtV9P
Cp3qCA67OOHQKYdJpml8LB6d5f8+Qs0sJwXdSwUonjckOJl8xtlhzsgO3BQdQtxeqj6cKqOveijV
jBYnzDtOMHGYVMr4cFPTJV4uyosbr/Pr6gw7ha6xyXj2UuGvfgD5m4kt6NtCfDnmUWBeSn3KmKcs
/xU4dpGia35cvxbUiuoERtgzJkdx1ZMrOH1FV4x4SlvReh3ZVGLA3RGQAjUIYE9hZtTOII1/w/ck
/J/tF5i3e4Fl2sGoFxncfr9WjvsupTGGgMZszJSSHjvRFk7CuKkdIIkriZ/TjEE8lcl7mxKZonVe
kpm1i/wRW8gf5ELuOoTa5Y4uiYpWLln2UIyhLwRHB6m2apCJZEwU8xqCtZ0+eyGVp8QM+wjh+3fi
HhEQryaITlssJ9yyVfoKsip6BTiGHoS2oK7xtJMLUQz31YRNck3F5nWYrkMnCFi7XMxIR5FvrrZ0
mxPsmPuy8KA4yLHsRmuigkwphx5LiNkuT0EpwCUOQAmsSkZBVmcHvjlEpSVC+U2CNC2Sp8H8+u2W
kg+As7j6Gdoe9RroJ9/jsZ0SXt6+UxPg12AsYswz/jlO4+7Hb0iou/3H2wixOy6T8z5D0EsqdDub
jDY+/vKFKAAZIWa/lJD9NN8BbL8kHL8gNlp3nmpH6mDRhAH9QDoj5sm8Gi+jBsJqdRyRSZ3IMz5A
VSZgtryUmfrMomKcdvGSu021kyxx1Bxq3lAnTrDvp1zXY9/+GdfIxZx6Li/NPG1AB3ivmewlfyd1
ZjXp60B5MKbZDvvOQI7z+PXigTi+puiryCkYR1E7LQ3b8YMdr94IdQG4ilVQH+kt/bpIi1OYsTyR
v4DS5Y98IGkmP8D1gpgXsndZUpZ2kpqSi+u3I81Ln3eABPSgjGBIcjLKzcEzNfpIUY8bDCncy8Mj
WdnVBnW59D/7wG0uiZM7Hj6vNVGdSyvKiaHnoEXwmY8XPRz1bXcfqLDTRf2sBG+Cyap41xy3+Aqx
xRR4nQuBomBQw3MRxARHwsndb4d7Lr8ofmzcv3SC2rOtITcyxIYJpMFrjIzMTmJHTl39XZeWC4dN
d/sCnfITgcZUyBep8CbvBsouTrf7u0+yrxT06TityNH7ffH6U82XTZwfwXivXe54cMDx1+QcyHDI
qOp2Ug64OxXAIMJr8QM3fNIDJnai92HqU4zA5+681oBdt0igz35tt37l89YiOEe0+ZUNj8B7TWBR
RImMI98iubajcg0N59pCsoygF2SmUaG2DzdQzkgUQRlPqqfIoa191DvVqwAOdD+NmYcLG9vdzsC0
vE4ad20clc5TF55aaU79dJUUSmL0HkQMMk0hJKGeyeAB/GZMLP1YSyPVnYW8sUzi8iDdqFKhmG5V
9z5UUjA8FMSYJKp51BdMO0MP+KQ2/zhg1oVEOWjDZMl7DM3N4IKW7J+kBBeyTVjrPeJt1Y6bjyca
NAop9AuNd9iq3Ku7XwXnOvFa+sHTwgrlzZWXjzwja3WOpnQqnwimuOR+GmrbAhnH20fR24ZLr0QS
GG21ZitNWH8J68RBQkQQrBuHx5pkyVDcuSVynKRwdikiH0VJxhvqZ3scxDrXUMtc289A/KMrHPHe
ZeQxbQvoGdgrFqbjpe38O6GJQsku4L7cQh6nMR4+1YOqi9sFboVI+T6+gtQFs2ZjmfeW2KAvscRy
KZM8b5Uf6fObJw8qosiTGQYOIWJzXRzzIRfVpFUXdkARlPlLOHtyKIPn1IUcM1qsamFCZLxc+DIt
8fXXikH6PZilXVxcx2fEL//dfHvYcjbgXp4fFgMdikJuEowjTVwjHkob1+jnEfC4mxEWpH/gU8iK
B4B+U7pKsdtxifnVTHHQo98MxEKSV2uxFNOjnGX2EgAzXeuJgc733rltJzz6flz9LxnP2BOZRbif
GLaSbRUrME1vYJjr9T+km54qNOcigEBLV6jB/EDDgGZmoJq5XELMu085fIgUVkkCM8WMVNm3PsYV
0esrhjKd4VqHHuvJ86tZGCu/Y3ct184q7pN8A1hji3c6abINR6ZN6vRjyOJPZHBz6DqAS7myJNrr
JonfrvAHdFFPcCXTAd57fOSKgl/6L9EAetLbugAyDiCnv53K22jmMXwcZBWWaKEgtBdyjC+TcTmN
d41nmbGFhq1MUIcI16p8iUUMon5RqW2wlLRyltedggRFOTNaiDG7lcwg+MVd0FAuoNleplG/9paA
TdA7SvrooRmXCbnNahA8YZOOeCtDfFgj2OsnMkt+dXSciMk0v4dGJa2kUMs9+UnzDcUF01ODpl2m
DdA5T2xTagFnEljpH/LIrVCbI3Vlecy498qNc5h2ihe43sF3cPOeJgykMQ57fgWJmcio50oa0MMH
TlEtAJlvoyXJx6GEx64iaxVJ80m05aHZgXsCKrF0B5zi6ZVVTjmeW8cwl9TFKtXitI+HRQwca7Q6
4NIHUGtTdjHpUVXD8XUpOixz8/zjIRloFlYfKfeHXQ+5ofehdIZbKQPxBjc+AfdlFS7HRHgTRO8f
UENntYTGGCG2lnskPRiqhWCz53VDOelb9GeT+TuecGkGnMBelswV+few+hINlU88wGuQ7aPs2EtC
xz26rvsIddKvGFdSKb8bMxY7kb9Y5VURtm7OHo/bOIbk22lCLw4Az+Ww/VJJNl3AolKvvm8r4CMA
wKs0uUdRX3pLBJI0gkoMJAWgh+2WT2wdZQYFWHYcdXtqenaKUwrV232285habNmhp8HfTM54bCiC
6KuXo9dCTMgrrepsNPzO7WmCW0LpIthEYGXKa/nYRx1lcKxamTvzkLeaFOXbTV6EarPy0fXHqNg3
jRXTb5NdhxuQeGbcj2/SJDap80PN+1b8xfsJD020Rn0UaN0CFq4XwubEMNJIbRQsm+JjF1enr/TC
bhcvDxGrAhfCeMBVT1T0qdYdQu/sceeGWKdqmr+ehVsIh1QCGou0/dF9/1hBJrL5awUNJbdm2GqI
1YX0O2loyLPqtr58MEZ95WvdttBwX5LhCuxqaqWJ4fkm5OFcsy+UPvJh05aa2pMZ3PLGbkymHRb1
S2BM1bZSf5BomaeLyzkKefrEWEKOvq557Nn0Rj+KFDJxCazvN+lZ4ZU4/QP2vlD/uxdGlXxMzXOZ
v4gYTQPcIju92geBwT1uo53OozcTnBluNmzFqFqvH5O/AUs9co/8DBfiO9aYeA5UbMmm4tbbz7Er
anM22YEfKwbHRX7a9hzVfNnkmqSwOBUcaQy8OOWQOlRsAYws2wgpu3YWfwEmIoPSs5otM2N99eQa
STf5aB4gplNXTeQCg56/J9CVd5j1kiEEuba7oJzcWf4RrrkYSJMTZ7POxybV36ABzghAiP7Yt9C8
7V44RbvH6F+IzJMnxvj6l4EwHv9Y5GKdk2KRqaXLLL7xPx5fXfmChPbL6m4kpDCp5qxI9ySELmPW
9WCUt6FWwlzgGe61JGBsSkhF9Q8A6R4gTJJxUCOzVpqsB8HZ1K2E4ER4iwFpmqW+2Hamhn3/pzXr
lYOx9YRBUqY9B5B9osdBTvZ/H5fz0jlpq2RoMRsb+wjSIuN584VhXMuVJlh7nMmWSCF/MrJDXRPr
XfcXofHQNZSfGmqr/w3Va7EGWIm24hxzh/zydCd0+WAOsZpfN42CuYWsLZ8OPRoWWZ0r4RQEniy3
JVgK2LeL2+AhNYn2q7aEXZNlRt6IYgwvDXuqZLOQijbstFxpTNOKic+xBOKOLeaFMA9XF751CWub
rQd1dhzRK6nHRZ3KcK9dxw7PrcufV87DYkoyywd9DRKcLQ/UBns1CW0qT5rr73ilmqw8Twuemq+3
TZSUw2xeT4nZlVnKM65/ngBOzzseNZI9bWu2DLD8zgJ/jxgHvl7rANPARxAhmD0bmYPcDbwe7CVt
Pp9YZft+qcrydEzRX263/Rc4i5z5D9FpbijuKjOJY2Y+ybt9he1upP0FDbsIK9eE+ib/azXF/KVc
355RbGb0m+KgzYHlg4W6Vrb7V8ZfBf8+1+qslQrBe3o8h1ml5V/ssy8+FRrbrmZwldcJz05IN7Cd
+28PshAkfdWViJSeiSa/7oRACCjB7KGJLE45Bz7CPi1nFwPviSWE/yAhs85p9y8C26urnUI99zVo
wELoJ5faU+5I/Xc0fk+gWnmVdIvcwljaF/4pFWLy/TeZAnsiADKNx6Z/5bebn5TkvyWOZxwGyl+i
ziP2gBBH3MEN8dNUSWUD+z4VMx6IhcvVzsRStud79zi5cxhXT/iJ2L7S0N0ythqgbRavZoNhRJgO
wCJXocH8GtqQzkxBYiki9HWRwAEvBTL8lS2cdu3Fpqv2ibWfXrZkMv66REZMrzq2Xom2qhM18Avn
XoKJTJNJJ+W7DcM1wR5VEtBzh3thg3AdVrdIyULrETq1be49n1Gb5I9j9nxWE3NJ1mHyadnK2DQb
HP3q6pQIzobxJUSoLojjMeU/Qg0nBVJO/Tzhb8qOkNaN9bH+/Ov8YvVMXA1JFSCbV0TglQDm2gMv
AyVuVdlBijEiDM1g0e24mCQ01gJ+b760y25vOF/0lzobAFMzXLxy3YBfJU6UEdHs/brC5033QDmO
9L+Lxnn14etaHnXK7a0SBvEYnVNW21DfCJwxvKb51eH2mjCDR6OCTHku5iIz7XhWeeEbzjzpjzY4
YYRLZQfZ6jEvKaDlKB7vMIaQr7MHTACTKVeghNgXDAScudGRrIqOi7f29+ClzdxujDioa9iTou4F
6Hr5dDdMAsmFQBtVpuJY/FFMOM47pTiUCIlOe+X07GNJs0PS5aBPPe4KMNqmcYemKkMzlJpvmsCA
/Q6X4Z57i35PgT9GKraH5/9B5L9zXTi9yoZSdTJGQBtxBwKIk6ynlhdri0ROVqLFfwU3jS5vrbfU
k6x5uM1he2jVtCpBvZuBcULvuM5ICFYbdE/x0JJu1T9vLZsmwoMQr7iqKgymGrlOpFsSHIfjHo5a
eUvmQRD17YUsHrMefxejlcQICoUsaD2d188luzdux3+sw8PNbGd7sa1QJgW0XL/7rR9KKyEm1AtG
iquw7zIuX//Ede6dFEUs4JsD9wSXazLtqBw12giApY+6YuIsTVrh/+Bcrg3PcF/CIKKVJSTdWr52
em3hDpLxJzbi/OoNeUnPJyMpKAgvVNhpYPSZhIzchdwWQiAc3nsM0NhA/nsJ5+rD6Jcs6d6w/RNo
QJIHkY4orAAfETCfy6I4Y0JxRfaOhpGFhL2maUPuzD4gxDZGYUma8J8oZE6X6ge/Lgns2uKCv1EM
gokx0jEJO/BeaHwLs0IFJj9PFyQP8hJk5q1kYyBSvCjc5kyDnLOHMAjYw5vkxp8ai1DywUhQ4f7I
okWO/kebMnFuynOSrOst3HPmxwZsyG9h8yjrStWP0XVgWXNiawx2JmpJNtELUmSr85Da4Tq+gDC5
Ij44Ya7eAB6JNuasYOcy5ZlDySwKiIPZa5UuRfmicVrPkAGrdfggqECh7gnZfuQr/1YeVBWx9OgD
wjQZgzDg5uE08dX9PpHUEX6mzkezCIMKXLofzdE/+5yXMJXejHQSVOdzDW2I4xzKNBe+jO913h4f
s/TjCZ12wy5BjSq5foQkb4mYSRHClBu3LRFPaQKKSlmih9tlsC+wJBoEwjIvF9zTjr3myLtK8IOO
DCgreHNaBUY/J8lZUlBaRmoor0QdjzvQj6XFf9cjpEhoJ1LXUVDrErH4xwZmnEQD5hF6pew0xDSr
Bw+rc9egzM9qTWAo4z83Rti6Yd18dKDfOkD9WmPbctVvz50lvsdMtF9s/MGhsg4NGVaTy+Qac14n
kwRWxbOYlaAJSR63VpKBn0GccP4h4j7OEpuA0rCwkrlmE+c5Ve1a/INsVV3jLKhqgLIOGNyQJhQH
c9lDxUBE1ZoorqTIJe3YaWr+avI1Wi9Ot0VT+RDKDfcuAIRJZJgRVkhmgHJL384clcPMuxs+YfCf
/KItNT2uy8DYU9ap93G3jPqRbbuypq0ydwEh0xOJC8tAIVsnTmu3EDOklm2YE231b56JWB3a9lZD
cfLnf0Ta765y/EW6IpIoIqJ5NYxG6o5H/WVfeGcwPPf4Vmuoa7MliYi7udijRt7rmz4c6L7xpHjA
8nuiUcP3pTK1MtkhtbEfuhVbaTf9RWQHPAhjbuelGzLgy40F8sZ3SkwbShDuJkjEhuRHOMcmwYfD
ervyTQ+4WtxbkpQg+dBzmavrpuOu53QDVglTLaaezg/vZin4G9E0cCkFdTueucmOi+Tyn/D8EPNi
XvDfk4dLT9rs07KVXWDTZqmsvOR3hZFmx6QPWLjJYluhom7ErUSbmMCiIURqMffN0X4KUDIFpnbe
dXKQdY9NOe2R4J6upVZeUWa3cRyPhloa5RV3iP5Zhp/b54ODdvvJ+TxjcVM0bz2ah+wGw8fUkmm2
/aLtvLQXXi0mksff/ayid77NDLEkJu70S6fq1JVml8tVZnfW+WUxhYlFEWnuKeUVFojQvaxm8ylp
V7YV5noYpxYR2P8K1acGxEiRmQW7EPuo5XBex2bW+oFYJP3pRzFbOW9k2z8/0pM52jBoD0OLIo9C
oTe50AV2iNQadmcR8fsle/qs4l78k+6VQZPcBz8EImFA4Akh3oEf9nkgvA5nX6EaDzHyU4kX0uyk
gDPgU+DcXYjDWKvH4h2U4NL5UqtzfOyC61dZIuOIHDzPmuq1huSjieiIzYkezgEIIow7dx1WAsmU
4/lUB/0K89P/VWqP+utX23QMNJfVHbznzejgzRdZduOfi8ctx+47ggQBGI//JV+t2W8zEpYbx9MP
Cphq2nD2qsXFMJKHrAemV7oOFygedMJZ3NAjxJxLdW9kj1inS3JVeFhaq6Sn0dTrmKCeb1MbuKiu
scxxizcsbllkU0FuUJfLOMNHDbzvHw5wrZsr+hb3raxKPwc0+mLkcEK4FklOeyS48Xer1KUtGegG
YND2mEzOAJ3fE1Lz9uRfMdnTL5TFKbHRkMaE56JbDrVmX3rZB0pr3eUg51aEVyG0MhdklblN8I8a
TNM205H+FKiF5cAe7WBtfmOBFJrm1hrNdmByE31hmA1n/er4O9gW28luZoOWwPgZSI9jTT5whar7
ctaeS8f5hZr3yJmP2uUEkFcOGMPQhXyInHHzMtjRWBpXqhBZvus61OlDq9TTYBEhb1McRXykUcdg
p4kzKsgX+CA8gNtzM2a2YWCSre39nPjK5pFKTClWgraywh6ovtAb3TC+c2man/+9mwBRW8RahUpF
32vOYKTJgOI1Qd1e0vKfCSMQmd30euBfunikri1NC+cBSXQxb1lSfKE8eTQSGtrOcJb96+4JLrP6
ke02zGU2BPzBRaUDdtaDdFANKbJo4dkbTPvcdVYEkJagjul28CT/x4/53BwCw6hCNxCdIGkCBiIE
P9Cti9RE12a4pmB75zQP4nyj6h8t0aLudhLMYqsxGIkEqUqgqzQvDzCqdXHg70HZp+a6WaZt58WQ
hyMx/r854e2KuPcAFYb+si9R1IVYsZIuU6smy1GrV2/mjSsXD1qjmPzUC6LobaLEvKGTvw/PEy4z
A8cj6rGpaV8ALCoWUNvKWutpncrx0eYeFsmbwpPqakf1tnroW9KKdvM7wwIKmmKySFSc1VKDXwiX
po4ACA9GTcQu9l12Z7xkpk908KvJoUUxb1+Yt45T3d+MeHV1nyVrAvMltiQ614I3LXO1iO42CjR1
kOxasJS+P+Tc+Y0XOJ8zVgaqjFWlyhMax1YvFxw2hz2ScB9mTO0UTWOTyWRWKz+HQ1VGabBh0qiR
ETTACaj7zoNu06gh6qEwPgfLG4qbA/XLXI7zh7YD5p3CltgVmCEkxNharOOCK1jKfw64+9cKFASu
Z2syX3AkTNEuaVBpvyvC6B8OyOCbDNkENRwFPomhEu3jQNyku20RAREDrGWctPwZS3W8u5ssU2mH
l1//U8OplQtfqZMpPxphPWIJ0wPfoOhVgPlBfdqOyXxI7QjhWi/yyIlAS0qMQmxEClGaEGMGXJWa
H3Jxh1fu/ssJ1n9DGh/Z8Q3XEUf7pL27tT6ZAjKe68H6ykU8Jgdrc16webptu0zBpLMU7tRPelSP
rXdW0G8/qfZb/vLUdixQncq8wjI8CGmIiSBgfkBJFta8dIBa2hY6yqFKNgbLFR58hbGy9JHTnJeT
i0lvfnLMHJJ/w/BQprY74lr1diSE+x916Fp7hBkHYPRwsmk5Ulq0nFoC2jznwxPeFFbX08nXd2Fg
W9Xd7YHQFnOk5sKYm7yXFv6ObaCXcHiXklAFCDK1q6vftXdhX4DhZ7SnFNn3LSavcTwFBfGfl5cm
48hS2ooeuuBHbJ5utkQkU0nmlQV8I1X/SXQdnwYiKQ1tmM0icPNKNGsWDSeKDgwBxcvOEBXSpgc7
nks76gAxogd4p0PeTBGNICNCfbKz6uS1SJE1cDEUJlZI/zOT9w6+b3IdnyhDKLVZENRY+KeO4wms
fTe2+8Ffv9KmPMkrk7uVo2SHHXSAXV21XZ21i7OMKU0gXt4isPpdrEHpeTO2C5LVKW2bAo0fUUSP
+NLw8Dg/d+aNqKoGLuPvXLy2cIKR1CF5eHwuwV8FLl/YsDsPBT8fNqA9AZwo+887dxc/5WQGygn4
U/c3F5nWbkjQWA4Qx3P6tPPtdPruNk9uQ6VH9G4B1bXvH0juLzuqKlGQIVd1G85UVeGbsEuWp6Qf
/UAVufWqWQLZjyHBKGqJHMxRjETqo2BRWcOzr8CNnRZ16dQQ+SjpZBvFkAtZHXiMoKMj0xFudmn/
qTpGHyTRfTyXkQfsfGFW3CsxsXx5CPKEAJvMH4ckUr0LC2WFNq/Hd5f/AGEbx+mdri8wv357jaGK
qvdGgXEuNEWn7Z1eJHCuwksITzznCPvAFd9mxMzcebUZRiVI82OVsxqLzkijLPfzdTLUjJczS+i3
zu3SgoElm9y9395FsF8waZIGeuC/lJH7FzEPPE9YA/1G36teCE4Z4bB/VVrXP0f0YnOSpOoyocSR
n6qRdsM5btGkvMIr2z394Tw2mKkxU/7GlQNKwk/UjmboLFyj5lmQzwYcR3n/S8dDMytSw2sR/bt1
vg6Ca4DHxaVqlfqrtu4hZV3HoIJb9u1kMmS2O60rDkcfF/ZczbwZl1sFIwzoYKCq7/9VmnQi7he6
+bFU8X2MH5Ncvpri9cmeiFsN+UqjK0F7F5pd0vc/TVloIUOrag2IOT0KGMmAMFFdtytcw0Dw1wKn
I19Lccei6G8xdFLwQ9TFTvJ+0y2OcgaHrgEVoJ1InS4amrFvVZof+Azovvd550jNuxxrxTBYV5Tc
ZU/fcmD6Yqy35Ul+4WYQ1UUIDNNkb/FKFJWMDkyjsmp5WYO2p1N69fCTM8RhrlHs5JHfTpNwebfW
aPapUzmXfBKO3fOWObgdDsCPYqiUA4MNMfmQGTOeriFoU2JzGRqN2QKm29zofrxgbpQdEVD2e1d/
kYR27i2gSslezrffltTmqBI8Gwcumoj226UMduZJ79GKl3pg+CYr5a/6+Sg8qDX+0NnCxCgyz6dq
atvlup/HyksAyZR88GpWSkOtdBeIlLCwAoLSCyqfePsHMrO25s88/UTBK1XWhAoOgf/MRN+CBxYv
gz7Y8wUN8CMKegWBNXTYIlgVRpWnkljEe54S56CGZpH4tmdDjDkxK/5mSNTK1X5HinnF1kV0XzsT
q3P/uAFgiUNCLaxp10fJFhstlQDX8UYn9o73QgePJMfaNpL0G7t9vJ3lkhOgc6Tbe1kpJOFlrMPV
k2zuO4X6zhdCofH6OeMTcGj7w0kf97zi94tSQunkeRq1t8d2ztF84rgWUQvYHdqeIVTuygwho/Km
PIA8WGBmgI+56b3/pkkST+YgjQhX2q4oNoO90F6mg7sTHdj+fb+UXphjA+IT3033+d1WF/thhTXp
0ulQmg78LTpnafode1TgIS/+fzKr0Q9K+ZNbkI0LN8n+N+3D+1UK7HLixNs75qAg1x/o5Us/9m1/
YoMsofuwO38MMdV+KN4fB1IQKr6a4Ww42AjGL+tmEq4nRL2BGGNd16Qb9KXScrTtPSETR/Ohyzwo
Ol6y8vkwj+xrCFf/4zzzW7umxzB/FkKA6moH/KvtnAq+pW7vDQHfHYhMdOLbv5t4dIoZwLmK4e/G
Bg4D3nyw0Fgb3DKpJQrp7ArX4dPVYi1H6inehsk3HlZXRVbo0IMw+CAXcQWI9AeudXILRzI+/wR7
DniL5rUzaJtdoJBooamU4CmsiROF8MegDylgfw3GR0/On0z5/2RFhFH3eg4QA53Z3c+SYTmh25zh
lK3A7yr1V5Pejkq+E0bApmvBgFTDHbPrnMQNivExAe1tAoWvBM13ht4vU9q4A/D1QCAms/YEMQ8T
ZzNbXZEsqBbKQG1OxoBqXJ1QOeJ3/rdICASci6/0FJm7lqJ4jD/03Nk7HRvmV53fK1jBKhYoNjHi
TsiXFbJo2V2S58VNhO06y7N7W0S1rR8oe2/sLMfxnwrwuAfdpYRoF0TjdW7RuhaqVWJI+lB72PjW
F+YzMV83D1+4snjVHfHCTdrCUcT0pbp0zT/1W4xl9CakOy3lcsj23WwwjZOKx91lFV3KekWUonqg
5edRQP9wMINApxh+AMi/eEjZvPQowpGLGO02z9Ftixai+1VGxshROlVE3N+RieCPYzyOgvfSWHhy
+Gfkggaj/2vT9wL7hj09KPRZXJ157WLISToz76lktauwRCQmwzZv5XikA2cFHegny3OSOh8FiLB8
ZcAnnubiyM9k3Wax4yldDz8xIuG9GYXxXXQlKVnNhD1jUBu/Cfbl/3MfXAlnZ/9ZAjVKYJhC3wwc
Iqr9S7LQMqT6MpUnOCltcTzC51ksggAePkTSmj9pXQlRV7UBM7OtgRoQ6fb3Ieh0Hn9W7yKdK8aq
Vyjyu7V6AFUW3O2On/VoYgHjNv6L4cSCGsLsFQ09b6GDKwZP5nk7Opw7Ih+4RcgF3z9+FryX0592
7ZpeN0x8d2UOVMmSDV/ZCFsrsvDwabc7jfFnJKGTniM5izXYoQAFWSx2qn3uH1ytE+WHZqMJv3Wh
KSpfM6QyQNYGkMd/2g+OMzaQc0OYfj6dcRrVFdZrFV2ikn6T5nj4v9HRQFaRmM1xCW+rERL1Abjd
8Y3hY1xBHKw6DYyy+SqCg082v8aiyg0cQGdATswde969fNbJvA7ZmManuWwTrh92RupkxOUFPHCs
Sq6SBMrVsdg1PnMfFe8XkZN0S7i5oixlatAHYYM+IzqJNdT8bhW7qvXELHkbOV8IzbbzNs9p7WZ4
t+kO1j8rK+mpdp8hrSJ5hK1hwEBilb3qyyHbXiUSgB99klK1f9wHGzXsT812ue+wDzl1gpYNmR5J
4tJsIyNvyycD5lWFWBbAN9u2SlsG1/K1MAVhkEwEPrl/q3wSTE3crbnEJ2AV45fGj+Bw27H8+oLO
9N06nQAOsTv3H8zTr+fCf+yKA4IK0VeBe1tnnFI5kje1+X+0kd7Z/VEjaIUrhmjhPTgaFfjP6bQl
/zW2WbnwSV2eqB5sNyfKv7iIMGn6I5bUAC8dZLluBjy4CCG24ml8E/VejBBP3unh5mobZVSz0a37
+QFtBw7WzapPo3yZAt++dVY66BCYXbQaFdKe50yifKntfdauabVuyJQpFhsX5wJT4yELZNPScKhm
D8ftbtnsWBIX/Li+A72cHgHyi08X4wI+Hbv10HbJezf1hSR4XA2CErrSzz6uHVI71sKrbzPqOcR0
7Mp1HhkzqvYu6d7XGfbk9tnuzni5synx74pQWx1XycQtdbjxjdkR0AIfeHo5cepCsq1IBSkNJQt/
+DKD3BdMD5J2LuNoXNtRUqZSw/FIb2eX/ZKniV/w2MUaBQ7+0oV9XNd7RWxg83rXepH1Nk1HiR7l
kUG6t3EtxI1tgRtYrEjYGIk2nm6Isnbgj0CJvboU/BKqOGvxzky+/ka21sPrRQfA73iXAYvrV/yc
1jUyxrURG6sG57i0hIw4SIeYpG/PBlYz89JcEOScbXiVrIyZTPe/y7PfFDaMvaZH40AF/4efRwio
Y+QaSsSlnMBu194+d0IH0KvjU/vdNZogTaed2gTxx6hktwOcvEmW/RZv600oK+EFB8xzpPXj6rf8
Sv5Yq1ujFfjVuYJzTc3tQHx8snZ2r8+WayCur181yWTpmRnQhAvfyvVTVZ6q4VgOhO5yaZgqV1K/
72DiJf8zn5+m+/uBxLR1vYkKIQBpcUSPQKPmY0igrn8PSjo6+XJQgYm4JVaD8cGIoy3J6zDPA3xm
2xnBGUxOz8ilWXzG+17LjOKPwyeEbKWuBmII7T/juVnS8Cv8+LYlfk8f6zZ5/Mb3dZqJrwvNr7KD
572Y8zpp15sPSn7XTFFYzkqtA0LBYjvbokYz5ZKZQvBSFfFAGhyHjvxX+CWsNv5Nekkozzd9HO/i
TQmtD7bwyT6ccEY/jle3W6QbYSch59FTjCFqsUBJD3alNrjvmqUS5BfIBUkIOkeNIllZgdFtNp2p
2N7sYi8wRl2lFr7q/0XobMNLJcUjdBph/o6NSdi/azNJLaiKUhKOOMZd+pyliga7CpNA9MCUkzor
6g30Tt0mMwQ9Cy9NVUZJCNCV0nm58J/GfGzKdoTKklRNSrmCxtEL4k+e7cjREiizOGqsgvaoOk4v
5lKMT9cdZXFPZRSKGBEEbbLZLbBLghdnjlXql1MiLoZEsNNJRLIWWi8R04NhnGkD6foNS68VS1To
TQLcne3oFC7qQ2tMUvItn53WM5I23pCGFYVLrU1WVszi39ojINBooXX6BiXr/yTzN1ZHNDynzzsD
0GLoDZPG/U5Ax81G0IWr8d+hjI4+FrWdVp53xCXNEsVEx97EoCt1zOS2H/Or/gubmeHAFf9gdtNZ
nsUVqD0LPiwUkwHfbi0XPSC5bo7tx5pH7j92lmNDn68xNqhsXUX7iWP86X+aBQW7jj2kp694Mdqa
mdrRhCDQRkk+s/DBOXIJjAaWkI5xanCRI1I/x0ACA4FX4p0vUj0Df2TeRM8nM4j9SQk0KA8KQkX3
nzpQdBtOAr4BZqzhYkIddSjaJEYRX1FYjJg+mZk0+iQ1/FMHN+qioXjLnmU1g1oSQIO3VupCd56u
4m/Gk+4bLhv4dpT5OqxpWFohQBC3GBGGSzSWwJRPIrRg7Nbknt78vwP1UX9WSkNUsPr9Ys97T2CM
OQckh/KtcP4nYOPaF0v5qqRXCTyidm51cb7gTilVS1LJk1WJAbsOrKFF47XeASBlyM+m21J+JSMF
CddxNU7u0i5FDHUiEQq+D4Yz2Ag34VA7LDRisNd2Ma/4oSP7kz3o9bjXhbU9qmRyGRdjWsO0i42A
nSUWCKEw6Vwk9ULvQVL6fFGtRaRgqS34xNVWweyFXCYkdSf/Kc08hXdKKORJ2OXbBWsj47HijhzX
J+VnvBv2zvsJqyUM3F4bfES23kjDJOidpRHR2xwpqEqnv2n45AUMMNSQt+0Ttur+TCtnVEfjVaAh
kLdJLLbWQNJUtJyW3GDAmMhy4ozo0Yw//0zoz3LQvsnP1vSopyz28Gnf4npK/9z/Wv15JSUSaLSc
ORABQLXqGAehmCgSACDe98O1bE2sgdu0ckOX5G3qQ90tUpIPNttkHB0V1cGZ9Xjw4OhbwoWKyDQP
sPitpcKy+C+VEk7FwewcH24msbpowM2pWNeOo9cJ9nnsEVeMy1BT3n98vzfUAuzmx57Le2un9l+7
LDovEcDH+aOmBhZkpMXSEo/pmCPCMw9y4wQdIfYUDTf6l6UFwmAvfIukdBfJE8JLDV4/Ou8Y3vz3
rXVrvGYSjS6KoCNGZ1IM89YicJYczr8twWTZ2QfFp/2FPvbqRuVltWs5/4rhgum/P184Uw3pnFZ+
yBQsQeJCRfYJJj/91OLickszFWblRAeCBKBo8wBLzbR4SFslKLD6nO9Ckdh3v0MqWnm681/+gCLF
SY8kwHqbKK4ZuZeuJzLt+qGlCg6XM4KftOsMJ6HUvc94hhozGwNJIF3CbUG1vVedc9iAaainJZuM
09AbsaAvuie06o1/0piziX0RAel8lObES4pZhdIjRierL1sBEnCGmTUxlss2SRV0xMK7icA8xNYT
W/7ikFjvymXtyLbIJdEwsY6ixX31AP7A6ndXE87GCjhRT7RqoIVmCmDZvRzqJjrY01vDSJeZfUHA
+8k6sa6F21rBbTVcx5v8jVsSoHeCaiZTiL10WKJi2M3ypxRQvifKyvT6jzPh06h6IqgZlNSpBKD/
FE/e35N1DtpaP8phldBNvu7iuQiUG+A5VLk7FWpcLWaViZUlMPpFIEVwe/4M2XzJ5hDCNmjwVDpB
0iSyYlIV34eE9E1lx8/TjF/8K6GfvsKkvJv98UwGETZ8WmZwDqpzuS48F1uSW1RjuW+2B6Z0Jy9X
RApowJ6sOHkfwUGRPc51OqzdL31IGDo5t2gHgroCxYYVAZtcihHBwwJAO9VA7lnwjh4a0q7ba1cL
rOEkid+jlIZPlqmCUt6ORaIDO2Zq7oLHcSfOO8cTq8yEFUIAqZ2asxnL350GS2BVmPEE+9GD+c/W
pAXqTs8bZctk3g1Yfqo/KkDnGACjeOcHdyk3a7nGAprm0ItjynqRBJiXxE0DZvB9vUUN09YdH13K
u8f9ghX4xGwcgcIY8LQBjXVIR/fej33w32ja2nBaRBmtO6ZbUNFkkbOMPMNNUGS/zghiq2urouFj
PSn955EoaYsa6HkFlFlBYutu95QSv3A8NlC6T+5QYgAZ/ay/daMEylzQa5wGs9wUtiKjBw5XyJKn
i22FuVynMm9Y4T+wE+ZTWMY/nnbZQ/3hxr7rfxnbAi8JeScpUErbCmBvA6qQ85RkeqzylfNvT4m6
1jQOZu3CjTfjNtX8qWLGnXtSHc/mF0MbSRMMlrRPVRPIySiJkWGDXCJ1KS94t0j0wZEGtchWV9iM
GiHSyEyz3VR0Y6nKzp5/lDRv3SJawwAm2asUZe6fwXsvSEGLxvv9aOP/1S16O4OwEsWa8K/LK2m2
bigtDqyNVrWXT+cCZG6jqMl65wzW1jB9AyKxoTD5gTfkzvr2BF/XgJn/R5Qmc8FyEftZ6SfW6pXY
nJQTmW71AAB31UX4Lmqw1Ng+J1Y+qoATsA9VWW0FJSurZLof2ul1r6N0Ka/hkvJiDpF7t06pWiGL
46jEC8+PJa96YtkDQi4+tUeD9kqa6xCIvCg7pR4RUZVWqtnvNOvpK/ucQjRU6cn486l0YjHqmjwl
lL7uLQdh2Nqwq+f2YMBhsNuL2bWYpL0oFENKGRil/xAxaPD+g+bl5HUPpJmf1RRs2merkfOVDwmJ
reiHzp041UF/JDq4SFYhI3q1smuHZJJ5ONPay+yMYRbTmme+8ZpHB0FPYjg4Bnamql2PKQYyw0v7
Nhnf0asMs/cSCz1Sb2ETMGNoUXMyr9czXN8Py9/wyAZqDEBooiSvs/xSmJL1mjc4bOirAoDLvD3J
VcHyRrteE3LupdS/DZGAtlAa5d0b6jkjsSN4kN2jrA3OEqFrK5EVZSX79x6tAFAZgXgMAyqYvFcD
yIoJu8lz9tQf3fox7/E3ZsaJLavDFH5M+X7az5mHQ4EhpAcX7gy2zipJMskjBxc7JGPn9xYfN2zy
boaE2o4y7W4N1KL4QWhOunX08vPuGWIMJ3ajavxAYkVt1pgGTbW3OAcnMNl9V2S9UZrN+OhXCbsn
TZ092KRXkvppSKCNMSqMRCIUaEroUPjyTG6527CIPQPSb7n203PK4SrCnhi+n+TwTyE2yKWyb6wg
mF+ao7zcs3P2depxFHVyF8vnlUDbX5WLUT3QV/qr8kHTZ1/kkOqjzo/FkBZ4+veSJLQ6iiLekS2P
lBZFPGLWJUtXdgHT0yb1PoqL8lt825aLYLtBbcr2B3M/t7JClVReJWp4Wujwpq6vrzF7H8t5qKlL
p0wh/u0WhbBa4WCm3ymUuMMEVNrp/8tE42QdJcrkSR/chaEAugUEGk335CH4HEvjYFHuiudxhOep
DIXyUfUtybCC2rcYMhc1Z9fEBdiEXwFxTuKEyCuz/ElGuc1AVQE94dh11O57nCsP1xMdGDNgIcje
51aAs3NARjEWS7gZtNAW1lUZJ07pB4ccQ5h62KKBfo/YxPoVNi3oJyS00QewO0PPk6iA+R7PB6DD
AlIJb5R0SpsPQfS2CgPAzQNu8iv1acp12UBuqRLGj1o6zrqUbIS6GehZfIOZQi6qexAABXoBiMdS
2DlEKP14NrVRJiIXCyOzlI220emKzZzJzi3D7OIAykxP0FfpG7JNni72T5vN4WAQ0v/uyeOVPWED
e0snmOc84AS5rU7O93JfRRyQhNvWr44wxdaeB0N6gnNuUcYpKkC5SEofR3a9dZ4vstUjiFMVlAms
u6SpWAtozt9iFzhA8hlyRjxtGCNltAM4e3XeUIWeJYHDwEQransGkqtoSAE1FB7TsrXTkeLtE2PQ
Bgs5jKrFynrceKluK98Gnr2/ZRAtFtYLm/gFduj1OFaTG53Dmccqfsyxq6DpvtY/KucmCbkNbxvg
dJwCYO2vQkxeFisJJ9N59AIX74f+iuSJT8hX/6cHczCW7Ct26/kpfp/7SsYhMxJGGHm/mtrF5j3u
w8B1QOiNaVijqAGFfhKiW67pfmrGKaoWG6nqEuRh2Rrpeb9e0YCNC1y9GPXsc3zUGJr7Q33sZXoK
weqgLA5BF/bci1Vxb744brOlBFMJuDwgBf37fkpO7GiQAtuVmnK/uo9peErKH0nKCuqVk3gbxUhr
34VzIv4bJa4z/uxAVMRqJ6IRWh/p0NKgWJ29Dv1U5GlXGiQx2LSYIUCTCQc9AYVNd4Q3BiIfNGF8
6/0q3rkTQkJuPSRpAC96IcVU5Dr4N6wDmI1nWlBAkV0aql1WC0TlGsXV+S2Y+xpGOXl4BtOc6uHB
4DQLhu4Z7d44VFPT6dffsn8pBE20amDrqKnS6zgXI3F3s4l0SuQLs3u1+ewVqKjrAjDrrME4dvA5
6exTZJMxSV5Wh3WFXnGn7JhTjqv7F7ULDHx3wBfOJzb6UzJMFrREBjPrQbXHcatWZigK4phK5K6h
3ZKVablqb0gAHl+a8HlCGdq1NaAHEdg/wfy8YBIlpqNInzuD+RwOeMH0wWNn/PjcZwkwkTt2PzG2
huywvG6eOKVbi8xe3NZz5Tgaf8EFL7nhxPMS2jXlELa1vfaqbf0aHRxk4wUZtL8Kk8ig5kXivXmr
mcbzNf4m5tjXneyh41BHJR+hekw0jsyDX/s5q5YyGNXj/23FhRF9SEktsqJ4FNX6qYdXq8aKNiDM
ILQ7gcmK3flC7ODCPVjjWgXos0dgQc0GnZS75imfkGHbcY2+ajtce92StIT22sFr/B9YS4NXuYOa
+gpxmEoyU1FL9ZKZl4vgjc5t6VK6+iS+VkR2m0CIzQgRZEvycF8jMqzb4NJh3EZs10R3iYZdSpz6
pfEKbVvFj0lGqT/h0CEBu3YqhBHoK1MWlhsN6vXuaJMy7m4nXeCHrn16+WTmTasRtWhQY79PLrVP
tEc/rbTTNujn5hoBOmcCqA2e+YX25lZ5u8e4nThpS+owFbUzzv7BtfNaB2UZNPFiIf+BzC5Jqye5
bNgd6IQiJbuZbwHBZ62nPk1V/xzE5qMZJAH8IVK/iCZhpZVWOMekWXAHfJiHzx2DYCALexQNe46s
OvPdScAqXEK306SDuvGILBmcOGEElxsXC+R0RNw5vCpz4PG/XsEtotuloh3QAAmTTmPvNxRQ6bLm
2QNNuCcBizlnQjXWykvD6MbHGOJd3/x00Gl56d5x8f6tyJRjBBv9boFrVRav3CKAq4hsv6svnfNM
7Y3bQmlTCGK7P3pfWyWzKBZKbwmJHoWo9DOBwEZQOsfU0ZBtv4htCFeXha5t1lroMEaSduwCS0kN
HoBmAXfeSVBUJHnyD6Zhzk4GCPxmWuvWic6Dnl54oLp9sG8qXdkClH5NdRw46ekbpbKTyGiyHp7p
BAjJjLCbDaGHT9N8rWLTtZxN5luWoHyyFABFqu6ZkB12e4c3hWb6NNwxXVRY/naFFUPmxSFSPd5L
sp7ZZl0TNlYhyYPv13n9HgKcDRkLRdfz2DvBMDlEMT7XdXT4zJDHlqAR2Qre2DrSAxKctTCiCBBp
OT/C8WiCTDHZkeBPhZWERdhFJD/ytG7soI9c0+XLEF76C0xp+MYyjVulLARUtKYR0f2K85QDqgYt
mkrQObQ/kHwn9wq9Eohw5MPLHoqiei1mVfHg4RQZKfpDr7y1fuU2ym+xWYklX26KF3dLlPIdKsfw
ZbeowgazgnPMQ3V456D6JyySoJ2i7bKlaf+U+i6FPqztxUX2QeOsQryz6xLsIZiBedYnwut2CyKo
/S2hGrE2s5+0r5RiJpf2c0jo9ZZs2mhkhlw7ivN3BUBogvBeQ4mvQBZNvTxl97VPKARCml7IilHg
xakPcsE8oR6/z3Jl/M+qp2qZPH7pUBRL7Zzev/18vYuSZVKkA8jIDZgQoSktJ9r6wdsczgDKk8XB
YlQ89vXLd3bnzsLjCZLLm3nje5v1ycBtTIY8P9Gu8ju5nV5A8xWSsTabtzujh1LrZPsIlCl5f7on
vORp3HLFewfLeKwKLe5bCwgJqN23yh8SOCEZi46G9ZlnEOrF8jybL5vFYZ3vXp+gzHxxwF4I2RIy
kYXYfbTm4RfSQcOsxj1CRuqAzo5RFK5tYPdOZelxarFX73Cbs/oaQx+HmNqMrMvjgtLvQcWZ85RT
vyK8CODVPhXjQd1eEgoLZiepFByIVMf1IdJ633hAUN+avr001f8anVsP6pWs5atd65+PMGJQJCI+
w8UFi7xUqO/LqIzKYdYfraGF6XMaIE5GbOYvaEIKESG8o/bmmDMw1ZLpFMT25kpbdFElPnHMoydx
eSiU1QIflA7IbWAjpbTZzGNb4rMCeTmBHhBm1dxP3TmeuFhmvXzfvZC+TZju/V/d0EHfHB12/W8J
X/kk8vJbNq1Vm7DCRgoCmBu6WtQVgyoi3WVHraEermLcys7dxuHeT90kpU2NehV9Hduy0HQiyZwK
oH1BYqIu3e9qdTkD3SfAu0w7dPqG56FZRPPcj8HBnFMKUG4uINMVqEbqjE9apmQFwTtdxOsW4Yqt
5cvwi0lc6WE1p9dDRVA1gAXriGgfYkTsCEGesk+ZIjvy3n5YoQyxkXtx1/dFOV/Q0eHfgptjkipg
sldi7/I4yN5uZnLI14hlaa/It7vf+gEpoMdZmFBDrYDrybPDUZjBKBffF2I6tYf7QiIwdswYZOXp
DG3ZG4CDAYNdIU/bSzJdlHqinejxYEw2fZbzDggzw3ookb1sMyCFfzXiHor2jej9xDojOAWMRBQH
NEXs8VX/bgolJab1lBBhxwMuBmbod3Qp1mekVV/V2W7niBZKO22f1th5aj8N/EcV57UQgsY5ht97
Q5hPZsjANbdGwyzdgaOP9rMWVU5SE+Caim46+gHWmuw+8zwwU/m7QarjYmbDipS1cPlUadgvdJXH
B/CXMONSjfJ8/6rpLa3rXP1j8r427GsKEcSoa4Y+9gyHoIiBzO82wdvA0i5zDC/IOnLIPtcA3dq3
w00LuJPs96Tb1eFRPNMmfZLGWJeYAAj3/ina0F7N/JjGMFxtujCoN+z5ZNtM0vsFC9SqSbvLRsX8
C3VLmkf++AFz+6bqUapY6z4dacPHfIve+747Xm3ijt6rg19lTnFKqO5/MwlyaIlnrSt786db1gwm
q5FPvcGR9oxybiA5keKbjiPqIpvBH/Hg1UA/yuJIxIVb1ijXsNcb6QNkYtfLgzGBqTaeBn4MMNoe
fhwrZPVOla8RmRpSJUv4MsYZNnRKmHPdNAMeTOh6EMFVPmIpqvrqQJd9i1LX7r2CtOqNkXoO7NOi
2DB6bmHbKwqgSVNvfpi4lf1nhBM/c8v2ItI1WtlfXN7iZ8WljbJHFaBq7nA6s0SKTc4A/ddgY62W
kOOiyg57QtLwBzZC/q4u95f/ACIJW9ZpLEyLSQsSh37kwMTIWNN0kr41BkXmV1hHMzauarBQ/HNt
gXxec10xKEEkTh9uzt5zQ8T3xK9xADARus6W7OZ6A6Ev7pzyo89fNTs7yIDNl2zHdh+6a3TeWDsF
XyQHb4MJKQs2bv6tJRUQ51XUbAxzw9LgqWvR6IN6koEj21dFga574hJ2dIZAXjosOGtTmzpWQvJG
Ob/w2hZdo8TgvMKVizdE/H8XZAeZDYD0hSRjUow/9LwIvNLCnian6rL10B51SeoqzXcFIQv8bqBD
7J8EButuhwQuNITy+lvEuj0cKBVcXKuq+Iv/c0GutQHYOSvdbUC0BnoHFV2uRWowj4+bIZCS4M+6
sMn79Qv9fkZtNzx+KM13UzpSRRKklyOcROb38oxncs/9zTt0sJwL0oIbnNfA5DXesFQp46KIGUkT
wbgfbnKSfVda0oWmVNOIloq5j8WYAF8xh1nZVqdaaahhFOLmGmPsh18xae2SJjqBCowP8ftRZMKU
vpFxMIXWzC8sDkRTlu7eZ9jBiUFAbUmpKNLPw6dh/uwAuppVz8c8g9u1Pc7hCUp3hCHAu0Oj8xMt
wj494E2zT9bheO4KCk78nuvrwH5Lvxiwa9niB84qnfCZxiLZqdls09jChBc0jtAs7cLANO0lYzeA
4Lnkhsd56u8EYy07HlbN4/ZtEh6glrt5kRGzthmqKyR9i+t/hycemCMkB+F5iqiCDtARNhLXn0c8
9Vyi9JLjb/84+8i9Q+22psnjKUqktUPHZArtVapeYhkaC9PwPb0BclbqmSccWjtvlZ/ydoDiLPGI
/KXXL9955ia9QKynsq00XNN+5vcCkoOPYWcfIdp+U3hilaeKZKSyKQTv6KSDw2G72fZul5hSl41V
JPxcbXiOsDBBqLy4VlgxLe4/ZHyHXZ0kUGSjfZyU0B6iRwL5t0KBpuse/w/3xf3H+Iy5VLRdXH7a
rLsBskjYIQOKdkjaPSEc1Esx1xjE6NkEPBBc1iTzYIAbw2meyoQaND4lPyd1rbPR2pY9IJNgmmP/
F+2iHQqUdHSrKvjrY0F3xgKZnuWUtIl4aDteIWYiSZib4fT3zp4oZesSEhSUD1056m0z3CYm7MXK
BRisdPnBNgLT+YcfuRjZ5PVnZD74zzg2IuKFZ+vVA0Of9hks0f7qm5pJTv9C3reYjgBwce2u+s92
+Zman9Y7SPDqWDUdNGpBl3w1rRPCryR9uHmNlt3KR5HFTnPTM6RZXq/VFERtSulVBV/AgLuvILNU
Ocy/N5FSheNVkrUOQ5CUViiiMDsw0zR/6x5gij0KMRykmdfh0uieO61KibfbiIHDK4yBkDLoYKdZ
P0JI53g7giOP+nRotEWxkDSktbsONCkHg8in76FMA+qkUcrh4rKo2d2jtoneZAHmjzJ1b3SGYFtn
E1Ir76ksDR/RxC6NBkxZxXXEr4uwQl4lOCdltLCdbGk1jjLNv6d/D5v4mtY+nFP7m0GIHXIr9y80
nr8pli2qvPCge03BQCN+O3oeNy+/AbXZUU2m/nBhvQkAJsxtABze1DCpFGvC0Arz6ejTnRR+RInQ
4cbqUgg+/oEtDOVkgNzaaZYYbrlpAcMh2mkr/nw9CiI7Iav0QyBzDuqXE/6T5nUDS4I53K/rFdxy
aue4shaMEv3teuDzADfc68qYCSJ+sl2C8gfXUFE4yPZyJk9CE6gajTjHZy75lEvJcsH+UvyzSPVI
zn5kJIMpg9cjk+B+0+EcY1FVGinwQmbiouAg1aLsIPeDGBKwGndGjsy1SPWIVXWcYEQc1E8lyooP
pWjTkoZnrH0A2gw7c8HOYJ9KECkm0pfyIn6AvP1c9aXj7ePbJo6Gzl6IF6DnR5BIZMW83VKoqAhI
zsrmC+AHZgxDJWI0gbLW9Ree5YBlBtzEufQtDJbrJrnyqTgovSI7bI2gTk4LGFFmIhKRV+e89A0N
T+jbgta3YaUFdczVtKU5XjcnDlutPpJzWVTF3g1n2AazXNBXYZUtgBHFXLWvG6XEAjcT8jkiiaE6
nuWv9c46QVdvAwakTma9R1kFUL40DFZwZ6qc+eGnOXQVmEFDdTH4EIyDh7fYKFG4vuRMEvP3LD7A
SHfCbuOjtTJ21V47FGVaxyxrzRk45ZOH0k/ioX9knZeCkvB/kBPbUPSR5ToV5QsJIlPgFi63+biM
krWCAc4ipKXBkc+G1Jmv/6Dt5BZLgIawCZHJ3w7VwOBOJExBVC7jY4uVoj7rbNKdjkm7Jwybr4Mn
zmEufJb6uAR0LYDS/rcRT8QXmXYn40AceV2fGUY7q12Pkpf5OsRzFCrAl7ucqJw2BDigtdzvYFKR
icm5tyYP4iwRIvkYMN5SzLuExF2EvpI6XSyZ2SAszwe+17kwbiBsOh9OwhywFyJqvZ/WM7oxfNeh
vPfVUcat1DMRDTh9FtVFnurIe63tkwI1W7ChVM3wH5M3POBbILsdHel6xxygQjvWUzy15q5BDKb4
ugQ2WtxfGwcPH/2/amLOEF8RXh+XWbXX5FjYI1jHQDWWkvyGQWFNMWQMCVpt2CHwcCgq+RP8fuN2
0pGNPui5w7U/c/+iyocfyPHzYYpBtjvKrsuenWMoM1LfcF9f00f7bZrg31tHlfrC84JapcAQdfww
gOwKhGDJAbTENJNbtoG+SLSea+ti4vpE4vTVpvgPeqBlzoZkrbE32SBgfzU/L/Cm23Z2R3yso9fM
XYoAgr9jAehGyBQBF+/0EUDUzwuvpgPXBWUixFurYY93jTh0vtaUEGq87A40yacds4HAS5yFK87c
3P+hFAlWuVnFe1j/E11rr1VPAhnZfaAYXjZkAC/qM9f3BhTN6fofcJQhR2iSM5a6dKCAC92CatNK
fkZhqyg8gUR2xI8+DTEZj0DO8g7nBwhlujmPzsqVDXcoTgc9Rb2gHMSPzN0lQW1tskEg8lOKSDzi
bUiskMs/YROMVk/Kfc1IZ9Ex0rxu78l8pXtH/w3o2RFYCpmbX22DjElMeiLIvn+d96ncngY7DKdR
B4gc0J/aThIirZgXrm2SOmlWMlVVCZoI4oDbupKtIXxIl8tGF0YdVEQNOsprW1jn0yo18U6dLNJm
YkOyPd4BOuidKrwiDlThMx8u1gjKTLw/pogCPzniXinZk+IiUrHpdwlh/0AY9v1kG2oBh0ssChk2
AK41BEDy4BZSnG0IElYVSaYepTk+WnvK00Tk/LWvjQSV+3VsgHt9/ij7zA+mxaCqOt81u9DH2UO3
EmDy11Q8eV45t7qpe+cQ1ky41AW7i7tHPqz9va2oa0XXTgE8czS0JLUZdv+omF/xLLXV27G7mh9L
RC2vkEgJZEzapT2iWXlwJGBP4ZKbV/6GvoqpaVgnAzH2fXfoSMLm2VzdDY3d9tW+nuCXejAJbkYg
7f2fRRbHXb+YhxoGNrzuj6i51lzAm8ByyJNlsG+zbCKi5duQL2lmIj26nTUqvjFRpreY+ZhN7sQk
aWY9iJyQGzQMk5zekmvHiJnErPvB4Pyjpyzsd/SXUiDIDzzxH2K1B1cO6Zm2LNAp0+SVmxW94+CP
huiPeNTuszzDS4sCjJtr14Cm7PU6hqnyTos7ItvFwwTcGIgbl8u0pFrd/GeFOMkTDlKkZxO2osH2
5euiSJyOtJQ6qM2LG6uUJCtIaTvKjDAB0UPj5QqTOUu8XIdrnygL9VHuE4QZpwR1EQ+40x3mXMtJ
vatMXv2wRnweUPqVlozNO0mDj+/eLaD2j1mRwhgqv2Gvev7wPeooXsE5sdoRuqwl5Nw4hH+IhYXz
WTcJ9p8kmbU04WISsiACr+6gvbyHIwc+860yI28921BR3+tyV8nAo2rNfB1VE4ffBQg8LFLJY2yu
6XBG+xyqmpE4P+N8MSpyIBNqYU88oNXbxlLOsPCZ0kxD4aIQCyBjE0dYS3EvbS1Qp+oRUlY/mpJV
NE5AOQIGkf45+hof0S+W3YLjxNWkxlP+rF2DGfl2DIlhDzLtzK6Y6bbNVY0DWPQVe9GxlCBNzQHo
Vq2HDjwI6CRQVE1MdHDGWTbOTKj6Yfmw6Dw6cjRX0MnYUduOnq2BTmfLcqYBID6DXRKlVZxQblnx
+fB6yhqViT8dKQ/RlyyiCkFrOKEj03AoIAVUtfLsLgHB2FGNgbDrH4v+EN/B4e8ArRcJe56J0KxS
LIRoBLP1jeUjPPeF6TwarSm5PfNfDKwqlf0pF1+6GsFEkFkRsFozBrKH4veuoJhW8dgKnA1kZJTN
0+sxT+1o7X7ZlltHPCQ5ND/EG9jx91xRq87i6eF2fcTtebwwonmQoajFAjXiEe0pcAMi3gFD1Yjr
6hWjignGjhiUmp88XTzusKsoCYKkhEtPzMUPCIdv4Fa63AfhsmQql2UMyEzAz+eHP8IuFUx8iljf
ZRM9X3zACSjjm9QmEHeioktAYumm564ddVducVHqW0wXMu2+yF7kPnIo3BPi8zfNDzlBMdVTfSAi
i3rQ+RhumheBtzfsK0LF4U26m9fXE6lY8tDJzb5Jhpo0ziYMawUrDApAyKa8nwPc4+tsx31Vm3hF
5I+nB73GV48fXWDUBfqvAVXkxWzYK9DBrRSA4JbuySaLCFGRPizbV3k3jh3vxuYT/6sJoYZUk/no
1dwmmgjDcnPCkB+KKkvr/B12cZVO5AadLrYaoX6ZmiGuVNuyInUjzp/rknBA9Yr+ahMNf/McQsvY
GQo8RgcYVJF56vgYS1A08jL/+S70NrnBYN8U9eoK+piijDfKyfSwj3yBKnMGcY2pUuHULdeaWV73
JWr0SaMpbxiUYD2S8uRDGTE1PZpLYtmg8azdn/F736QV3Zjyq+AHtVCclAVrKy9aSpen6BGD+wY4
wYeY2ZlgkKdgUH3UuBbri5JvXVx+TZzpVjaMceGG63sW1ssYmhVON46Lavhzi+99TlQOVa5SW6hg
/HI1LoiWrPdlY3xYju6PsxHCiVY4FtOJh2H3kiJ5H1q2wuBACFUX444mS+f/jRDHAkWDyDtmVAhf
NI4/nZDdw/SqtF+JgyDiqFiJSfzVbrvSZ1SsqLswEkUlnokV8Kw7xjAdFIuylEbXKu5DWGWs7e2A
m9JRjnctfNqF2btYZftTlTSJOY+ZyuE5YwL4gTShi0uX8irOxkKdhMLjUY6vJNEKz3Eo5O8z48TZ
QWQ9oVtzaPUJ7HODW4QGs+V8DdHHjUDuJ6BK6txHtN7/OQy1AEtOn+nGplTPDye1AQ0XCSmA+ST2
fd4P4g6Q2WSDVzVwtvP6EEYE5uOprjNwPvkT+dPVSqqwDzWxIiADKJZJ0cEszwPa2xLn4Jcedc7j
20ZNZOnLiVI0NQyOPzJvW6Rt5Btl3XnA95+ryrSdOicIHPSMGkD/0MV1cUxBt8sRzEhAr7HGCvFw
sB5NWFgpXws3GsegIhUdDu5kdEyXILog5t3D+EFQkKYToAyT4qG4Yo2PeT7TpNOVL6Oo43vcc5te
UybqpfDmh2CgTqM4M107x/287vCcCQQLRbMPYG5BaBUwmyLAEvRz6Yk7IImfd7Z9fli7FcXJ34r6
EHMh/Pm4otw3PnS3uy/3SjBdO9WJNUc/CZi7qV0DCfcUiXqenR1SHU8MKiJI3a/e9vdsMCfrex9H
oIqn9Qg6cBM1AMf/HNkhOMPmiSG+whzLfxFaQwBVFMgDr/ZEnXPwBFerOnVazKM3WjIVxRL2SLh0
BhTltAbTmRTRDRdF0/E0FpaRQQ1rzckqqy++6mbecASNMjiEkBSMGkhy7TVBb+6DyEqk33FE/yPy
ay0d9fNJC3cfm8t6Kv2m2bCoIB/KqI1pcLHMhLFYO7uV+uk3v0s9vnDaxgMiStKxUzDQmzCv/Dls
bddXdNwnjYqlFytOYHgZ4AtbPUqeQGgryWo7aJiSfvOQAFo5rVKtICa+lrrFp6z+jx5SFdinNIn9
+J/NoKoNrKVyqZfYsa02KlQIwmN44ROu0OtyI3/MQ/6QJ7RvNcIwXBZGYGfNNP97m4kfzFkm7+r9
vmXMKLe6zubBP1ZcXm2QQB3aX+ORra8EcO37ByuCR/hVEka20y3N5xuF20yv73IFKJiMsWzl3/gt
HXiy6vFaKRds5C2+ClBKP/bBe8QMGHPYKfMeLUQRh2PmmESjxOAS+DIbcefK+4WG8ytqTBB4ACig
JaKSYVDbuVoActEas2hl08XHqiCnwG9W7HwYu/tPM7xZb0QnBQlkQqfk3u9VBZNEtglmtVfDZPHH
LtfUQ+Xz4xX9AJfVK+jzMRtrSx9IUbCM7IaP6FbwKe67/Q9pKteVpPWSY+kJsYwhw35829BCc6AJ
vbncq1zrZrirF4FQTnR6/CVdGQKgGg5Dn2PfvQOisCVnkzHSz0ZHh1DVVDcVbZLLxFHITjqJi6PA
7gjGNC9qHIM9OHuQoAL1NWdM4/96eIVprWEqwhqXkvGTg0qBHRGiPayAb0WYDcSfSwdszrbVBh61
VO+Qba/m+A1OB3VZIVZf4F7Wd/uWJqcVhCN1/WTKI74WFwWfpLXzwEQvpDMMZUBwn/QpzHvvj7kM
G/chGAOUay5p1Q/o64zZLTGDcQVUlmtGB4U3oqI2WOnK5PnoOxg3UtBhtc8B2UMiGL+O5Q7bavIC
TZb9U3upwPIxBZFb6rHMPlBZsMrHJO3uWp5h/n/sAi8o2GxcjlCNqFzRvMsro38mjp/JecwZIgxp
rjGVR4Z+sQIbEuV6ZyefAIHHokH46UDN9AaMdxSA8oca0AwyPmdQYPUqNcPhqg4rzaDDmO0mq86P
+2qyiQ77YjQTilXDu6Ld84CaffqBcCAW2MyJMTnriIv07dWC3thq4+FXSqK1tk3MnukZM3ZQaaas
Cy8e0QVIxXl63ZFVNi8BXFpmEqRRvxHQcxeenSPp2KmImaexWi//CT9cFldYGSp+SuizdLas7/mF
irmqgg8tDeXgwJOERKnKI0jHegZrkZjUaPeOO5KpxHnkN8nb4ieT71x/nnLK4IehHqxBwDnEpy5J
z6m/1MKwPxOMWfnia8SY9ej+jzem8H8380AZRqJYVNlASbaz4OVQ9y6refJBLgXlXAfmgVyFi3pj
La8CTM5y41z7wLL6+jucdt2olDON0bEilpeEy4UWnk5LKiPejqLhCKt75nbO3S+mQalTPdmnBxIa
Yc/PwAizTf66LrZmb9qA6dXGJAfXW0kk4Werl5Ng2SQn0rMQWorCcz9HslVKIb3tennjUSerQ2Ej
m5tO/n91cpCZ93lujS3Umvs3ZuqM2Va8bTq/X1kUZvy9+eocFquVfHSQrCYirSMqvKXCQy7HGUQY
CVjk3FQbi6958YP5eGElIrsFVOaufsRLWSfMIDwZqp1gEjcdLfyYOXA43298HsWcxKxDW2KgbJhg
9d0n+lsf9PTTc64Wpgew3//9qleJdJyWpm+zPnDiaT9D5/17kMYMI4X2W6Gq6P5+1j71D3oeiAQp
6Cp2fp/QZC6gC3ZErLefctN5V9kKop8bFC22D2qiaK7RBanGAtlXWwenfD7vclXzq0g1KGl53BuQ
lJKNIsf8a0Qkxc2YqkM0VastfCYNB3xLrbWAZ/LlJgYyE+aMrcmQuAsIuMdJLnNCfjloEDQ14SrA
GS5xnfXv0uvUpeMepKfEqe4hgE2s1P7AsUvcmENaejcNURY6O6zS7cWQCb6zLLUVU73ZjaQm6gJ7
Gpsji44wltcNYFk6QrxSZG08v+8o66ZTBzWNlDQYUcZppkx7HLJ9IumIg3acSOF/9ku/oI4xfeB8
8IGtWRGTGntZ4zyJaP6CRW45TroFL0AhRGCzm+b/b16KHAU4NeOrlqpleDWdIQQJ8LpWh/TKZzvq
SCppLBclbeEzmQ7Ukebe3foJou7gaj/UQY1iIzjPLjWR3jx9CIml8IJZNH1ocnXw+aZG7Q/pAEfy
r827yb0sexmWf/IelIXVo4agzHSkJd5ArHA2du7wjSNnYycXVTuRSQYlkEq1KJNjR5v7eVSTA02r
PZySZVwC+0/WrkLmbQ8KrljW1wPecxkPR9NKOjxQLMhxDa5ADpGzXka8MrHJGWRGINnOrieK+4hN
Z/svvUpgCW40pGuaJ8kel6jiT8I+vEo+hdRgPO1s/jd3TeNp5QHDfypjRRELXJLqgdVefoSIlXo3
OIk+8X9RdyQYOOMmcQPk0smt6nG+tMXaFmJR27nM3wlQz+JT4Z7te+ArHtfjNvu5fBMzHabCZNhG
48eAYC/suMtak5r8NWN+QSrNOVLG/+oFRtvZg3W5BpXeCWZokdeh48QXO3+dJ2HnkDTsJPdmtL1e
tH8quVFFKNTMpkQ+0NNqFC6jvWrFvVLzJ0lIYtGSsi6FC455dulukib9Sn8t1kYdHF0Ho5yD1MSo
OapDTMhLqmH2fvRVQBW/gn5xJ8x58aCFiLz2a0R5zkmWDJtg9w5yu7/G/WmO8VcDAnyJe4OzJJBV
FLpNPJofyYQRTp8U5rnwy3MKMeHi3XT5R3KMCAP+iEfUEfFhBRXUR/sndH7eSjvKfMeEm+O68Dai
tB5Sm/scgGE8h+sD64Psv/jrB3kgJZRc92IZAzOcEC4FbckA2FKsi0bBIBYwbAZLvJrq1OGOWf5D
qhixk7stoMcrsNtV7aIZUM0pd/zhJQ9d/gwFjqLn+G/QJwaGNdwq906y51FvPvqRgPK/P1F+AYer
J+xIc6p1O/NZV3JG+DYFPim96310e8iEdU7wxyfGzsqsAyYA1/wILGkBnVJzLRv7bsAAt2Ggteil
3pE14vRMPLxgI2/QxmPwq9u7hBJFUbaIXq+UUz6R/y3tO0sbr3jU+DTptQRasXOBFjTTxmHYYxd7
3tmIAQPEmJD9I4lyaYpSDmXykWx6yzQgq9JSaJn7AUzgZtCGkEYSlO421cG4qUzbTuYuwbFnLhch
x5cXljkO++XjLfK661LWqH5pNvh+QQDSP1aXEal/Uz5JO0rDXhqCt/wgW7AcQD2pas08ZKb1Z8kC
QZ9cvjEZAy21a6stGosLGvjiuWDpg1tW02qRgbvgBOUve1V2sEq80Vd+TeUC5+c9LW9kzHJsL1yu
n6zBczlXPSIXLhAbzktpEIegehkrZ6DQNGst9P8ziTY47xe7qlI5SFUh+xrvTuGglHAbeYCOuy95
hPLXVJb6od+QfDZiD0hJdC6c5zESAoVGrJlfueVrIJ5uFGTVslsSX277z+M6fBIhw1lohUssgaIa
0ENAzb7PDtWhEmcu3f/V3km/XLACdbKkEcn4GZOsLyglxalfIdxv7JCl1Pq1FkoLvGRdUYvoXsRW
QwahxlKGen5UZ5bwRx/Rn6FOLNWJUmvtDMZwCfBBLpa5jbeu/RQQcs50LBcz1UhBCr/MW7P7PhcU
Nl8mkw9wAFbNWKx9bZLUFLeokAH+d8X+6afeWK19iUqTj4XWkASG742MonBIpWzbu85IYqB+wQrs
6tP1YmrB14ihS8nS8V+FDfoAZoif+eS/rnO6va1GCqBiyTLv6atv4HfE/38IDmYg3EDH74NCJAnU
DwgVZaqs2sCo3aN01xKRFDcHLLAm7Lu0d0F99JtqwU5c6GJbtIx9ZV0BuKcwEYYKr07mweIm59/W
uditf1qXk3wX9b/HLUXzPi1zO3zT62b0yD4a8YhmfE8i8tK6cF+Pyo2N7t30fgC2EEmgt1g6GlE1
ZxUGorDrUN3epz4tVxHJ3WMS1LUhMsvx7XIx9OO7KZ300p7jPcH9Yz8lHiCcgsy/mcwc7y8lRbkQ
RPbeV294Sdo7xan8dcXmymEyRDcVGgy+z+42ww5HN9yfXPo+VtzV6M5CL/GpjzjbfNgE+M2TKpsd
Mt64Oyu2fmXXJFdPMQrS1KGDnAAijw84JdNuzrOAzlKF7sZmf8sCjncekA/d3Z+cO7I8DFqGRn3E
6KwFJMKjId+lNlHgpbJopcBjCDa2V2SxD6zlhjNGcQ0ViWDe8Iqt1LmYG1jsQ77M0uHqLHZcm1b7
DufDl/vMx15YdiIrUFyhN+rJJBwIj4i9L2Gjg0LCgSXTaQVQiMW5fthxBJQrCr7zcHjkOewp64WA
njJP/7rBNkFbWLABY8NgoTBKPGQ7fiL7iBtmx4KLVc0z6jMCLbxKaOThsJL1bOklOCaMQhC/NxAH
2JYLlgghBjUO8YwsUdHw4HjEcxjGN0rVJh1VQajgYobbyv+u/xTzwcNDybnQy6TEvOrPWue6/v81
iwPmilqMqdSimQn+eqal5Fhd0lLfC3wyPlM0kZTKAkEgz1P6UwvfZCZ0eLC0vMimP93QxT6ngqHI
S3FxxCW5W4vcx2qziFC8buuJbXboPvfF2LOJTsfPbL0ANasAbljKTEeCOLVacAGMemZMbUm/L2er
yXaKu1UxoHh9kxiGoAhFV8gscIREq/hodsNxH3sgU5j9AIO2UldgFzj/tqOS0zhAMQTZ0xiJqO/R
NlAuVu5M2yS60//y0QKWX/m0RHIOZzyH7dUMFzCPAt2nfMF1Fg2kUikjnuqkVH4V5BEhxRQgpVjv
ei2iPXU8aXc5NjiwvnDsskLhAuAdGiyMrUf1+cRaVD/6GsfGP/wgE/1RhCWkcM/g6eRQ7vG6l/A3
JdOxI+saglP0pGAsw6uvWM37hPSpNizTHX+46KIkOdUg6fj+ncc+SlTbpuk7SxHruw4Fhw7D6V+n
mlOTSl1E5UPzAXsA8CkuPQ10QOYR+TZwa9JzE3ahYIsIHq2GmXBMqNegDTC+Qsh1yQcDjhaBe0TN
zVu0BWaRBJkXwJ1Cxa3sY+eXStspJaFDfWL+zjtgx2SnbWzIF5qCLaGz08hyFPJY62HSdkAAS3/2
x+eflfsZgIAKwyxmyvDvy6MuSAIleSCfYxFIigTp3WAbmXy5SPoTMMbdxIxl7FYDM2nuZBAoQ+YC
q5biEkkK59wy2uoOkSPcgsPaddsydFibz9ZgZOvuniycpM2cJaDrUQWNLDYkw6dwP1HlFPbycyqz
qEvMIODs9dd3/YHjzJdLBoWrj9oyuXTh5jXDdUdRs4NnCK6CQnaHfbOk25EgFiHzG19oZt7HmG2T
W5gd74d+bOKGheBDr1mXz+1aTkiSHIopiNZmL6+/HmWUrcHYHVnH/0/TB156NNBUKp6bdoug1IMS
8Vfh0K154SWGU6cYc5YxePXQPBhSnC5stezGVkNd2P+8atEVYOBSrTN3D55/B6z54dqFFEn8GKUK
YqqyBDHElktmyzy04OEdy1C6/818dru0mQ4JQ6WzXYEcT2ZVLkSXcAizElGrI5RgVvhYJ6KQFIEq
eVB6SzBbLYJDdgvUMJaIAtg90gWKZVr/oh2u+ILLNtlu2mR+Oz7vT0o72M7m7cS202FKlS44VjEQ
PumPUXFv4nPhDkN5K9nGpIyrJ77Qzz+aJtNbnXOjCS0cOqURMPcrM+Ayp/1emazMixoFiwUIrDhb
B6tKVecSqRhWcxDR1w+u7EYawz2UUymmSMTbLQe4y1kO8NL38RpQ+QhjMPCjeQYQUm1u4E4R86dm
fw6slJuQ/e6zntMdo0oZJnBb1OqEpYfwbqG+xVTY8YWt405cZjFEKWaIsiN43NYaNh3XhCbZWv8m
DobdJ96jUXLem7HmGBpyevFS2/1h5iQXO53wFqISzb5F7TgKs0sXVT35u37pVSdKlPVgNhxSQMOJ
hE9pLJ6G2ZJlC/U4dI5ZdYiCA9Ly83kVZiR7kfjx1Mz/xR3u5fCHqy/xaj1uQQiPQpmwqcGOdw6y
cPHgqXOK4FBo9kazluT/NpMdfySNh8B0DtgPK5iikLPZYUI7QE4HKuANSwjpFES7pecqYCotvZwm
s/aZFdO4J0+EnuI8xtH7VjVQYjiCG+oCA7+jPKmu2bB5DfiRd0rrENYde+NWfZao1VGrDjXR+rBJ
g3xLXHobUZHCVKUWNDeqv1y7mVb7nkpxXsOkZJHEUyFlEqtNr9XWdbIFbG4u2e05qyNeQM8HOLsY
uhX671YxdDwI46ZM6CBTQe8EEPFu6+s0LcU/28+tjSDRxfIGebrgtl/a2Wp9HvfhIXVx+c6HIKWF
9xSRdZ6H/J0ssGKWV3LrPCAsXGv6iZo8ksiHwrLCNrdf77ARS8iUcGnr2F9dgo4/6WYk0WidPa8L
ExDvoDceEUVRWR06GJgDDpDrDqeDkuB+c85SOK1HlbaZpunZI7kk/hL6VLsiSezt/ytefouqt2dO
uy7Tk0btA57MvbnaTNo6Gy6KTZaphpaYH4WyAtI4HrcQUxh2Ra4iA5SRkxWX16PO4ewgTgvBM6Ca
qSQ4oIawTk8D/7Gu9YuO2HiBUvDQ2xd5hF5PPdD1R0HKZC/DhVuwr+yVM9rYQOV82JpstbiDb4Ry
KxNxFHManG12V4Z3saipVYuG8lPkAlExHAXDDI6uxHIlvffcw0WjO7RFQ0AgYBUA8ZKv5Kg54xxO
Y1RZQQBzKRUoqCo672Nc0r6r7Q3D95RS/stABOXANpTj2RttALpYp+1YHLrRqAZ2LuSYLUkKDVGI
y566i/nHJLrxFC4gRfNVW4Nq1yK2jQllbxw3w1tKjz6wkI37n61VEH/8YwgltfPFcK7SRWXWSVU5
lPVspKp1yOegLYFwDqiik2Lx64hgvY3bA3nyAuwmoS/xG6oTRAxME1CL38pOLjZO5MZGVZxShbOj
2lKflePXQdeg7/crx4jMMXp/U5+Fw1FHRDitCEJ3mJ82qNoi/xx4x5itFW5BsCCYJI9ai/pkts48
eccbMeNMMyOT+0L9/NeekpHfDdsgtQhtVEMqLhOmxycD1qRNkvPfMg1/ZTETWPt8ljeIOZcPHTTV
gpF3kn5GcY73WXCqeYvwhJtudkWmsJ2OJPBSwwgAZUMGFzYoL1aniqk8TsdIbCRGMPGpu202crB+
qmSCsOhvEIbo1Vvgu58CnIrbW6U0i/4jiOYlypJApG9YndFpu8VFaJGoU8C/oUZoEnKjTRaPAK3n
UxQStRe7/mxOSlqKptC1GEALka9smuTeOy0WzZWd9jmPRxfvEi3uWDWWs7IjS14gsXCMlXPqxbeK
qK7u4gqDR2xViHz14N7Yw2dM/6RGX6jjoms7ShvCK5av5Ekv4v6R2MrueFNf5pyh8LriMdCuyhNx
Cu6J1C70/GXIgGQBuoRSom11vb5iRwpSgP4G2d8a1SoLrYY5ZRHZXIubNKHMUyrPVbWPSa23sKm0
HMuvR3+ZaEPkC1jFy51zeDyEfwTw+7qv/gv3Ee6p7UNYyKbzjvtqgGxLQT5ylqpSiko4Jsi99gmS
xg4eHI+Bo8U2347CBYM+CZkI8ReaUjY3yp+fyMeHLiZ56zSLu/wYDTY07NimPLbE3KspuN6cJ1nl
DBgqx2uFxOCQ8DQ63YldQhaBkH0J8W5jL99FG/NCtYFAzdlR1xRDjrqBjz6fRVjjX1oi9Ibc5SNB
4a8m+1HIEfE8K4SWB9WdawT4/hOl0Ax2gNt2YkVapclVPMs5WSzwx/ljs7IQ4Y9HCzrCXYTrdeU+
/pkWqs+tEYlKHjrSEe+iASytCDuat4RJmq8JTk1P8l9/RN/PradPEN+8G9RmE8g1Nk/uybhAbmDP
8qZFSS1k96aX9707s+1l2LVB6PukVhq4gv7uUOaY2BlhdAaY1LRJHqLh/uuMLo8wjYlSo0dF8YjM
Bq0X+EZDTedwV4O4KuO2hZON0oFWkXBHFsW/Q8WddgTSpvfybzinHuNXkzEjZkKr7kitIIwmwQ4c
pT+hlvSmSOy/l2bPcxywzKCK4L+gJfmv0gcJf8C51H7XVd7LxzZ5mik51DwN4KJ7n7R6jOONC/xj
UHQL2AKaAYLnLGgOe2sE719KU0XJDSv/8Y+foJkLvC666oURxgyh7ip6NJOs5NOG6np7Fxlh2nAA
JNw88ys58sdIEkLuP/9eRIfDceeaGHal9VW6qAM5TVZPb+aHFlAzJ9vYVkQWrEv/fuQhyJpP98tC
/uhFyKwhQVrTmlKNVcZNDqq9lZITcrXUBnTF2v4qiyNJiFu9t6zMPIryZaq4Vp62fBgBH1316oR1
1PWsQ0d1vd9fMgaQvbr4XqfVHlF7qfuxBKm/10ADpnG5N52OyrG17rtp95p3MMqrvJmdvjL3qHBP
+SFFXnxb530D+4CuKjFQrnqbTFw7M/R+frOyZinojCKR3553f9rsyDdHmooy9A1btCM8do1aiNJT
xthzYdegVWYbiBOz6gEhLh/Y+8r2GKah1YNeSV7Id6YjKaDMR1rQE6Sbimz+gRofI/HE+w9DsAh2
j7wI1ph/hK7VXXf/X5oXng4obr0H7Bsx/eKTjofFRZD9wtIxHT9pGjC1rBEj1EPUgxcOScgN/FbC
BPP9qLpCj42xuFBHKrgpDatH5Rz0GsAtw5EUcnyOU95WMxnvJYLBxUQPA6jBqHI0yQo53z8T1/+r
O/UPOqT+6wFuWtHlVDkBJo/MvK00IR1RxYgA3JhID+vFZS9YWYmL4l6aWOJbEqEqf3Dw06sdEtc8
rOH3XuUH73ti5xtAGLQJ7TzOolfQ8siLDwSHoqy2fMp59kxZuurDRkYdXN7Cxn5iE30NjbgyMigf
BE1DUyS2yhC8Acvk7Q2y+U4U8yFhFGbF2ZDECUC/29iRlAb+MODZybFA6vE7hHfSwPT2wqvP1nZi
ImjLwa4Ije+XHRWuO5KgyaQxKN73WgWSbsC5zueIDp+BatHQ/m3sdJNQgJ/7/Vv4A9oFGDmqLmTa
uQvnunqCa6rBkGpjOKyPRHZEOT6oij6aY9ifj40/eH1+iGO8QGIJkpEZkDnTooJsNb/VuITLAwtk
aPYTLsWupBJSp+h9SH+Sx+m8piXpDPLLXF7aUfGctruvr9CpC6Q6V5XxDLaAoeOjLrzAjmqGR9C4
uopk5hI8Qa9YT1nGRcoPrPdOO6sLhB/EnawdHxYGsXI02GLHyinZLJGU3LKcEhV5KpwM1lmn+SqR
p3+LZWSHH34jhJZkCPmte5H0biTlpRS6JaQWUUPXOERK/xDcLKImDevHPbYZM/UStwegmVJt6G1Y
jvpwTYEPpRpw3sbzuj4Fk2YEum195DtDq9PUvOjMQDPDf1EvFLCPlqgj+1hRo5iy0HBm2pP7Rtuj
21bsy2kJaJR6bE+zpjNwX9Osnx4ISCI5sOQxzxefQsm+MNvtnqs7xYkV1adznLVCi77O7ZttsVHo
bK5GvnwjHE89NrfIISg3p+FncwF0uVFT6C0cRNeH9L669pykgE5y8w0uw+NmFDDwu5pZdTQ5uD7g
AfZ0zdBB62EKE1rbgjVoiOzmaCq/S13etuuIPjCXbCENL4bG5oNGnNE6yz3/xyyIVyewShpXezyQ
lNmVn3GV78yJ+C8FASJY6l3VZIbz5wDZx28BbkvgZcEdVxc6CGWeb2COBhk6xuuOGdLLfwEOh4dW
04OeGwVIRuzxlrjoq2WalYwP0lLz8j3ElM4Ho+ofQjiSs9HG3peCo25LXifk/qJS1xAgoKwTzWsb
RTjhFJvFPSt85S0PRHOEu6AJZHj8n/YCE8BFTq6KlMjirjVIKWPSeI9DpVJeOm2qsTppzXaoemgp
mZn7P+zwviuTsk+Bq0OY9gj9/CtsWCz7c3B/9XGkFHrKykbG2fnC4Go+G22syYgchYYRx+Z4rIjB
Q7jRPrOdCXGU0QnhKPQ/lk2JDXySrh5UgMs1SweFpFtPIoFf7Ky2iEb4ORLW4ZPUyier/rHY7Xnw
sb24ComvxKUYJrX0Q1Tn9aNOK15gBLTsWg6cRj/6phNkCFWiSjtf9X5UqS2/9K4xmEBQuN6QawNd
u9wtX2JC5xUMiXSMvU1gxyoq7xBuCbINGO2SCJ3EgZvrL804HAzAdVGlWCJv0y8NV57oJmBdS+6N
LWuLoPOu6D3VuAvyloxDgfCFGcL/ujSoBcsGqtzM2oNd0gnTe+D1gv9uaMLIi1/XdNHPTYrTO43o
3Ma/ZurwyPux3QrXu6o78FmkYcE2bL+r6HPxyt3Ygo3kg91cigFHdq3scoGdPO/NIstBcVqsDAlU
Ao+MHtWRtBl/IfSvkaq58qSyoB92boEsDC93U/+E4iZKzhlOzbwUWgmMW/5UY/jMMkhAYuXNYLMm
TPtzot6FSI6Z1ubgfVnWH8HFYNMM6XRK+2I/9G9RNNwxM9yVEnr3nQq51kKezWZglQaopFmA4h8D
yYaMOx+cC13G7c3ocXuv71jVbEo/B/8DLFPDioeVhWa2t+89t7znHVXZ9eWJhF/hnbhOw5pSmOfS
r+Sd1s33+SpfDkMLwVyJnTxK6htUHAlZAPCx/0hO9Z5tFmNyovyHYd2YqxQmgOP3KzNiGGNCvWpz
Ay2tpTnwC+EIG2UePk/JBQjlHcdkXUDlKTMdLrR61Q/NO2caY3hGmV97n8y5toiBLJsUN2oB4UdE
2B4riJUYE1gHPw5nuFqzeCCmZmJGtUF0gGfqoiMlWSBx01vhNQODwmMuJ4Zb3bsYK+aMMF7dDKWB
fR3pJB49XvFyy07EiWMs9uNeNKbrL19TPcyoVNfKlVQ/JHLL1I6b0suFFWqaTUk0dNk37y8E9SRg
pGOm/TBTl2ppVM6+bVISti/XBXYDMPAmncr250OLL5yFYRsdZ2B6YSZnbVD/pdqTaK2eFZ/Z1l9Z
Y5LZwCd6UqY4wjjCKov30qcCDhpziRBbvynBPWYClpWsWx1cnzSPSACkq/hu/amp/+ChzaM8dsNm
1+5htnVekDUBYZeZSniHlizRcug8QMtTOIiiApw8r/q/RUUNWadJn15/wKerW+ZR2Z2c7dqgT8Hu
ASPj7wlKElQ83WkYLXdFNjENm+F2rtthBU6UDAoNviD759vhviId+0h/guT5u2VvesGd0LoO5HJo
cNoVxFmlMRixzqa0MIeZDGkFoenBJltrnvDAROf3RYh1U490zhfA8Dg096/nQW6Jn4a0a0xRevpP
sCFKE8CQXk7ikRx2vcOLbNohoN6kLFH4XEmzPj7WWaUjRoJH8YE/DRV6UCkRuN8wWGMUbDL2F9DS
SJR3lu2bjYY3wloL/GfGyEycGMC9LFKHYxsfWjj3QJGxmfQsd6FjQ851B/Smye8zbVvkJnEV0/Ct
9ZtXuvpK2o6GInw6OUMEzQFyJinRZv8h0D/nxWXG9TfpNojIswHl+55VsfW1Fu6lqCvwAi3/xEuN
VLQ/FaR4pWtQ4gEh037kTTwg3rR41g4VE01ib2qyspFr7Z08Vhl2BQYHQ2VawGEjoireKa5nhNRe
yyGrISAWRAtxiFW/i3Ph9JT5/JHV850RMoLhXdLyiV4wNcrtnxDouf261gUCxyadgkuKroFdIqQq
1Prr+VF/FjFROjWI3Mv1Sc6aUJ6+7rEhhln2xHZzR7mYxs70J2xQm+2lID0tM+jyT+QS38pRvHVN
5c2iHe8doHu+eE8cC6m3G3b/xUO/SxTF9lHQSqgZpo8EPh/w2UlZiT4x94BghJ/ItDVOeeAcSMtu
ONNiShN36Q7ezkFdjs6ZzByP0LiaGvefdLUHn7JZHkHes7ygiwWjVUBvmUitZalBWyMZcJ7gptc9
xIJ3RY7d+iV7FLtaUPw9bBd/p1iVtq4DNeSX/eVK0aG4ETVIwWkIW6O1s9yeNKJK/7nYgVZHRF7a
6N8QCTPUa8DcayYOSsPpBIegMzupM4mThjZfQWfvQDsuN4ngE73NuRktudUEdRRTq/QVsCYxS+I3
KdmETkWztrxQWcRNS07q7/VVVYsidutP+OCbEEaR2n28zpEOMQTTgg+N/9VT4nszf/24iB8woRgx
/ueVAwRYTazbUjyh3936GSE6MIHTgcNZp+2TZgIsMMHulFOjw9E+kllBrhlbpolsR94EIf6LIPhe
Rkz/AR+1nm9z+pSYCJjEwYu6uAFAW2hsO45TFJCXB5+t7MJaqwu9HDCrcNz1kTxM/+ezbMayvO9H
rcIRGfh7uo1wApoLZRjv1vDbuW6hjhOaHByzAUcNvu5H6Cv4j1YMSbHyFkjYzC6VL6wc5A1rMh/r
u067MLHRSDXS4uMg2S6n+N0lOq3Mxau35bXfnmgojrafD9Wd7v4ST8/mLUzZIQ2jAdYMajyzgXoN
TbibYO/bAHjq34+gIU+5PNRVJXZNLtQoSY9VU8mtVdC9j0Nosbhm3hrLH8e6CbEr5tiV/PCJ/KDv
MTQVxyTZV+98mR1NROIrIk+L0s+ZGBTUNi3Utsq5fqDbS4w0t77gXhdYm+nOn+5GtU+nOVl1uMnc
Rfvn1O+lsicA+TI980JISUdCr3m0yD7k65LZ3em9w4UrNWREEYR8Wf22dMsUVVvP7d7Z+c7AMkRr
x9oMEnrL9oxKY7/L3Uln0Y+FbKyeLfVDDhtMUqvvZHd0rGHEnjrk5TREKFCuT4sRcQ3cfXXC/Uq1
o8Hos+sTePx0P/c5gWunN+XYXrXGZJhH119cN43yQ6GBuqiWU5sU+tws2wlEn2jpatvHKLTv+MdF
wIqXCYeE9I+Gg5oxwDkhz3BJxJZ8vufu3fb/x2K4dpLciTfMORM5P03x/vUCgcppKFJOLYdiks/h
PSyNkle1xn4LcgB2YOgjq3OhP8mpIgkCjiVtMSE7pZJU0cyx2Z8xRAaX6roBRcBLzNv6G3BhCe7w
fDjDq5mlGMBkq35iqJwEdPn6MXsDWkwgQpFKNyVNCFd+MmNFbkP8yYR902TDftR+QZf5XIFNQ70m
7zX/6UUFo0z3goLK67KELNsz3EZUBDsmY9oM8/5GYmDSTjMZ91qod2mKxae7OSFdhreWi28d5YS3
zIJkJfdsAadcdVyVIiw+WaYYpbESd/z4AyIqZB9PJ8Ur5n8i0ImKJNENbngpl3NpEHFR0dME4J72
sXy2AQP6npfxDwrr9Dl/YYxhJNwUqE+TJZG+/Tt5KQ5//swyYo6zqk53qTDcaiSw5APw8MLQoQ8q
QBDLa013rOM1qKKDJfAg2isquDjdppiOD0XH9NrrKpoI5f4pzBBq/oF2qB0D56Cc5XSmkxJq51n6
NClw2LvcKUHxDRdm61UaVRG4kL6RNUluJkx2v4i8K9fjFmgJ4QFkO8CTz2y2C0IBx/GDFNzx9M9D
Q4YAdxIkN/96/nXma5erwHV4wDw6dVKuiYSynSlN6VLMMAJobm1AkB9NlUxTz5mQCS9ooxCPKcaW
fnfFQ7oBXi6tfaCmJjh9EcwNscbsCrCxT2osm+0ZCGx3WoO4xVqcuRv3Xh0oy5uNuZcnkegKT/lN
fKLFBgfrEhkrqfd1e7K9bjRgtNS5a0aJF8E2Bo13OBHOfX3uMLQBRA3oTKSzF1rtgHmtQ0Ml19iT
xIi1KdrhqRl+iMp+N9dOlywFMghd/f5UOZYZQPwuh2qpP9spT8Sq8GsKS7Adey5VCGJip3qfRwTw
kL+yldaecpNIwd9Daqm1uNkqTOFbQyAWTyH4KBJi26UlMndXv2ka927oD6EYlzmIQwQ6106SLIuh
agH5l+v5kc4f6XVwzi0T3TVaTQyreIgqjLYp01mbdj2VyGQ4fn6EmrPUjnhazvHBVBbSYfAaO52A
DuZ25DP8oPV97VdOYXu0BfahPMs4qHMoFmwmfgQmkAupnHWVbtgabotMgAvSrB0ArzcjUT/7Bgeq
6MOHYnJHbSwCAuHPdYBr2DwO8pLpOiuKc2DmTPtTelrsjGUx3XNbOrn7zFYUGDs3kThfTdD3jDRp
7t75kVt+25RYLzuBeOJEwgYa4eTuBfn1Ucdr38E/Ae0/m1FjpWFkx27Y92joW6MRksklogf3VOHS
JQg7gJeAat6rSJC8Lb9w+7WQ3ii8tWdq8hVibkR/hJ1qlluN3+qv/eMNFbo11PzHG+tFUFJaWpXk
yc7e88exrWZljiD6QSP5cW/dAuQiOlY9DYcPHRrbGD9WLf07MkU6zKcVovZ+FOP7LUrOnxIff4+s
TJ/dj9p6IGjYRnf7d6ZBRwYF/c4nLZMWU3T4Dirt17p19Y5+J7oW9KliAmWKXuMD0UggqkLfvkXC
4MbXnBSUJ4T1/zYH7sPajzXEcM8bM5VusQxEEWioCOLr7l2pQ3AIhgLNizW4kj62UaO7+fv8cQ/F
mjtyfiUCxEQQe3QanlkWBfRezGLhqO9dyOGHXaL+Cu8TgwJ4/D7KbSWVgxHq/ZcSEtG3bpyMpOFO
2ebwq9lz8FyHxM2supkolx7Vrn3Rwr+LOQ5iD2luwmxF4Tea/7PytlCb8w90U7YUQN9dubgbCZf1
Bab231TPl2xdDkMOzAyU8iRdkGsQEus3hlB336Z8Zo3DjZxY1gyTpeEZM8JDb1k2sNWwfkkQXPe/
LxEPobyltOwN22L61LkA/F1Qk+zZ+hswHbZ1dNUBci3Tn1abKyv5dcoqBnc8Z5347K4/1nCxXJ2F
pYvQ3B0QqD9FRnVQrheS+oh97Av95YhrTbf/sr+9bI7OvhK8ceHR4kG1xrceOYHCQIYpWB/3kw8c
8uQA76WJ1Q1fmiSHUHbhLDd6uyVLR1JOE2ukwU42GgCccMxBsS5nzprIHPJENb08JCCqDWQDDmaj
Ka0cdmbf0YbzUqOAihxlKAZyMh0Xbov/BBWSU87LTISJzvL8qYzu3TURKMw2A3rH/P5fKksP7kau
vkxG1fgN/6vhIqhIJBZuity00o4ovRWE6beIEChxgnDpnfFnhv8vXh+Sw7IICSAXAPNDgxukvupH
HIjHhZvjnlj+vjTlWBm0BwKuWU+5N5XiCFkgVxakvocBfPbUOrgdfHUsPf+DKfUh5VopDTpZ/u96
hDSOJOMKZenXnBZf5hZBWkgqUehooYbpWBtJ5cYMxCk09YWykM722DIXQiQXeCANpSMKhXx4qxSw
B3vgeNw+jVO1wt9v5zsczY7CjdhteA35OANglPrNeovbrlDxH8JBc27ubpR/IO0OoyjTuo/1+WPi
YiXziCcH9tjwoFB7ZvG5EDZ7I0g6sQgm6F6N+hc1mRULGIbVZ0t6Z/8qZgJmotwOomFqEs+NPqj8
CsPgNhZrPWe7NXD8UdwSlYjNw9GSLxy4Ih/N3mcBIkFClOv/yPlsvytXkbOvdgRMy5tSmZHYFI3A
oZc19snSH9+q/ptGIhY1n89f5SVeGpYa0Zz/YO31XCHBTh4v9uLl0lTj/TqvhVejR8lOhyth7Yo4
h9hgzMYtsZTo8VyuZXifNxetLm/xW5kfxAy6CoCm/3FOuAXlKFts9RLCg+vXplTbt7UNFXCEgIW5
MGEb+QmRTcXB+ryXbHLmKVAwgkhXKM+ZZSgZJRCr+Yiyu+pfIKFm7ysukOMWwJCXcLU3C93ZQhDf
Nz5je9nkVWTtHAvm40s27bEfm6dJRkiHQRIb/3px0/ZDnjbcDwtF0wTSZoYz0vF5MLqjPEhlxm/E
6o5+pGxv+Bx1+UCYYCqyCDxmD56Wgjd7CH1Xl2AZqEOhg/4rcOPYf/JePgRc5qivkacMZqtN+v+t
ul2xjCBHnLdVEmGrA0DYpJ1iwF/Z0cOiJdIdNghh4BOMGjqJF2EIrtG5FCL5g/XCx0mNgfoktCVm
XVonfOxjmhkqqqladnAIqTKV9KLbB/G2Zne9BKTAUPpu1F4PUwQLIPOxjy5F4qAy22yYSwjY4Mww
jKpoW/nK4BYgneIU641y5yKQ7rpkV1W4IzAPIkbNbe1ckScBXRrQMUXjb4RKZlzU6CF8V4BJP9CS
QA3MwXAlXcDxT9DsY8j43LstFGosKAWfjSS3dlVA8nVFzkF2rgJq+05ROPbiN6tqFNPrFKGGAkP0
WQB4l4wxXSNrAm553WotUPW0AHofEEt03vEv0mC0tndKPPX7AhSK1wBgorFQBl4sdJXIuaBth1fR
jrkelt1uGjbNvtOH40vA6IG05p4enqu7Oerj+JbfRpvQDthrBGI5nt5PVnQ4U7gr8wLO7sxs8KNB
+vn7YRd6aJ3aahFpb6zJh7CXeVTPSvPvtDs+XiCTWzOW7nsF1COkIsqcpvO69mt8VgEw7OmdFXdP
t+jCY2mP89QoYxQvs6ud6LPbjSjJGazNM0+LQgACzNdi5p20UKEkM157C29r2NRIpcHP79rUDNq3
DGOMXL/xYPRo0zoLpusUu0m7hY9RqVwLlMhEIkhAr0rUmquKz5KB821tLW/0RGr9SPcb1Lb24Ojp
BRqrE+uMDMS5WZD8c7KEmM6xVfpu4ILHlB2sQAhqL0ZqX35ModJvRXofRCvalGs/xfpoKljHXHdu
MdxCgM3DNURLKd1VOUUjQ5K+ouOvP45L/xYA4RmuTy1Zx+D7X6UdAdeHb6z3+nGAWs1j7+2kdt4u
nCR7ApRL8JGtoFgfus1uIjeKXImLDlcFUt5aXqjHAYalPBMwlt8MIIoWA2sND5jbaCkPyCTaDo4K
vcFDWf75CtaLJ8qyugdpy+tQrELMavtTG2ZxigF2yUtJFg98aOSVblR0stOBIfkEjr3/YvFFsUhz
7opInyrnjoxA5+jg3/fbcUkeVONHg768nIPna5t6RDNOipt00aNphx1veUsNFOB6atq51aW8eE+0
MAUIipir9wSqNVlPblaplSCbdlCxnYmMHkKRe1hRiBo3guJd8jEJSxh/AgxLGu8UHLyjXSmNP5ts
qIh/q9ljt3jp0nFf3t3+GCY+uN4KF49dEv+rTDi0AWYbq/OKylM9uSuwt2bSCgXo7R8anOVNgVLN
qBHRK8d5Z87yQF/+xcKVPOmTZ87PL9UyZzH1Z/wpcDB+K5ccAoDgLEYB4oDp4KpqtK2shRf9ecrv
ZTjgWLxlNMvB9h/xuWelpFIQeoYvrKNIqasn/v/q8EHis9db0Ig0aE5dwp0Wp2Z6LKM9DJG48LRj
xHyqRoLFYE4Ee+ckoZZzn/qnyGlb/EoI+fpBOZJVpNUzPQ1dG1XQ2EfFb/MMcQrOtAUd0Ruawi6u
9DZM2GE2UrzMNj9Qqj6RDgE/amvb70/Gle/drVh1NTdTlGk6uP5/NiImbkCCb8PLtEc/kvoMVDcY
t/IkjW7wrayj3I0T+YYmQXAE3AnnQ53cz6zjfuf//sOJtoSKT3Cl2HyRQgkeY94WmAawAhqYkiup
tLGZOXEVA7lFzpKlQOFdJ0r2Qa1Fxc3dFSOFSO/VhWbqXlAR7aKp7fjSc8DMuOYySmZpeRp3Dt2g
PNPYfXjdkkiCFyEZsgCJ15UR/28ovzwLLJTDQ/9vJ9FH1xseDzeHE+EWYE0NovsW9hKHGGfsqbvr
eh/tK9gxx8liPGUUJ3ADd4u7MJQU8rPM5eT0ECrxReU3OLM2YQipvLy0zYyF2+nSNIwu0/kEV6i8
LDS9hI/pBBrdYi4sX6mMbDLCEGym+CbrlqJbKg27xb2hOj6VFPqJVCQV7eNXEpglBadQW0IeW9D5
9n3yJgp2KvyTcrMTmwJNaMo95Nw6wJEmxlViCkG7iThP9t5Pg50tKT8pBjRbaeRZHKiAXJGePLLr
epyTrLwv9LHemmHTyp0dnGf80G3Qu608cZ2jEOIK08VYidLllEa3Jgny5OUQ8puj+TW5pveqFJKn
BFfOI2SfqJXBaxxeM4X/22ab/ozl9WDATCuNWXPzekClqOlXZmV4OwPEHzwSpYUkjBb1aryP+DoX
JcBDwAoApZOzFPJx6OVcfH/sKZE6EyXZh/gTcMJOwSZ6aovFapZ1SSqgvWCdx9gSfBOFAR2cwYAE
bvqwhvsGGzM7q9n+69T2ji4PvkjkrvgaK6zUbQdE2Sm4acFiGLQLRjKUYb95pwjeDyfj0Ni+H5gR
rKv1/LYjzjxvHINbcPf/CfezKglC9CHkPugBK0L1O2XFyIDT7e8peTJVnfKQIRugairqOkNvSeWY
2BAx7JmSZMczulJDsn/Lu1GYielVp/pvJwh57wafrf7xTgfx24eHxCUWo9X5roc/YOg2ysRV5Ji2
XrOQ2oPmSxqGDLQ8LhMgw3hpz8fK2au/3ksWJUM1pQWjJYSG62Doi8ET5iQYJ9BUG2CTFBxXHx3S
MmPCcdDk5azVYuhAT+TypCzTV4+JWV3BC5VTZ8CZHOBG051+W3j1r3QbhyyYj5Zeq6WE3p4qFbhQ
7cglZJV3yHxUa+tv6WG3WD/8xbQJ2yAAtUcpSevNIgTikv8LYms1EZ1J0G1kdsjQgjQeXoo6186O
o7VqrgOLqAhW/tneoKoGBlvc8Qcby4awmRQBx9jvAy40ChlInFQua/Vt55dZbIf0MJ87wAaiaTGP
uUPgL4B5H3qtw4hNLIqtjg/ZSoMJlcyfi6nJs91UaICJ6KkRDFP+ykfGjJWNB1jaAeU1/p/QHRyx
nElXMr3MpwtCeVsfFCUYcjKOO0BHbWMFjiOr4u7wGA/2hiEckzNAHTRFW9/gXs9LMvm8E5e0T1sr
MPV9FvkTRVSe3a1WRa8Z7Z+MdU3Xd4EytknWxYokuPFWOZKLx2zDEU4gqA0QGxT1w689+MDKiSqk
TsTFb2dcGt6z5CChJK8jqPYZdWp46D3WvDi9ZtUDu/ANz8p8z0Z+ReT+L40zf/js1yNwQa/ngrLs
QMJkpZf9/BnKzDUUDRPM4nvKubMWI+yFc1MV8NqF4e4brTr/N7iN8cIIfPWyxO/pRfTMudHRq+XD
v8thXAJYTykJQlgVHJMLJVpD+lI0U1qw5zjul8Yga73EkbR5lZaHpYVt47hDSI1zdldshArDrmHK
DeM5z7SU9drHcVEEtl4rqvbWLO9JKzIzsgSLfiKtPvbjf1k9yn1E8Lfl5524J3Iq+A8+cX13LimV
0zEBbMjr5DNEv6E0a+E1tPP1HEpaeTXCx+9s9lIS3uHZmVXzEDzN2XQM9DbgII3S5+qb6bNzzqbS
PsSbQJEOWDMAA5KvPFtWbwJOMPIhCbw7ZWHnOAuL6ymrjVb06zv69xHA7emDjZL76g2hdh4ohCzV
zC7e+sFNIDXbRnavqXRTWNiZ6xwrIcNyoKE1pWVW1FwlRzYMQTmDsQIdsK64CHjpqJetnglj/vt4
y4efT8AEZXneO1hFI1696l9Dqu47QVIEkvT4ihhtBvNi6B1eRa34ZUOB4Vw5qxSeSpn3XW+Y6kcn
WNOo8GiOvRoFiVHEjkLa69dxKjqxr6R3w33BuxOiuB+Poe+ihYLyYwONSm0lBHBAQH6PzwAN6Sdw
I5tlshw1EFpBQWa6PQWWOS2mBhCpGkK97WcQ7v4u04MjE5RVpD9EtZhDRe3f2SWuctOiw31smClm
wd+RkGxDCSiX7fI82qf0uHQx0q0oHtWtfD55LuGfSujgENXu/9fuqXm9x2HFj0+2aa63LrTyG5hN
uQc0vDOq/A2q0fus4hWIoYh7h8JAeFMcAVAxt9jzJ3rwz+YPH4gl+ujCszt2pNSwAaPObs//0Cd1
mGyJbZJKl0QygxbatbN0YhHwlATCyYJR8GirRe6dDY/waX+6fALhRGkcXIDdHp8WesKJPQTJJYZH
pVb0RfSoB7nBUTOywocrwkvabaDJlfus81IPW0Hn4TPE9QqsfqsWBS3DongTaDjevHmx40S6KOS9
cf64yG5afhonQU1CgwX31v4N6W/xMTrxak4LA+aEa8VTQ/BbS+pSXPbXf1MUdHXR9Fl2u8j/G9pk
i93uFzwp2mRyXUmB/9jrGv/7iLX8BwL/WfrUIpsaijKIDJTrGBU3FnBTOMvo9iNqj8Uh6PYIKvOD
CuYNJsJlZ0aniGSGnfV+l5rsT0ax3e1bedwwdB25a3ycKYzyywsZFec6TsbP2359yOGk5v83WhMo
c42bDtzA177WM0UPBgSxdaSRY3hefwqBKcFCK2rpEULzZ33T7h8Mfr2XpDy3SY49lulikn48UbME
Bp+7y8z6qSWT/vCCwJma3+eaZTbdI15I8Z9WHHBZWB165s91e55VP/6ZI1IWLt/fg/MO42yr2bQI
JTtJF1IvwGPcC0d5jDomYihnPjKM3+c9gZCuA9Aik97Hbj9lALuvJ+N+TS14//46+QVWtyIK/pBp
7eduX7+sLIG64KKTY315vpaBkGf8BSLFcbhDBoE6/l9kqsXr42+u9migo0lUQJguUHRBgFf6WUPr
izGM02tAhHi/wQ1C++70+SHOdfAOGrHxvhmzgshpTRcnQyeDaYtOXgW9tYj0R+9ow3qV2BcB9sUq
ZnnLXGsc0ohwEQ5VfJmYArdHAzowId4UZZrvSbLKg2rGHV/VeRPeTC/KfXOOQCJC/rj63Hx0DNzl
8EGSNbG/8VtrN0GhgcSNLhUa87PAs4X/VcdpheLz/wRq01Q9lb10+wI+rxdtRnA9YsqkqzcsnYT+
1rQzFqUMY3RTFg90yVRgN6wCthHWpZz2gP/Ck/OL2x/EptcZ3nIW4TCnRvB8xTbAE5FLRFNIyakk
uWpJDnYfR5mOb/qeDzs9VmlYd1YPfVjsUBrrBoUcHpuof4O1/9dLZeF8yNueYPnaBVqj6dhcwpoP
UDsV+Xu3lXwB0PrgphBVUitzvCY3TrvBrDS/0PN1QVRsHLfumfZAhjjs+IL5+yK1fmM1Um7Sac9T
wMgWnOW0HZ8ZC12C5BiLKJ50CYfN1gzYyZKr3Q0+VAIJxYk/hvgNYXphiETIwdYnYtbjgMGGyuY1
a+1fllGgrJgjCkgolllE7TVI3p/Tt0YFDhx0tkV8LVk8FouKtrOXS6bqELayDMnirddO39c+bWZq
DQ5sCFJXcsQ21rQzPwEcP9fI8uzlDvKAcbqLLU7ZxQn9JMz/cKJMMvzF0P0S2001WhE+PAi6T/LD
D7GgTSrG8WUgpnK3YoWlPkMLt/c8rBMz9D3kXiD4dQz5YnMVzRh3oN1yJwT7Qs9ZILS5HtWqoCbW
3yY+WnP5v4ubzmftU/FwQDMN/8XJ4RUQ0ZmA3feh5kdFT05rHwsZB8Sk7ztkjYMqNRWdjtK+7U6B
JterRSxNCNyRItnrBb0sSFktTSZ2X0Nw+B8ScHtdztjlSfr/oGkKcfJB2p92YYgKoe2CzfcKos1e
6jj8/hQ5jqoTWrUQcMoqjg9k1+X+Mqzxavtqom2DmGCymakYTC7ymQo/vNLdkHAskH3GxQSP/Shs
4cm1mwzVGiEzvAgGmu+JhoKm/WANZLY7cIdvbFUzKcjLxD+8a7eqhrwh2TnRRHYUuyq3si64KosC
a13qj5OXvmQbhu0vzUz7q8hzoubbYNgEc8mM1/2PyNWLaWiDw/3OGiCSyNZtqTWMXOB9kHcPrqzx
B+w3mzBeDXR0JEhzmzIQeS3LG+xL++sYm00oDoMOBVBxSGF0yaeYiR4Y7RWtdrVvdtobOQ8Tta7/
4dl+1x9GyoQCDXfK5f+iU9ZzrIou77FgNkO54zPXKJvWQ2BA0o8TXfKqw+Pz+E/xBRabuUrg9/nR
kUvF/tJgAVaJhEqxyMyJVHmzppHhSw0Tv3NlrVdJiZ0NeNBwP8gkOJSGe2K7kGJ/ETZJW4z3pfl+
HvkQ7AamBBuu7Dr3zs47FObIeRE+TUlwcqqxt0slSbk7dPusE2qo6VAkbqCeiAwdRGyMkfbk7CkV
zCpePGcYVG7puZHEmmtvhcIjflrbRWUkArEdO7UWQ5og3esWRD56qg3K32UpFe8NPhKIsNZK5Cs2
hJdwb0dB8BRSQenhWFtDdNhUL3tobiq+MapY6fX7Jm18VQisIso7nBYl+mNVgEvY/k5IoCvKNXSY
Al8pz3jQl/qLB5kDICFP7e3oCHasPNTNbvLmNhFsdv7XnY5b8KALvEwXZeY6rHZhTNe14ngL/FJC
UkEDXk4vUZNFWFQkTFqm8+x72+OXkK9zvxuEZfMshSI1b1/BBtw79OuDoyVQOxOQKWN5+MJNBPr/
kfceuArFjIIQxEkfMA56eu8f6J+gkz72s6q8OBRYO3n3ikSSUzDxOarH8OmpXrkI7rPMHOECmllr
oWP25TMlvyJ68HSAOfRYKJB/qmYu9p7PEZ31uU59K4Xb1olscPDz4yU7Me3Ce70vWLNZzM9UPmcH
F1hFwWAju5T1VJcgFXdj6BhkVl20T8iXA/cvWWQeMC6ZkHAPpfmihOCt3nPAZfRa/WC01zQzcq9D
28o4LM61VKcvi38/sUMOlHuLOdyQ0YB4twNSYGL9X6shy0nYbqjW+q0IVH7cl1EfrydEcFYsbXY/
I8CMtItZhMO7M1KPvgZQiFJYDuIAv+urQEizi9L6WCMqgJKXPvbzlZsGBpHkrgboPMZh1mRTV8r1
neymnN8qhwlq96K9do2LvocogdduBoTOyDQoD8Sor1um20KENf33pk0TB7nbwIX6jenqRzzqwhnf
R35ezr2mhyE4bpyTa6KBy0KC6up1KTg8IyTKAx1R2q/+LkbJ4Zwjqau4dcUojxVb8iMePwyMvMC5
aj/h/geP36kqAWaFVtI+ZLMW62zbbm1G5N6jyoQLAh9FubqnOl81UpX7hS7ZMGKS4r6WUGQ9es1b
UR9dSeC7Sb3shXXLS2eBvgbHrEFumiD/c3FJKwPvJy5F7dfTYh/9dxsgQjYBeIW3L7xrYCnyStpX
wYXfro3JyAak9+y6oVv4V18ELDa0xSxpyyYyTNf4joIkkX7NPSYS3H+5imywQI5sCJvAJWAiLGPR
qPoqr1CVQmb/HpYKctrJEb/SFiq0nH66l8+IFcUowrhmkrYXpbKXwBWr9HukypDaxu/wXpsLQ3ew
5VE+l1cEbV74p673stMSX0zzEF9lDeUgrIJFGcD9UkbSWuDtSEaMZTikER1LBeLREgFB18sNMl/A
lNoABqVVOB1xN7iTXxSIbxaHaNIjCr77Sh0jpWZW+40+0orcpjT006jFPw1vPgY+cELXP7WWOGZE
Kr8DC33SdSALfme/U4M9NJP97I3hJ4r8QAKIrmbskLNiQ5BWzrTELHu3/IxwP1d1F1THDo/AWY8X
9mRDoBaYBekZ0+u2HnQRcbUv9t9hfuHDbIU2ckdG9K61+HNg2BpUPH5GLUlsue7M0RX1Y0spG7j7
8MT+pZgVPT6jJ3Ex4J1lmdXeV3hN/pYs5ldKqsHaYvGCQk8aqy0ucygNH91VmBiRIeUJ/0aIEJmE
albNVnvqyezUrJUTuCdTrj76WhpQPdmuw4kmjTCbY9wgiNm3oMtCB5VxyQpNrLY1iVk/V947B15h
CC3UQO6wYaMkqDSATrA+em9eMHKnTvdlZzkS1MgJxed1B9uOi/aN28EjRybQglsxzIM6Hdtuai/B
K2+9HdAUyM+1dIFH1Jnl10qCGKXdFiul8khoMw1OMjLnF60piZF6Cdo7dtxG12p1u9BVIZDPI36m
h1CB1GB1QiJgzni9dTbIaVpP70lETtBMP5lPo+5J/DUjSjYlp7GCGAh3XCbHujEhLmc8RrjZNTM2
FWdjKsnBzJitj1CyBu/0vt1ob6rT1wVIBCOQqX0iBUzDv5hiNvnTnfKOxreKFInq1gF0x1F6cFv6
5hmZl5I2n6usdYLEqeBBnC6THvzwYVkvx/RpwYFzVt3OzwBGxDj1WPKGmq4PCE4iTplRLRRn6XgR
WRCqEOMOCNmikel2XeybKNOwv5PvObLYsQuWuY64hEMoN3cFosFDk7N5QLUJxpS+XV2WWjUOsBKN
k2mwCZndeqHQUVCTy6TCxYs9wmh9HzVfz/cqYvDMra/xKJw8rxdhWnjwbsfnEJtCOC3LIV5CBhU5
TubTrXQQ2nkj4SGjZ1GKN7SABMg0y9QpYn+/LPtxDO+HMNoqWUJwZITaKNl9C9rpITQX5rvJC3Mf
wmIrFrgAv9PwKYP2Ytl4pK3Asu2eJ/wWqlgMdRzbwaGqb09lwNwfSqjxVFLtqnhkRGnqtCAmdc3F
2s2Q/QFHMi0OwiqiXKIjZ1rkiPmjDjSyun/qXHNu1ftDgMALmtp3pzu0Lw1VOEz3Bhldb4jkKnZd
7q366k53I7DXw9VCb3119we3ybZTwapWyJtqYrXH8JmfFKrzJsBZexfVS0lVEny2h948B0npdbMN
HKnvezuSqTla43S7HdSuSehWZFfvXIRth/Ny6FanSPSH70WIH2XJlHi2TAJwVVb4QUBh8opfi8g3
UiB+VpUeNyjKM8Vc1ssWaRRqywF872IzOXN8EBus8HqM4dgRbiYL+ujMtpzrKyRuDRmQCiqhTeOK
E3ZRn3HPGRuX7i1V0vYiDj53K7hbgS6iCKDdR24EPf+1f1SI+e1QkxYmSsk0KBfMtPZtL71ZWEmi
e15J1zQL+yS+1bWy4KboeM7X1Om/bitFl04Ub89c9+CtnlCW+O6rL1mu8lG0jF4vvv6VyjTB1QW0
+kDE6eXDLyuzWY81E+gExsIf9yw0b3Gl0AJLn3rSxdpC7D3yl9nX39XuoifjARFoy5/yVQolGda7
zxpTEGJyMHDcmo+zpHobYEHVUn0u0HOtLnKtXTS4L81V1BHK7ZxyZv65BjAzu+YJRSyKKQ20Sr6n
zfBLiyZ3RML3+9X4GxTSSLT3QeOqgGvg+upyOFKzg13tFR+jJpxlQSQmme5Pk68AsjJ6Vvu1fg22
AEEpumGt+1hsYBERmOsflw92mtkoMx48/EOjqkQxefQEYutytiNuEZ/w7qKSLbK3KrYtjzSIEAPt
MoiMrfuu/5YXKzfTbdMaisDTTJ9KXIHtGEEn4MSz8jXJFVVuQR2PWp7NXM8cUctfTFRVJ6J07ZIV
PFOGPmXyB52kZFRcJC7wSmFT/9BpBOaz62AyhZwyjWj19irXBQ9J3jD6bgRjmUPc5ymBtc43Af+e
p7WGWg/V2Xm2asLIwFdHVNoMElqsZUbCw2FRl/iXjBtSKce9ovObGxyV/DzUxUWg2tv6aa2lhq1Y
YHE1bRBH4Mtn/41lt48ra3GutAWeZ0rrT/5lBrWosNiIBlbWlWblwbtrnGmGonXmzzqN9gKoMVke
+tMLpruGXUz8mq0ni4UgXIYLFtwxrcdQi59AA1f9JDwg/w+NHJ0qm8mvSYpNi3cKS+rCeXmaasLS
45Jeam08AHuUkGa3M+GSH6QkM7h0pg35OemiCc/BJyae9N9h3Hpqt2+hiwTXo7gs44Hn6mlX1kua
zuLBv5rc4FwRjEv0g+XUDtY3miZGqWJpAMgdODjgT7Uwage0h8ZnbRfmtuGLxJHh+U1KcWsbyFS5
PwfpSN7XZ6N0gOsf6A6P0L8DtaTqd9a9O/BkBe2H3Sh0CwzAbMtASv/jPAgkiAJVON52oMXlXRKU
aKNKFZ0dZcu2aWeu6Ep8nIS6pO/TASaHKoORMTfMkzPhcMta7r7Qg9zYZ5R6D5VXvqNMl4KY9/4s
xgaJXoxEiYn6K6wo1VxeIwyWel0fZ2vsKexAy4d2s1NcditkPLc5JZYV6q7+vGBOyYKWSxmzfY78
86CmkIHsjWXhUkfQVBstXcHe+2fHm/1U5COOUjvXipWXLsOyKmhkDxgjHeAhton7GhFu9yr5F2Qt
FUtKFU/CnQ2GAr+V+EyiJp5VwFzbK7qht/8GB+uRByK/tWSsbhTH1jG5c0qkJLXTyQT+Ra7rD6ng
PQBPEUYoGaeSRzkrpefeCFt7hURROfHTDsOiER+7qpNuqXuWcZjqIVqF74IMq7tNzoPMSEAb2d9a
lrw7N/ElPn/eKW1gXOfMRWbQ8sS3pywNujt/IxqocZQxMj3KTA4upTnyz66cSrcFXGgTrBuNiD84
kjlVcfh0u7yA/2MgvaiAZRP2WchawmmpK21EpO113IZ2p2jQLZ/s30u3U+mwhAl81blqADcLHjA8
vvrKkVX+lPcXGYvYbkJcMhBV+f3ETc/av7B2eM6Vp6/HhyZXkUKAEZMF9vmKrFvuW1F4p83TioE6
7TleAOpuM0rfWSmjxKD5p6CoORsYPl33GE8jlGkg1hqdgV4Bgvxds8hF7dj2EaDEkfNCKJbrlJp1
/TWRjoHBoLs3WFAGfBPf/vd1SOhHYvk1xFuaRODpwQuKPHjrDkk9zwXxOisptdsIXpISNLH7DDvJ
JqekT9uyufnUUKb9bkpqRpn+qtTf5hnO6MG1hlx1/eQjNaz2MJkLS34s1G5WvsMtQNlxRRiLNFGV
79Dx2K3LRlOcdkspbklt1BMCNETauf/yzJINFaGfoBb9WAAPXn6tdBeCKNm/U2o17RZl6mFKRvEw
zc56m52CB3oQ3+33TZOwBJyWO9jzgA3SI3vrGYH+xU1g1GuRNAyJMIPyKqZM5BmSURoHBzJhXaH0
8aLTjXn0sKpUBPk+MWH9MQeUxIm4NLY1fncmrj9eR0xhd0WEHqdBhzzD/f8sta7ub5qUuN4/Fdvl
IPEj6AZFW0IVtV5v8lvQTTTEL87xsvYUpnKRYPfUxIsiBY7akVdIbEdSGwTapDDZOKm+j9Uc6OYu
9eFcjJOx/9IeDt3JWZ3zLm+e9w8Vol3wIj8m6MEs8aX0ulquFJvpYstlbGhVb+n3dKW81zQ+XdMy
Vx0QQRbbTI7v46ofKdMiZFlJpO2LoZ5pES3Et5KBrl7QM6E1hEmXWoq4gJbKtuwIIGdekydFcCd5
tneF+I3a1yCr+mx0BCym3rM3fCSc4zFY78tRfS6tQdjVpKCDJ6KFYVmsD+H76TuGBZC6LmsG91sI
hzKueO43+h7G4N84JiRub88PUeP4xWQTtKhUxvTGQzqCpzjod1rWKE6yj+OgXuyK5TnDUlfJ6OsD
f1yIBnz/E7Eeca4HWCaraoKyLSbe0TTUah/iT2Ie0llQ/EmBLubfQfE/VLm/DgcZxGavnJdPg7R6
GD4J/kTChFJbCW1KV4i7/8/IReQiCSzcACs4nFa+edoZzhhC/s2ExcxOb8aVNMcDOhZ0+I4ju9uY
WXHZa7XDQoOJxL8CnIGcfIHmYO7ZU06IdQDaK4AfDKiWLj35wPThtX3CkqN+cAT0onllmj+HGKN2
u9FtlqDPz+SlyCBv81Z3q/In86T6qfZT8azyllzVtJJOe0mvxCqHCu4lQTLCBggNN5XlWWuj9C2C
/62iBsr9GOUykwWFt0DquK3FL/y5ARn3wTbdxujyUG/LlNHeVgSxXKvaJ+/rS5vuO79AFiip490X
T1bOnrWjcjYM1tGsHJrkJK9QWHl8W/K32fUlrNOjZJnIZk6cA0kT7VFznlTzf1TdP7zhwQ66WR20
qslcO3OQNtIBsypHW1iN3v9TtLXsaouV0LHwVMFVA6QA6tHsc/GhhhPclsyLvhk93nWsJWYJQw+T
IuF/0mTUYo/4jQDRlE8ej5LsftIK1uwZwKskcrP2PyGkLEmqryv3NVmgUNCHawqfWBPjdjaC/XIc
BHHkahZuxa7ZRAhqn9kTJY3rLivlR9FVv6ad/GCENqs5mUA7F1a6A6iYcXiNHVVf1TSwLPLLTx6o
jClwcry1UJ8EEGlXzynMsORikR/Y7XHyugZycWVaq0zkfDhYbV5VDS69VnvHgMO/PCwvhEScO9pd
TrPDNZBlggDBr0LRg3atoAxwPQMcu38XrLuW45i+l9WqC4DNbtk1x103zO+mHiWM8mx8ueVv6mEv
VQ7YYP/vRCZp7BBZ8c6KzpvJEmbCEWUIw3u4usMZOPwP68TLKXByNZZOjnmzJA1n7wImPegAxQXk
ScJBac+Lb5Y/7hmpU4XVZ7uKfG/hDlLGFezdiiV+vlHs0dwUlgxRLERH1C9gGJKrah3oqIN1qKaa
PIA06c+X1lfRn5huV6sOcv1Idc8lGMlxul1GgQu0N5JGuP7vdY3SM+T53B80a4x1gGJhfNefrQvf
9k6MSPtUttwoWsm4ZCjbIfom4pw/I81jTRReA8+rKiBFi7UavWgiJnljOAj9cz+W41NWEhBdZCnT
/zD67VtMosRJ6IAQrqJG93R0j3lWUe9sJXZ8nT7QzkOYYnB3eQk9GtHwLyNJy+cWJq8CVJfXxe73
6o2Jer9neX9DCIb3mDgUqP58kY1ZO2TejLlZRUpdviqWDP6dGXicm5HYdsYJG8FMXmst0iNto74o
KQi7euoczrMnsgE16PWYwQ+Rzg5UZGJTZkCbjHwiBHGKJQdUsOxKLSyKCnA3eY+oYOvg854KngZQ
aeM0PYafbeoRfNZTMRSYciUBG7M63biJtgWu+pthg2OfVDNwgtastiqeOEn8Go2pKeRuuCsiGMpa
vLxp4hZF3Qf7CawnpgAMZF5ionzr2+vX6r941rHNJcnm9ybFn0HC9SX6ue39oQHFOPj52cks4DZd
Uy4G9MvoIqx4L9sbXBbUdhhGODQwH1Bj2PFVphIJIIzGn8qHUv2Q2QEIjwDJ3DLN2oKAAoLn1pAV
HkujWSNj3Qf1+D//fiDeuLWVwgjo+HgHUJZCcqs7YvB4afwuVziJUCM4Jv2PLsQjAB3dALOQrYRR
/TLmEPMHPsMHyMeUR8Tn5gFuaSeRgr8k0XssKf4WbpDBU5MYqDZ/S4iTXjlgGzcBRwVDeMmZv8bx
yqwobXOk8vSGgzfg/uQrtBqICaZ0hDKGsIwyovhNUnRdE9ZuplQmJpHkmRnyM5LVV5pzqYNFTBl2
drCDI7v1SRt9eQ9yE/LwzUxjan389rAlsROm997HDgWfazeUtKAdGP4VCFLST312dtUnRbCFJB7g
c/TO3UBjrNdfHPwRmrjZ5JtzO+1nUzcc31xYhQTeXwhN8stuZltgO68XoZg35nIZnRiY7H3/8gmm
30pNLYiHbMupsOEKCzBt7DpdAji9YmaBObicXk3hscXUA4yeW4SrvQkrcqdVX27jAmwvSoOZeQBj
Kem4F7nRpGK+IuYKoBO4nNbXMT9X1aPnSNSWzUgWNXpRYia/laumT5NmnZELcENY6Dr3jaMbVi9I
LisYZZ4Q7gdayYFXdU7snulvaXcOo+7XcMtYWT7pzv7o8gr72uH2JVyql5HedNQ+9CV6LtHfRvqK
N5eEhn/LrRL7mZ8n578FCl+NEx7DnFL4yKpmIauBXcWzno03dCQvxlv1L4sNhiWuZP/1Q31F0g1A
W7yXs8wTeSVBoiA8Q0qzAD9ds7x/jR/+Rxl8+BIpT68vvFIRnZXdSyHXgBmp6CoYQoGCAodSbOmC
R00DDaNLwllVotXCnRhuOhQ9JKoX8Il/98auawLFCfS9vPlKlJtmGuk228HirOc/1rpDByiIiEIC
ZWj8tvpfNS7rVzNsVHJFNCZ7EsGD85zmZb1KVdb/qQYFU+u0uvxdu5dLkdlzId1mhB8Gf89cx8nC
L5kAz7AOekV0F4xb5DY9g/vapTooWZOX9Vsyko46PytN07+4v5+EnE/uhs1IF0g17SiFE//XIA3d
NphJBjLLnnBoRh7ru6xO9A0y2CncO04WumFcOIuy2ZRlAOKhFhideKgfyyVKQVahD5/ujaewHjzm
U9MJjReFP0Nm8UQb/gLQdvynONdCEEZiRkZbZhsWYVRsA76d534xoryI5ssSRa0wLm5TvelgbCTG
Xr8BQwos9G79Fh7HYP3rgffJRhkn2ozbkXPPBR5frVjpDzeFPNe13kBjsIIOcTEGXT7I0L25iegO
ZSypE6f9MSS3WYvFJjok57WEb+R13qhgQh7S5DWdIWu2zWBOCp9xGHunEEzIBX/qWKTXzHFEJq15
BTfTolC+vEN5dck/FStrjCuimczoZzQt7PCV7V7e8zkPxOtxblKB6mhw3Bq69cfAHMvfm8+DgsVx
dzOigNCSo0RqhRXyQl+N7m1c2radkOfEor4Nda+wwz3tm0qXD5Z8CUWXn0OtFenxz5Mxqrzj89cQ
kZ5aWGJdLdIS0pAs68osjujBhA6Ig4uRCroqTC5SI6UsarHHZUAwszxOsINlSLchI5NOo2z+FDiE
6a2z9AisMBunpOi0ettd/HfnmQQF+9NrwSdcfBBkRpz1qmNt2rSoJhshtClPiEet1AMUkeOVrQ2c
3reoyN+KE99tlKsqBqKw9xHi6mXxbhZPryHxheLMAUNZn5b9KRBCnDGWEsKK6Si7RFDCpZFkjnX1
yjZKis0aAFePc0LZDjsBh/Y+uIeu/69MYBDVzzZxjQWl8O6BgSe4GBzLF7WezQeeU1wtZMaVXV3M
DBxj0F7WUnyu0iq6I3dAx+VD/q/sDUvYLSm08kZRfJe5/01xa99QLxrMb7LAOK/Df0wuOC5Twi4m
cZfQIZ+rV70q1EfUUDMfhzq6/gcJpya2kvz+YfCZcQyBWNMf/AveMy3lkyc13mWJHSAXu+cosFGb
ClZB7cR5sHSqmn/eLG6W+oKQ6T43yKcd5270hxtSX8/Zy2d8DS8p+NLjqQn/jUopg0sxNSqvZHiN
thYuNg/ZGdscA64REAAoioxMQWRyOOhELIthzpacCiEh67pWX10GbpHdfpmq/M8vkdnMF2eQM8l2
1nPGybxMlaHqMPCT+t6jFllsGDddZMWFF5qlhwN/l7+ba5sN9idADMPeBXl+YH/3K6eF3VMhUJtY
TdqF/2fhx8J/AP2AQfglVdkiEUsgLXmAubmUSCk8iWhMADApNPuCukR7YeqlPMDRweeyPnqwH43Y
BODBPKwoSZFGE4QxHKJqwUWfH50bkhH6dJcBp3zxKkNzeKHodtMS3AXGCN3O6zBhppHLKX7pldjg
Fx9PpEe2Zu0BmKpmgQxCa+uSOn2J9CM5HNkZ7qFiQekOuP6q703/AVlK0ZE1X84KcYOLVOcQtZAk
J7QSQ6QyZj+zDQszeEtHrzsH18JvngleXiJE4kUmCrckSaiKv7eONthkYirrYnsz1V+0c+cxe5pA
kFfaLryTlEQ5AcefvU0+9AgBspsmZFQaABgv23KDQDgI0HZEYlOxyZF7eLe3lKSKe0a2QSyLPhjz
zUPHHHcUYJWYW0AXFkVbSg35D8AWmiFkNjQsFQY6w55ZEFndgmw6Cm1Cmktrx2ZQcGJr6rbDLnJI
HG2rvFnwIXyY83hFQBj3mzUpmQ55fkzTJXkjUOiyHBmYeYamVBJT5HezTEL72YUw03liZe4B0/9H
vFIQ9b7KnatrxnP2HA/I/gVBuT51VoWo0SmIMusdPUmMaq06wjkB2++IQXdZA/Jb+Qhtfmmk29hX
GjOHJPhtLI8tk5hjbuM/DMquTIZ11W9MSS7kB2syvJwttLaMi1sLQ8yiRvSI5kFAQ3w8AmegH/yW
x3VnNS5yLNdBv2qoWBcw9UMBCQyB6PwlXRlyKABX3S6aLT85wYrD4A2lVIyaEbbHtwTmv5J8qXaR
v2ZHJHAPCUWkmF9szn0X/VMh3QCdW4o97noYYZjn82A/XN7/DaaCq2DtYyzv82ECS2xf2dVOFgg4
aK9piyp0rncyqHOkPu4jIXPFSj6GDKtJo72QLZ2xaYutbJgdM+ok05Niv9vWey0W99coxZLEqWVv
jcYSZ5Lyw52cNAyCfH8y5cr9GLz60HtMI2M960dO2DB4xms9YPDlpMIrIWrjRD6b7o12lrxZT+7p
7R94AA7c3vHCFhvlVsN86XByiIs84kyZbtHVn+auVVTar9xVysG5lCE5A+zeKoAR13JHUfikP+ZW
kzrqgFEbAJHe5H02CMgffTHT3JmAfcjAjMM9atgiuFDbuIt1NW9uBccVinrzk82UkSmXVUPuTW11
WGyzdf6l7rdkzi3Ytmz4IsheaYfRkKEnVrndmO40tQke+AXq/OqdBVq9UoOY35ZZXWuz1Wdnli06
XiTG9LCjqdwQBZDFvELostO4Swbw1Oa9W+4MrKsMMMtEF5xCQ0NicS+XIvM9A3VfbKauOiSk7Dlz
It1iRuLSMsnj9gsximM0T2Z4qwJeQcTqwC0OiCtGLeU4lPJO3pbl6A2igL7xpBV/0GYPGSWUKA0G
Rjw2ZS96Ve+4nR9K/1PNjFXYzEFXxHlvdo7j45lPOwXMIum67z5M6U73Zy/6ObmkRFL0r/ka12WA
rhjiphHlMCBq36mJEFDbjR1edOWHNq+NInw1OqONmrp9w9b6Y4efDQ4pe0TnvTxmn6Cx2BpGdIps
ISO0ZsF2Hum3mDOT48tsUJq/U6j2B03FgP0PqTz8+BgK+V/qrG1lZT3c0mLzEK9MHuPp/zYfwJjY
AlWCOOkXM7GVeKX0cRw/mgP/BM+9X1Akknxrp+g8O2rBJO561wrmnZVE5e10AaTCZdIXPqhrGPSd
p759xsH4Srvfwb93o5derSLeilWt9al2gp1lDHA8e3j4Ur7sjU+YC2+sLl/v5/EGO5nGQ7KK67UR
qqDf7iwyaPDEK4UxmnouSDRg2OLMeG6fSxo0N+r9Ys5qesIvwV92cuNcbpS10zdHBaxUPypK/Blt
vjfUV/Lp6R+NhToYUgNywOsJi+lDGWX+Gllnbr0DwJUhv1zZo6rrNpgCqgSv5oCVoUf0/aw84VJ1
3uehA6VVkZVUEEJat2VRt1Vdg+vDHYDXcyVFmP/sxrF45P6uVmf9zhL/IrJU/TYmpF5knFWQ5z3+
h7xb9mSGyQPX7OAriksUhMab5VZQu6G9Z/U0yFnPhiJCYr2BSj0uFIEpTM9kHzSbyTPlKdclPwEc
Beq6KT/R2+ZTHJ83wic3B3/NFDJjBbFArYpQ7qIz6Ghta6zKoraUgNMkYwkKb8NjGbKWBKFWSD6J
Kk8sesEoFg45+P5cjswNQcLI616LZUxyTizCKt189zOdv9x0LuaM0eAgPcmEhGc4gDznIz4co8/4
uBKelhFiEp1TgdW5d8klIdNjIi1vvZuQDY1BH4PPWArLoehPpHKHxbfnpSav6UTDC9w0y/2elYJw
AQ3e3OOZVH20pdm+SNMPYuThxUa5VmSqKK5+QhemMIwTHPfSw8hIFcd9ioEU1GJNbGuF4ynepwJX
FTGkhlN993Ehp4pt3eMgvCUiSXq+v8iYlOJrVNVGfoD5G5pTR/S/vqdYbXTrlbiVSxpy9n0j/t+V
gJXFNm5LUb4NfVYHMxwsVqs0QNEShDa21NkjYz4TbsLlB8Fbe4q2cltVzU7hG0TrPdTGHbjnt+Xf
EJbFYkR1HGx0Q8U9orhGntikktZOYr7qlRm5KGWH7/E6tyl1dnLbiHXIHyQYkJIOHUBK9+lm0OJt
nfGcI1POGvFHim2Kdrd5elnLsPVLJPCo0vvDugIRJSePLGIVoNZFVHVwZ0EKtq4ydFj62FScMCW2
zZWBKi+mwqB0+KFxjp/opjpas7iVtxSg8/+mCakAKUfJNxdv2b+GDKMvA6/JhakUUeA7dFHYgxQZ
U5KRn6UKj8LkIrgE/dTSXk0HyCU4Tm69gtKKCbF51bNNhmPyKPDj4nLrdQoLU1Blm34JYjMpUAEE
Lld7wyx6fKFDSBhb7Z7TVzCXXOTZwY1LCLUnZBgSDjC45alPBh0gSHg35fouEJpGshl1g5DLs03Z
PRmmGlHaLWPA4cnGTKuluPJKbIT3XPgxjUGKVS0ag/ovVHcjDj4kn1cfSqs3S2nT0GCuy/hyzXZt
cjl3TKmG2Hnpk5efia1hcuFwBNeycV3I4+JHa755CuRoMr1dkJIl5xHjVd0U4FxhIuv0EAea0VZK
FPTIPMWY5UEP9ES+QWEGA48Y1K3z691mP2tVsRtPJ+IDlOIga/dLDJSd1dDJPuRfYEMOTkjku+6S
vtSzX4UTPNkgpEDyykV1PF+p7dNTprd1mxQ7QoEmReEi+z8u684MGIDu1PxOKr2AVOFTeutIoqMV
4cA/D5yKiutR13g3CUMw5lcs+dostIB0gcemnwIEQfGWM5GxuXLdaJcabuBfOaaoSRmMWYbiXk4u
acaNkB+AOj1LBpxuH11ccJ5j36jtBqvCm1L4UoxTL/jfU2aZXp4XAcJebn3bN1OwIFAyjwEF65n3
BCXrtr7L82EbkQeYnJX7Q1Jfwj45alq/YopepGpzvRqnKu9hyo8XOvqkb1SOxhG4aX2nPwuqZxM7
UKaoJyrdk/ZUurQ+WvYyAiQRp0ePQHFRcdoh/UZIf9pxTMIWQOueHur65oliXDqqBrD2CJtzKazA
WbZcQ3HHpg/iJd4wITmXkjcweGyFHK59XSyKez6BL80Z5hisHKXvAQ3WsFc0mwB6ug4RHgLXEOzM
Rv+ARy5cFEYJdsy1R4gUdCYvuHhSLlM6IXMSVg40HVwbfQVGzQmh4VeOoVcNYuKvhrdN0+1rmylL
7OFLyarVDvZYBH8/k80epRntfrlbmxFys++xxCrA2genfFpAS2Z0Y23CV5VNs0+6+5+hkVAaCWaq
ocEVhEcH/LiSQ6/i2LnizaOl3W6Z1+Q2vYNpHLV5iSzsqb3l5lkD5mBmTwfgLOi5u3yqQAvAqvMp
ypmlczTuOAfQec98Moudj/v83RPwhM+ezPtHzQqKlnncwGEcLC84PDvO6b9g+CuaCurDl4jOuPzq
/fXhX7WJFTzOyBF1tKd2NcFK/SgtxnjdPWk05ChhQrslYGVgyXf/7ubf9r0hLjmoQpKrYSxD0Vuq
N6AumBMyqx8DUADboPwcuVBzSb9O3fSvy3CekrlpCjQBk4hgpRMlnvJdD64/j7prqOBRMtAsHaZj
wBPSPvjkxkPj10Pk7t/h3DnVihON471djEPTWxPJTEPirbv206gcFNW6MR3jYijA3ZaFvkvbBg7N
NdwRpAuFx0hRUxlRAY/192TSQGH97ihrAtwZ+mrm3YoEUkqWEPYW8s2Wt4erkfcyLxoa2vrfEef/
efFbbe2A7r2yYibh2djrNBCQ+mVLkpdYa8zWI2jdk0npFqS7k4nFOZc0pq+uScbGFuFUrUXxA37o
RmCFjuccBl+GEVj6tcya48JJr21cU7xXTP9mOKaOTZU2QcISQVm8/VIKcjEVa1lI8SSTaZ9HAQGU
70psaKLh2a6ejnc07FwKHBoziFEpVutUnZ1q6PYTrNlkFhwZuX3ISi9+ecHCxz1aSCL521RZ5IAa
yoaTLbTwiTxJ53OwZepYg38p6+p1WI/iEqTC/zofW+IabeQBlGTF4g3jkOtCt7uQgyONxNdj6HiM
WLKwrYvikQP7cYDbk3gdKUELY2gL/XdvNS797R+fQLIzx6Gd2R03Tm/mbkGMiPAifTW2igYOGS+p
61qTIYpTet/HtCngLmYb9940BxgL8E02FgoKQjF+ktJBiagkv8IYrREJdlz7M8TM9Ym+E7HiS/R6
c9MthppNSRhGOgClCW/cfHlQetLLK9GyMECNzXhHT0pYaYoyZMP7bha9kuotOAuxRrMlmtT47nnS
PP4Gf9ZoAwb6sFQsslvd0GKA3GA+0WOrMoZCxCf35IcGLQhqVdjqePHXOsUmuIFedidG9MbSSc7r
uGcRiatKhxIOf46DtUh9GXcnTCh3By1zhJtLCoVYrP2YRhqKK56p3DrMvm3/TE1IqdvQbxZxgN1r
vx0BkSDZk5e77AB4+OaR1EzzWCMwcvNhFPcc0/2eBD/ZBN4HxkhBRBKNTXZa1IgqUE+Ak29djfsb
eWgWZmnyNxSeACVTl7W6jgSJB5WJMlbafwcPtJ2wCvPobQFbR4J0Nj1iV3tjMZFriXq13S/Z2G3a
Tdo/OmPZ8yfr79trPPc9aiVfCs+0ycVOKqV4zDKAigHBkWMUqIae6ZCOb0d7/RoxPW6oeY3DwddU
BuL86J+mbHrV7eg+897YbJpSFBoArRFLPbcEPbqA36QNZZKvhw23kVyqQEUngbH4IqCkn+Sr7324
DBdppNzTiHDBiCHM7imyu1B7P8GKL3cYAZ4jQldiFwGp4FVnjilhNTT3h7k0glOSSnUjBU8Tvzd2
JP9fQ/WQbWKpe8AlQBiLUZS1QMjdyj3wrWRvf6uXu3bDbBVKbd5YXaKqK3eaPH8xq9A8GYmLJ+ln
AGL2fpeoM1GC8gX8qj8kA9VbAm7EIhuAyaarUCiZUK/v+zVyCKy/53DNEMVBd/OaHNoF5st7xZli
2ZoXj3wLCI40Qg4Mx1C7RLM8LbS6CJ49xArD4kF/i/Y6bbE6lis6lWKk6Eixjt0dIVdKd6m/lUgY
ZcsoSVzJVf9NJo7D2AayygfkajAho1s6CqLFjpOgXEY6PYyTgtCJ3j1ykDi2YtCHEgq3ZyGFN1Lw
WQ7lZXZfb4CMWra7X+E+JpWCRnL/yhNW5+TiiNOVBMwnlhf/GOH7KxOjuobQuSnyuMqHA1/PM+QJ
r8HAEJY3tY/3QjiBZOTUGihs/EPWsZenz9pG/Vyc/OunRTi15GdK5Xi3kxZKXEGkCBSbs41epLas
TRqsYIpwLF6mDiq2SINglP3C5eJK5GrTZLHx4vc18mOQ4pdom+Cv9f4+piDSa5JKK5UmW6wRf7CI
A0YkQrCL2RjJrQ9yffHu6vBqZJjeYfZmtzVZ8WsE8iprcN1etbbdt+pr/z0Nb65wnrdM5X6gWWqD
ZeRVrm/Z/RjggR1hmgpBUXOvQAWFhaJ6qOsY/uJ/L2yd7eZ2KRWibZb0qRCiTMxsJdwJJuOG6uEH
Us2ISPXrf0s3PoDaL57+HuMRD1eH1wf+Qg2eIQdgEAzpjDEEywBOEyJ37CuGwUlowHc7olWwYrgL
u+QFrBFLbTmfbxT1uL4e8oMHPFbQyTYw9i/PJ1OivRTqagcm00jmeD+dmoNippVgEm3A1gv0RfgH
LbPgoEElGpvQTpZ4nrUTTRX0+VHV00S7kYDya4QSINfI34uLz/3UuTQeZhYEodXeUerDbnRSEw+m
QPJQ1IswW+4MndW5VWuVUtQGVsrRTN7TeIdu9vwD6TO/3ZKc0SJa2M2578WEgPY897hE4skyL9Mg
K1AP0ha2OYk9wBvbiNGZVG9+cBim9FE981NJH+59GJ6dQcSVDZh5zz18oQYYwvH11KbFtQlvxCdx
+oxIJG77hSmas2Vyy4UOhd2dwJU5UuMfdcTZxgJxFOi4maENuma30fHN2DBQhNH0iUjd+KtoW8iZ
kbiqOsm6MBkFkaenm9Ab0D5jlPnZtoXTTANKZFy0NNOWZd9ZuPtEkaLcG3zDbnQxap/e35stwRJJ
VU4mXPyiEPXL9XfB4JLGUPMuucXtjJocJRIASX6gtw1lVqrvzN8OZMDwgXtUnvQmmKoxSkqKlu2q
oywY37ODlBgJnN376pD/Ojoa2jX09jzXvoSB846uUjvFME2Z/c5q2Dupj1pZaVFn4w9fRTi1PWI+
FQgvDnyXmHtDsPhiHDkDK2jo5nUkuMqY1j3Lp1BFvY5W9T8yWgDFYyMs2IuLIdUhEFTBd80KXXVB
DSKq2kuuIPwn9CdvjT0k+1vVKadFIdtjRcDKp+TibAPw98vZs92dLhTo0gDq4Zf9+nbgRs2amjDu
7r5Gjhx0KlsoXs8o/GqnCV7MAEiTX6fKwgVSZXDdyOCmUs38F8dUXMcwyhwk6zNyVoriZWlCfDO2
eytVVxqOPLpxuSL5GwOzhd3sugbr+QWVbwPG/IIdfctDHxlQw56KCrcBnHhtAhNhJAJmnFEpkHPe
lYO5S4hbOMt1wmMs31qa6NeH6tgUfwbbIdZbC8kCaqAGvdXmfrDZ+wzr80W77Bx8mCwiEx9v0pPT
YjH+gfkZpyt7N942MtDtjjiyOUMfHKnRTkxJxIn8o0epaAnk8CSLZ8qKjRLYlz381ISA1G9UFoq5
DWzo1fi6ZOxBmakEAzxZSoQBC+wPg8amhiwOoBTZWzLVDZJxpKwJDveTdDN5GSjXjwVD4KJsZOKX
YM50Fl9E52NTKAqvN79L+JuU1z2gM7WSSdNzPFAmq27kEek3sxenJN2W453JcZWxgIAdiH7CSU2/
+gopKbEUZ9bnAw9rV7No/e9MVjDInQz+YSUFNxi9v9IACEzx7nHRrXoNTepp1O7wsdafnHKt2JDv
OM9uLoLIvT2+cUpNGdqF4LrVFuD0qw/wo99JOnDoSU1xoQ+++IIfysd7Jz0J0QCMaUFJHGZEhrVi
70oylj+2wLEktROJhX2/SVcczeZ1stAv0ySRqu+iRt4P5o+/4lMY00OqPIVPjsu5XU0xTNVopQYo
wi2+mzhbtk4+ICYvYvpaG4A7wdbOYo6V5i8OLCtrytgAArUKe7eKu+DczCJVYo2wTLqgrNZWGGN/
WLhCoAuG8urvYkX+CzRgw5n1MZSlLpOJvQCGwxcVJJMn+tX/hhqx7DV41r/9nwAYFSW1F43ABDbc
KZZVKbTNBIuI+zgd87JqhNHM+yJH5Er0rMAmwGI5Ae5bwkklR/giePgCuS/zi7VKPpyG9sysUf7u
VQczLUvOmfsOttkFVODF19oOwsO09Kg+F8+fbS5WH68tVdDKXmJDIJCwXgHVMDpR84ltUp84zGgG
kF0C3dX2oLbzttcijLi1IdioM68YPF71iudvD/dIkSn+9jupauQIerfKWEXi4tLE/me9y283zVvB
0Gd/BUZ5EGnJQN0Kuf0Nlyt+h2P7t/iYQsPeL8UUMCpVSkzR82cZhmHnCzAKLZtyjs8Cu2iG0lVk
3Hc05GpmL08CnWsD5HGEUm5UuDvvtwLBC+Vwr1wlntFo0OiuFKeg+lIv0J63yLf8Aq/5XbshKmyA
rAB6b4+jU0R12IA9eLhvxtBBNRo61XuQsh+U8I+2oOcplUo/Eai5Qx/KMCjKAY44JQIUcZI4bTH9
ATTzKyY/693tfRiJB5TasUPs+irBr608Qv5pKkIVJOpuBXE5QT1ZDkAljeZhsQ31Oer9xRbqoKrM
XlYM86eVrb9qHv2XSWNumYmlnHSxArxMdoeg+wgP16zYwHfSAuzHa/DUJTpBmz2c/QwJ02JSj2Dl
Tfs06UEzWoXQwcmlX+vi/JtY2aHs0Id5uNt8mLN8Ce8ZYzP2kFGe6uqZzOOGhkzBZ+aAcyKfus6T
FBVWPnaxl9GByXdVCzNHIQNuw0pU6t1TYPxWUIu++eqgSt9W49+o16GvEdCvn61ePyDqM4OHwUmb
HD7JalDe5cwktiXbR/KDag06/u4KHPED4BWeqn1CeV3dqsiUKn1R0Jfu+OP01UtPgBkcMOghZLP4
6YcBcpQL6pTrfT7Y011pXuTGw1z3Ik0jaAnPbUgkkTK9ADcMFSrd6OlXvdGONeHKuAZZIRe1SGyh
EJN/CbQYSDmqKTx9agxVxHhVIb2Tq3mWckU4qddVQzFAyhuztkrLNvb2xjsqQQjGLqzQJVUEiz9s
+jaHxsCOXCn2onCnFV6lRPyFNfvo8TJD9+RbXjQ/NOpsgQ2Ge67T9vyqozDrwuOk6r5r7pgxMXBZ
Wzquatv/QJrEo/4ZsOWOCOJW3sZIxVuXMcYSiHFmGdvLmWYH3vdhXgEpFcZhYThBL2oNKktZAPKw
mrmMs0z32loFpwsrWq2yN80XqIEkhNyzivjYo7ocq+Fa8ooPARHMHPIVu3BDVRtweA57yc3yGKPK
tKnQOsGidjUWlc3neM/z9DdoAjp10/DJPD/YPnKoECAuVsh3nAyWjAERusahhSYiZKC3yl20Ds7B
xMvMtc3KDcjkfN3Cf03qZcSUvuzH1Krs0yuJoP+p0O0CIhltql7PZRr7OUCylOuA5HlwQ7W7bziq
fLAwuRHAF/dpvHxREa0RLAtcQe/qZ16kCsA/5iIRundZoBYs1VF20g0SmqclX6VYfZU8ZV9HAk0u
9uHl8wuTUqGib+gTZrlEO/S5KBHv3Wwe0DibqZO8mXx6/JsPTLJLL1b9y0pHJ/CkvibWIq9r4a8u
3x5hIIa9JrRB5qoCE0eRpMt4gZEBjOH2Wt7jESYWWUTiiiSPVcwgysK7/QnGxpevhIvfeR7ag9i9
mwBNQR2zMscU3RGTP91laT7e2U/S9UOFToXfEDhySLVS30hPN5U6NePsdj69TgLsfGA7zM+zYwsA
GUOxKPHzrbP01as4RddkP4bfSkDUcAwkOBdWYoEKlVvA4dt6/lwinZqF+R9OXZg9S0rTMQUvccUr
7HmAUR2uEXf/DM5//yjWQ3O/LZyf2W2TLD3WEABh0p23bpWN27irPUYpMvyfqmFkAh01pC3wPk55
Rtzbu2GSgonlBifq5ep26CdLmdpAVdfZUEvHpIxz5MwlZGPAq+hB3d6INIn0pAkcFAk3Py5+SdmU
F+KVoGlyGYl027JX8RYGlhilt3VUKE9achkqwuzcUpn5YE7xQDGOHgmGH5CRrcS5Lpgf8PdzEMvE
8CdtLN+9atdB9gJCw6U8tauZd3AXJT/H+Q7zR4sUQeqU2Eh4Uy0hbJBKT01311Aa3A2QIGx1K+yk
HafMdgrA4Afomzpuyw70hRu7yYZy5dR05gKupxS4mtrab7mrkYYUARsxh5yPj0FSKd0v472ZyXqM
4xYneV5r/rl0ddNyXHytWD6uYh8kaTXR+DAwDtwYF2DBo1E1WJ3cz8iQyVOyP9hbnTMwXu8glEZz
ZEul8C3yNRKlFRz1zAbCrRvcj79EId5nlsS4mkU4VF++RJNkqlxnYHp0OVwngsqrAoJ6nRBe9S5a
6xaBeMnMuiJ/HJJqo6KpB/oSOxZr1nVe3Uv6JnSjD3hYrumkBLfnjFaWXHOj5oAD8sYqyZBanZda
HcO4cmfn41Ep3Ol6DXn+EIKiQs1idCcwgCBXofD+qI/qmNbNjNMuPAmAQhArSUH8roC2Jd9PY4Mv
uPl8P/6SaBA03t0nnXGM6lpnOB/+isB/uXcrefYGRNoK4YPS+BXfah1aQ5/x7Wza1RIdxvam5Stm
QfInpl+ZkpRdp1tcBscOcGi+HCU2OPunG+mUYrCDh/Y1Sds6hrLL+eBLEnNe1zicQC5Bbu+gMrpU
uaIix7Lkp2eSvtSrV4MHboknCzMH+yoXOzvNifEjpDp/e0VcsMdhJi1NdqRNUbsszE0hCHCHjTNY
K+wI09JkRQ3j6ZTBD6N7D2K39QCjo9P+SNG2TU91Bdup8+hAQ8fPcZlrUtOOC+6CjnnsW1XeJGl+
i4pRxrBhJIooYzMdqlShPXLcK8p0DoAQme59MBBxygN8POil2DNMLXgA4vZnwhoDFYsICz+qTJyV
AS7k8PWuNS6gaOc8VXK5mx6pBBhNHY52nlVdp3MOg7NCAO2nWb0sID0SqAbKWidF0lnn5LQkp6of
WcIRfcuGXuG/YhYLS5yLnHZB3ndNLOm7Qy51t7+SzxTX3UmPDgRjOazv0sa9bvk4OGOQzw0c5B+b
n+xl8vV1wNA446afjtQdi5GE3rFVFoqEPyiZfuSf/gh/tU7oGJ/Au8vOP0rvJFnIhKZUCczEQlVT
QlCy+4+F+LivNXvvZGbw3sAhyySCXKOyuQV4+2ENc6is+WweZbQjxGqA0EL4PhmQ4WsmTJPsn4R1
jLDc2PkzNHoyV8s2UggRUhP4EAQXyqyUnkqZX2ugiQw1zWTyXrdkCs+Fz+fohQBUM86s+XyHYH6Z
2v6bCjF1/Nj0aDoFxIGVuSrZG//x7mA8fqY5wJteRKW4/zHI3cWWMolNcxFkaGnuJVB+le73RXSm
CQMwtaILEZ5QfxH+oIHQlaQ/S4eIgh2MyTlrpYS1AJ3pK7kTQnflSs0KHcBZyQ+sF6vqrnp5J1t+
QRt9nnRh7T277YNCiKk3xKvajE+ouDv8OuQSxAV1pKLXvqgUIqg2uEhAlDvF1pUZKIDAUIepw/Zf
5C5P9e/sD7js1Mln2/rF1bUKbJSYeASiPlSThYfA/OsjuP5rRTUk2Hx+tsnxlNkK0h7fdCSZjcvx
FLqmKWDdHiWJQkV877kWZKXT2H0sb+CMUj1x76p/bRK8ALo1Mp7W8fij0d8+U/pFdJxOYCGpB1N1
Px8kZcPFF3HG3PIDM2x3hdoe9vkAkViXjNVIKCsmAAooaKpiVm9qd5jRsb+b90pHsDzDLBDllhij
iZ8AhHqWN2QLsio61P6fHUL7rPnqNv3c+25AhABkfnpFbwpiI0deIH7So1JQF57t4uSngtswqhY/
xVNmnrvUhSIUfOqzC0Zm5nUvJKlSvEmgiB2jt8rzD6qSTYgJpSJqQwJkX47PMZbsbt93C/T/uASE
c+66xmlmawoqraiGDWCag6O4cvxbA7HlApI20IsCdmWyCtJ7cmK79yU1z9sXduNj1I8shWyWg40N
3oQFE0UFlbTrbOKTy5PjaLVss6kxVkM1rRvZf/YfkkQY2gYTPb257RBWseqvazhebIbPyYWmz3OX
V7V1D25njuBGtTy98tIdRa21vKWJpUWeYE+En+EOPYe81m84XAr4gBzBJ2l3rSt66Lm5lPdADRZT
F5e+Q9+IoI1mY101WC1Cjksev5rxeI1eDNMKTWoiukdugGshBZC9gv1Zd/FNvHkiLqGKVszMEaUM
w5K6HFBMnVlL6oSK1sxMemvaFa9xnzVMalcdQ016QL1TNw+p6vt0sIvba2/BbiIfAq/3iOKezdDW
FjbEGkxl07n+XryC53Z8fKd8rGjzjXA5KcNCZNACYTpueqlXMW5KH4/LpGAG1Eu48fScnUGFKdes
3r/KQ2vmFZapcOBrL4bKEtWx4jxc9v5ynzH5gySGmw1OP10bxO6gXU0W2ZFkFgwzqKfyuy1Vr25+
pMiZCGSYd+0utwHJogIiNo/Bb4D51F/c1ahin28JracIPBWXUs1ncyEbSnYF6AoxNRQwZjSZ91Vx
TprwD7AaVh6A87/y30ynj7rVC6CnTQBeL7Z89aNrceQlEGdyZh1qA8P5qaP6lBqqlM41N1yUXfWv
RpcaWSZaVkm83CFVW+bmkGUFZBr8Y7LJbzaAxiZxE+uP+DrQtZ/oE/oZnHm5B4y3qfJ8Y6WEIO2O
/ITGlMvdh0RwoaUwysLeqojN4HaaFZC8CzaVmSAtzPwU1LMGH0COnR5oKkLcG4aDF4qwjLHnVgO5
FFy5Ssv9hC//6pAXVENalmO/v5b8wyV3q5MwTvv3ciGkhhNyFIY8VBBSFUwHdvIOIE3GRBlyuYxo
VyGrxhbPh0+0WvdsB3QInlL5IfONdpFzYJgQHy12GD9jRslAGETJ7T+ElLgqx305/ld8R8fM8kh9
AJaxMafRgIGHZn2Hy2K0njfe8ctNxXJL/r6pGzOM0sXT/Jk0HsRZS4BoYyp2fbJsXdNmgLDcQnjs
IzvO02xCCE5Cs0Qizr2HmB0TXNMConYwJQuYXh/z7i43/t4K0zaNfkx9YDylk/Hex8ORLsNSU80H
jUAJhItzK5PjyWBkZB2Di3ftPCXHRxMkPNqvpoVSKW7fBRwYWOS1aY//iwTbIm27QVSm0nrVqQQL
yB1HFkCN6pMIMXxhCR8Hajr6JdbGZYLRzRVRusV8mRVXm6s4P1VspFhSYupB25qdHnc+L8nez8An
yKsqy7qt8+VlnoDuRlwpNv2mSjrcUro5ZVkrb+7igIyuM2MrkoofPehx0sBp92LeGdKZ3kGrU2H8
e6lYXw3VJt9cvmS7FOhHv+ULy4JK/UhoWXWAiACByvsrqii5e6Q/u8Ua3MdVIycldOyX61DOemVG
AJIOZk/AYIABwJzw/Cq/NMPccY/74gkcvPDTQqx7piIfoEFPICKk8+TyUnPPjBVYDFsidpGVPCq+
2YrygcXT/qVMvodQtnpL4H11XOGjqQ3ua/SL4OToH3WbaUV+lxVPn3rUh3vB05BUtpIwhSe4LZm4
EY7yUBa/ObN6zm+u1Yb0xMw51HqqkjuIZQTVaXQ9ZEm8l6x8TWp5i3lbSG1Tknwxvl/SaHRkcEZn
pF4PSnveW6jw4dyLchCCWKPvN3CQdp1KOfAjcTDQoy+HqQvbG7+SbZozJsrN4l5MDzZ1/d4but8n
ko4ixPRgLNWEr0//TX+50oJEV0NZjF9WNurXT+FhzeG4ghSTCbD3hC3nUjd1vxwLEO7SH+fCDtOK
6aaFHgd5RmiZBpn/RN4gS5lHTgkLIQFMJrczncWoj8ocPv9ezlPPddy8n/OKzOaMk9tPwy5bLJ0Y
r6cN76BvxhaE3Y3YYnISnnCfMQyYZrUFp6HbQPWNNtz36n9KhiVld68RVntbNds46UlJHe+scFkV
pKHKcSDNvBf/9LJgftEcuvSgLtiFNJo52rrDpytgcPXsxvNnBbKSRX2yGoXxmIq//Xip1esSYe6N
TcRctMMibMwjP6X4mMXkv8mesFradhowPkSmj0olaCjYj/1noybCtp17+eqGP8SDRKgwTijzcMdz
l2Wl9cIaL1mZj7xoxoyClW0Top18PWimrVCe4wQ70vQuNavhBXNht8G86u80JK0lH7cyFcEgOK2g
kC9QWMOibGcGKBLMTQKCe7Ux5npceRK/pqZyeMfIlVIOLCEcB7O63A1mzQaZKc85YCcpF4l/5gXV
87AG5SDMTPGEAWymkprhApCx+sWRg98wbsWdNGIsRIla9tr6JPf7Yn+HlGeyJCcMmobDWo2dUEwD
xRuMeknMPjHkVoMEQ/fFr7OWJnhld4GkXSOMlpc8UmcK+PQ0rbdVpwandkeKhmcJl7zokZtkEyXf
FAGAccJMKTuqTgkcLHT+KNY7WBWcE9iGVuNlb8pK1oUAPKktgpnTMJIHD0ZqaWYUzeDrenuXOtj/
ObRbtBVmUCKPp3WxuduIJLEauPGZHwZuaKszrdB8V5xDZRFf7pf8Ef+0BPviOReRdJQf/u7mdzC3
hNpLMss5zbAQRtSCzWTTbXHcuZAI8JQa+BW7YEMwVMBgySSYm78TU5QvF+lGucLUVCnAu3bvEcuq
UC2ilcFSlCL0zbUXG/3Irg+zZ5+ju7pmmRoNwaC6VfwTwfmbB1aD6glbLBrkbcVzk1wGDub62fxC
R/zPMYleXgYC4rrrgzWwks9jjqjYWr8nQlXqz+tnj/+gQzqp392/Hf1JfjaEEKVBaU//62Dh5O5x
KSENA6Z/eZwP6QanO5kJeYqPtEU4XZn/Rg/QhWVrJD1VDk3BJc+se3LGKtJByEhrTh7SnHmk6/2R
rPHUEOobnsowlIs+2x0Zj2CrXuYSNyxUboflRKjSYGNXbMQDygTl4UZ2j8hhvyl9KFgvhhh5SiNP
yh8GuVspTBt72Wnuv9VVfCwaVg8NM00EhgslR/g3bye8LCkraSlEVoymbxORefmmODY850RsURv8
wHu877nXgq4IO6g1JhfJPOObHgxDA6uMaHr7nmPIe1Bkk0ITzd0O7dzw8vGEHAnJ5YaD3E8gS6ug
7VGuHYMZugxODz1JHYwajTEPuQwS7C9QUPXtN1KZCVwUV+6I+q7mhqanykSshNhW2qnDPoZvi1BS
tGJJB+ikmvYvN0wNg+4a/ckL3/Rmb699SqhNaZ7cLLIGRDera0PunEs5yJ79J3MzulBy0Yu5zA17
qHl9/3eBooiV9mbATK4a/alP7daIB5NELogSLn7U5RAj3eZ0IoNiDuFI7czROm+Q4jHaTNkbocZs
b7C6JT+ddXzaHPw3+TF2/9JWr+m0SwbLTIzCDXnRNKSN9l2u/ecS4cP9W11p7rr8FNwhauwnHqDL
XnS7gm6dgkwVI7bZksFGULBdVu3H7ZAZ/gLuuFj17C7bHnnVQx7F7jDIW7Wa8zucoh68qiqkUuny
ugk+gQkGy0+C+iy/53QsIw9dPDYyax+H1/kl102fcQmSwX83gx1dgnwpbcXxEJoYAjy5H9kELxMV
VJhCJGNcju5GTbaZB9142KqnxR9EysWNH2eytHKCrS8YISwoU6cQB8KQfS8HvI96SrukR3YYilDX
4ldjiJVBHAQYzRqSUtmkV+9SeYB6QOsscakNynLFn56ABp885lXmnrO+qN0GsyGnSV+YDSKHMIPD
EbsP3ZkKyT0lD1bMwfGrl1yKWasvm++qqKXBKyV5uvL44+agK8Rn4tnhFXAQJ44D5wHI21G+kyAa
qj0V3OJlbNKnqH9L23mJPFbdf1cY67pMD2chWPG0UDBOCvRRMjO/geE+qMe7vmG3V950/Fscmm0e
XC0PUH6i0M3KT/nGIDP6UdNlEs7qsPTIbj+iETtdYPpY/0tYR8rloYqMAqN2o03GXZlYX2XX579s
phac6J1mVB2fa1qCl9liovxnrlunwqqwi8LRFuylKbCywWgNEjs94qTy4yyJUsl/x2l4nYDWcIbf
bFZDwU7OLLde9KT0EqfYAzw9BeETlvom843aVXP9Jp7XHNVVCXrltTbEfjg8Eg81/iJu+aCRg2bf
giVvdslX1GcrwGjgQYSLrGooqZSYkUziNt2t/uCEtDuCQdoSJWK9vJ8KKVWXem5c53jpySrlk45v
YumuBTI4sWIABTmRawat3JXY5IdKeK/7xzUGVCOtnNWKdsmMh/oFEevHbtC4mpfhB4T19vZPRGoG
jJJ9CXeVfT/Wopx9e6whmXuYFVGXRuxLw2ySptm2Bhe2Hhriflqv1x74jj6t9aYba3+OAgPEw2Pj
nobxCnqhQQ1Od6mzdvS6u7T8fYSI9jaOe/V96Xj5/W3EFqL63xvA79OWuCLnn6dH5b6P7tMbAzZ3
mG484ReF2BXuOzSTtCajBG+Z2eLhCCHyWa3EfdPCqsd2ROuMUkbMQIo7WnpO23KEZslfLf6YyF+a
yhRbKoVMUUdMLL0hB6FnL/LBm5XZF52J2cjGXJEOnytWGpqBuy4dKQgU/35ngGCmEUd1gafRF2Po
7slvnd2xHzfWFhnRoQQWM3RKMDTtbt4u+eKkGoyQRC8XQdod3ff0Xxrm9E+Oq36qhYGt8B8GIAGb
rg8iJfm/8O5mr6YM6cTHP7GKI9zGL+3r2Xh7NoceXbxNwAA/TB6p16EQSSUlSitLcCRy+LZGXlYv
+qVQ5vfuZOGi11BE02kNFdo+pqzLxUHj1g6ofSNXeOctGeVoEBBQ8vJ07YrwpYz5gONQLibUxgxJ
sjGS358MUaxKW047nbkJkC5LW9HwNbhbFXZTbbd9xpZO6IWZXI+/nc9NwzefQID+IRtoawImQtkK
6oaKBkYbZxEKtg15/215zmGvd09hxIdsqEFyhczAga02miNByDe6j187lIeg4Ojk11UAiRH2dCJ1
Exo+zEyKhvayCUco5AsCVnRdXKPfFuzxgJF2ru2XG7KO5x7+OXhcYkYC64bxNijPTd8BMq31nb6a
WLuAR82qXbjfblf0MtXP04IFr2Yjqhyp8WHp5vKxJBlhrfpR4l3bOuSl8JdTKXemXVjJUt4f02B+
IrdoXviRhHOsYZuarnHccLCBEuHgqcBgJVI54AA5iT6JfMbMKXoyBfshXCPxBci5/BN+zuSWQaPL
o/9+AJkZdl5+DahHoiFXTlthSL7/HwpInDM4/q5IqqFC8L2jXsxGa9/dAPDOl9FXwKPLJOP9Tu6s
k/rfwREg5qSACfmEAUyZo+uhXIJaCmDpD0oFo9Rif7yOk3lJjWIu1opn3Y+8BcAmS+73SJPrcilM
HpOsHLe83oMDddeMkqE90uzJor53b/HeBybpuM58VUoDoGUjIKGDn9wnymk0O8YkNRZuqNAbz12G
pTbYRkBLJAq2KQmvresaFU0lmwVT1kfxTyH7ZDw1ehUoTMKi5OiJE/mu11YLPGwID/HBuLrX2EBw
DT8CBB8zEb1ma1rRcjAK9PtF1W/1Jc/fKAY4+MQgY9yX1n6jNmf/QNVZVJx+X4/XAbnjRRpvbuJD
gUe5yaaWLP4fTbO+9HU9bvMOCUdorSSKxS2CRiCfTENMOvNb1pDgj0iUsdm93E5xne3XnBB7efWZ
7o3stwHI5uUumAjta0gMLYX+8Zl4J7nFDjb+JrP8a5/52y/Lo9dokbt8wYYe0/558EN1kP0LVAPs
j1kJCGtFmaH39DtbbQ1Iqaraa0MyuuSfvhuwdjXIFFhwHffH9tnfCBklsxk/ZE+aqLFiJHlSRblh
W65w4RmQeGyW+PlGsaxz9A+N5bImRb36Pqay8V+0gpYYcUO+/nW0N5JhcHC5zRaMmZHpWfV/ve1W
4ZTiCVCYfOjx2iU25PFAfZtzmhjO3fUFu0tLbfepjKkXEDGphnSrx7Ovf8m9sRLlL4ff1+2R7aUy
+hAXKbL0H14perOFzTler3AnP8wJi1etkh+ZK/pgfRzIHfah/N/X/dbnqsfguxNxZTN91lI71WFh
NTn2UMJ/VdA1RGjZi9NfcyjZYbE7ePz9Ah+0aoILQlvfbGsg7lRm/t+lQWF5gmnCIv6Dh/2PNXMh
hTWiAd8u73HZI+294cs8v4Bd+8VtRmDnU2/tEWh28PunPQTaWOq6iuw9Er4l713PsGTnHCbGHAd6
RaRE/ugA49N0G/Bi8Ha9LKBRd+pwAFMAG4nLnQFO+t7oTMEYAI0iirOazd9niRP84gz+si7BvkFG
pN8daP9umC3yQo//M/7LVBZzf5BD+4XKuJ+31fKGq5CG41OFd3sRKmj4v6th7q5PUMmZ38PmTlKh
oib7iByItYBWn6ftjEyNcIsg5o+G88hIOobc8tcc/DWs90hWvkfyMMX306twZmhB2m3B6wIk3BfR
3CaiIOB18eVU8bDefPLkIU9WgzdPOk4lrCOryGMqGkfekpLD2BG6CCrEeZrKasogVtuxDYcn7or5
QiBgTjXQg3ItqNO5wwu9kwKcJ2S9BjaC5h/Ae3OGDE22Sl200UnFmKidQ/qin/Jk1Jj0HZPDYUFE
f8oBIiLGiv+pVAXarYoaPRzCagec/xjoecyvFOsGKCf2eCMt94PU+xvXpHuNxjiR9WBYpjsyqUfE
g5fqWwpSCBOBnEEFIDr8Te4PSIaW0OWAte2/eEr4+0GwKX68dEw4QEhMxneJfENgBezG+e5nIy7i
hqFUlK7XkiGGW/rl/LqT+kteZ5MC7LX9XE9R5EubmIELddMetfxRvCEnKL6F6eaoIV8MKQlvVUoW
PM/4sGWw9K/N+qQ7uqbOjU4IZ0QF4ZWh/p1Ua6xsyeWPIWkFLobsZgh48HYxY7R/+DKnZ7ZT2kM9
6sgMvzvM71qwHzoZpRshUxxaBQ46fWvzGi9V0GdU6gx7hli+Er5dUuzUX+5QZe4+B+6Vt+hOFOrQ
+MoqmluaZdjYZu3LCybWuHRJlFU6WMySs9EM+nkbYJGJGDLu0QR/HqQ/MO0KPRohsIJWhLkEP1kB
W/dpHGeEUbLfRi1ANFMhxXuCkivD1L8gL4K0MMsllsdUO5V8br+J61prpFq24yRqKAM9KfOrL/bK
KYK94BVddkkaJDyICSWVBbRPH5ohExAEJuvCAd3vexYWkF79EMdOjf4xGkIMr9QYdjdstKVqYhlI
Q81kHY0no4llzFNNutiE0K14InT2amm60/21isIE98f8lqqoz7ehmw+8ah60pjv9dYMk4QP432nj
n26FgZkdodAregZ10bRCuyMJHrySZi4SjThLOD6T5N/1YSdKSt8QRaO4jvlsGpa3bXOMTEX2CX5r
wnSHVDpEpFJ+S+kE7MqFBxU+4NXOwrMb+uSsdObRprvAau1ANMTvasstAnfegoQsLW8JNF+nLk6I
GuWWF6pk3GNZ7xLQ5nN09fu409edbq20cR/sJl4vPtJj+EumAXFswCyzG5BCqYfAquHGD2ogV6Nk
zeOeozzBqnPyLtIMVL/RNxpWxFjaB9dUAxfJjnTNRcMWnCa7gMQXhjHqOJvkKzam3DsZ+hHovPHf
rzkl6+uThU8l3SGMAzcxdBE7GTYQsUAuCdle9F6oEbqnbzFCobzFRkx9HbiVXRs4bFETz47rLonI
xklXtMJO3KtjLeT7dgY/c2r/ATVcXUPFSMj7CQ4WIZaGDnVCE7JV57AisDSdOAU89I+Ka8IqyMY6
iyjwSoTl6SJdT3YAo23C9NUVzQ6qAiAiofK/hGcVc/vbQpivKxUPRgjzT40ULDy3qyJvLJt67x5F
HftDPuJgCjpZHNOB2JbRQBxDBUO1KVsZB+HhoW2ZJp2SxxWw8vk/mYc868LH12utiBaxzgyZ8VRM
tAndtaCR0kD7sjy+alM8dofc0BACH8F29Ev+ic9f/ebkfcUp4IlupWOPQk4h+iK8Nds/WWdzqfK8
lf4CNXz2Edux7usdY345V1bJv2gIUf318LIZnE5pZ/g2YVBomFD77z/kHH5t1s3rAfBbq0wIDEyu
EP7sgbkP3bK00h7YQoEROFo0bekG4B31/6A3e+xBtHHsCBGKbhVexrQ4veVQfj6GNWjGIXQxu0sR
yOKCNkNVQetKS3JKmqUpQ0mVqHLvHCmfKqswrPN8yxYlIw9ort77yfm7bYXHkT8eOesM7hQbMQcn
gX+6jKtQ2x/xCxGkPS40p475SNzUpzMwmzLhnJwWXnJ9Mu4U5EX/0z+KNx02vh8E4og4Kv4qQeb1
1Njmd+YEMD8yNd1psB1AN/J2pNqTAwihtgda8wpyWLjvW04/SDJSMgKRAHDRQPfZ2XypBluPuC99
evba2tQOJoGJcj+SFTvH0hQ3B7fjiqaeRxYAqQf69ATuYJkjIXBj0z4BaGxFoVlNlO5Tazk64DPl
o2ifoxyW2ABLB0OJ1hLEnvMyVfyEq4sBF56fGjNsuAny7rttUd20IH9iPEwmuvSYdT+Ow20ohwyt
t4k+EHHAXrzVAg39FJ0TkEH11xvh5IcBJDlOwRJcHCAakTjef3sG/1QMfuQrf4zhhud28KzUVh77
e4eDPNNQr4TzvTqMc2CKOgAzwtQWcaFjjWn1ss7Cjm89QK4sv6YldGT2CSrsUrMztIpsC9P/I0D3
+xh2bWRZkoC59t6G7ND9Utro/mAB46APfzYLno+JXeO6Rm2ty28rkJWbMh/h7exhcTH2KWn9VGcA
/MDjJXJ2w+r2uz3coe8ClDgPa+lym0Ye4kYK8ZKa5I0Fm6KEmI99HNJDl2mmrUGvDe/dcFNHB4Ly
1uC3p/HMua4oI+lrppWrTKgMxRokIB1Ch2UQ1S1ChcdkuahWVldNEIGGE4z9kZBrtoP/kPbTV442
bOZFLWbsQ5Tm0wy+OV6SQBy+agxac1KnM7ZWzhqvmN9pOxGaMwMv2gfA3trg58JmkPsed8XNofXu
WNd8hg0UidfKgq//xwgWb8GrZB1LEustznygvGer02htm0brX3gjuzp3b26h23Fcet5L+HsP6lEI
GW98HYCA28f7/DU/p0aN6DAfwMw9PSziT/yQDARt6T+RbiciVI4pCGZUJfiQ/B7YG8gUCE0BJ2sa
yGihzARdiBdHGam7BlpNuQK2TdY8fQw3zANhlz9pFyGPa5phevSrguOQPaPyaWgsqBD7La1z10dN
UiKIrCEDihmUSOK2gNOVeSgmcvsXLLNepJTaSw42pEFTMekfjXevD7TaKKTgALwTZxEIYtyqlExw
WY7087SkBR/RtvyE0fc0wSvK7fsIWLaBjEy/QPWqELaRL8OQby+O6NYEzrlkS4dppeNHEdIdSac+
ExAHt+E+qblM0ITT6ULCYvz+TdAYM6KQE6DENn2DIyqqeEpBG0a9cPkQUzpD/+p58vdFX7iLFy6V
6iG36YNDrEnzHx5hws9M0DCHRr13rlejulo0l3egVsoP0hQtdvZQkiNoj+mGEAlxg1RjOZcGnbZU
Dfee1jWiyjFvep6bUb7gzbAWD3X+0HmBE1GNW35wTcl7Lr81ckvextMByA6TscnI+6+3Z/TTWHim
NK+GaZMSrJKKhXW5hTCed6cxx7vOhoi7K9RrJEoaRNSMGcLD2SPMrZAZ8lRX53I0Xi8LO0UCyKJl
SP/3TuhNpxXG/+AYfGD4x5UNBjEBKX7t8axvul/nVrJu3TNrh7E69DBpK1ov8LHyWTmLgsza/sJ6
u4ZzdYW3O4RqQRZ/OwLBByvVUBFO2cKJLj9Wc8KSi8kyz73Eg+jrYIKcbK1tYOMgzElP0GmB2J5z
TVgVpGUwZZJAsLrEiC5S4gL1KkTXM7aWqs+a1iQBAhHKVks1MKrGcrKzMaj8IEi9FBj4ZAHIwo6x
IonrP6Yn52MY+aTD0+ompA2V3kcPqhtFcsQR2/ERCPXyVU97WcLYf0mctH6dtwRfpvA+FPLPqmiM
C544reUdvdfahSFYNtmSX8ZX7sDL9uIqhVE5KtLU4OIBpqZfFXSgUWU7XWEf3UuseqOIkLrkTFKf
7F6JgJUH+r5a4lhdlkgNpG0znkpU1OAh+TJZ8uGCG1US0Uy8XWhOg1rUfx5P+RR4A17VoZcFgFMc
Oz8lz2ksN1wrwAAEN8TGvJdZCj4bltVZa/EBNrFd6VKdXP//VUgVubV/s2mbINE+PB4R+W38eOtr
QUTzQuAIBcuyLV7+Guf3YlIkW0H4wn/x4/nhsEd/mTBpMoByjPteW7yVNZAs2IdlXyDdWc1ueCk+
jXUXkh9M2v7rlkLDe1a3xxiyfhDwA7NEEaGZkK7Ut1n2Sq9DcJJJfpPR/V25or7M0fVMRZjeJjUt
NQrcHqVCW7fu08kJH61c6VuqFjiWhlSjOLZ+Jxg2z6I51iFnkjsKJ0X7Zw5ZGkyT0fX96k3SAXzP
aB0nrKL0VcQRtldz3q8/hFcolK1RPel1qcsQMCEhYDHuWQjdur/3wdizFeKLMfnT0a5aIlajSuov
f6q7XME+gAm0cPiDi3AJe5HFnGYbvX2RiaRAmlBQJRlSiDpNGsL6sLsJf+zj9zaYXXVXfZDC7IQ5
8+VoyayNT7CSrVmbcx0SoMNbef+xzvGkZxBoplt+Ix8Zt9yeKwHPSvTyd/CnFbOOPD2JLEWARGv4
XsAPmybKGtqW3eAfl+YpsFFEQsP89MzLsRWa26rtzCzSbY2mf/6fpAl2XW1g012PhJtRDCTPsb+U
aouvDAxV39QMNzWKWp7u/e1rwyzcDcBpliaY0y2omVLJZHdv6hKdpv92sRo63LwhpEKWmnunHAT0
zot4aZazdP5yIPgysxolI5xXR41UUEx2zbXlaEMpvv9I8ARKHqTfSTRnizjWoyaMUxjn/QjLpr8f
zvZxbAD/KmyEhw1qP3OagVNv9SKIebWRn56h9y9HeOjz0PhiLwdimb3kDNCQ2E2OHO26oVMBoRb9
J+SCNtEMVimYSom5tnF03sy1OTI01oB6vEHMzjCoGjF1lr7klMxi4XmCAtKTpzzXi0wh8K+IZFOV
miqaSjxU3+Myah4C4LwxtKHDUwMpU7qUdfDwJQwce4Z0jhYzy0CtDMCIfX3JXxwT0LAc++m477Fp
UitX9oUqzhm/N+bUAKmlSGhUcqa9xErPenQZ3ZtawUNCZtFQgjgjReCqfC+FTMrBJcTdjIIHPAqC
Mfu4e5ywCPF6195PeqH22rEJO0KjH+uaUDOKYum8sO0WploiekJUb2+wjVSsQX6hILRwPYlErbDj
5dEnbSmJvWnn73sJcBpGtODvpMAi8OAamo6bXXHynLbQGz4+Kl6jSr22ZUn2X3plNLfTR/pesjYK
wpqKzHR+1GDOjyvgXYNZOpfInBAfy85+lz6OkcrYzM/pSqKx4ElldqPeKTRLi3OFRK+2LyAuGan5
oU/VAO/4WwsWwgHIfcZJHPOTgEuVxX8NTlOWl1lfd0aGNqK6S/CcRIhx24H7/xmhozV8ktfproT0
7JCTShAYLNJU6VjZDceu6uAoNYRnCEsfxgW8imMRyTmSvIkHMVipw/NQ1TBxxdLQPNU9V4FbUXog
IzCymQAgWJemI9QNT9BVhpgN5gZiYw28Y5ro7vSAOCW1Q2Tx8HODSNZhVYGZe1kChbhM8H+xsfWN
taV0W/A+B+4Ag/v1/CsTYCuJhGAniAtmPNydT5vU9gFsp/W1CntA4wMJ3nacaUYRMrJiU1HgSbRc
niBoP6fp0rg7YYB2tvXp5rGOviJzQIeE58AtY1qpIafxsPic6Ghxb7zWetRRx3oE3OfNVahoSJCM
X5scJHd2g5Ce65FGTU+90a6vHUEEswEIOL28TolIUfz9lJc43qovgV/az1/gJ1QMZ+g9MEmw2E2S
nIQDv1Dmb3FZb9WBHEHzEUNFPMAJJFq+6itZUbSNmT0X04Z1Wt3WlvucIgsXEJTMLG1V4NxPTUfD
URXxUHkhKVf0uv4D4N4QmrY+U1RxBwzgd2wVI6HdTI/cIMufEa55fLeJDyskWfxcvAVdrWuIGE94
ysuDbXfYsBltYNi+vC/YI9yDalKGrQYwhh5sh2SCuj78ta/D2NhBmz/n1/njYrGHiFZ10cfbQovZ
ewM3aYvGT5mAMcRbl0imac/bHob/VGj1/EP+BoNLbht6SlJ7PT1IcNJtP3VKBdVGk7AEEIzC/SsP
hUfmvkrqegtYQinPKQYSH4Oop+b2l0p4X36O2JeNDGLXcLx9AEI/TxxrE0n8YXb0XrPJ1fiyWNxq
9Aj1J/NmsvmvKGmrVJ7StiRIG0ADmCqbqN0zpggENDvJjyaJvGfs9nYpOrQyUZkVbYjIi4Vgt/5p
FfTHPJ4T4N3FJ+MtiKRiQkuBDMPEEJPY4QhcAiKZTm8evogJXSLFmJMduvRm3Bpdjk3JhPLuwnuA
5z3N/dnMMcrWPpICpqTL4DGcNOF58lfLRqsFC7Dc+brytMD95iwnGh7/dUd7zScE7/NJZh19VWCG
shx5cWgjiwnGjcGlkyGjHgPWpiKBmvO1P2vZiUeR+zsvmjn+lSUkjZ/ns6g2qdv3HHEdDN+XudEN
4cbzkUG33OAMA0tcCZKQOP+A7FObKLu8flZw++oLCrOAHwb+Qxf8HMsxKeBB/flG8JoLGhTP6MMe
LfiDL1NAzlCm3gw73w1D1UjU6x3Vx+3AqKgSXBACZhkwxPtjrQu185OYGxKoDMNIkOjtR+x4QMJ6
hXb72QecaQ+XtER1N9Cl3pm0HgMY0Cx/4wXsUrihtBhduJEPCXzYHWOmy24XAZ//0zu2O16Y6T1Z
mTnnI+pYDquFAXOMmwA62LMt/puOIKY3o46sGs89TkgcwPnjFSPcXkKXNSua5u3VSKm6ovu9AIAq
xvRMDIgSaDlUDQ1dKvuBAcjs4IuhTjNBFwO92/gIV3WNSG61nLS1L++7bGsS3+tBpxrWp9Q42BG9
DhQu/lzdptZt52RXOhv8bfRPoX1oywQD9JHF/ljOIACZmz5Qc0UKNSjKFhpVOdhJEMJmT1MwCmcN
71MLJZi26u1q69wv5QmjXqg+YT9sY8uwZMBbh9nB0AVpAGlxZ/9AsG7MQTCSMst5FXGwp1TcKQGc
DSOsPDkqKzpHR6nBneUJ1McnJ/+XH/0tD6zptQajGeN8gyENsLIz2lX9CGUUpbJ/qxuMOaj6WxOZ
afyqph3ZtDtkbSZQk3O0AB4Q00gG9GOybe57ZsvdoMV4HEiwtZl9AY3DJa6i4LT0pz8UpSsEwDFx
lgSsNOSbpUYNAw+rTyaaL1Q6HWNwGrMZ3sRcOiehXGV/11GesqNPjbOaFWyJr5cEbWz2gZxSxPnr
P4uEbuMQmLYt3jMFIWeaIKUmygjYZaajb2kAAzOBHA34Or49nJivFW5A4rpnsvmr8h9z2VemFJ7+
8GzfWTPS592KZVC6zBJhPQt2fFcxml3m6QpIufPOc8nV2BHklLjZKdCSDJR8C1UoUuA3PEUfFVPF
MwM2NF+/xRveM5E6DIwmaBDQP3fIntQCWe5EdHAWCPtE9VyqwhfCN3BUicdlJhB5WyTCCwoKhznH
DiqpcrsFEgBCX8FTO2kMDEY4JhRkAa/JewWPq404/vUhJ73PQzaQikxw7JItWeh0iQm/l0M8M0Bq
Sik1Z3RF7YDCMjthohYl6S9ufPJwN9pLuBbO+79FzDPXhQk297ZroKaUH2gUrUHvl8bI8VZEcLhB
JHncYeSi5mCG9835u90g4c1P24MKZYibhVLZGjlZOJzCBmE3xeamHniiHlVJjo7IDILKjtzjbXv/
xRkmb6WQ4cbLcaodqyE8oioW+YP4uSJWfvy3rtD9SmeJHC+JRQXH/SWrEyLOfmr5UZLGfPiFowcn
z7xh2yUr7jHM76YF8gZh/SlKJXS+b31+7AJ4dqgCzkgOLhSJf5we52NIyISgAttF1rqkDXyuuAi5
VOGM3kbnPfWUV3ErgzDfCCEElB8R/vGZGzvTrmNA6/rKRw0DT3BcraFAPLo5WK0GQKAvzYKyei9i
sUFnfR9tERfIpS2vy207P5d5Iq3Zi0eZiXtnY5hMraAjlgqLIi9hltdyG7qkxuOzN2w3b2VVH0J4
EVqFCA7s3AV0GKu/gBrkrh+bDbUPlwm/S93SLlCiggGOi2Hf7PA/XMbm24w8YHrprEbIbgeWp/Lz
dxO4JIc5+ObzeAZqGjkv00YLbEPfSim6wc3NkG3/5q/p8smX82j0xd49fz0MwcqNNCmpa6J/pYwD
8J4LqMB/agvDU1Q01ZjOgC4oUPrEwYy5/3PpvRKP8D1SvmXVmv1eVnqTZaF7D5ZaTceliDUNWRmN
Ba1PdNKtSX8p3dmvIbkd0t2IH5cKGBn5UI3/LOz83exrh58tOVfW1Lrd1yT/lCS79furj2bWjoin
Mrkn0Vsq2vX1slqZhv3XQny1QhBSBubIYgZ6nu5nHuQHOgf2l4fO+Pa49lmDW87EL6LctOa4/1Gw
LbGIfkpIdIxOE99pu+0HjJ7qMwDetvergqkH2WE2HTG+nYfNyuy6NhXfGM8wm4BhADn7B/vWZ2qv
+5PC1GZ8WTvw54yoPBwmgHWTMuLROlV9R/lfb2/AT5NiISvzoH25uD6hdUzyby4IB+Q84t+YLBY2
xXvpuqoLTxh7GOVjIYXPjdrRxau7hXtXyCCH6mqNS/L6XPM9VRGyckSIlKR1rxZCDIAqhLiB78V4
ZuoUoqHqmF+yzu0kudx6n6bCuy9Mj4sGdUrVtS6KAweLYasIBJXlUx0jO7+RUxQc1LRxMbRBKfes
TMlAg9Y8DdS/jK3DAdp9vEDU70YeoNA9u8qNuBuHpi2L6W8/NoLSy2+6NukT79TxSn+CO0FaDcj8
k4X6zH7XswfHjsYr4iXjd2QBE1rVl0Y1UpSdUlArIgH0UPiHDGNONbib54rOqassahvmJGhu0Mh1
df/u4JSI4gezcy3vHC99gBgBkshASOKBl+WleVgd+pz3ZHn/CCqazIKtFwHgnG0f7X5SncGtR94e
S2lcm76Hx7i9KETDjrRI5FduO7fqergfXd6YPrZYv2xqlIcg+6W65vMDBb7NvjqAXKplMzD1GIWx
uILWVK4sUxaYEzUolMGV0gBzSO4YZTRSKyfvUUrd32BCXbgP21hNVcK0NkG4MiO7/jTXbd/CetYi
pVSqeh9t6y7rZFyKx7OMfmHi0YAz13JUkkSrHabqNieRJzAimuX6kst35T6N/BzmAejfBwMOgANv
yP7gRbhBhDGRgnLLxyRbdOesyieEgbOrnOFw5ix1z4gTTBKw7D1mLyEG7Numnd/1dcoFQZ5PK2RN
+ua3GyKAbWn5ifgAuqBmATmp1C0NMa/wi2oTqfwhx+I0Veb+WSrd86zNVESXrH53JKadcq7SugpS
OeELLleMCZfapF5CXAJRpYgu56ZCVbcEXtFY/C9YniUAbvq8/IgO7HNajEtEyXbdabjeZCd8TnBE
rgjM1STr96/HQ5FExrjn//WllzqHXikwq1iG0rexjXDDT+rpbrvjO5izCP9PAGHrP3oAC3S6Sftr
jc6lJzYeOUb4Cn9nUEyjHMph5pVieh8WH/OGqed36mWsgAokh8UCRd5SzP5jhKg0SQMIofqLc3kP
aO9UtUYVY+Tiz9stc3Zgc8SbtJPBEiNlk+aID+0Bh65oEg1NB5aFPGnVVCY7/CaGu17LR72BSzyJ
pkT7iGTi1z6tz/XNBhgyIbua3BVeUbS7VYsmTd/JSU9V3/Mg5LHMkh6ndPzCRhOGpbTbD+fEhsbY
EIHKYqKJy5YOGwTH/J8jvAXL6z0uD7Er7j04vUOyHIWToYV1na9Fn5DF/XXbgFNqmUx9/ebEKGsk
0P2RH/ghqXvN6C+/mbfuKkB3zW1S4f4oNYkWNy/g60DcJSDaTYOrlTFHldrYUfGX/X5g1xO0E7qU
K1xkVlSxk3iqCld2iSJERVylylHnEbSiqc2Pn2zg7yXnah3pdTrMkxJjLw4uNh3jl2uvr95DiDJ4
godF634VjsfOHQ/t9bgEXY6L/ZkeBGrdZW2OARnNkdijjxRIrL2P5k41zPrvFzafnJbvxh2PdEgn
/mDZqSOQcabZkvo1h8ks/iZ2pMdVD5PTO8fVzYf6yGMsOkmLYJ11HRNL3YkBNi39Fcj9qNPTGouj
jY2IuUhlsfdQlXII9nXTqMeaKEhH9w+q4z9wRp62mT70NwHOIqaqE4gIQ1VLjpiGSXzKU9pVuydq
qUHDxnz9MwgOtKiBmFiwTNkb0W4nq59nzSE3RUffkRuNHMQr2CW9AbfGuxOKPLY1R3vZEwXs1iNg
vSlBjUuVuvSG1lxq7FjW02BHDWkiSJGWALJSofWmaLZhX+4eb1q+7VgwOI5lbK1AY3FSYijC98qe
ZmKdjM7GlkJG/RSaF9hZRjD7Y17XOFCE1mimULXBoU82U9HoSIzWobjw9Fsd8Z0vWLBTASFnU65z
l72ae2irCYEWnP3m07c0UPlfklCD6/ldKTjUnr0yDsWq8L0Hc2kdqvJNcvsZA+im6CbIMvwCLOWZ
ImDBeWMP8NPeLvBAJGW2HX/ml29wrZ9S77dvR/t+l2jM+KEWj1b6NMDuSSqkxWgYT6OPZQQoAblH
jh8KEFvYgUjv4fL3SBtYZ184UPp2sWjDzPFLaU+8DBki54jQedYRBCuIB6dyg9HbXURM+MbqhQj6
cJSQsPYVpAobUdU7muDxj/fLTSSZANr6p5FIBLy8xUNXO8JLexnBOe2iAvlkrbS4Ycsp5LYvc3iA
qp9+cS9aUcNVFvr1ZDJPG9wz+XYxZ8dHAZ8+DsvwkoYK3vMu8YSXXgeX0WKn8c0cKvtxKD90LkUV
ss2Aw+mpFDsaWk0W19LmkzISuLcSQtkeZBsuU863mgXhLcm7LvAELSRD6TuDu6QK3tEmMl/W1ndk
j7tOu07ziIxtsApqxkIj+NJxbKAnnBMjjEdkrQ+0z1fJUBxWCJbMUTaiJ4BPTYv7MR6ky1NuSkK6
3kFLSO/UV8H19FcjKpxlg9AvA5+CNdmgYBDts9BvMYJkBxRZE7SFlo5+ngyZk6dj5D5mSMfpWmoE
m90jh5dV2BbRcNg+SyEycuDdCzHuHK3USuO3Y9zj4P/h0izKu4UT63Zx0TOudIKnD5sELTE9GgGr
HdtJIR20xO/oSpsRd0xRT9+0WtNw/SZSH5EOmXeiFJFvY9nax+SlA8io5gMbO+F9sWyPGzqZm8tJ
yk/gjIMirYbwxKYSoYShJPJ4MFp5UamkIl+ZsdEGcy1JumadjTMrNRWuAR621sovFzPeM1CSRq3Q
tSK58BAugqD0HYBc8saG7pp0pho0WvTSAG5bhO1By+jx4B/GLn9r5lPU4x7iVUtLYiKFnb54ZTP+
vVeq7zKwPxR8S0NKcfWjOQUV4DO1cKQs3ySia8eyZ1nA8Mb+7fCBJHiGF1fdzLnJj+mABNYtPBte
rk4kvQc4uWIL9fAQqYKAy1RSgoUZ0/s/KkrXLi58Thlf3bU/s45rxXKLYHM2YscNm6VpioXIgC6F
ppM9TMWr8vY3RyKTy8ruLGV2YZG53Z1G+553nU2skG0hhS0l+R4npkrGu5QuRSaHI2WlG0hsaIXd
KXOx/mBMeNt093GN5HIrgNbOHOndKt80t9wWLsB68zdRHrYTHtL1N1jGz2Sd4pod/LdaPrZjcRXh
WJYuctwd1+8lW0WP1lqIoycC+rmPIkMhX1p/qLvMeVR0awZBbTcglcZeSm6igCFyjR27hEA2wA+W
SzBBVPdShcr56kVEniI80ZL8iWe39EEyyG9dYRMvRezbaSI2n+6mjbqaIQngtibQ5QyRJqEMEq6k
cLDBBkY/cRhTwPr4Yps5nZ0SU8fEqNZYk1esEx+d1nezI3QqEykIDZnOEOW7VmNosUyhHXy7oIAT
54u0BCmUOmgGV1XEvUGH/trgJ+/FhtEk6EVmMw5XAU8vMwfqthSWtbHNbZMtoErRy7jBtX+9FDVq
a0IcpxSBj5YWEAApGObPt1OC3bbUl/6TaigjZWLzioHnDewm3NaFqRlBnvH9f6Di2q8uacvNfQOK
SQ145tcv/34V41yNhuAGymwmx8Q8tywZhTcbWw0vFAs+0brvPkVxTSEp8IaPjWDslpXn7yEFIUHE
JXECHrYCJTM06BodE54rD+RjZNBgaY2oFT00SDMuJA17KOmE0gGYXdhpRgVRjxjeV/q2zJp77xs4
aQ/wNfGbg6EHuZsRvJhgEZbmp9qZpUFn127/sheABoIp4ESGuCZeftRIWM04EO4yhSz+oQMMTVc+
6stagFXD0Ol+0bLE+Rct3/reVNsvK9ydjc+aqwnVdP9JbwxnqtbXyeKB8heYoHeyJh6QD/VS5PKg
Qvun3mgreiQMv/wSz3DiXJY6PUWKDM12mf9FdCQwo0mXiYrgL/l3GKoL8tqUw5UT2zb6UQRoWDSH
YErHgEg3FqZohbdJis+DrGRg9mXwGENnrQDdT+VyP1Zo9wYTxhA008A+e0y2Zj1edWKQOrpCDx8B
Jq8bzMHK/CiqVlpj1lId+PurlcvdQdK45/+FRD3Adz5rlhnK+bRRngGkNU1Wmhhh6hBIlWcON7EU
FH3XtolB+dNPVQPySkRdiFFOCAo22mGXhhE9OpuR1Tpzga7flDwecKB2Mp9IhIZQjeLySQ9ZlYI8
sxqEJt/IFKD8Tebi8fanFM073SILaJ/efRydcPEjevs0i728qPwfPPral1Sc9Fd8aAV1g/SUUQ4q
Lku59pAtH/XQdqkPZSqzlJv0IxKyh0UEJ35lFol9NLQLgITX90/fbluQpC+LyOGeeV7+DaUQMHxt
eeZD04+sEbv56OtiCdp+tq5bDbm3cN2XfBX4ObjaIuCN3A6DlsDem0xdKf2eAttgniLRco7JN3oI
Y4QuFQo4oxxcbKc4DJsUFUhHBO28NKjtNXbnPt5L9CcUwbLyEkdCSt5MVGM8oWD3Iqd4tKkWiLL1
X0sJwEeyBSkABU+HKhLnuqax8wMON6m/OwEDRul9upXRcCid/4m5a6byRjrJaiaVHvPVr504WrGZ
ye48Ya3yDJxj9wYhQ5VsVLfaB9kmq05IKxqYDt0lnZeeyvFVGInnLEm3ukvEfdLUka9TxnmNgk8a
Ju2DW5zR5ZiYm4inVmaGs68dnokL85ZZUtxXwldkSiEEth6W6qKa3XGl3PiOk9gsYZlmcXmEYyXN
6qi3ZWRZWacDCS3/838zzG7c6ofNH2UA3JntmOMbqlebv8j84k88SY1YUinde9McpQG/P3TOEZy2
2AAAANRTvcyzrZWAY0i1m/FZWXxk3atI4Z+MeyAR3Ynla7JvqgvMgs3KaUZpXzNI3aEjZ2sKrRET
wSjLqXCV+7keHR88sfjkMU/87QWnPCWSgUvwBfGs4/sPa8UUt7POpmfrY6xQJM/q/CQuuv7I4k4/
c6Ktm7szsl/cCoa7VuDkns2+9ANeFTClWAChmc9ZFdKXp6YAP8nMXJ0jVCT98T+/Zqh/sriZ/SaQ
F6yim+qTd0mcaGkC2A/lHzdjEbNw83uFGfav9FLinTynmwqHLoYc3fFyUm1JAQ0RXmV8FQbjNlNJ
C2g0u9Jb7SiJWTKEez9UCJeX5Ju0WddoC27ox1lUpvltgaeZzNXoyzelsS2CShM2zHN9JHFaLW+4
PINrGCV3bro3u/96MBvneLUwIMCKYbQNEYmbeqTV/mlCNQTkt4pSpszOWeiVY1JFMl1DpsEe7wsZ
w1DrKZEuCLWmkhQWf/GX058lwJH0L1AwxJcU/g8AJa/Nqud35OxjlrmArzoqq/avn28zXxvp7/RE
698U2GlunmwUPAmJuZ+beepMjOx/HgV7c+P4Q5V5gXrRy0U1oMzqn8zovwWx+clRsUFHsqSN0u5Y
uzGo52VJjvpZy4F6bkfj9E8dLrB+cEuBFIjryqI9yKhcBxWKi1Tlm++LkLVSZl3sYTdN8CZ0h5hg
BNTgMEmUfRGOt+lN0oSyTnAalPDCdrSNMDNk6S6oW/racoWYZ+KscSYDT8guF47ToY5TH1X23J3A
7mVdkyp603lKjoxIXk2/uMNlhL57NQ218Jvq2z6p7Yoy08r2zGBkk+Ex2+1yJ5HaDOA+ZUI8ztX1
oI9sQ3b2Lcktf4skdr9vxzGjh7/qDMG10jNOGaP0ImzDfNze1ZksIMM3rcJSnWwXU/RVU0ivcWSG
bgx9eid14fH9Em/kLLsD3TFDN+bbt1rEfngB9ox6rOCgX73qcn92V4rqOgHkENQhUQutj+NfWWdg
Fok/s0MlmZPL/Q4hw14n3IbhWU/pk66yFr5L+NuoqvMVRaZfcfwXBy6Yl3fWEU6epyj3S2l8doqJ
P55OIjya8uWLuuXe2iZWNWdhP2XK/t1Wudw6fDYm2vy3PXYe9f40wS8poDhdYjixPgsTZcr1UEki
k/aH5PL99aUsNMHowkZgxQwE9ZUOkfYdqWlvezo4hLmCibp/wfLVOdDIvgtV6T/s9eROTMlzxG0m
lPVJK5KHbGjKFNO5NeIZv1EXpOASj4ZIlhsWPDHVHbXG5eTv3Ea7rFHf54Fb9fn2rZhkiAV0iD2a
KDbaQWhlUiut2GyXqwC8Yq80f7+Oa+lK/4VU59A15l5+0T13g/fqebp0F8ZsjsFiTAnarWL73fU/
ooPNxKDvSg8EctsEZAgeLgpL8y7IAuvFqIH74B9C6c5dwqeJLI854bMqvm1fEtn8+6KguA49xWU6
8JxtDNVyRRPLyHfimFlJfR9rLYozX4gtcZSvUWeZVePetV3GUAEexPHnhstfRmaG2fNTmlWosW0p
kpzoG1gt7iCKLH1msZyvoMCNYKm8pEeUWktmqwWlV4piJCBjteQ0h5Tr6vR+vFY63jvpyFvakE1J
a0DpiifXNlC7pJY/PCwaGSfmytDgWbKKqdk0VfkiS0THNpXMiMqqvH2b8+1t+0WCwkSQLZqFKrH3
BZ83ZLEGP8558KU7bHxrVcJw7m9tIThRu4Zx/hhiFWAhkP1IQf5rCfgCN7nSfEW96vA4jSscE9nG
i3L3bf5hhZVi2MvYirDu8y435nv9KPEvx4YDUt7vP7dgCk+lWOpppQak90hKqp5d9IK9bLtjf3aX
MXBnv51dEjQzssOcKfgci1i01sKGGvd8VSZWY5g92KUlb+abSwaML1Fe5GzhYuEulfRp3xgjgiPp
oNPyo6BMaz81KaLcNSfneyK2kneEyc2P+7XicGjUM2fOYmfcoaDmxrLDGcDn8osRBCTm6/tFzLSC
oVlpjjJ1iZ2VtDA0jjSjnRzRB0iJ6uJQIgc6Xj5OmuS/ToCYurWj80OK/FzL3o5vRLWr4TazNVWQ
psADT6vHocY1pOqf0fpR9Hqcp21MIjaiTwl85pIt9bZKiXNzU2DLWFhd1Hc9Jd2NIYQ8R3+XbMGf
MBr56Tgxo920Lwga3CMC+ob7lwPkVKJgoZodgwRSEsM32WR4JjNgcF229feifm2SvCbwa7eppr0x
W0SsKpm0hjmdqgyJCp3id3OwwXqcp+9M/KueeRrsYxv+N4mp3JGuncfWIFNTRsM+/GxOtGuejlSW
tGEMLAqXTN4LDgaKUYxdIXX2BIa6iRkc+9toRD1xx8dLlQTMBxP+zOwsDAvh9BC6QJmR24m9Eb1m
pJlXYWyAn9+qKoLbMBSIYE5V2yVZfANqcJFGNDonqt0y6Y07sV7E1o28qjPTf9X/BYICZjS3cp6h
3qqTNSyQFaWOo6epIB98tL2l6fvpQcF6EhNnqY9A7BCrFGe3y1jPmm3mW27o3V6owIYNhcQ6x9WF
m3pFyUQizk/OO50j/2sq2jVd+vNPR28y8cy4XIPLJDBuqLohsqfyh13xpuVT1FIby5qJU6g/stz7
qCCiAmoU4WopVeZj3VaiJH8Z93vrHTxNx1x86LJt8CqKyJ7ND0JXtYDTxEHaNeOI2pa+r0y6RWP4
VhZhTX3HR3+5sznnG6jQrnTtWivxitSsbSrVCqnQWkEGEKKLNLW7K0wHcYU4c/fVL8kU5pMdNWJd
aZCZsosS7+fREsRS1iPyQWzwIyU2tLahL0x4Mmd5o1Ncc9mpal8ObXDyyiZzOIYxAp3Mu8fyQ5ge
YwXiynOwkZVv550+levfdfd34QdwSAhPRyBXa+rrpxWooNZYbMCiUR53NBqAuauYFr7oO/Fh4KyK
RTxPSIa2FP3B831s09wgvgWgovhn4TKPgPHzkaiRfz8Plj6T62gCLahstd1cK7vdm/Zv/lweVVGr
K/cYSonu9coUeh7oGFHplJ6bupSdro52JHTZJbxgARTu5cf3na1L4KpC+BpvuP71Hy6kdgAmm13u
jGnfYVR1LChcm2mdzhL75+23RlpwVH9By4sxQ/RCK3rr0nN+1LS0qKvt/uCUPm6oJ54irL4hEUIE
sYtH/Pv++Fj1kmoiV+NKwAS4AEF7sb/yLDMihyagVV/UryAS3dLLYCljlRNWORgls4EOQf8C8Mo4
GJ2bfhk/HDNkxfOIU9L/7UsKHefuPCHxBw84KAHtSmdnPqiXAeRgfaREd6Iutb81ugZq/vgC8bxR
F6VQqzAXXu67MRMA2Qmbh6RpBf+K6CUCEPzNpI8ezTlVhWKDb3V5pJm3ByvepWo7/odNrFxhAn/g
xFedRSl6+PHEBMkQr3TkA+tpDAMiymb4y4WunSc/llJR+74UmXQAzBoLgFJKOSR/lpadbWB7UXw8
ANT6dCYOP6uRsRX+3GgwZOockQ1hfai65y8Khhkecd4KyEHuhGvT63hY7wSfmhl69ke3zB/ZYwfX
4bIPXmynx3qsBF78dsv/GZUrvuyJ7P92/TNRbK1AcvFplqbp53JUDxwfE2KUFrTeGqhKGB+Jq+fc
RNa2lERreUJ7S/1C68fsfuFRnSHHqfnVuObaGqo7KaSSafaUtLgF5f0gamf6INDHtd0D2ufNiCdm
xF1CkpspZZH7O2U8YG69vT0jWQ6BHNYZgTH+fRCysryerxJa3u9ouMIKIXkOtfDsmEmxPGuOt74i
pUV5VtdTlyu+bOVjWXlUFMVOE74jRUpasxqDlj2Aa7RO0Oh62Y3/Do5DahQ9f4BFdY2A8nYxImTy
YmbY2GdNC7ULlySbDVs5M/lPjUwYfDKu8LkOIX6qQ24cZ5w2fVfki8b8qvETnXHEk118THRFHlHc
u8wWI7PJr+XOe4nPfuklvJoTRBAfzJxIG0Z22ecbSwuyktcm06i5CgHCoJYHpWVUmO4CZo26giQd
6fpkCBQ3fsMd0l1SrYdwHCPEmckvzDw0p9SkX+HGSUYjdMhYrqZ9BzPblYxxGsgWePtHJM+adzA3
HTSPqsQOC5Zvmzm8KVhsb7xKjDY8gwHPePFc7Q7JnToW8ZVKadH8flcFW+VnNbn3i2cktjvFEyaf
uxHKLW+f1tAbP08YMVR8bLxwDLNp+u/KQc3H33VynCE6mB5jrLoNJ5TOW+QileQe3K6QZ4YsjtAj
UwJcQgQkUCJ2nx77pgP1ad6s6JjqfC3gYzcP/3FBMy8yh5Cc1yNd6wbXuBvcKPxZ5o1lKA7e9P7F
fHzR/63R75JQk01d5AIIPgghwnXYiIVZRH34y0PZV8+QO2Y0FAewsp0VBHVdJX3EwPPPIVJrWO0M
6+5I9SFMWGrut//qMk2j9kiD3O80ZjEsofG11Lvo5o9MWVX2QBBtVzF5fEGQkfp1qPcbPAm2LsXf
kVTpcFJV7rjAcjzTbySSqglWJ5ko/SxqZ9j8vwdscU0monMbOMQDGXnvok/3aUbUCFfb/Ha+fxMS
bp7p07mPp3xjr1POjghlS/riON4yUHzqC2Ao3GsAuJFtxwEMZ0Fn0fia1RRiYbePNnIDKBLH3bnA
K6U2sdIpGWT5lPCzZ8AKsoni/fA7oVlhRx2ZDp0HnY1j0ER/K0qf4DTas0GEl0QBm5v4rQjS/DMO
yPK+0jQOclPwKfdHYMPgf6KcRipH5D0Ci1OOPEXZ6zdHD0dxbQW+PbNPLl7FOULSBPO40mygVFHM
pM2q6XPX0hdrasWu+kd/0bcU+I7B9MLuft7ENkcSR29/T60ebV2x0+L7e+vhLMrxTyiGO8pg95pT
ITBFqOAKgAsk6t2FMYzt4QPkaHtA6BgJSK9kprK1dyQy1O/0lTGPKLOt1zmVQxYdaARSKwooV6Lc
XTgoKXcNLlvZ1CW72cncTEKto03o8ZPITgQh831qdkfpGCkPG8F8sC/2WEr3hUv6XN1ElNs0Wqjm
GGDJi0rab0AMZNFFHENDPUeip9GRBsq5uAOPFwpBuEHDNdONjazvxVVUPR50QN3l6xpxySgvo3gW
BvwKZ827RX9MyQwljFZBz8UpJPgPVJvUsGsic0JPt6sBs+9pYdo7z3gYrn42Kqy1WOVyboJxCJBm
QEow7BCzBxExUHO0po1L5Hne+J6j6trFg9QNWVTPyQvD0drcEWJ9Ho+instIBH6Ofj74C2FzHCx1
XW43ILgg9wzVGjcEoVyXP5qNpZxe3CbylUJfNpKABwvhcaXbX/auh0XPSW4fbzqKt01+7hFVns/b
ek2ByoLbJGSAJC+WaO8HT1SI25/iCWbUqcGHaHHoXn0aqy/SDjXOywCnLxk7X0NFgnE49VFyUu/l
MVNHYKiecOg5JG6/Um5W0oRNA8kW1IBChcI5sl3ccRWmsHY3dU5ZE6v4nst7vmA8RwzGAdiHvgQy
9mt404RN+rShxcpVkMDsVbawBohBHkuDQWBzepEsG2hEa9jZ+TKllawXpZn2d/oNDtCvsJjTMUbA
d3uAerRpmOGHVJeMig0oWkynpqjmZq1U3jZBFtq4oMwKEqqYra+5lrhaR7/ipz69ALKmHhoaRRcp
gKsBXhFAJTExr4sx1+e7Bjmq7tOjo9HUQp+VOTc6dxBAMqXSMjlwZQl3RWluPr9BiVz9RJvUTeAX
lfRmqX4KcSmbWbMwoFjv570/65F9jsBkfVYuXTuc7ej2SVekrCyFoWZx0oMcv02hIOp784oqKb+x
yeQU6kp+QRRQGPMpX4prFL7rttNvx6oIrXa64GRQ0a8GNtZaM+SbMKHqFPytiNYZRh1niPqilXwP
HfWmBJi2kbHlyFAx/QKQvmq3KDgBkP2T5UzjGCmcFMQPvkd9sNwUsSv/LjyXkBz/JUg10N27H1W5
6ZMelbOzk92kYdQr1lKxl0oU8r9/pOq4+lGtOTdl5YTPCvrwDdOwbWW2+1e+kUlMgQ8BLEIveLxL
hXuJBE2HPuadu80KhnjxGgVuZ+OqUaP8DVo1rRd8fYQPMv4ew1gYqIA2Vqq0vhdk1bI9lYz4b3Ae
Ns3t4srReUEe7kuTmv8fe0Nc1s61KarYBx4c0a/EULAqSAgUmRHcYAFiHxsi94dIycR9YA7GMv1D
UoEndbzxPlcpxNPAuGJGBA850zcQJZ3fJJIwS27adFkM4zO+9xL6LGt2D4VgBiCg0VCXTi9vBxu5
YB4nbaLeY46gZTopeIxMLk+xx1RTn2ewIK/Z2RsFvJF+tsJ8aljz6gFPLb39EQGXjVPxNE7h/+rg
1ZYGXs2G+hH3q9QpRPcCVb141WW/2kzqUDDsV52AADqK1PeB+O306TEV4FHuy+MHV9GGTlx20pLs
imzj4ncz5hMRF9bYUSvjMWEPf4aUKP6s8f4qKELdIudl+dGY5m8yhiL1hyMnHiywoIP/wo1KYHcF
olEEYtktlF+JUppOQwfMQLo/DCaWL+29sQMaHhsS+kZtHsdHhr6BO/ZzjVvNbtKhCDk6Q9eENZfX
YMX9sIMVI8UsuQMJUop+ZDA/c4QiK1JxNsr23FRHsdsYCrrG7sn3RX9UJ38vnjvb/A+o7u/awjri
i6uNBd1cLRRDTJf7OyybXBKeznVkF0OKdAIQ19PA33c15IM/lXo6mhRqm6wISVsh8xISHmCSLTGZ
pb20Zkeignx0DhDOnKQnyOJW8rZheK8OwVe1q3p9Sznvmc+S330ys9ql6+w9Ksp8OYdPW6Hg40xN
Bh462fUahWgK6y95M7VhyD2hYYTsaZBsIvdLI4tGhLPycx3LPnyXWEMf6CO1lFW5h5HXzXJ7Y1ml
cFtnVZs0NRKcdlTPK1bMeofQh7mQVbDtTEnZz9Og+e2saVtypHXI+MORf/ebs9q0LdDtaKAN7rgE
k7vPpq4aOG/r0Amv0j6nhgHft3xH/qwSGymHgccvsDey9Bk3ySs+gukeMsXSM8wcvonlsW1aSkRh
ogHan6CwjO/CLTC8ilQFlKt/cvrv88LjJQDK3O4MvG1uuY19Jv//zqIh8BFAka8d3GemWkKjZJF4
RGscSphzSJ8I3jcnbz1ZagOsXImg7QEOxO7bGc+1l/bpzNHIvyuHSrRLv6rJytXQdCcdNCqEn04K
9USdXrvllb13MVEX7xIO55DMq3BkjsjwZKTPkq0cbifqtfOKFeFQ7o1YKGbvRLKXK6BI44gWQBAv
+uW3RZ+w7I2F9mSzEk9JclfjxIuRViFyngCPcSUIvVif/zY/x5erp/Rn8NXW14KQxh06YsX1gh2O
RuMDw+IS+5EsuROkhuYtQ4Il5+cTR/8L9LK1mcCE7ZrGbOzEnIoDy1JcgD3EIyHIEe6BXbzV5K4H
dNrLDmIusYn8yfoD4ciL4GUA+D+/wYeqVxvfM4tB06Kz/rnd8IGxu3XoWEJRjFvuHC9J0wF2QlYI
wXW6+jbCVyKNBZZUl+oOIOUp6UOP4nxkrr58qodk0DS6WH08qMueUKEB4gBY73JAwGCeNNRtCDrY
mnAnxyNQh3aDtHIiPRKV3qJuEr1Aucg8qJAULxWY8eIhrxRNHl4/RuICIaqqw0qdYG7xCKgM3N8y
Wt+EmM5JTbOzDYCpLnUazRaWgCetq41r6L7B7F+891zmKyEKFda3ybQoUqx2bnqrudLqnvfbihZv
G+5s0yma3VTelFu0i0D+2yE04SfJFLzrcRLN8VCpoMnltAFH8dS2SJ/qkKy8KjJGp3DOhH9kNRZr
DEJP/YAGXahkicXt1v1hxOaNbnX8DId54eK5ctM5UVfzAA6nqY4jVa/WFsJHG83hD2TVM3l5K3Jg
Xd6l8daHbmHfErHkd58qkHOl6vPz1rvxF/DSXHDh2xiaflFh31oWkD8/u8G17eqOuW/OaKMEDUIi
mLrW4q+vFWm44vYxVMlzRzIzmd78YsZEXDvbli6QpoamACfRtwsoRRBCeRXN6l2kO9K8mhBMEQw3
ZLtJBq8NYsQGzjOjDkA91UWwX+xxHiNbr9owRfmFnMQs57oul0V5YyX3YBA4p6pu2tYvlbeVSL7y
QlOfv3Xji7jTBhcQaAwsrqSY1vMo9EvKfKkgfgL30p53B50wgd5T2cLehhSx82u4Z8rPVoIjun+l
LSS7FI0O8sgkdC521ME+gvfuZi0WGrGRLRtwnGyFvwqakL1FzuOxQkrqHrXQo1JXa8aRUOTzVks+
EvNbtHsngbQRzwH1Ug6ebAoyVkgNH4XefduUtr5i/e8+S616hLFLDuImLBits6o5yAYfN+UVc96R
JpqBN8CpxUi3Lmiw0TTxD3Byzc5Jx1eNgQefGZiDK4QdhU5KOtcmPbKwBg8tLN+p8Ht+qFLetPJx
X36mdiy1tRtQyOGwIn5hgH54XXyUpbWtUsFpZ07um+x/HdBCOKsd0DWdm+RpRuUUiT4jdobya2Mv
mT7RwHS4TKfdykI7JfkVDPiO9B7kB+SL9Ogkc6kE3/g8efMmytz2ToJ2vAhr2l+qX81Jzoaq3KLk
ubMadFj1RnvUJGHIw4mFSxliRLaPDhpZn/XjmNbwazJKv1Y3aCzfCkAMgs7KdNXU6qYYWKB5HUJC
aPSem9XfPYA96gqRfwFlf2a+t/kzyj4gq76Hc1Gl/wKTO8CLVVK69aKWlmuLrr4r0DscT70saWlc
AQq2TbNZDbnidbmtG6G3wBFRtovhITpouA3rpb/7ONiPrxaqWcpNazCN8/ufVGR6x9JqKv3WQQ4s
aWc8+7ha0RRH/xMj5DgTezwRp+x2rg2laKzJHk3wDLEiVjGhIA0OIcjqcmHJFK9GasR9O6QBgIB7
8TSe2pUiAQWreKGdk7XckrOnAOUQGtUTLMiyYpcXEiW5SfnT0c3BaIa1Akcf3jeBMXxpZGQEn9xb
VaC+SZvxXvYnd4cdayr0Nfz/2vKezEoXRSFjeRUevk2pfcqP87egN/ptWJqPlG5vV+rXyczm+eRE
qxGt19U1CF48vAkOe+M+92WsIOFcDav2K7g7W6sQPVVGs70buyEZqUpCL0RzbFGRATBYCujxjHD7
77vKRCWV/5K/OdZtFTBrAbZ4QYsipn04uUPYnD5b76HTbTt5Wa53yso3Wzzz+sY9rh0ckaaGUJW1
Y0xB9Tg+tLtbRkaFcL735b91qcStlnAedTSwEQxwu/gvip1VcVy2XpN+1IlHkCoiqoB7WnQgu/uO
uY6nrl5ETt9ud3m4ecyxTWrkcE8Jkx/IzJaq6Tv3zIgvjohLIOU66dd5+QpLzyPmFmKlFb4qGGTG
sMsKnZ82HMcudWJ/IuzYJusUPjXXEd/7jpWVl2cYWmXcL1z+IfRqrmKxID4oBwen7H3LYGUy17OB
uNNU6q873wE6WGIQfrfofAvhJJyjEm+AAs8JEFETJmn3mvGcwb7DIHTILtz/3rhtXiXnrSqn86pO
z/njSfM9J/4N1FYeTyzrOhhANVEpzx468TlU3rUWtyX0fnEb0lo+dy3uSlSRG0TqeLqLvSRTQAcF
UlF4/GIEPJJ+5sGRol2kVFPROrZrMQPMcCBE2jqKI4WPcsIvMSGRHWR9Mxlx52RZBYjSZL1X2eLz
/GiZqDrZmjJ6QSFzpcDd5tbCmGVXPLonSvt1p7/Ktu7v9IYz943CRR0com7edc3dC34/ahkeKnku
g23oreU5DAcoNpDfvNidxoZFWE4Ov9cTqnWxg/sloxbqVSwqm8klG9v2Hn98vsHZKwSerCO0hWXb
SNYWBfjZcwCdP5k6E2L3MUqnMS/UQsjgN2klRtfjnHgGdDvAql0nRJX58p9aHCIW5Bw1MUGmC7US
g9LsEhyKKnZHpFYFqehPCMvXodHYsT5WG7sB/pjkCCFGz3bGNk5zYmd6QjClSdLexRPKAiYzRmTd
IKDUs3rXg/5Y5OZ8vFyRzfrDQuLCwe9f0lWI8rmvOyqUnWx00MpqgK/NjypcniRv6uiGBiPADqiK
TuaTiatBCPequ3s/ph01X6GZ/bAvuNk59rjqvht1W8NWWLIFYtn9auwC0DsOoILc65jAvIpLZ3hb
nhgji9/lZYOt0I/YWKh4k7BRGyqWBQNwtgLw/0a6zMtzCnqcBTkQyi5uevyhDfdFjBxaCQ3sOdWr
+wwt+rMuFhdCf4PRdmDjkgSOnnszwe7QLhOCyUZaKuMFmudi19+zps4MxAWksk8dK0pVDWDrNwub
5aKXDn1WHU/7+8FzJGuwFIIAhU3jt5T4aEiITztpgHsJnrE2eO9IHgm3eKYqQdZORI40dxZ67Qmr
MeSsXXmcdWoNJtUpEgE9fztvS+wCM0YRGBHEdloVa+uKg0uzF34qRXPJGtVnYurDJfsMsaJA8M0U
UkAE+FraRhjURODT+41NvEOg9rBL3UDlXdcAUaGwl+O67SQCDY18Z6mQ1iX+50gc+mTiKVETolLj
rDANdgMndymRHVJKQM6UL77KqydCcICDFcv4vpEx6cn6WV8ffpl1Kt0uWyVdgCgCKk91TIwUekea
WkFq7lIoukxnA0M7K6HNgjhK5pPg8fRZ30iSa5MRTewagOYa+Ee3wlZbuc/0XfjxOlIj01CAvefO
+XKbjmlvtqdegZfytHO8I5FwD2q/V5wQJYrFbJCfhWXawf6fjpR+IbrldPA5vUVykH+Wj2RIZj3L
g4S6Kr9S53lNN2VRF9+8gWWA9XHkcvimYUsIp7mUOobNuaKkeKjbzCCNa2huLk4DVfxLS5qDFPFv
24TQ6x3x/c4N26eOoj3PXSklGXZDejA4jT4QGb2KuEXin4zG3Fw8/docHvri90d12s1ZllGilqve
Er5oZy4VKcyGBsL0DZDF7XH7wIqOMfiCNzlnZravrbeKNh0GkESPUj5Qlq87hnJW9nB88vqdqgKt
FleiqM/mqrnTgMj5lxwnJHez2k+TteSccIjrgZzMxnYs/WBpLjcKrLKAHOhrPERG6UmZnlTjM4G+
TbXfoCm5w6sN64mAO/gzi5fKur3KwnUUnoCa/RlMGTSR2LVxumsG1W7zFd7tpWAHC5ypd9/7Tiun
jy5c/g7UGpKq0o8Cyxo8bUAtYyWJfDd6ftUJSczl9VTn2FK2I58AfAfahEExCKLs797nfJANAo5C
UdY2FweCIZioE3pnZCtSc/QAkfbW3ZBH3QaIvb1Bg8k33bCzYvqrJSEbB8auED9mwP/MyPzurOAf
a7+5EPZIk3t8v87GWE5L4zt8d0grZ68EUNfmFG8ojxGN3nZVpCG2ezbwQXtwHLmwW+sHMWAgENbA
DDLitqMfNXkVTC1Vba81NvIbtRDSXYVaXsk184ddsL2cjz5DMmslvR1uUl94DIf9b10M5Z0kbDsl
h7uLwlHTzxYXC/XdbJgOzL+3bdPbhOD1lmuRCL1fREcWanw1Oth1vPSOw8Xuoqp+hwXClm9MK3fD
jSaK5gbs6cp8j3Ldag1AoqQiJ4KJ7QN4s+kYLHMZUYCKyJ31KU23ulEAJVkpkMZho1CPY+zEkfgG
e/z52NNiCr3QW0z4fbS4BtxIfOLTrd13p9v3ks0mU4SRSVW2NSjG2I+QD0gopb/dNwo6nyFwQTpw
1Zq7WnYHBG5WTN8lreA4aYU6iKdPSsqcV3ZjUm22g4Hk8+keKN4bfFGSobzeaU2OSoCZYt94ym8P
lMgQFlxNT5/cREsKWrZ5dTlqZR4Ugw7R55Q3l6eL8ZcxIhKN7iQK2xbAECEHbgPMf0J3YBoAK/AY
B3UDFJ8Lzxe8TiHGLYKcC0cIREL/A2/tRSmlSoWsfMTqFpFCoXT23AQGkw15XYOWPavcED0aRqZj
EjfPgLP1zItdS9sQmw9kMU+IpcwRFCdSMeplk1KXHxQgu2A5nqPFf3ZWKa22pgtf0CyS1Fj9TXOh
RwoMwCLaCQlGIFut89Kob2iEZuLnh+jlUD1aGjHj95bSo39qLUHI6uB3LK2DhJidrgFFKN807rBY
VvXAo7ErcWWInU7yka7AaaWk+CCL1af8VunjBWWNFINdmTZEZQCbXN9he1At3HoyPYzHzmvQDAUj
JvK4Bpcl6mkisRiLCwskLiXUL8HBTStTOeS3A+atHbQuihQ4v4XURPiKo4l+ftxTv7Le9FnTi76c
nHhx16/5u/1dCl5nE5v+FITjnOKb/2biQ/+iW3Hp4eS+ZNXYpxkHGOIE8hRASaZ6D9Pns+y5u12t
5dyOe6Cpm9mu+isxTJ+z292aYyT9h6JsFZ7c+WxEcgXvgh+NF4oCeZyVizuVA7z9poMA+fu9vWNE
bxdVkIxrBQObtEvk/wy3AU+UMm5t8rrmhcBzJJmh6yOjZkXO3eGmMgDKp4cUSBOqUQieORWiWJLG
xC0/eza3yUmXA5ts+0aoV0iAId5yYVeq42OWCB9QXLwGdPJWJTXFQmm62dp4m7v+ZVQyZzUA9nUY
awjLru3fLTltvWkA/L0ZXJd2/O7vVW99k7yYgu1dtvljYKrp6xm3Ic3fIn+B7jBNx/RqcfaUKqHl
Ei2LafEanqO6x2zjbI/3qvAE/Z8HqAARVBiBb0oiD3W5+8NKErofZbqc1HZrHvHosHjaI8zhWSJH
8QIC0JSw/x5UAl0tjd4pzhXCR+2ru0SICpm1yqDoBGv5bRFINDjkmSv5OMjc4cLVqOfo2Cox4I7o
EO8rLkUNv9KMiyyLaYNDOhomeiIMMDmJUf3hSd8fiwVpH3kuoZeyB+M45DWLd1EsqW7v3B+KJvN/
Wkw0TRIx7e49t1cPfZGh2rr8uI8sWJwBCyOGQjnX3W2aSxEWku0VYQQV3fP+Ata3jsjdJvN4WPb1
HCjN2T+xxFEmvHWcDU33+n7iyrnaCIAaYcm57FTwr2nB3QS9nJecEKJXbdS1LeCSjxaCzh+vI7iU
NMIgX+6j/bsLNohogDHlcL+2263l39Qx60uhXGXGJYteSrqQPAEvMKWb4hto4IAEFHjlbPOdUz+K
e6wJO4p6XJErwhjiZPrEWrUqnuSO94xobIN+Sq1PDwv04WcK1ldmZk+rqMHJjpVsK6uoC4xSb9xb
ngF+RrImpjt5DXSYwS8TGfS9Qhx3hQKnyhANTmVw1Cl/KIJbyFmATIIhBLBgs93n/sDjM+MDjTPr
4lnLcecEt3EVzSESOX6UtGL8PAMD0K92jQPNfU9bkDR2mIqb2gg2vZgDMvdhiNOR4dNWy488PyYh
HQ981Wp6U4yQb0TEoBaeYpr0+Cp9Mo4MIxe5QU/oWgdD0r12dwnHlOPMHNIZknANmM8+Xh1Uv9Gs
9MZfmCssPwXHneaS96JSOJOQI4OE7uBApiksjssi1nyW8BxmnmhbEtGUs4bWAT0nlnUxV26RH6p3
Ll3mQThKShA2UlxBc+yUsL5NJsRBcatuaI1zQVTW47pV1B+P3QKTYWFzot7HjWIN+vPtwpe6yd5F
77/K3uv/Vgt9zZVKx9CNGyyKaNP8DpFZU5eB2Nj/1xkNRwV183iyO6j2QIKn8KGjjwiWVNj1yCsp
bPDxwzsj5bX4qODfZznN01yE2UgdgLWYsGgRyvUmvRbFG/LA3oLXdOFZQsT10/OEYY3cCQ2ANB00
iSBxhhqKT6gtacEYl1GO3cvJHSMN51B1riYIPO6MwsFK+hoiS99H/C4cch8di2H6AVMHFXisZnfp
0SA3l+Y9vO5z4RTWHACCf6EIjTbt+Pz2i81QOHeLsxYxlbm5Ui8i5kLBFcgcV1DykG0zJHdL+OUA
Y/zweUDM+GpFD8iD30T5iABbl5hS/x/wYC6KvCjoMm9lnOwZCilPr0X0tc/i5wIRVSTPZhqcoqxA
8WfcZXtCvFhHdi5WHZmTfMXrIbIUTbXLeXb7XNAWrFANyz7jXgv6s/su24rRNLgXONS/XxSEvqQR
C3MvVNU+RImDi95EZeXaC+5B+tBt4yilXITmBtzvCL6auSyeQ12yAs4ticb/VFD/XH8d7WS3uJua
VDtZAGYKAQfZ5RttdZ1P4nJnFXRCF4S1A2yb1LiFrFh5ZhIWEh5XNCSrHA2IUR1dPp5j3TIPkXlE
Ca1+ZJquJ9OOCRU96jKvq09keuZH1At5K+g+DiI73beoe5EmhFniWGtcZWsWaV2zi5ttPSAW1rP5
IwuR86Ujk/Fv6Bxlp8rBy8MAFBz958WGLkY+jeuaoqxXP+n7D2sP9UJh/hwVeem4qHkf6RCc3bfg
n9hqQMmCSmxOI37ijvmc38mfwidpVtUZXhCar3+aAOV0DZpDj+B4CTzO91bcX7s66JlmzbspF+N4
D0tHGvAP+ya9OTiAVTjSADTEB6jTpbv1WeYloTAOudoo0dDQoKt7dIDOo1/OhyzETcZWTNEFVbx8
zITzbCVXmj9gLUBEokx4xxXKA7aX/cIWQDu6LJudT29hLZsKu1nRiWiCh7s6xXf6RgKeOHlU+e4k
8FFs7qZmpKn6Wzt2Jq249bHds5KzQbqmk6lYcYgHl2xgsn0ElxJm/dMw3nS8tn2/7yZIfFxuBHR3
WphJe3b30E8JG8AVgK+qN3X0APzWDTaug088zEGns9UJNvUDGDfJXMhvVauO+MXHjNFAdD0yP0cW
Fin/AGQjx9ZzIwah1BX9KgxQDR+6n909K0edStLMHSexsfIumZdQqUr3a7NDJ7ejq1642YNE31Dd
xz8fDJfflL1lpQiO2N/AOwBSX28cPOz2/jI1bZla81Ixni9GuiyPSIWOLpTS2wCrwlAbnZXbwFNz
rfq+IJNecxKf/VOXLxGlwxRpSF23yhZNZOoQriM/qf+qSkx2EyghzKkJaNQHAn2RdUOG/9gkSerE
XSEvRoV4reuwPdaz0ZdA+LZdi98c5EJT3CzNQzqJGYNHqsCbqdW+xmDdqa6W35pNxN1nCSN9jvwz
WBjeIG+NRrs/sVBBEkgfqfN8fX58ahJKg31jU84lgajwtn/pXpbV3jLF1zfVTf5vGKPRzfvuYCaF
+wfjNlnk7qncv6pT63AYbyJzo5Zjb3KCkiSfUGZirqlsEk2gjoAmysH6osmApdROIRW1qFvhxJx/
xfVLR35/ZALT/Y9zlg9VOT4aTrgUeMKlEuFJykxh/KDTatmHN2gRLMc9Wn1df0yvvmJPVt7iBVU5
L3EKrKAE6MkBZEPtFF3B6zNp2otbxyDe0rmLLOQ8yRJh2ZFJ3XRmo9VO2yVrxBIVGlwaJJ29fgRa
uAYUsALuEZSZTyPybLwI56fT7leMPGYWFDXyUORF9UUUd/qKBhLm9mXyRVUT+2k5xZCtN3YLsl4B
YfeN09DFSggx2x64VEd/nYLYEmAYEoA0z5oS9JjyyQ/K67HS+n5Q6tlAHcOco8DB9pDOGN3xeqWq
Ym38s5PTpQHIrbHYD858sfZwQ61LRDRrPQ1iruhsKfTA61P0RFBwI36r11s+aVhzPWrA66U2qKQP
UgdOF+RhBirDzOdvsqJPpVj19ZfvjOmlhTjQyukqDnrLj/FTIbHMSJOwdlZegvqbSLbppayJt0eV
+3uBiicQ+y4TitrYO5Ny+LBd11hfw9xUtpyfIeExNdXE2E19w/qgRe7uboNEKAu0uC4WEe6mRDx6
PueeSxW7Zj4qoJSF8oaQqsgcVbUOw2JoXaqf1eQbBoTTdN/WxlBIC5GMuKUkwp3dXKgSDcisOEOW
IUW0s6e0iTU1dHKnyRcNbI0KU6KaDhMjN067t9Ckbabnu2BSXCKUNoieQTmRV/DZaWK7DHLzM17l
ZTRc/XRkZOctx6LXrLERpDFf5R4sVndJYjLY4ErufbN54E1UYAcp1bLEY2aACtqQWPHO4xWxDU7g
QnZ6To5TTMWroscf0Ul10aC+tENmtgab+hZJf4dlki1E8tSSoZ+e2QX/HS7UaFPmS8aqljmpQbWa
nL6kVs4Dt+cwv/r9rYCZa6yc/umHOFXvuEb9Du8ToHTtKjTfuXI1OoZXdIcO+2gGZbiElme6VjzQ
RopS8U/VF5L5KgVPCwdgm+C2zFdRq+xM9w+31K88ycRv5v4foeGeHon2U7fMHLHfO462J2bnGnw6
/yRQ+NSSactY+g8OV7fypIopEHvKYWwUKe9Fh/IwseZivmrtJKdOrFYH5wto0aCcmFRk8/N8Ddm7
kFtROtSLMHyGDrpmW3I9RRL8w2BM6A2G4BbxjelZzm2/aS49Dhe9mAN5PKj8xYGNsrTqviwDnrAJ
YLHHEiys63TUmiZ5bS6bv8DctlbvVCOQAEnE5UDjER5prt3ldgC3/LAaJU33RfZwZuvkwFSdNV9E
hsTawl+GY6Ti3E7xwSfMC6uEdSCt4Lu7v5NPE2Tyzk/wc/5P1ln16GTGweyUQhcPcE4Pp9W4JjpX
uqGheSEDsAvGQmv6FxK4I1jL3RrgSWzWobDfE8S4O2QyKVqATXOxkSoJAQ2gE1FZHRF9VS02leNn
IEvFnlcV/7N4mnL22987Oab7FFjlFrX56Y8HBa+2BRRRkJ9ee8Xe/rqDzS4LthoTYvS7uHpJgYFW
MEeBTXrsYIXvjxl+6WdV5vhQ5ajZijfvjcnEl63eBcpJn9cWQhxPxX+S2UBn47LdqWviWFcct0WZ
xdV2vkPy/Mq2vDqKqlIfymkh+pXqKdMtvdUxIOAa6lIe9keUKg8oClEMK7bTeRxxu+JAzAmI7Yvy
I7q64V9Aaog8zgewuzSkiD044G6Ks7Ws5NHyTAA8n2OYCsmtL3z8szK5q0oxfTi//LxWP4mZFIZg
RORx34yCX1WLb1gvCPyDUvYpAjmVXcmxqThYpXVKifrZ+Q3GMXhR8F8/SmuujLWR3gDVEiWht1SW
RcCfVp4z7F15RhJ5wEHT4oS4LI3U1jKg3y7pdA3gvNSQFuUZlU5vfwZeHmGE1nW5Qxnpkm5V4WNX
0qRRSeqrEmbNuGXIgOJPhVq3shKZY761bL7cbOJcrtAVhlqUWFCkQftD6S4cewM/HQwFPX5bNY0O
fFqrRhv9gHeWZdymMKsTkqL10fEIgIYjoE+qJc2eYCsRlXIhCX89r4tsHXI19O97CsiXbGFImHWI
zhkmnwnUyatjwiaGFesmKo45CLRHkM2FOb+9t7sUwbiC04NzEyKf2mst6Xkwb6FBA3EiqUGiT/6p
iPj9aQWMWSIHSCg63boFuQneyyugulhltzpCNxhj3LrqUD1+2Se6gy6hsvwGp0Sm3Vbreh0foaBF
zW0Af5Ogv7v/PVZpbaL7v/Pc7tXuuOwGvue2qVkvZUjaM3FnQBICbRaF4iglDYFug8IRjT2rqbnO
J7khq+lLm12VdfVs5XOcUR/mujs2m0eS0EwWCt57q0CHrYBPe51cOTT9btNA9dUidXZqDFhUGVnw
9OTDwypBCQY0uXvXmF9WSYoY+9zrUIUqXShmWa8obRug1OAxedNZcwm8+H/FfpK/m97LgcwC0yWk
wULKSa9OSXz2TIGNBKdIlTbcJJgG6zeEH2s4wpQFq/s9ucNsUYfhcYvYKZu0qTWnmf6O+SQoxdU2
gqHl/yywuA85JRiAeq4bvZ+VdhShs/JR70qMlaLRJXGYvtQwiLlzW3kc2lhLabw39hCAOndZak2H
eYcee4YoP4ywbgmkc5CzJaNOPQ7thi/4LyE8ZW8WP2sMtZpjgKwo61ONmNXd9PthzI0EaxDGPVFk
wH6vuDR31XdCJOnJoca8hgqcSG4/lc769su1icZIDIkBa+YFfjF3RMqNK8ODJ0J3RKlDdzw3r+Ei
km6Vdqox/AbgpEldQv/+B2DlkIWC8+PmHTRujiW4oRLABtPTyYSWwWCd57U3uzGkq5l1vDrIlH29
K/Sg399NsfUqyzGW4ZBP/Q4KHAQ3MsLGpGp6+/3R8qW3IwGNuK2ger/6YqAmLXwqBbVcsf2T/o+A
/j+cJvAiNfylZCgxEH++LsyIRB3PL1Knt2QXNIY2DFgP+IuhKcdregbgK8sCeLp4vBPThBCSUhEj
tkscyYb9O/BNm0cBICkyUnxe714Epw79J2i+Iz7WbgyoAOu86Er6jBZTEPT3BL1Efhp0WerF92Tr
/D7DHVEWkvAwoBd1YlUynU4cu8ewav8SmDNpoY+9ldmjLAu48wIsnyiOoX2izD5QRkjHjZZ6/pID
gki/yvX8spvq6JYpEKiL6quMGPuppUYMkfkoZST4wqOzMKyXOUANdgpD0diODuKoa/gpW38JQit+
YqzjrWVd12n6kXYjAKpFq+k8j66gUm6B3Rq+9ut/4w+cSeh1yRzuXGiba9wsSdRem74HN2uIGUCS
i5/RpFoeMy199FVL114Nn+Z06ppa/RhP8ovqWDpY7j1th+U6VIn+EWWA8qWdcOVtvO6QuJ8qTrWi
OYJPwBwzNC0Uyz0ewqXWprPq90QcpNZrAEBH5hVwyaxr8zFIMDG9/y7s1PkykjWuJwUTT4sC/MMI
3ssWuIWJBudE/7TpDB8R69FVFJWg9UxrjaAqsH1xpnQ9zJBPVqPjZOlv8CPGPqv0pOgGZ4DXhjQU
4+xgpGw1x+2rn0JO8WfY/M8OhoF7SAg5HwOwhsuIOV8dEwfbmmuUcjmQQPgCYKXGvaIFl3iMo6/3
iuD1ivSjJTILqsEY+46o+wUXCnrB/KaFp4POYSsJEmchYL06VYf101KCuVpJFiJ31uNoBqU2h7CW
mjCz2i6sLTbfXtAK1GbSHr2PtVb7/v/Q/PnLzMAVR9aY/LOWSKB/4b1M8g5XT6bM9n8JO+wTJurF
14aF1RUYcopOEQt6Ni9C9MOUmg3VJ7QGYxGD84jqtyZiNf7wCaxRJ/11TftaQw60TKvyyvILDwyC
jJFBtSHAwtZzPch03LnW8Y1gNhcL1S3M2oMr6SVKHw6UgVh97mNfj6dhTHkG0IrNvI5OkWeSUfOz
DUQnADucxGw+UcMcAbUWwWUOPsKGySzgCkGY20lt4DJyh8ej3LiK4+p6YzKER6Btg4F6a7mJCeaO
mOnOASYgzcIksx1q818yWAR2isKXhZCD/f4iKaE9CgJAuT5Nl0e/BgsWy063PanJXhsTMW9GO+Dr
NEnNOuizgid/dKTWGamNl7X6YrVjzt4oMpVDWmJSOMqc11U3CwjbX6wrik0bLdoI9GOaMPBoiz1A
i2eNRJwbM+gwGrjVoVETaoyaTaK11yi/ZKNLlxrFuzKBtBByXa+wDf7MjjZ9zCpC88Xnsu5OVopY
BOS2lSfmjaqPUM+VJHSbbIH5lB/+iK3uPhq+EXYiUUOZHBmsKwZjdDqUp2tkz7ezMF6znygl/eln
xfsuIxWTSOoXIdtNNNN2YJX3/Qu+zPGxOyY1Y9e0g8lg5TNWg0HB3Hw8xzKAsT0IbuqSfiNASXLV
WdGVpnBml7kN5CDUpkHjVWNPkZdkUXnH6Zb5vcYROkFkbK04c9VbnQ40F5yuJ8Z5oiNvXKDAtdHF
qSW++zvX4BRNZWMeh7wQDPTVbi1wAYzWVjnHXnVh5ArW8E+MyO4IpXiGzY2qYb/RuMOKETtGv2Gf
FPEtsHr+jWibs3twOGLo3BtT4FgkxLGOgqszJB4UXj5KLqatMBcdTK2VPFYKMVWlx+HDObcZvCP8
S0/Y0G2dYY94PVavQSupMUcU7HuNAwZsLv1ZXTb52aLsyPIgpuiRzGOW4Njw1mVBzGoh9qBodTpG
nR9KcCmig0D59ZsI0LzQB/xt4o/7PMKUpYtiuiF9f1VPNiGHZxLrBC490HcySkmuNuSdDHOglxxI
Sz9pzSMnmP9xSHKsDXC81/akx6mwCnLQkMm+xwUikkSjAZImZEI9DbMWGcdXQHiwfWFbOEngnyhL
k0fbBpwU54w+5RYtkmgoWMqAtnIeoIqlF349A9Isg5SWPDSPtN5BLx+9FrBmAbFjVtOtpoEOgq79
OwEmUB+ODFov3EMTmY5Ldqeb3LRpuZCciqXXluawH8ursdqUL7+vr+QB5cTT30rF30/JVGUYV+Tn
4c1dW0gSJ5zdbxUHICA2cCJtEjlKsTQJF1FYtKtiD8pcM/Aj9D99B4XmIe6E3vcXy71dKJvRaVm3
+bGlTcS1oWcnCOqg3njrlv3NTcnlMuX3lrQtOB//tV5nqq7vrhrO1eCQcCqvQ90QB8J3dN7tXTJU
YBY8iqR99Rnzp7PiGUFhyBqlY56FlCrrLQanwYuQsdeHZzPMqdiI4uQR3tVXozbRtmYdYQGLmSN/
FMdbz2C+qAG1BPdX39UY+Mb00HnFx1u+OhXv67E3/4DrkAVldYXtAl+AywaZ6/ucw63paSzEK7jT
+EzH29Wtr/OQGiy318WiQYU/B1DBmLTjuR4Iw13lCe0ba+1Bh3kuX91I9zPZleLOHTp2ohDYBw0W
4SybZjH4AXhSXXNu6v34lWp0SjGp5indt1rCxFMsalB8GNjm36V2YYOBcZupm9t6TmW2yWaAA6UI
kSG3VN6TnTA+KyDsrJu9dsTYJc8UPNPK8uQtR26FGuCJJosii6N2zs1ejUb8H+wQ1ODjg9JY+WdA
O23NnwnLh+zWmCWGp/fMs0NX8HOUxBE60hDzsZokCknYzIID9Try4f7EZjaEF0BYzzfnYUrOvejC
DiWodi9kkUFsGaO/Svddc+0jLcOHZkyKyprz1KQpSsR5RWoNGfIO1GjkW3tPXlkIdqvkBMyVYxHX
9qEqH/I4AeKRu+ad3cP7AURB5fY4/GckOhIZcjyGYqjolr+XRvTXEcJtqEx2aSpK5q+9k9oQmjdv
5dUsZmQuI09mFgMpV8iwlgi1OD6+L0q6LV+OUokEUUtjdoRdRTNbBYA57/Tf5Lp9e9GohpjxBIdN
KGVGhBHS4KqXW63boaSw0hL7pW1sjCIQTvgbWBIKm86vFKWAbUbarvTjF3KqSR2zpYXsCC3oTxZ0
3M6BPQJD257YorO2AZ6N7sckFMPPNODz59gN8YH8EzS1aK9xOc1uwNFKaagedv34mgG/PPZVMwFK
NkQzv8jezBZgj5RrDmhQwS5OFyXIicyFp/hj7FU4EQmh3kiBydNmcaCsM6fbT6zqxopJnCrWnaO5
6ioQ9mQYOv/POtxDmKgPxyQ5jRwyzPvsVxGVRSxoB94FMjDyTHIsthgS6FnAIBXuVC/Lxm+oAQzh
bKXhJSsBfGRjNj74qleEVmxumu4rEbZPnNss4ZQJY59R4fgtiu2DiLi5OGL3satAaZQw5K7jY27k
jGwN3FwkxhsLPjtcNWwCpJME7jzrZwyZI7flx1qre0Q+MZnUf1k8nPWft8Qt+4H+1UgHaajx9DlA
ggnQ7LmtV6ln5rGR/hQVHhKINXC2ULo+5y1x2bgFpJ/tvtK7sjpjp+Ir4ckxJw0dE2oNVbPgL+F7
tFisD/w2GTn4ILhkzP7b0kkeD1q5ajk9J/omVWkNXQ8t6fHXPTB33vCWT5uAw0kyvpEt5nb8DdHV
WOSRElqRTU5m2Y8R4wYjfaCmiA8LGIO1r+db/61DH1IR6CY0KbA8St7hJWIDPHqG9/T9Mh+n+Xue
WnKtNNGN+gaKQRBhdIxMmL1MSmTW7itcvbkDHSpc10rDxTzlBK2B529kE5TGO6ftivMprGnwz+AC
LndN2QXfMX3STIzb48pssqW0Fz4+FQSzWqtzCaP8bvKqPT61RVwVXOmKlOrIfEQp9lh1xfiukOWs
tF8Eo0DloluFN01k6LogslEOEDRNVHYZt92sNr+AsVDp7GPkx5zpCBzoRlbSzfs3/Y9DqNY5T+/u
IExibSaWVvvGoxvCuJXEtIsn7qeLPdEmif2YTyaVJ7n0ffrJqG3/GE6Zat4Wb6LUPhRHI28hBlBW
NsntcCX/tgxCORko0UzwGvTaL+gkuuBGgQdqI6YdNLNxAkGTLddBqXxShBRz5v4isnYrYAnx8f1a
tNINh2VTGjRcOxZoPxXcMUVfCfHd4/3MDKjhSRdaS6SanfJFrIX1ztQmv+gsy47UKTiwFYkA66Xf
1CDeZwQRW4VimzxvFzVBSybC2VZANdOql01LMEAme0AKep7zed8aCeqw9NwVJTznpy+uYICCzlBG
WBMRj+NSzwKBLqSEobiMeMIJUHnrHH5JS3nILog/OVppqO1RNactg6QwOsXXkbJ1SwlzhmxCeyMK
VCBkh2zT3QdpGbxfR0RvY2KwCmgaLnCMp+aHd6JfrVBs3Hfgpcc+80jEJrMqE4Kzhtw+hdSUAf2x
LfwpAk5+0IR3bp306+xTf+oYhFNvBIX5eAS/MwAY6JtQ3TvoPrdCDwLMsWNny4AMQdft035z8zK+
70HtDsiUN9v4kk34HKCWQ5L2s2gGofZJkQhy0yqFlyJNzpRCEGBJkdSyCK/6g1+Cse6lJtrJrcoK
G86pkQd6E9IulP0O4rnp/F5Y6+oxUz4iD2Xtukvh+zMQACPh8TfxWMwWdsl3l9OxnUESw07G3pHA
/Bl0Vu+yXpvaXFYVGXtsqUq85xF9w+NWSK8eDuI3DtD+8DiGDgjnxaR0VNYjKuMys+/hOKjt05dv
Cc+YsCUYhLVZE6V7xkDO9BKynpl49BhRmm3qstvv5tk1VSuxF7paTTVkX3h/YI1P0JdRdyju0Dmv
80at8laMlxXbLySbBhyaZdwxp9PtdPuWLHHEaPJURhb+8BiugbLyTbDc6tpGFmKNIy3OyMd/GqbQ
M57msbZp1iNJeLadmgmx/mJteiASf0MVaXXdybLbxNNcj3oB1BDU2of806QG2TLy/iwjRJ0l3N5U
1a+nuTwd1xt8IEZd29DzknWmqK13qrZgclL/AZicFkTGrxBnzNtBJk1dB6jncIT2S4m7atPKOLn3
NgLMe/zX+BoerJ4ToiRelgwDqYQ9Ytz6++bUAkv7il+jATSbPbdcooGBbhadlBg5htlid3bhHN4B
9ebrChDkENQMKfw3bDZoAevkbYNPUGGqbS/xNEOCITC47uUQzYJlRR/7Z1xOtZcybcWHXiMaMR+h
48sy3uuJT7kgwE+LpJB7Gt0bO69Et/eAhVYHshQ4zJkVqCZPSRZOY3xOTFBtymvI7/D6kA3shdTn
N+5iE1DLsaQlRnQMz6xJ9O7mTGHTwBJJjHsydZF4DRgWuuyHnxbT7e6O4IfLdODd8PK806IQYcMF
82wcAts5VlvqC0B5OmvTxUaj5+CfPQ52Lu9AWbKBDvCrbIMR+Ir9MDg4kgZMCqU5Cp+TwB8GXZtd
ofvpTe4UjWLYSi4nW/XA0zsmQEQkJEUslqfxKGzV2XKxJUt9sXV9K9Arg6EYLu64kKXg7KgzNV+W
Ew8zn+Cmy4cDA2d3BcICWrjPPDhkTF6b2FVh//g4ccmscWuS0K/fZX8pzKmtzbwcQ3117cwJpyKk
1JAuWotIAW6ovoRnFgJagxPvceGk2/clZQN0vWT88siR5EQUsXLicrlnU5J7tUxg5+FkIj5tDZ8r
JG+j0g3wNyDQEDZyqFWEiNZ+APkOCBAI0NQOeqf1XN6UQojXkft2K3JJKOGfrS0BN6lGFKLJXBJL
G6+1aMwnKD+6jgUPZZbpdQxdzRi45DFYdb2XNQVZL5FtLf5D0l+y85F8EJa0hyv/pFvFkujfsV1O
NdZf37y4LWqasJCNFZUVWZlIMLv3PHoFCoi/e33sgLNw6nvXEULTqp7wYsw47Q5BpLTqqFGrjsdE
OqnEZMh+GupKNzuG9rVZcjEp+Ql9aPOkv7dYzNkDkIRI2dJGVF/T077pb4wBs42RmF5NfIkveHL4
a6H3oOz/OOLCxp5dZln+NrzjWCbPO8aLchhBCBvafRIj1Jt9Xy6kOtnfmQ8/c1FaGBNXqQLuBdap
2HQaGvdmxiX2Ps9Jv/KkvtGRc3ihHoG6sdtatHMiD2faYMMzC4AKs8CCPRnLARHC/CTSvKhL9Xu9
fphcxsJQgmJaHEh8BfXtwnszqTRmMDKKWU06bc9ZinNJDieNGx3kwY6fXdDOzxRdczT1jx4yXVxs
4fY/GnTZ9MyrS3Q9ynbERWif3n7pKnYWxhHXn9lfSkHEu2JnEf77bR0ZFklkSNhBP9CktXc4i34h
r4EZ2JX4c5+jk5hpsjIsGgMY9MLeucaCsvID7uuHum/5IcbindbibDjqRsDx3yMbkEEKrM/4KZo6
Psqa3bHfNSyEi9ovUK2hgyeZd4rNgv5nA1o7f5VQOvrdWzqP6qUlGG5D5VyXbIyMLcxpG3wKHuxi
X+cFmxjUcxj5H4xk8kJp/SQaFCR1o5hCp6aKol56lIEWhVDRBYK4SS0ATps9qr8wXDRELPyKhKwR
aM+NB6d4OyGW+cwyNj2dpxSM+3pYnPBt1hH5Hl/jHHDpyaXklL7qE6nPWzaCYUOY58SZH2DejCAc
yZtILUNvwpni++VWApjkSheVH0U6OhW/wSRasT9jEeyPIh98FzU6OsNuaD0ST+JZPGcw6HoTXCTE
A/lj9OeNOYupExT7fbdLLGoumZG2hse2QEayZ+JGfV8VgXyq3XPjci/6jp1iB8VEnWcSpS9RS7dJ
f0Mo0SFwXdzHYCPcAelUMx3RNYZS46mwTRj5eONrQv9BoCp62loRk9qj/DIEuc/3sLeRFMYky74V
ICCbO1JIZaGMw7hG1ibJvZvSBuA6tDkODGGf6DCjXDqGX3R8YxqVfqPP0A9+LuZvAd6ZPvcHsfNi
QRIIO36Mw7yO/C2dnWLU/JlMUZBv+k9Vv6AOlEC9Z8CZGfpO5GYldReddqCthgSwg7rpbR8bc5ed
u24gKdbcYN0vnppLTj9UCpYCOTfhhfLMXD7ZS2w5LajtuFpuB5jD2pXxwR/AH+caS5aKl7k1oWvX
zpPUxWivGRF9kuH0QpoYf3HFQahUGmVth90EMeGOD2YfC1XoX8NAkLzVx2+LlDhs7Ba3SV8PIHpk
o5cQ8mskfBvxWp5yzjGpUr+zuUA0VYrWDYO969DETsfVAS/UrvurVeCqhGmeObG9oyGSHqLNMCTe
4nVlGA10LzxcvKL03eKr5HsIeYnJZ6eAlvjvNLathRAc+EWTgzjuuh50LVyg4MoXkg26FZuG8oKa
6H0OxSqViPipT0sIopMVLYCKtvVHQLxjSXCf8QmXtGxEDLXeAQ556LevZ1ia6QoPxMCs4lSppw3/
tNP6DIa8h53oP67vZyzp7mHEzGewqUHSeTi3rg0PFDnmgAY6Ybw0J8SyXfDfyBnyesfKpciQgFE9
oiPXld/ZIXgxNji8mGXyAa5KZDlP+FnBXuYSlull8cycF+vDA5XNnledi5HTFA8KLR/EOxSpwC39
arVNbGh1MLN1uYmnqGhA0Yislid5bbEMCuBHAuvbuXKNStVTZzu2A0TLtIMvr+wfhLX3JVoKM/2P
0nZL7g6Ki2OE2mYDzXld0Fm+pitAViIyn75L+2Ds3NTR7/LrT/J0mNgt5UNqA0hKfI6DyJ+kGZin
L6Gav8O8UHzGa6f7KQE/wMBQB5Z7a3n3RDVjEyFdxJMU0beydXHziZtzSrZ4uzAoOOVw9iFpK/hq
bP9H1iS4INyVIQLnxP+clw45UaNONgNug0eepdCA2NdaMhGY/gmsw8N89iDbe3J5XflLx5mFULh3
RcGyS1vjy5cvytMpVWDXdvUSKLZH9/FAEcOlugxsQVTWSb8DxkHtg3nghuMvdrqX10qF3KHl1GW8
OJGXSML6gwNyohBuwI6qItNx575Rt4Sjs9pzNACJ1e9xiasVhKXDIzhp/dcEAQiJGL0bxWmwpfgH
TGTOn6wI5cUjIt39O6rylu3krnNe1uDbyaxCHK++PfoST3KSirKjICBn2SiP7xsNTv3cBuMn5NAF
b155yP4khuJC2slkwW2grvVYvUkbaYfKse5lDnKRGk9vcybk8wm+k3lPQyWpm5tUmipKOfvSh3oz
Ho10JodD8u2rIKwR7htUKyZWl/2VPDHUA8GzcR1geetVkLO3ttb1PbgnDPmJA6F9kX0FBMGyg6dI
OCr3baHS3GMWwBwPpIwbXVPi1dJGdOfkgxbYsXab2ejRKk+vGpkjwbLcJ/U5TYozhspFSXgQ1hgw
00UcjGOTacOG8FtKBJYhTXxuGsQhl6lyxKl+E9iU4xpKJ/LV/6mQ8WJnSa/L7+ED1+WYmLBLzMOq
T/9o5759QswYFNQ2PY0Lc8xHCnDrDaJtJBHJ/SyF5eqAQBM57vuPJYwt8avd8htznpxba6Yyepub
OCxXYgrKdDwLN+clytb2ZGHN+cWmm2GcioEOC18zHLU1HUr8ITsHRIfXcyvSZE5RdXQlcDpsal43
vwkWwEvlePskslowK+Q8IER788Ae5Jh3De14MGyJqVXb31dLhNCVLE12f/iXSW9T/c1lswV5gXoI
pzHZdJ+Jq0Jn9Gma8aF9IOdVkdTL1wmIYf5WZ4RMvvDVR9bQrCt/HtbJbqg5QsEV1K+oQjPVyXm4
b3Gum5F257Ye4RsHsRqHIX2TSW82NsVxjF7awkdn7pExN3c3yClJnWGQwiddFmiiF9bhp9jNb5tg
INDyTa61tmHck226Lxo4z043m6Dm43CwIMEXqVR3gO5Qtj3QuTv7eTLCl9ZjKBSprFVjAYyLoKxD
8i5lgBZUtqm97omM1c5f3DpFIIzZ9LqvI2wJ9vgmz4JikbflXpJCbEAbXA3ez/BjNMTrjbS00/ui
eY/cmRP4Dj+MQmwNKEFVFeVpUdZ9PiD2BTOuKPvso2ABY6q5z4Z0+Vv65iJkKnymDWAn5uuprvHC
lGi/fQYxZTEjOVdwsoyosY5CM2nzR4K+nfpLyS5u0unLhHZQ4t5zH1kvjy6CKM78iDkVh5AVkfN9
Zq0zTtQb9bZu81GPXJEDc7o7XY1XjNDkwq9XNHogDI9mpdb3a4lH4WGSjM+5nSdiKIlnueWq+Ffy
2Oy1mSyFeAfKLtS7vVz86t+5MfQxnXjmCr7sAsMqOZiF/+YPvBBSBUg6zzuYd+6NQH5/tc2gm8aN
oPFuit9BdsbW+/jXuEKfbI5FGD9ySXqpiOf11bT6RQc2P5B44hzyc4kwxlFr3h4qktIS1yKXc808
va98nuKUK8fhFyqExGALyu8IjvHFtWfSXtD5UllVqT6AoXYz240UA9YF0xIMwLcoEDPFpIgFccv9
q5KOU8QEAuR/Gn4a23+i7TrPxZo3WqLwHCe/it/S3f2oLL39g6FeP+ablM9izX3MP3tMUwV0B+Yr
BPEPEmAGcmvZmHpAWQFlSwvvjRYoeHdEk5pSHA3JMqTtRt3ChmcgrvGKwZTAk+7PH6zH2EaRHuk2
KoOwD48eySskw1H1uEsVFCNnIVIT8k+4r0vDMR3KSzaWQrDDWEOF1JQdydTuwXvlHHqlr99aZJma
AYZvfvqeGfMMWm3+Ak0Z2DyALrxq8eIh4AMcmc0nQ91JPZtK1DXq+bWiivRKEp6ZDS+OWrEC7zgS
bl6qK6VWF+zHLi7iqq9bb99t789jzJo10glqsLiRwP53NAE8low4n0skrwNnvK4npn2bFUb88Kkd
ffcR/ornxRBrlj4TSyAXWV1QEFmsJEkIrFrAsoKrgo+DUi2CJ3wylqtjHWzcGMzD8ZH5+0wMbWJ4
FX5KxQhv+sZx9F4Kblj+SDGlKwrLoBhGhSgyNd0XJ9+l2fjFwD52sVRwbakWQ4ERtNyYQOqOxkDj
vGGfESELZ4yOZdkJdQf3GOs9IHGEv++BBxd4PYFs4rlU5yEnytR0ArtTfJ+m2Y9u4ivjPzPuhslY
xezxS+TaCvmdqVjidE91LBUBRwGqvY22uA9zucbm95Tw5X2/P95itrcOLoErsLFiFdSnz6Lwr3rx
bGFD97QyK8s80WxSfghTdMRgidc4X5ZnQNCZ1DVd6h8mCW9ZOgdUM7w2OcBeeK9QphJw53+cdHWG
R972c1VOYeSbIoY03k/3bKtjDveTaptyx7leB0fxOGFTZ1NvcNxUNtnvX3UdfQfjzZFXRdnE4Quc
0TYOgIWVbxmAg8bF0R6tOipPo0p+OPzA8K2RQOYp11+Ht/NnoXgzO32gPQge4T+8aiI9Ar8wajEg
3M4WXm3JyYan2W/zrNe4PGCOlx4rzrZu28mwlKKcoq67OxUdHIGH+DK5JOPrzxJ85YQ/2vTUwDTp
JS9oGg7D66VMOeMFaelab2DP3yheJdMoCKG5sSDhHEhWUN+iEUxMnxrHA0X5D6hbiJiHD83IfsK2
IX60qHQP/u4lQfhufpl56qwRAaReLHyMiZFLBIjJ5/uPVIrOKwAHizLSDqq+yuAKKEBDtf6xWQPk
ZJMqlr5O/NUuqFj35y+GtrYc1Et5EtFIV22MDq6SQ1vyzFtiWN4wyvzU1ubNdbykgtUkYgAN+wXK
+dAhcI4GxnS52vQXNh6jYI4cSibnWcrHVI0fU0Q3+xl7+Pu6/4Oq+x/uvO0flTF1qIPQ3znyZaI4
alTG1y/VzLB2PgwxyuzVjbtC3FXPvlEQbpFV3BSTovqCsIdu7e1ioRdHI+A11Euqllgr6yQFi4C9
ouhdAGtQG8nSFo2uLpbKO+/RcA4VEV1SfffbblZv+iN9Yigp2qAfLHSp8KsGk8Rqng9KgK55gzSb
qw9l1jU8Ja5IRPEyoSszRi9a6PSxdyv8VOEmSkJusazopEBL98/bfLUs3sw/LJNkAfy0q1SxVUbR
TJ1BIgbpfZLeBh++1ZhpUkfMboNvH++JqHX1X7XCr4eJE2p6jdH59ShDINQy9ebi/BwE/hXSOW7l
UOnk08IvgO9tvHq9ZWQ2AJOiJe4jyrnedWVcllvGWQgqNUnbVLbB2F0wTaEYKxjAabGp0uGbdYOu
b0h5ChYin7WoVgnndz1ADxy6fUUneljD5OlMOssRiW0tzvpt9o3du08MqKrb1EIcyMcbVD0TOfce
snSPpHNf8R4Aoe7CXEZFshsdFSoX4t4jorHtG6KDtza9IR1BEqecP8INEmIV3WwOifq1fda1ppU6
rksGxC5Yk/mK1FUYM/ms6/7Wr8gqim4YHNP3wxjzeCBAh9LoOX/njma70nzI6A8FqEWansGfEKGT
2jhyHICzUrRlun6jLDscsY85gdIAJoVCor9jmgLUh2lK9CW8K61aiMTbIM0PBm5E2YSP27QP/lS7
YvP1vp83/zktiqT9A0XYoznAd9qRXtAsCQistdKi+fNUGUEXd1ZHiFTRs40A9zSGmP89qTEXdDud
IjAo1g7svyVmiCFVHdhSST0QEkPGzTpBzh0u39XrRG/lAKbpzA8ZcIB/YIS3Cl4sv81AAhI+ftT2
iXZCG7pAEJ/4MdV417cBidtc8FZq/iuB4OwB8Ds94oWxUh4yes7y15XegxS8AjVmWbMWvvCLLkBV
+MXJL1vkEGThydeCqPEDCfTf9jdCEZRb3fDjy9cqb8p+lSFGBRY5+aKVPND5Y1vOy1hZlIFwJP1d
mzBWf8Pqa74xrTJCLVlOZYmnUQV15y36/1tFRmnblom6f10Zxww9j4/Z5mTkUYuYcnDvPjrgV7g8
VQk8mS6JsXaRbKYtEB+0Q88/tP/LXCGMrLg3rq/jRezzj/jJH4BPhUcmCtPY0DJtzC2axCGFsjic
t73dZJr5yj25qA3Bx6fTdQIwm0islVMfNTE/hWqbzpeQdaJGPPVOgwD9BJqcpH1MeDMs/rjd+AtU
mVG593fiMJmndZNo9ukO3kEqfnsMj6cyasUuAk+MuPVLlWpZlynXitPr82R3mGF/vbQIzTLVBtp1
ATiT+Gsp5kuFNmJK6wJCjq8kO5a3YrSzdVmHBKiohLIMsoyJo2mC3iVQiAe41JYaHo8uLe7pxt6O
GCjvc7riTJcqNfRB29tc6Hyuk7oz/u/mrtcnsxFP9hy5PD8PEr5matwpa/SZDJ1BXdpTc8C2svdH
fHepHo3IJoSl4GN1qD1J0YZfepPo1LRWJceQ6freBy3YL3HdCYo+9LgVvH//0vPZAVvAO71rAYAG
MX+g/OYa7MmX1U4+jlfHHlTf3G+nmAfh5swv8UScsNcbUyIgS6oPBxypE2RRE7HgW7tG+XtM1tsp
sqZw2z8J/OuneDezTvi9pMIsashy0aUnzCKWiPvPBySfsEVbiFvCP7gUEy9jXSTlF09aHWKOEbFa
06JeX1Ml6/PkgAsal90TniaQwnrzrg8Bx/4LKapRvhCnvRIZLsB7g+Cor7U1xMkL4SCrk9+5kW7d
Naz5kZFZxUHdG7bgrASkE6slmFbrihDNPiX8bCmI1ubdczoNjHn6gM8CA1oTwQakTZYvaptALKuj
n/uH5h6bMCRba46HLQVIJ2RpVc8llQJPTRHTToLathYf8pwJwr0nTPRF+K6rMZ3Bn36dil+19Ory
5LJol+QrUkYvqUkY5xDiibu4f1RDbMJD5DpisGdF28ZoaiERjRRw54gcquA1l/36NIWXdGlyRmJR
la1jSwjcDuKmpDSaGzwkPDg0y/89zd+/iZDQ3TPXAuiXZcoBL3S1rUvfXyRfWe5vSsO0pockkvzb
IMqC+YJIHluTIyXmzVAJfHN6QBFn/sJav0DxY6w1kN4JDcUVSZOezghsJxeM23mhtJDzsdx1UVnE
cbJOvrJH7YEKPOrwsmDVKSeZp5NEL5q2397ZeR+Ccz58FLjYA6gN1nk/Qd0JvILvaFgBfLFwPr7B
oeHVqiTYxk+VJtcIkXbRKVhM41I1bDUxllmaLJisj2SbEbaCO5llTSykx1e7tvvIOSLpg+18/D6G
3F9FxMjzW8FU9xdsz2zt1wc1BoIRviW6sHr5ebxAqTxpp5a1OTg8DqO3vn9Sf1n50u5Os7W5S1jh
MdyXcsHi7HXpOcz21hEgr/2XcRwI/05uf5V+lOGu9l6+uohXqcjlgNYOvsT9KKpUIiRPcV6Yfcq1
Bpqi++nSLZoSTx+590Jec/rj1bPVu8NNVT6GQ7ICnI2D5hkn/nVssahATjCsfIoF6m0eniF2b2vb
RcfRc5g9krNeWt68lUUiHgBqF7WPyPGxqL1zc8R8kOTU5OBsG20L59tzYX61PZgY3i5wVkpvY8Gz
MJRDLU+TRzx6tbHfxpEaTaE3FZC9bSKdF5V2I0Sx82bLjBmG2knp6/epGnROZ9OArVzMLyPn9Rao
unggj20QnJhTp28Ap6LZqtRs+ccM/YG4f2e4z6VV2KWhXYzTyZEqSuGVQFSzwDUgdAVc7Hnr5Byp
0tJ9UNcIouiGlRl3kQlkwi+Ded4Ad9wsOLmKL7wrokMHXIEuZIuAo7VkoX8TKihCtsUFK7kGeuER
A4B9cwWI7RJbFncYhuxXMTjAqR2cinVtrvzXPAEOv8W20aeDMG2y3gO3jWNmNydg64+K/wf36zis
7wOQJACiDltPYFXNuzsEfbOnNcaIlciPLNEPTq6Dy5F2NeOrwSJ/08xSthDcaEsmceINpqghoWMp
xwrYWMTo4Dp9PuHHQT+IwuaGemmBxgeyyEpRxWyW+55Bo0IlabGXn4B5dmxl03J/4CcGcmMWoZqj
ADos2UVto2yYDd8T+qEBwByK4eRVeUlRsxbkU5BM/9MSiYbesyYwbYPJwmB/ZyF2uY435Sd9+p4r
5s4Xcataxz1ZFL+9KpiMCQEzLMaoyWNCDqS5fT/4rk8PageaDWbrkBlQwi9hY1SnqI6pKVsEUO3Z
HLyrtfUmW6ImUJYzh/lWwmxLMa6Q3jXD3y4PMUF8h9S5/Q9Cds0cyVwSZWWt48q5fQzuzQ4/Bg2w
+gs7CXqLa7qvwnn5MRngUanStQg0orxEbeF+v6zmj25CQJ1EsubDIPyF8/ByUq+frYdBNQU7RlgM
fDgSpNP7sv432tbeUqbPz/aIPQIVMXfsJNZlOTK5uffbn+KBiPeIfq6gSex2GoMT33XcveU+Q1ZB
DWDgT/O775pxB+ltT6nSIyvjFXq0BbYZ3JZSS1TkHi5284sfEhOb6p3Mv663Xd9j+ok73s0rXh3A
pyPGYFYaNINKKe2T9ALhSSPdT9i+ajRSD7EY0/JCIRrmayLvrOciI5x+txCIBhYWOD0QIPcQaozd
zBqJd57coUftNe++nde9pdf6+0YT7itR3+Nl9PAW0qwoD+SBPV3ekGJonYP1hU7evblxpxVNLcUn
GqgIKHx/OtiJnDvXtEVHW5az3AHubuqBWRDwvNmbBVvYjb1r60PdXRrtHjFCt+GoyzAZQsK3Je1q
LVmgRA/4DgLUlGZEoZrEewBDesToehN43x7krkU2OMxPmgCB/SXWkWNHi1NERwa2qUdhtaWR1v2Y
a1W6Vj7+WjlUeZpE6Ol9OovfSCWiC0R5mU/ImCQM1rtm3hUhYfQYkTjIKh1Q8+seWxahkQ204T3m
o0bcbDvSKqY/ZT2KxixVVokaBbiL6aXoDXLkf+0Ax77nfmvg5icQoZbJyNZVdOFV33RS2xLkLeF/
GZXCUPsK0f6MhT1C+wdftm0JRaG9ApbGpUepjGzFWgSL8lghYJv2WtRdNF0L4i1J/5wCmg5B5iG8
GRDjvr+lJJf6DJwPpb47Z+0wubR0LyWcm2+eGzvkKONbf7x7ez/Fe3I6SzHYNvXo1iczIT+oacqI
zLwj7GwnLmolzKf31a4yDTxqfks/FGCYuH9SZHv7iRH0HXNp6eQ+Dv+JNTtKQZK3JZ63Szz6EEZ5
qP2wOaZjAm2a/m/BjQFxXlHdPUAhT7whEZM7WRP09DnL+Pyx8fCTVrtXwJh0vlT+Tsq7f7K5rc0x
pQkniFrN/7lq62hjC0zgniMFCX71HJSSGPqchvKA6jsfH+OQESpKfuXP1/yy/z9DgNssAfrxWn/D
9MIo5hghoYAohaqTOMaT2PzFmz38XGA+aarAeg3SPAfcq0nARnz1uLb/yt7BX4yye5j76UlghbWD
DxJlj9pe84LzahN+En4GJ9WvXIPvVFop9DsjygK5Ut0K/wI8X91rQtwR6NK4+5O5WK+201Cc7k/E
t0BwKo1bhp8K4KXivCdrhsn/KWxpYEdo+5YfrMBFGxiHmbxlgu5xE6cyF1S2FHXqDOc4a/xZNgsy
0NYkcGjWW4s8NGpKLEfjt0qJ8Tlb0ElB80T9jez/KohRwP0PeJGSWnhIEzMfVDAab4jVL6rqxYjJ
PnRNw/508KvrtwFAfDSwYKTWxy00gaEzcIrKW19pUnyG09VmQO++Ar9zBZABxj5+ui1RSqpFp5W1
ktTxb8HFjTADwsBl7HJ/ZsLTBZmpinpPKs3Mjd2Q+bX1kVEsDX8p0TquyZEGBJrydWqJ2Xj32nEG
xKC9KQIalm8l59Md8QYd3FMfL0qFzf8BwgTjdTNxY7/0Cj6JStqSIK3qZEb6eanGAfQoOfmh4ncc
x5pEmKr06YY0k3KDszoSSKAgqFPf/2fJbZg74FVoeFqsXsWyRhG/QPKo3Yju0FOlxu0iomsg259Z
LnQNMqh6VH5UKlywHon6nKp+2BEsGjjzjpZhz6SKn/rs3bicw+B42+HC+rLH3i8SSz2IhGAFl/qY
7NtK0YZaxoGvHsgLo1lGj36IlqJ4c4W2rWTn0DrhruNUoGC5TB8s+IdyHhMSASn+JzzFA7sgmnA3
hhzedmVCx64HDltXTgfNO5mb4HjzLQkWJDxgs0tSsjyiKnxGD4iC4eQuvEI4Y4W5vcOciSyXinA1
h3EkRl0ZFsKgMbFUHTEk0SWV7O9fmW2IAiAtW6vGrwHmXRWrP/z9loYoLxg6vFTfTf3kHyu+anxB
LQG4SLYzBKQ7GRpzoZ8zE0PxhkokrdUMoR5Ajd+8JJ60M38KbSlYwZxtj53M51bFnnUYB780uCWN
SnOz5j+DL3riaObcbZbg3ZQ5kjDQM45w3Ey/I2XldaRZpP3AHaL8DgO6CCB+TkUq5VZ4mjMwU8Nf
JQbpSA0FuJQ8AyNlM+apE9bZWuOdgYsC1SoAOUs6eKA9EuKlMfA1DYJFa2eOrrNSaODbK7yUM5kr
0GWeX/ffDBU9YzhNTzs/014dz8x4oJv7zcVrKJpbWdmxi1+decLacBSlzy1Hrwlhszy8F54DLbqU
uLtRrRR2KWucmhVIJYSbowvz+qJ82IYvGJsDVEG+KW5HZPu2EeZujRvd+P/CmyMwNIWZ7gRJHC9F
qBnC+Nm9Ka8Xb+nIio6dZyfnBGiDwIPyjUkIfIkMyayoO5TcQWVRFD64KLXUsrBUFGjKBOccOJrC
khEip9Rx2ZCgQ9RXkiGWcBcU1UCCRiXyBrVGGUhGEarl6NSlJiskkudv34HwKHkkAUNV9X/IHbPZ
NMMufIwlmekBGavSgEqz/npQGnQ6wrs8ePz06TOP3q3qxLAtVQq3lCz0Jwd66VSpaIZQ7xYjqWaG
ZH5M6cb83Pb+MiJWYODdidGDAOHR0CZTqtWuvf6fGFDqAUjCyixUitWu8gg5nQ9WFGB3G937ZbYD
mo9S/7iiOoqt2rbosuZe4DERf54GM+4daLHfdjfXkXck2Ti1vRt0bz5X+7jADSETXkpAbIc9j8yv
XCumIEl0CAekaIlXsj3gIaMUwIX6J8QPLViQNUS8YiUzZ8TlQfs4+Oq7DiVRcCz0EO/WEh0LFyR+
5MJTwoTmGsJbmFSaQ41Aychh+R4QIv42/aV56phzq82CdiMJJw2K8WzcC02lDgrqlkO5vrtIIyyT
vCFfg6mo+CLCKmgORgP6ivllcBHPpbZ9sf6zIwIQBSs/GoP6WmGPrZsTFUPta2xRMrRRuFb5FEXH
TDp71TWGA7IZxyVC/nI3tY4LM0Ehbo15qlEhEwl4ZP9G7pV9vRXtnFUbAlREmGvt0XrKFMGlUrzd
gBRGXg65XmVKrke2KBx+C1MyR4y2HILlsGYhvSYzqzb1+xYB4aqatDeYT9hZOKIEOEdJjO+UDfjf
WTiEXMw4iFR4BDDhF07H1ugZBuMvoHyLjsnUa6v86VPDXP+X2BbN8KioAtQuwwJJaAPgIWDeSMnX
NX+egXwrim6L+aZu+BetF8lKnbG98B2XjWbYayWsecpBu21mpPtGvdi8QeyXI6IiUINCF17OVqWF
a4D9CfL9Pjm0f+pZ9qWSle+tXmjIZ8nwjBb4T04KWleu0Gq8NKsUXnq2jvYs2i1gu+iTLiAq86WP
/gxQDJyOAborfphwCu4OUe+qB1QNTCX9tYkLSgx6C9BUuzxPtCxRobJy+X4X79ujhwSMqNzogXIP
x2mQ3jUIkkroOwCZTujams0/ZZ5RAflRm5iQIGSmI7mSYza7VeRoMgbhB6VJ39tfDBQukspwJBJ4
yLmt+tiyrYnIb9dv/JGJVsTHoEmbxSHSoVVdDH0R+x2ZE9jIN2ti9XqFPGvai9DvaUTLXo8UcwLZ
WM07pCI/0R7AkJzJP/aEvjexKCYbUbDUIqMtLv+uUGB4Ekm1gfovxsvSp72WP2PHYw1XR+Y3n3E/
Ryft5bMltXWDk5ECPlIE2a6ysZTo0hJdK7WU7oww4mptyOiKlcbswJOt0a9u1tIM5LLr8m0emFRD
tSzv+eDhmWUm4sfZoWClz5+6OqzvSj22s7OuAFUBjAPtZz6pH7RkRK8diPvAkR4e4LCLwdqBJrCa
KbIahWrcJqmgwSMIpQ5qAmtm9Y0NX+oNluhelLwkWx3W9WBvYoTzNbEx2EMfGmrjPIXTsmdaWR8Q
UlPmc5CNV64omv6XWLhdhOeTpp7i3T8MjjvLRVJI1vfjE3RT7cUHuEmHuwFW9G/oQR0z5oq5NnmC
U558y9s/fxLphYpOt/03FoeReqiAIQSSFbSuwCjyYrmj7QNZce2xy1RGCQbp6JMXU74dQFJDreSp
AIF/SsEXtNNF+O5fAxwIEG8PTRpATOb/Aj0OeRjIGOb7ke3Jlc8yiwazfJMm5NAjlWxHXBo2+tvr
/tKvLI0OAalasyC1qjXg9la81EcTbhgXv6eqGZ7Ap6f5cwFGPp0vN9PnUmx85ExzmkcRZy5Y8pXB
c2VgFFeAJdFkuC1B0IT3+fKLVRQF7SwyrRoXFB4lvhWUfY5y6halRE/3L4P3EzIaPzSFaqKp6Z5Y
cbSLqeKsOSMjsvfpSxGrun4+ONc3xYJFPZtaeUXkAPg6ugqrUNr7Z0Dz34y68kCJQqhi/ObBvMR5
4B1v+rxhD9KZel5G4jh0fprmTz+d4EXJZ4gKYybWQfBpT0JrhY5XMFELmEQC6cQbIQ8hUazflmPE
29v/K9vr+zdcn3qiisvv1N+KD6felqULkzi1JVpAnBeC21P3fKEl1qmK+G8kFoJYtVfZ4YbDDaM8
Fh0k0p1jK7lWEtRDb0+hKuqrlijihB5Jr/9ZNqFYcPhVb6/RgWNa8DobBFjD/YrlDqglUIrp0ClS
oS56RxBmqhRlJieDkApRcuizOIBi+QezyKO4gUa9uBTJVowfhafzw26NBCSpzNo5oEYbTFDPab2x
9kX+O6O3pnSJGR44c9vO1mhRw185oRxZGIZUyAIjQjEhOrX1uXBySvsraeU7LPJvEyyOKSO8HpE+
ckF/uuHUXUJVCEcv9Izh8NPbegiWSCAvVL/1bvgFT5f3IdNHrAHhNj9LP1CI7rAjftO8B6g5Pem7
VDV9dcq9tDCg6baJXj4ZwGdQ3SxaejGX5OAqsGeRjjjwSMih96x5Bc8LTOLrTkUe6uZfgIQ1KIjF
1qOdXA3CxZojOD8ZbpqLuq49xZNjZDMFT62OM5KW6ozapZnYI7em56RDaDbRDr0GJ7mn3Vi8pTVK
ph9tVOAP8zKl1pd9U1frjONiQYh5eXfTKXjffuuArF4pMZQhHO10rsjCQQYWlMfhsZYBpjyK3ifi
sNCMKYzg6wDrIzLX6WrDRueNCdbHQCGqsYavPqocOTt9cog6tlszoBZ47PHOvUc/Lkgw/V0/bMhp
awdWwP6cxSJ8CBcg8Tz59IMbKbwa6HKH+GdpYnDSesCGNCTWrbWUveC80sbKmBQorcoqwXqzEe2/
+fq8VqsAAv3W4Zu0+Oly7i2XgRBO8LRwZBwM+eyp3T85h3TUOLknrlstX/tyUm6nl5pQd37ujAzH
1stmmbxDb63wx3XUq8IJbUHbhsIYiX2VAHyR0NrZwK7wP972IYFqjqtadI4jYvKeQi5KprhALIR4
HHBfgIHmlCMVwPrZXkZWHi5jUMt+G2KKM1yqpk/m2PTpVOGZB/xvEnkn+vcS28JdDojocEw/j6Qy
t2sO2G+DYDm0pPD/6lhcoxKKbAtKeq5BH9a0OV1zr4cvWW3S9qLkncBCCh/xTklb2IsIrJv+gJ/j
DdKGjSZNAkqCWalWqVupNbtpCGoBrIJST/XLPe6lOS+O5Mtbed6esen34lnvy9e57Wkl6BmoHp/W
XKtZObRVChC8NF7KPa6WtZ6XcnqOMpUz/f03ko6G8qbxtgwuKDCtqsy1IQBO/0qsVdJmlZL31UDK
fMY5Vq6kFHmlaTLDSET7T5HEMhUSk3L+kHO3Dn5jYOXqLQ7QXV9P5WfDw/Jj70qZkjmIDsd0s4PY
ExyYwsR9j/dpTvA4mfChUk8nGFq5cL0yV5XGZI+zFyeDxZTp9C7aKcQvjrobs3kkzYpT/R04Psmj
/uHknFHTuoL4RFGzrDre/cdvVrjiYaJeiXBb8/qGAbPp9xCXtp4bARrA9MfrJkxsnXDvg1a7R9Ip
K7B7zgOrjlaVE3nGApz+49cUa6Ab0P/5Gfyikg6vKujBtlqyrRbEE/Y65T8XgzkEK87P4z0O57lv
pseX7wygpEJfc6YAAOxELxZr0TLqDpJcUVckH6+HJEh7esR6t0oQdbOJxQq/wE6Yycn/Sx62PeYO
CoGjgZokinRU6lhBDwG8xwXxaSKHSoNr3pe3uyUgysEkQLk8hR3ylp5ihuDdiu1yxHZ/29qHG0u3
QbXpgeYSGc8Je5nhqJEUhVimJrj0EYrZiMIfNvhA6wTPtNHc1ax89Q1tzJuV7xGWD12YSWTzcxqH
zaBRjM1rQXYG9YWukXlmxz/hNfJJcv2hy3kBUoH5pKywaQG94G1XETuRMICwm2IL4EAV83Tade2q
Onx1P4beKkjZzAJ5lp/PfYX/XYDt6Je7hkgxfSB59woPfTaOrCukSA36pvpLXFu36BVKmE1iHB6P
GCRCDKODqmPyymIdZQiQKZ90nsjJOLvUiubMMNBtWyUVyyp/Kbrb0mr63n5ZHKWeYQiPEYYdnpFJ
DteWnelaMNjgNXhEK7pps1HNAvmN1kmYiairQVPpHhRaWHbAV0GTZyENu+saMlMQo/avnoI3xdJV
kvYcz+6k6Q3DYg+07b/VQIckWtpQK6z1TNWEX2O5zUcnRI2So1MWjWBilP1IkiyJ4hoZ4E4Scqui
NpGQleKFwivIoOrXU9cfqt6Tx8U4gjuW7JHeJAA8n5BSgppX1AMZbr2o4DL7adqfUbFnSfeTQKrQ
N5UxU9UK0jGAMQr3dDP8R+c3ee79ahRcnVQU07UGAQc8dRnoHv9jRueCeBF9h/AET8CS2dltHPU6
R4NlCTQOok9lw/oC8fNIysT+Zenrsmc+JgdjWgCP09na8WUpHwU77I6K47hdt4+tTZJlsQaR+Z5i
jXyGL+EBvhWQsEOfVFoBChmn3a1yI5rR8Fckx/0mstA5icK+vF1l9ek8Ij3dxZpFCy6lVMt2468W
iBzWNNDSnzbbf7b553P71Sqv942uRD0g5IKuPyzgeqHVRSidaIT6Ai6tBzoX6hKmU+8RtM13L0EB
qkm+ZT2Puz1M7nbQ6xiETsEcSyCgsC9x3OEvIjKK6wPI+6tp6BE6jadohYR728phqEV6nLp80k1f
tCsqa8kgLYAvsinVMaNWh5dhVQ67lniEA6ytgAbJ5X29senDKH+2HzWnfaC9KkmOzvyxqkALWEeU
/+9WVDWislRsip/N3Z5sND3wpXkUjPhe5DZ8QP5/yp/w0s2lzGDk51F3HvYzuEsDACQuemWYAWQp
VE31l7rZNn1NLBzHePxv6knzoXc/FiAfnOWI8GH9fVknf9RWqL5O4vJcGuCBQ5uDUoECzu9dqpfP
YLUdP4ajxZFstPQ6cHUfPD5gMzxEz/On2WuqJqPeeLNniLQwBmQ+xD/buH7nIWTt7gS+yexcwbW6
+r7knGGO+eTa7+LQcnJq7I9ARFc7hpas9Fbf8EGG03PBejHnmai6PWRyDKpuYPe+JiSglHJorxa8
w7whHPK2dKhdengx1bVUuXvAMvr+Ce2tWQOXGJZHsXN2r9CXp5fsnYm6LdInzOyANxjp3yUGRXz+
XTvSPivpLUPt9qmI/j/oB74HcSsPYvIo6zomQsFnC/S0Mzd9+qGfe61MlS4xSGcQKGjOyXq2HnSf
EzFg12MskN7UbKVvuuI+YTVWOM/5Ybtn4TLk50XkwY9zd4PmLTuMZcUVazB98YZglosuVMT4zX7D
k2oTcojYyIpm73EZn6ELOFiY/VLDgbnyh6JiGGIkp5oC4IVsIkcXj1+DA3+JnTIo4G2OD7UiSWks
o7NdDcM0qNbICXut4fpRak9hEVtWOYIiUSkZ1lLoOnJfWWwlNfi7ariMm+5ofYINlzVP4J7Y7WqH
IgMeYpRtufvPHYHyU3acgMG4x0knJYj0QPZmqSKCURGprTzkKfsMNTZVxqgryluFhTsfe4tn/3b8
Blrk/QKphE3aWgWdCpekymfe82BMneyL49bnvI/la8nqvM29oRj3tQM0pQx0knqN/q4HPUZv/DSV
2PkMZc+eJcgp55ZkSu89Gwj4oFtBkfXINUPIiyPSb+qOeE+RiJK5IokEwXx2uzKtNelOg1shsKIZ
2Po3+2VoovrLA7bXVgdDMvhjZDqHmt5I6gQ8ocpkCKPRSRz7iOw0qGqfSfVGCTuGbcNf7E0hHwV2
ENCXNoBkaq0YxTkDt7NKs+1vU+BiSs2rcCyDrRUqdbq/DKiGTLhAC5Jy+1JYw38VLhgEmC5e8N8g
pf0N8y0/DNPRcU5T9TefbYuNEnXHdz5T7kzk+wTalJC/YEA7J0FnFP7OaWHF+4sBPHUNcwRzwxE4
e1MAJOiOpZjzTtG3v/cIhtofuCZYBTbtM24tXsfaxkJoRVesquArtTV0M9rn4Wg0+wR2LITe2faZ
r8iuIja//kd3NEz+DO18Dj7H1HFbwtloJW0qS0RFEz1ckKTncCviRDCE5jmdlyoXSX7BwiwMLj2L
qMJWm5IcXin6YeQGTWI/sC4d2KIJw8Ptbpnb21fcAy/eZ+WPCi5rm/AoOCbrbz5dFP7gBXhotk+A
ElqL0R+iq6ZELpmuWQINRjSv8SeOcyM5On1tO2B2QYJbnjyihSbYO2U5knSZ+J63oyGFVBq6kBw7
VPoWr+Q9HYtYhGFtCy8aiKmpwub7xDuzFuf0tY+QALqFi/GB6PlhNQcXDLLSBZ74BUhnpLVnWeNW
jNUoVWvzIFUT8foYbj0ZaqqO3pfXDg3AnJg1UPxcRvEec3bXZ+tHuek+P7cLfFtxfjeo08o6QMXF
ZsprQ/mHrJLeGkTg4vbR30KCTdHyjph4HeSNoqN+ZcOI3MUbOjA8lJtgZBZoPPEtVYCEC36zcVrl
l8AJZvn878tMwyb4eOmRP9JZcwrIiCqhAXG5SaUmfwChNRbLftCp60zb1HlrdoCoKJUCZW5pTRUt
cDDC/YF5v5V45/iuxEGsyPlD0K2Z1jvZx9k1eBFugJdTQ8CUJl/XQjxVmJ/MBX7HorBd8o+SrhjZ
K9MVkOFvwDTVD7asJAofqDM9QHFIl5OK7t+/gCZDGpMbsaeukqBb3puYwUoSl+AQQVDH33h7JqZ4
fEGUiKKZ3QcuAe+VsfYVysHQxkSxyZY1voLwR/JkUF27RXLhSAkRleKhu+5k32GYexq8MO64Kl1N
qSwHDsJqM64zqOURZmOEWvpdz5FnYYnz6SZ+VrNNja9GAgO8EQpmb5V/wKyov9SnDVGmlACUWe+B
oBLLwcuispLXiJnXCYOQKyUHYHW58OqT5JdCQuVlOKZUN6VzeEihHDmzmLyGVsCUaH8N5NsAV1/O
dzZfezSWldBJyeJliRYL3hDdmFGagGj6ieFRW5W4iwwn7K/x/pp4qPjcjk+xu/NX8CfluBoOk35e
DpReheV4DvX3B3SQTg1ksxQ8ITVwpEcGvMOiS/nUNB5HXfRGAFw47eD7tf2dDsS8fVEk5USy2S/f
GsVkQ4U+R6tlyhfKBN6ehTgReLWudkulw174yrP8X1vauJ/KYwAJkRG9ROn+Uew1OZrs341H41Sy
rkG5lLpeIAxdZEpjzqixpMLhc6k7R8gly2OKnh8riVhmm/GfovBEe9hfkHdtay1VV6cByPrSxDeU
1b4KcuvNKw/6w//HbXyRffqKaojJ52Eck8CABpES5MsF9rXfl+1dRDlAlEU53rjnJ+UAAQzFiEnc
3dicLQjEyUge1i/GY5DujHPB/5dYieDOWKccfAdEJTaHqQ0snUS3DAPVICu5ByoLdf0GoTS8iOnT
DB9spqAdACNOpMv7Yv+Eg7bUZ+RE6NrTr22lrUNdT0pzuElWY7E2cDOZxALD0VyUkRC013fLsb/u
4MpfBM4am+nH66bSjx/14XKFYHJSl0u7BwHnRJ+Yj4SpdhGZVhc7RBnC0NoisEIgMTl0hLzbRydS
XK7gj6xyv/TRSQNvftVDQie97ISTniXsbVTncr2wi/CWk0SWyx/pbh6GbIUBM47xTf2rmQq72bGp
xESBWdAJ3JrhpH3T5tMxDEm0W83w2vTDAr8RipWrrev9qXu/cJheevSFxqk2YQPtvZNYx78552UK
4GZbNBwAYsdSNChovvG2HQ4MwGKWOtli072eSDdoKK43ATZQj92lioap2fHZyzwQ9yepbboKBMKk
Zw6Mm6Q3lYqsLrEda6CMbrarRqMZ3IJUZzj5SjxRVPZlaRo+7tw5R8ezHGTIgeTrMxMnaqiZ4vpK
RF82PWIo78zMzr6ayOhTxN6NTPUWiZujDr7ItKqD6uPKrSiEdnpQf96YyseXdJJp+tLH69RfeygC
pVvS/KC7z9wPwCSFGgIU4ozczq8V/fWlqXHvwGjVhjFBBMZ39pSNz6udAqty18ApINfbyBewZK0K
KPwd0T7TL8bljcro3X61Qopnxej3R3Tzg2FDjI3RWSP/Y26Y+gPB8mIXemo1BGH5RtzdAwIYVgt4
clr4fj9hhVHwHgCRzwv7eVhc+CrwCxlvjGp3BPCK7+AhqZ3QXifrJcwjZkaYzfd45jsqjOONKnZo
Qwl6mz74SbREgu5IpbiAbBERENoze3s6k092TnrT7MvZj77pQx+syblRXgLsm+KTFW0hKAzeCVHV
dmE+wZtefa/lbM6TcD1UBlvBNo6LOT09c0T34Bf9iDKi/4YPiwcxFJ60Lo8v+v1lpl9tL8nIvImh
geUW8Pb+SlyVxcnV1dgG2S4HsT0kLv38bl/kvp8ShfASAVoSxnlJCCtEEAaBCc/s4D3HP2PeLmZe
tFhNmxWWB0JOB5YlKgTsi/WjLOJbKsN3yY+0JgHHa39OIemPkaCH3pCpIbEtrXRh5Psu6Jjr+k2f
nHpqpzkPuyHeGSW6E87SC5pa8jEi+RsK8gDw/d7VAqVzHnMmYPuTwoyMpbMpb7S5lb0Fcq85Pvlr
RTahb98Hd+xlwOO5q9YLgBu7ZGcDHN162ZHMQ1NZi6u7iAXj+y8yIErMb7zKWHB+LNbQfMyp1zN2
xoLxQXmqCx67uo0JcCRFzaJ/UcNThk1vggTiZPOlswrkGpB/52KZ7mwxxBk/yj9QYSd0NQTAyzOg
p16H+rmDp++ocfuP2Z2AF8xKJFJMn08adJUXb9dRAh5btKW+xAifRHQiVQrGqY+EcEs4zxfZRsdS
BU3KxUulne3DgYnqO6QfjwyXo1vbZXXTtTY+5FYIDMNX9qhGbLPHda0HH8P9rjb4KKMaFfReyCiv
Mzfslxi6UdqUvgZjyvtE02XYP8VPDSCpv3o0xbE8OLGqQSi2hW0mf9tHCDnVOFC5rP01q4Js5bDT
TH70UjYCbCi0zgP/nsJ4cJExiSty+z3PHdvoMZkMyA+oOCskmkOrNCOz29bEXq/SBtWttFgTyH4g
xQNPutFWLx2X5XUWs5ltpoGEzBtTJnk4kmezKdIBT+NnxGhjE3gd5MzIM0KrbZufgjm/DFeriW4B
FjBj4zrxwz5O2TZoetdbd8/mrj3ler9Md9VYXrZ2p3BAk4zhu0NOe7RrtIwtv7dfJ5O2TTEOxBe9
Ps7LdyZ706RuQO+XoLoNgpxpzSVZDc80BD48DP3xaebG9r9wryzk9eT7c3kkMpEPV67flz134Po5
ggvWH7nwNDMU5S1wOBowzlgU1ET+DzOkjVaLdc1KUJXjvu96V4TZWYLFCOGTVn+gIvFuJgJvk3ky
cJwZo22dffnPLgG0m75q1zFSujeRK8vEaTnou1QgrejOae0T4+1jAacXRnmYzmfp0KmO16UWQzb/
RphcP7YBUVg16ocDbhencTJ7jYA9s0ynqPh5YOMd9URMROrLqdTGKNnOVdRLq5IN3dpmcXzWNy0N
aEL/U5LHOCPZTcmL6uRXWgHjv38l/zeemRsZ7W18jh8m57T3WclCusXNsp+ZhE+Uh8a1YaCfEc8K
0DN7qmRa0+Ul16ZkotYb/Cy1qTkgCi87W1turjdi7BgKAmA3SGdrFXwuNSfVMaKcHP9IEgslGb/4
sLeVRPu+jLPOxyooTCLqR3fgVPRAnaKS0QCoyvVjVnk7ay8TKbko57V3I7xq856o/gaX51MiknCY
1VD5fi/YwJ5tGM8syZtHbxIsT4DIwHI2h9k7dKOiMYEbEAZvDsD4/OZkAb0DvUEdMXnlEWPvnyX6
6RxsKUK1vhs1yaftI4SoSEfb+Lmt0bLuiU/uQyGQTMfGKiY9BB0LZ/l9OvhxDw3Kex94At8jQmcR
wupkjYYfgKAHHog1U1/EXxVfPy69lsiIhPWl5CD9n0sHb530GaDbnKcffE9I4LI9lM8CfG8Q9bQk
T/xAUQtNZhIxPTwLVLJD9BiZJ+ju9SRw+UH5xSeagKiADEvnYYf6h45yP07eADIhDF3jbqqPTU++
yhS7lFp3p0rZbeTUKECJ9+Z6SeT0DuQ+v8u4tSV+0ur0+tsNdcKdoXiChm0Xm7lYsMoBy/DX1XF0
r/cemMjFMoSGHa/43/5hKeByARybimAjiMQmCFs07YbK6oOpoIF5iobQsGHnFD1MMy4Uif7yowZU
jsjUPWYW9dnqAFF5j0HySSIK4KfqfsHmLBsezBr+IH7ASE8ZYYTrdUlBaO4UT0YG2uqgR2V0+f99
vxK4ny9kinH2jhHLnBeG7mg/4VjVAnM6R6uXPPvlIE+6mJpfeIO3SJsH3fmEhDhtF4zAyr7GSdwk
1+P1/vynmolD6Lx+tlTiO305sol7U1Mfw1b+K8/6imqRMmPLnCkhHDHkouOL5JaJ5jsjDMbGyOJa
VCXLpcHB1uNCCPzXzuZ62+AEI9iuHlT6ix0ZoD0K201lFbFjZFCvgdn07R74JQnnTejbsUU+4E18
18F3fSEYD2RSxEXxvvgqcP5E8bIzeXx0CmMkvMuoBWJKrJTrfIrvwrUO2oTr0rtCGGObLvH0eGx/
5wlLvTmNvrB1ez9V6RmAwQAJzyGNVXOWbjIYnt6+2jkgTuzOhMe+Ppt8OSiuaawMYZI86IeAG0+x
pgAHVWSpjdmaI38exiCXG3wi+LSse+MtlTOvaxySLQk1glKpPK5NPVRCOFKXoD5hECsKJwFBoNac
BMPHMFrPFRuYvGBb+WLc6ugkOx/pS4mMES42tjDw+JqAn3I/PNynSJ33Jl4jugfzZsbBNknc6Omm
4eMl/e+eeHtRRaNlabtrsMhLk9krZQvk8rHdcpKV8jVU6mlk8Y7FCLZ67bqzxVv/ORwjXK+AwuDm
HMFR6xiU5ln4LsjFURcZvEoiBq/GFxAuq85cxu+ryeD3K5pN8nTLTJHiccbMO8t70ltQfQwK0m42
59tWhA3nZigWoAAGIkcXldOkXDoXgubb6/TMeOmHlZsWnB1Qcstg+z71RO+Z3N3/4uVIWTomFzCb
ivbC9gvCsILwBdzrUxieTUaSpO5WhHIWVB7IgHJOTLiuKoAd7ZIxMTSghRr3607qtfyi2aE3+dLZ
KK4WUhH0Z3r1vSRSePP/qFlm5hxyPFV8YoqY19x3rlvW90t/zqaUF9u3uTtj7Ft5TKcA6AmZ+na4
QU28r159UEBpYtdDxaTIJ1e/CMa5EKEu76vMpRL1bbb0sSOZ9TRlmxd28sqrGFKKkIeySQqgLnQD
8g97dmMDyCz0A4UEqF5yksOyaOkSp1dAz3uyShWV2tmOdAvlHjFCqwSYoVSv6CvkE/4OH1BqQ9q/
xx/XbGTXu/6eLMXHChVA7e/n7+xjkdODgOuXU1kTOWNjzWhKvR+bZ32yohAklHFoSqciOLA9ATAw
fQQ3jyQaZjKd45d2xMQ3dhnecz0NTIcpLgttLOoBCJDPHHxisxWwR6+CUXMn+UvZmfiUcbmjsI79
bd4q7pTTqotnCog0dyrSUEf3btM+HgLKSuHQ0fRdF9ciNKKJ5lEHntVZ79P2LVEAcCOlmHAej1X8
WtQSLMImptWAPtAz79n6iauGrlBBYA/XSHGyfNKBpCZ4Kj/qSUaUMASebODlxdUIsvkNWNIelvye
/gX+mGQ/duEsvUPY95xAelfDoPMDStWeWc+BFpB11f6GLX6N/zzHUWWnb4l23mKgTTZ7iY4joxjP
QepwzVoiqNWQ11OokTIrMhc5fUX9nJsfM1LmCLPCRy6H4hR7Xm28za0Wzmpq7XqTVuv8hw8Qp75U
Oyz2MZIZUgu3oS/uYz9k8rSv38Jnr7WPDevp8bcYxQ4Pn/orVOg1gfC0GHqiwOvNtDVlBPjkK1fm
gqcVMDbdhPIjeWVykwQ7MN6krwNRcGlYJ4Hcg+68mMsqesUz9GfuAC3Fs21M7z2G2HCABYOZXWsc
F0hWbOkyYhmojEAA/Ux6m0nSAixGgdgTko2BnMtIY/CLQWWJfJTjHM/KgYs8NUt68ubpQGwBSv6W
Wn7ht+QdyqsAZNjP7i8cUYwQidpeev8edUB4t3ExJJ6ji6yjZWI7Tbsa7GIsBSqKGZA9I16+ZvF7
eqq5YhigOf2RPRtf+09hHoM55KTFoURHtNYbVaePFXvEG3MMaQvkOrc8IMdY1TOZbMciO2hdlfA6
POkMjTl+WLXmdBVx6IntSZTQv2+y2Cp1JMdWdhHhNqZRzzXO0jRfDAKMS8u819PIAnpbteiG1vrH
fBVwppxE+K7aAeEvql2YHVCVJxiEM0ubRc8OSjmVMX3zjpLOq1lwxAGkJxt/+G76OFcgbABIJxbe
1uH7iIXTkjF4Dk2sjsMnkeqVZBHGPpu1B6O5YWRV935vtQP/NEiyUVGTAR46Mr8qyDDI/WOZ/AR8
yvQi9x2Frg0wM2lCN9fg8rLSq4V8gpMsyH9RqRqvq78xMeU+V33AmUELhp0MYNT6UI/8SLKy6y5j
3+c+xefOvdx1eamsalpgCkrJnVGbGFSvaUzUEswD/8Yc9k1FKR+1WaNm8nJDBgZXJon+fBpaNpI1
tNCAoUv0HSwQEtOOOAnNg5HU1QMl27XkFckG7dcU2HE5My+p2TVnPrNxX+H6ocGEvnEy9zosV7YY
wTFUgij3o0KWnGDR7vIXmdTmtpnY/r61G36jgZGCBtWevpObujHGMuT1penDBVpjcixzdmAnEL3K
RNNBypWBxeCmhTNW8FzChCdixuvQ+QzwvNOfTSPIhrdsq9E9VIW21xB1QZjUAvl80uzzwK2LSjep
RdudKsRbVlUxDG0o41GcmC33VP+MHqBbWfX3C89UphJ8b7Ne76/ppCXBGnU4F/hZXT1iYM3JN+S1
0AeJxXrmkDD28PeD/E1r13YBMy24tPau+soWSGQaLMNyQpfz+TA3nSTp3cfEE/UyGgiERhv2leil
9xx0GX06STy4eYnltLaM0mf5PtlEQkpl5gS4SjKuppofmLBSzqWYGBtXc/Mx3PkGmuX0Jgldoc9+
WYzo29TOEIWARf30g/oiJKW6ThrZOPBelCvD/qXvVPj1+ngAh55fuJReRMK6Z4PFzNJ5j/6H+W7f
LuN2SgDHtbGvqUpcQtzxKVRUqHUguhLl8yOnzZCpswcrhAD47yt22q8tFamlxi3L4LeDbD5sLwI6
QDuuGYetZYDQHbxkNTXsrxIA4fzbA+xmCSUHQTn1a3X6WXvcqE2nRmGuCq40daMDt8GSCIHKJ4G/
skZNrcV7xq24m6MhV72HLwUCd74opk+61+DyJkZKo6HPmboxSiCPSJpOqnvTy0ytJudM5wvxcuYa
3eg8UgUHYLOIa4xvX2piK/t9il6IQ+HnPdLVt4vHN611MqoWwvpzDTzSW4pghYwmnNM7Fg4k8V8V
MTCXgGcRnxhvR9uRlxQjuO24kU1tE939ZUoccbcMbjinLlvvtqxiN4Kl0AwjDloYg7ru7InFdhiL
oZxYoKaO3ftUHUlB+Gjo5sngjGz5HVcxTPXcXS5zSiMmha1AvEbqQdofOHYuIHbE7xMMcuTns6gZ
NFIbZIU3cOrMVOkBDG0VgNWgM/LEH/Mu85dflOoWUbl/FmwJW9K7xk2qpe14pftbZLGcfLEX0ACr
1N6SjJJFlAXDgwoacY7OHbTt4uYMD5oDWpQpADjXSY1Wyk/u8T5+rPsSmsCSd4tR36wBqEzU2jVN
2sybb6lkFscJVmltQL6n0WI/GckSQ7zieDrYDheTZPvNDhMGjwVJvwUXx+lkKCAjjw6tPnLaEfGm
OZ33iUIV0ZupSV6BRSQrU1SDoWB/2cdIXzXORj8TYyxK+j9/20blhpfP/yrn6rVv0EcrGi4ExPIh
K1k7vwcBb4x42l21bY4qeBvfCh5bDQU5qOfWhbCzMHqKHnw5pGt4mLEnu0k1jlSLxHu/RRD/InmG
18tOMf1yR2t9vDRrU3haKSMsKGKeHEeXK9aeMQYL8HSTaa/eNyJ9XDt6OE27bED//y340sdvGl+R
G03BARFlJeG7f41j7DyGmJ7f7E9C3Plw/7PCR11efirHCISFI65cqoVW9T6HSd4iy4KOYoOQ0911
vyLJBzJOg9qGopXhP5aGJExRfRLOeZIKDv6/9nQIFq65UVwxH3vSUAdIW8oCDzGqtyhcJET/png/
dr1y3VujMDbrYSx+BjmMji/BX5Zs/dxYwZXcfhxF1eoYjQkSShWkxFxe6X+T08eU0GMQxYVLMCek
QcKRvPEZnG+MTWiFIswu6k3NmLR9jFTn1+c7ZqJgTLHOi/gw2HptMEKP6gzYmS4IFmZaf7H0qokj
WPBTf1JSZSOq2nZlPfQt24UkZ+7Jhe1L4LRvVZkpb4tmcBEgFAw9yk2BysUkTEgAwLy1Ze/8F4y1
vKGDpjKflja9v6zl0l8026kyQGkFBEc1ZauA90lpRTRYg36jH4z23zeR/ObNTh7s0gvZcgovRznv
H25IcCj1DHvONjcmWVAeD2sNXmpHeGos8Mn96bQnkCDt4430+xKd7Eo+a/Twk32d+mjJdG7IpEnc
CI54/8U/wAWFVa6vT4aJ7925Tj729UrTNsnhZbrLsa+QIoLPocmrJtoXEaXWYSsXAKbN2BAGdHX1
W/0xmIwSfQNr8rR1nQ/oO/0YcFSDdfdeiGNo5f7XwX7FzHUUc+d+uXbDr1eTLKv3l5vUUr3FeY1S
GBqyJzsKHU9VpBQy56Ra0jjc9J6wYyNVzAdx/bFUzr8vMN2xcP9NRlQGdQU1U6RRqF/a8QJv5cA4
P6mJhO/i80rrf26CYu2KU5FvzaN3YT3BzjsR82Gc13CzYEtrlNWnH9edp2xEV8sLv2ngABg6NfgQ
hPy40lFtNjKABxu0nnOQipndKntkMZBEtkjCBjw84FxQHJrfKZUMUXpvUNEzvV5/GdVYl86dDlrA
NRSpdkSjUzyToy1RIjGSsGajbcLV7zB7boLR6CWpIxHvjETs4EgE6T9S3LcFRKNOP3zGBlDIHXRv
EAGcj/0Zof8AYK2/UxFcES+hHn81xqwE+Cf+X2tYk1PLK202IaP4GM6UwUlm4K9WT/wQbEvYMFWp
kV5uTQ+FB2W66TnxkTYAXpF1VPCuPkaU1NTKZs5+BxCBXpwIa3tLzgnrsBibu5HIt9ELac+giTq2
vGiF+p7Q9ZR4L2xg5Yp+vR4WGxadeGqYzHlwjR8m7eek4uFwtay+qD3eF3FAhOd2f9Bap5RtdsUU
A1ompVt4Y0/gszlHLoUGn89SOX3Gi7jkVCjZcxrmrYKuFzlET1QcNTtiRkQV38oEAzlPeg+Wslex
Bn+of+HSEyg+R+oWu7ADftwCVSkPg7EAvVUOLD/sBE97b13mNlXLhl8NzlH8aAe3BhjY2QhOJpqY
YrRnwSBYlwuXRPfVTiavwDgSgsSfvTIMKpI9awNLLK7vdWmXSXF2Ib7/GE/FuiXNun8zLYJyKmuD
q967jvsIcKiTVMmpr/uHW0DoVzDSfSwljE0s1ZlU3HIOVUiZpR1SyUpbAudhk+XXsDhA1GzCqxsj
i/jo/WFFIV9sRqjHZPlanR47DQBz3haKpvTsAMCXlCuLrbhRa8rr0IGBvfzpM52+IThxDIP5SCRg
Dn+mQiHBPknmGJFGs/+OAMACWM4SwI6pciXZtFQuDhpFh4S8eqY6h797q0xbNmFtIfku+LnpsqzV
HbiafV2+pA1R/6iEBoI37gtW0LSUew9FNUUXFzGveRwTelIidBbljoICWmNf5PyNLpZJxKa+8liZ
ScWP/hNgbyZ3AYirc6m+8Ldo/Wr5ruGBDsNIRtbuvEFYEEyI36MrWk9DghH4GI/n/vC1/5Rz6RpS
t/kvVHrU3l+loJ5lQpFPSwUaVynyKGk6Nh/I0bB0KmJtIp44wKPssBTgT1cZ4B9IzxGnqsJTtLnc
STydthF24qGam1L9ovMIYBR0N78aXhGUPuRN/AzH5YPfQ50e9Cim6w3/rbfezaciCXnwEWoUL7T/
bmQsj/VAbiLI8N3akw8UEp5M5tJsIzI+YbdvPGY/TvAtZpnyFbMFFvX+1JlD/hNg3bSKAn7+HlTp
gOCHA0CtVxAqK024ZVdKyBDPo0H56d6wJ6RdUHwDJHLAw3pSs7Bb+j28hffC5E54TUvVTJsXy2fm
Lp9lO4jzCDVSmKfBOMJ7l+kGzJNfMuT6ha2VdmX7hmULO1kRc92Z1n7uIhTLXEx49/PX1oo04N/7
TissxJgBRlZMeib8ZudhRataG8sz1NG0RBpWdHrHabYA/wW/Sw7jrCztz7cvUOwc4TmjxT6YZcfT
4TNXnm7pv45WW7VhJQMQcGAi9SeMZmQs42UTVkWRHBf6h/FXa/RGdxNKzjeKFV1IP5JfwEHcwZhR
mu5CRgOey6Pblzl03/+06D1GnEmLsMLKgDp1Ld4m9GxtBGK4yd5RNhMulReABA8MTJ/+LudEeI3s
VV5+DsT2xsyTAbHGZiD9dTKmju1IsMuQkoN+8jctLhKWgU3ECUVo7oonUSdMDPfXUABrSizjB8fX
JVjNplC4afcr9uVTyiJoQxGLsz01qe6UgA9Ec4mpEYNVji6kwpfrMCejCXBg3xtTzTGgOHzGEhvH
BBQCFQJvkHVIV6fjzDCL62CrsR3MqyQrjrAjds7KNdFqkiM/L3Wbt3CCYs41SR437Wf4OgvS8/ei
eKPeaj0qyD7UgTtaAB69o3unRUmJ5WJGhBYjV5LQAQoX3/BCWcKyISn+2Ncp4L4WX41fJE67fK5T
LNvLWnROyS3LxUGe2gzOfRBC86U+OXdAc42LAJcxXS6izpaVF65rkNgh6GYoqApoULqOSpzCbkUi
oAt5dVMTawTsVo44rWWycxaYqZWC4rZMWPfXkJyUgvgKyRGYdgrFsafMA/DWKnlLwdv4nz88Pa/B
A2gG+nKv262bsHCPXSh+NUUKehaKWNtYUfEuNaASuzLao4iakFFrLs7TuGimKpLvvBEcaS3ribJ9
p++VHmR9/PCd+9Qn7GwHNqfqiY33XPwE+RehdkxV3YqKFt/FE4xNutqQDDjJ+gEyJDVourWxZmFl
3HGlo5VsO+Kb88FNdWCA+S8xoBrrvX4jHbmP+scB16ttry6I3YxjyFpImCLtJfIwA+DKkIbv7vT1
ZJZmmoLhyhMf6rpwnfK3iz4BxrPlKlHCnF1JD7B4Z/eAAtf+ScAOPgwPpxxevgIg7b4aO97AZotI
e7SQ+qOE95hoWju6axOM42AEmlr2e/IVbNvzPR1zVTWOqOYPWoxR0StcI1h9zVXgvezURmc9FxQ1
scbOeT2+XAlFWPS3osfMmPoAn0ptmPHasB2ys6ITqP5GFKvYn3dP9HsmOsBv+dvQaDr2Za2p7wLY
4eyOTRQ8DXrGFNDLKGii3sBPuWNRtKJdMUCibEvNEWDj7bkYZ2u6OQIeR3lQmKp4ez/OPyunSrSj
M2LC5eVZ7uqStkWBUy1teUIS5lRhpUXSSEpnlF57vNHVIxdeYThpwIk2Bc2flDu0TiuaU8mJBZQx
Z6OpFb9ySFrn3PH3yGdYN7bXo1+frfCf/8kAi6ZTpHDHXdYRsBcI4L/imw/58/HeA4vBftNjo4Ua
IuaVoujYVuYywIE4k2W0efiXrDIF+dqdlsRtGFLtc+x0tD/ClVddqnJEd5A6jJ1T5HoCO3nQ0OAa
NY1DJMGa46JSmrt2bnjFwZQyU8xcx171vHuxEgLGChY4RmKcMcbv4LsYeJKx1yL2Zb4hpafBZ/6r
hpKz62xq035l4N+ca/ZUdaWUOkR2rqdWmEW+szSF1nDHXOhwMVa/5KGbJy3FDt2QJd1zbVqLsevV
0YlAkVd+Sz/R8Icmb/6pZSAV1ma9oAE/Cy50QlGol5nXKQH3SENcrNf6+znjKlZyRZpN86KAy4MA
aokikSboMroIC0Z9cqN5S5geUkEF8nFg5TipJZ13naiQ+bJ1HhXBxMvUz3Os8vKWHp5QtSaAHn5H
bVkiCrfNmcLrsQfZypISoYlXfgmTuilYDLgV4kAZJ2pgzs4XTZqTAevEh4IvVRoqPC9virhwMyNL
XyK/Ov370kWPPAnzKmJx4vhKP1AaAYPNxY3EjYFnJ6pUpfBwKLVpTGSR7D3XWAV9pqkvUtaroAzD
PmK+s6ptO8+G4nfzDPOvcdQJmiTTT5SYR5mfRyKGbcPydM7JQATYHKdaDFbX2ig313QMz3cnzz1J
JQq8ReoBqCRkz3bwUEhbM6ToFc3kbqIm6D8NE6Tmlk1LiXdhhzZjilA+Ax/+iR0K7aioAX+JkC0N
w+twqZCzY7+bJRwvVL2r7gVhG9sxAqm+m5/hiekD3wRdxnwzqMPB0V11gg4V4/MJU5k84IVxUC/7
YyzQYSm0HZus0loNXJWHQkMHvgfyQ14/muuvLC7dQtQmAWYc74Dedo3EIWyhSobF0Eayxe7k+PLm
7fGr9U02h2xsNTUFCMym7wrENV/Y4MryutJxD4m93ei4aWD5e45mWb4Fmn7+7ltSwxirDdc5E4jx
cULe6bmIQeqxYUryw4fQ0+4F7OAsu0WpZ1KJcUzT4xIkpwrWgx+9gf6dGBi82eH3QzCyTd8I04fP
P5mfJQR0XjL/lmNyVWgx8lNOaW9F8UoTF5KwjA2o4yGxQSzeWB8TjqTDGlpXYcqDD4nxtgPIXSHr
3eOjfLfr4geekwz9GIBPF1/MET85bHvtB2+tP62bqyQXZqNAR7tRJmu1cRr4SI3mBM5l0XKNutUS
EECezdztq/GBfUsq8CROHK/AcsVetzXWXCDy5CKa/yg1+xTuYT6GSWatx03YRTW+mx1CCkyXHBRc
+vm0DPZ0QB6sSegtMdyxivdqiqNXD3DoivLWeYf7dV+HuN1r3JNGPC+INXq63mVeNNrSN8EUNti9
MwWHryq8PCs3Q3BI4yDkEEsvyo7DfdffP9+40ZLmCy3O+mUCIEI2ksSM1BraFuTAWwdU07nAkhCM
MRlqB2wjEzZSZbkS2lwK0VQ3sfsrhXGJwI5/ZT4MaIAvvyaqKQhWid9/FjcZc16+FdtaGtfBTm/M
jzVBt5J60AoUAd6t91noktchrvEeBE8PKi7o46FVzdQXIVghqcTBvWcASmptafR6VcKye762fkkR
xfA5Nop7FM1vEK2ROyuCTZ/vk1xz8cPX90lzGd9CaNhK8GjGYCSWiCQC5GEEmbshvG70FlnVYWil
RTo0gwxysNcac9UzzsA5FQpkHPcEcD+kU6wnzIdMPgDKflQjxHsVPr88G2xdB1GlPR96Qqox+m8A
sjKYEvOzWXist5SjhRCOgmVmCtAaQRs7WyH7uMfJf0xIBdcz5dypfGKE1eA2DZP8EcPw4hS9khju
hDY0MQOAL8NUpk+vXtQrVMpeIr9rfwsL2uAY2YiHwL+lLc/7U+kLAH7p02bOIF2wNTvwObAXFVHf
T2A/HQsKAOmw/9aNJ267nKrrWIpolgp/5BHsy+NRyM95pt3MK3Sze/Rpqs2bszQX0kpRNeF2IQO5
U32jPjd/39Ej31llXtvgHpi9X4a78VbNsvMDKBiTh2SiRzwg4YcA43cNcUoxuOw5Ex+s1X/IM7ca
cPpLr4Y7SqehaBVDfAG9DIeiNIUWzk9kXoiAtcTaQAyK/PwpTEaTYvM9dJiJFRH4kvYShP/Dc6iB
ZZzMAaq5u/iFyjgtP16kzFTa9nDrDw2cUR1ULMoxgHoBTBgGDu7AOHYtxcxj3IqqQQLN36i/kHd7
u9+tFKFVzr5oTSQ5nQvVsSGrjBeWjO4gr/22Vs9FE1NgKopuyFEB3izLiszSb2q2nAUPKGXBCHsj
uhfzS5xwltYaeovWddQTAbUTbhxLtrWjEQS3G0lA5jMqyaNUxBQ6GknS6XdKswvr5SNdI4iaYG9v
DXR2nTwDw7/+/KJXWUNa4l1TcUD//I8vPB783Z9a0OhYUnCFQ3YiVGq1lTZ98N/W6Se/n4Y3Qf+j
OaQzG2gp2M/t9ACXVuwyK2wM2otf7lU7CAyIjekViBXuXIWQaaMPDCSFjbkc4tEKmIZNTIn3siyA
CoXy1OIDn7WnP8xyxg5/cDT06oiUsfoNzqiDrRMj5riKRzn3CRqj6XGckOBmhqdJMWRpfpgPySiD
Z1bWI4rsYL6rSkafl97nQEvARQZxAo97+PxiNqS5QU1oYFDJ6HQt7lpBT7ogEureD1VHFZiz7LMR
SSDLSvzGeAr75JaHM/rT0qNohr2sy+qFu/lv14aeIGD0/oS0/mVILvILKHS/wG+/D/1Qvlxi2hYC
lbbZK8EaUg9r30QjgBUwAI+S8Y48cJLu2OOkh2oeCAFNjvM1bgMIb/Xr+SJaM2INHpEWfjbWu/24
d46a2usuzk3eMq3s5+gCAqbOUNEs+iLsau1Ctq5SKGr4H3jimzrV/QusVaIvS1U4ZoCxKlfAkmdo
EN1p3QIzhUouExDHMvawKCa6XHTo5zVGT0CQVQ2ac2+3q1+PHRk9mbfbNSVsu+02lDDoyOjpK2NQ
g6ZamUL6mFZArI7UNt+Etn4fF/l6kx0F3UH9IHPXyJ3s4UidS2HxkQH68wwcipVVXD0De01Bvm7j
//4dzETa4+CqZbgb9lsCtNh4D9jx7jvPasEjr8EKVbm0e1sklqtL6Oij6hbYbUY9N+UEXWT6Dqm7
PrZ9BAsxPLHR25HLB/uOkLD3fkX3vtxa5ssr9W6Qv9KKfl3FwT/P/Xc8XLEk1xqBT6Z8wxLcw9hJ
bZ+4C7gl+zOgdAWELRrWjD8PSE3ZchJA1/akM/93Sq4a3WB3dpgAgxqsAeIyZeXZv+vR1AOVtl4o
ul6mEZYiI1NPHxGlnHdL0gLv2/Gc3r4EUUUnjlyqaOs30z/3EDQZjeNnD/qp83mCPw+bzj8TyTMa
yDSmFa4lFN0oGxm+BclLARo6/Yd+9cGJeQUVrT3fN9A/U5nE/w1zlLJg+opGwMWEPfattxNysM8J
2GhV95V0tf7g2heWmUL/LOAP37qXn285UdG1+oW7uKad1mfjNbvV+EtFyBgTE7Gzn5Us0HotuNYL
4oRhPa5iIbV30HhCjsbVv7eCe2WrCctInvlG+W33XbcvOQ/GWBXrG1Wrg2on8ddgmxehNa5NlwQz
rgEHAQm9hx1T36E9SiJesOkrIvMSzCOGT0VCOSLYzqQExEjQLEEmhKkfgnnS+sHH2a9X5dwcNchP
GE4q9uTgeuirImUWvCJC6VhWyBK4CfdVCdjrhrcybkKwAFAZLbxMGXblO2kzr7zx3ymyJ5YuDwEz
E0Wu8GojvbYEXuQXrfBO4f0H4vlEkbVt3yQrvAlvSKBZlZLA36LvnboOBAaimz+SQtuQmAQ1/J5A
o24+F9H3DWWCPqBs+T1exxcBdR6Qwx2RhWpu85HZ+Tcwjx+w0N5E9otG6XoO/Ir5pkGvwzbopa3n
AFZhgWu1GsooLNSmOCf2jSTieEnuEdqkEv9ZoczEJFa3zOdyPRAQta9m/tDxfaRpB1DrAEIWdpWU
E1uMQ3sk1S12VaiKIe4bByNc0M3yUxrXKctV0VeC9K+QDXsyMYW61WUuYJ//dyFT3RudBVaUJ21q
c2FS2TMmzNkWajwcWkwciflehkfQw7ZQEGHn57k46rDsISCvDjDlpTo2xy1t79dM4dyN70t5ygLk
eB1V4uPHw3v7BthkjZMG+RTeQ9+sJj/wLJHXZWs5+W9OBNlH4W+2nX3vW1G3vCH67FArXZcmhfFA
N4mHTwQX07mTW9iy97+cW0akwzEPyQwx5HiNF7fBbShrT/0BZchnUQ1fAYA9V6Ghu+bBQ98EIt3f
cuZ0SOhOePtWIZ40yHTew+MWZlqgldKHh8Cq40xr95g2pxzE9xzCwzcdrtT9JZAYPbVlua4JIhNm
hmrGCYuzM6hhYeM8BFaDUBfMzqEtmjzmKNbiKjDOj3XF1nUrdfnFaJqr4lu3E3oEnETLxGTsS7Oq
OsRkIbbbW2dx2/qs95Bm8cGkN9miFRB6NaMN2FWH9r4WlrcLweT/JyqGi+iE4qXJ1ZptIOJqbdUv
tKLZFfyO8bL6s6MjFzO+xmR51EtwM309qVcIIiCooz3Ee02GbHhZhORjqekE5XMyX0VPff/UBAMu
PXaoCf6Zt9HxxpLdm6/v89W4pUse2V8NNG6mLr0TsL26fgyBF+nc8fJmwsu65KoE64pIvY5ysNJO
/zgO7OG2AxSiPJq4C65iV+5XS94FHd3IUmotzCSvMrmbwBNmuJpugBnb9FZLRNJYiAsc6gggLgHh
9DvVKqSX2A7aw94wQvH0ayywASyClF7AlYCGs1yvhyQ6Kbpxzsk2bRW61I99G5MOrjqo+CpX/LK2
fPUGLnyq3AQfcoCxAHfSHnLwGdBogwUpHxoR/CK3rtHS9M8CoShrr6I6OsRBWzz6YWNkLOdLyjNQ
lUzmY4mXcCNp5wWaP+mraachQa2xOhUHArUhqAs78XxBwhJySk8HnKhI7fWRCr1lElcJNnUqMY/c
rRK+CyboxnblWEydu7JHIRFfUGGTLdZTkIrcla6tbQkwRAgHdv/wbkIPf9JCMYoJjGaK/FIDr+KH
Vmj15+klYRyKOsbCMGzFrjZx/jjT+RWYJha21e6qiQd+ZP47PKUOrPrxlnQAFkpnJ3uZUmzdObyG
s10d6UJEfE0YyJativC2tTtmnpCtdvKT3qrCrHDx/FGAQ1LQ//3Xy0HdPi+czjLd0re1ucer0sPG
XHRPGvzOttgiodJRvtPxRN61r83QlyQofduba4grkRpBDNBCERVcxqVGM2Xvg4hilH3D1tuA0SMz
r/aHbchP6m4IJ65KUtgFdrzTgGJAnqy0hgU9mBsUxdfjllqV+MYaHc4Hh26JxISv7EnCbKcCxVm1
Uc2+Hk6MfTN55bfUrsxi2jJrwiBUqOEfC2jKcAuEtFjB3gzOOJrbuhG9BmoGLCCVczj5waUhfcmz
4LTayef4fw4f5Sm90Tt4NxNCzUVX9Y1VztkvggnqBV9PPagHEpZ6spmDyAQANMkZ4giBoVeXluou
GKZo10tFpN0XIiGnkifd6W+soY/wIDi3mPKMBU3y2lOOUs7H65E+tPA9ZXa23CVUxadu2E6aqIH4
gZB68XbQw5MzNNhfrf4i89thBDsGyr8f4FwJYwqfRs6bWhC0cE4xct+pTGktP9ggHXMnda/ScZeB
ld9wQhFQkxdy9UHGEe4MeXHzAtImcRSMnEv7V9L7vjLgFtOVZpP9i9x2r2/jTxmdKNBXq4DED4Ec
GAb3+dnQpjPk4MWmDOVpQQirSKha/+KxAM2amapEAJ0Xj0KTZHccM6ASSuyQ9g9dwk7R2tAEB3cc
FVSAzxJwcwrPMS7AdG6RUxD17fOCr1RkzND6/Ng+JDQsjces1jIJb0Uifa/JAyXBDPKQbAt0e2p3
LPg0NGW1OqqpdzeY0sbqqSQjNG2AW9WH+8JKIlVZxqb0HRw7s6w9zIUwRTx/3Ef98JI34fX2JcNX
7Jo5lRwk8UfMJq8GmATR+P3WTtzl0iKC5iorIQ0QGM24kPiGGCIztZByrYJmo3UGSxq8MZStWDGx
az4vNOfcegaT3Ofjs5HbpMDfW/MmjWsW4z0BmqWbKE8sf6baE2RSC5ienI3vk+dg8W4Eu+eGr9T2
bhYCMjTYhAhs3xSFHBh/3fOIoq7Pis+yiUhRLQ5DtB9JiEe5JrOTQZhXtgT6v/9V1Sd7CoFnvma0
c2J/3NVqbtiOQZw3UXf/eA/TnnWbko31eLkBGi9TgxZ9G4INT2Lua026B4B9Vido7uhDXOf4Jh/x
1esFX+SRCNauK2t1oY9aBWet030W0ODGectGXPTSbUhG12OSgQyXEDi0LE8X15FeEVJTAxlC4ggF
UF3raDEbWLKhQbYmLJme2zUQMiwMKvb5mgDd5Z0aEznO9Nfuhjq3LzMUEDBOY80xEZcHrWvnOBHe
ymcddpRM1AUT5t8idRGU4Fl2dND2SBKDvLdkubcu2fE/rEmIub5RBfmWWMlbyU8SLrtB3uPHj7ug
6pTPN4F6CldHIvUC1XjeANwRu3sWy10rrM0gFn/j1W3kO/0q9GCJGu0xliHomKJgZJvPZNfVkPUp
3H/vmHKywHaLoHrKu8uwr4dSUu1D8+mWbXAYjtmsWv9xsglgj/EgK3+RZ7UBMvOEdLAt3p5raW30
xBUnveEneFHkZRoa65A2GYI7UuECNLd+QAnC4ptZ5YU89mRDnVRPZ4RYQeaBEkkV/8ckROnfw+7N
4EeSdn8VvUC3fjGF100Xel7rzeZggoEj3jbaNEOtp93Xz9oNDcDKZqX+S6yD2C9tt6vXRdPAhcoh
bbChjLON/Rge7jIEciig106CCZo+2HrWUO9cjqfYu6n3rj5887RE1luGOPH4rSGhA7XMRpOD7nHg
pZ9iTyMgFKSiA3biU5qyt5Y4yB/+fcMXMZ1OCA/kRso1BicjSPbisIkawElLD+X34NNwl65y9fZt
Wjb7FCnqG6RXuxzy3y8BXl7KBpin1dldjFQHXaCBineMVT09ueyYmLQZKReEI4WDXeUzkK5zycrA
sFYsSzPEMmUgDOmmsGCYerhGcX5CG91398XePJIxXfv7kZ7Y8f7vmGnyVq4lNFAniM+bXY/cIhby
IcB2RQsyahNGs2oxRMXKZNJrYK9kBnzpUR7MpmMSjrHrYuayx7VjgLgnMMzNoKok5Stlz92xJWpS
xqUlqLkJpRUGLtkormBJ8OgcEfJZATCiC7FxD95ZZLI0WMgZw7BtTegCuxfW3Xp5XdZZ4tVC3/Mp
HEMY/M7ZbZaAaQh7aXiHTcsOgzfSz5f0sOA7VRV30oq541jLOBoIGeigX+1JegsGH0OZH6mtnFzl
NvOYsKzfPwJZYq/K0wanIxhn3Jy6KdzxahW5YEW7d2Q8/9gyoc2y8JvesyBEfolzwSnKP9KWz9PG
MfjJ3+7fLUfJptk9sD+kgwUKFN21joJ2ZPjDcHCC/uAP1vCiOoCc+48QGfYmfXa/858T/B3TpChG
GYYwWIG39e1eXHVoHOkpmp1rXWQCHDVFV3YaUG2yLC3gUPdjHZ7aBeJkbRa0F1qLV2HY2DVgMWWT
ckxT7fFgW3eXIv0RfYUYwPCTXGMImlUSDovICg0VsliK3xnc9JwYK8gjLX5ZzUOzFAiFbShmjlxS
0e3ZF449nMyKZOZtZeYIfGTPmLirUerrmEChDBieTwKKxhYj58pxv2+NQfK6fE5zoi+fVKKtWY9d
J6x4NPVkHMYR0iOQ+KjQgq7jJhTxZABn2TcV/IhtvFrsxY1QEwrwaAswhbZAs8B44LAtYZ2XKqa+
kup/qs39637F3hGavegrzHyPwIbRhx3modicLPe61h3bFotQCgSkHTbrNl8QFXeX2/3MdSHN9Fun
0YQFPyH0PtLQ0m84Ld2jzU3s8FhvxSUw1gnc9yNkhwYMigjep/+JruM8vbxIbJrbRye2eztuFuDH
0CWcMtOCzH7LYjwBiQCqs90/NXVAfZmhpZcVmfb/6J9Wxl1wIQCFkR7TQDuQuBLGW/tlNO0A2fKV
2zWsSR90qjZpJiNk+g53OFdh8PGScC0xzEv0S+4IS+NLQvgufufbT8minw3BKZBDO9bk73i/g9PT
QbATPd6pSTXSb0x+X4FVKCN9ETQ/bzBqynEXFDLKsB0Gy5dV6IxxH0vhnj0Rq2nX7tMu5qLz+71q
gDBVm4s0rAhvEUoOEGtcPJ3QMouYeAAxGHETFapa4atxf58gZBZQMEz45lldd4lthr2f4jAUPRsC
lFA0gqXUARM4A5SZbmBcnfXUyhEe/GQt1TB/uKaZc+50qeNnf41aQaeI0sfVsX/4DVzLiWvIwgKz
vov1PAxRg1Ll0sFFAiVe7v3QdL0dWrwdEUSmVHvVb0nM5P3da8XMv4g770/RUFlPtZgRb3iw3MDM
LtKcSaeZeLNP6GkHJ0wSjHJhENChJtetRXhBoTJzZrWN0+ZqmxsTPAve5gq+PGAeR0JUUUv5JBfj
k+MshYSkFuKY0TheQUT9dHB2kvRypp2X4h1hOiBOk+lkEkZGPnQGJtMKPgKXoJKUnMuxrRxP22+v
rY6MOK3suk/9h79U8qPqvjRzsRZ0eIgqj/J8zawKxAoQffRKBsoOS3nnb/WSzxDNl01tB5R6ISNc
CKgE+dpGz+QV1w51RtsoohaspFWdLvUEbI/8GOVWF7CUs2XRMAzWeWpB0NBLJUpoRs2ZS63YCjS1
J1/ybFaVTTom7C5lFUw4T7PTfg7z3uoMYqCsjsbR4YXs2I5oU7s2RWGndNiF0kmrTCkUeo2zPNWq
rHlle37zHSUd2NmU7w4XGsfgNOqvm2F5qsPTZ9fdp8zby6ugMwfPopdcEsF6Vi0xOxrdrs8lp+ud
aoHDvbbMpbF42D4SO+Bb2H0NrgvsA0+AXRYLQz1KL6Rd5EvdkFJzPVja91/M6zqtCqi14CE1PaJ5
UjmExfGgXpAc9BtUhDTC17b3QiqE1bA1u81npQ4ioIhmbyCcLghMJT7xhpy6MkW+/md1nxvhxLXO
eFIuj8WNmIQIRk2CCLdVV4NsNrXKKySum6izVTJZ96YI4P2nIDl8fCqnU3HOQaULz8ZjKtXIRadE
6VPN+iMVNrAoDDG85wGZjDOy+UQEMFwVWSiJ/jXmObeUXid1sdzUmm/nRTHYwQwHJKzD6j9yuF0a
7JVScwTnySBjzRSjjX2944Vm5S6L1iqZoZC/buVo6Dopt5psoUm65r9BP23mU8i6sPF3fdRwxvzL
9XI8mWjhnvGVKkP2qCIk6rEHvc21/Xx/H5d2cFTg3Hcp0O7Imv21Wi64TVJ+X1pfpEmkHOoe5ny+
5+v77f/0I+4IW6N/9xSdelWXt+gBrhB3GFFjtGOLG1P1zu5PfIeM1FPYYitFoeXyMvmuEjqmkrdy
oThH9el1NBPnt3YANEoV7lp02fjTG6+tLgmfNF53soQvyS27fb5rwLoAnKdcKI+/dd7Jv4zbEBm0
3uVD/ZW3Poprxf6wTeMFf0nn5YnT1GHkqSha0HGcfypxH6HF6jzlWh/o9NW9sMMtgpwcjCLSdb2l
7uz8JpW2ByfeHitYG1EjddJ5ahDJwiKQKr2/nPn1Y5MzFUE1uOm+zj4PKm5rCk8NTYBLIVdvXr1z
L1bs1OCHxft2sWvnkTKUU+HIeVjsWk3bdGp3Pm1YX+wJ/iI/M8oll3e4sPY59XIIqcpl3YLAvgPC
BWyXjCP7gI5ZAyvHK0W2MxPH0WNCD9TeRHdT02bqBsCZ1Wy3T0b9iS9ydI2ji/pB+VFZOPGHuBB8
cIEW2mVWj+1W6Uos53oLZ6mDEoFTdQZ4TG7hPbUkrvnZ7JJdSY1gfTcOZevoIgP7TAFzEKaebDfo
aCZUZ9g+LXzC0QJRxqa7lauv8yO9ryRze8ORjDg3Lc0wzyQrpjB2EuNzBR5NI5AS+XO6QWGIGN1d
hvK083tvGaJkNODhTTta7mvcN/kb6dzajvGpPx9Vgmbj01llvXxQqNoqtqZVtgcjGIMqyRZOfvMP
vMs6NAshPsQccmXC+K49aTK25vXsP+alIFA7PNZmZzfaM5IIvPPRHJMcbHAAdT7L42kT+1dY0a29
boj9fCelN11Q30Fajj1b72clZQINNl7meJmwzkgTQbAUrJC3uvDNm1wSBDlzNWaAx15ETrKkbmS+
btEh8gis0F7vSB1m8ZakHekEPGPIQUh0PBPnPEdWwhn7Yrsqb4cp+BJlPRnTwe/SheojE5B7AiXF
sN+L2YMFfRn8UyT5B90mnRY22sbnvUtc6Lkca6SGbjUwHFwd40fnOQadMsJWnVVUzMYI+C5DGKtG
ovL/mIPFRkjR+/Jkyeb/PWqigz2Lh7g1tTBtu6qaszYuplqyCozvvoTdOde7jsZpEar4zASYCVMv
9rQZ2XqgEvFiOG8/ifP2jFZXqdUmUek6iB4ElRMS6CMyi7JO7yzIwOQNHB0T2zbEwwdxTslttfnz
KiS8HXx9ExxCwY0h1FPckdHgaQiizvtU9si4m/hWjDneqlBH9JHPhUbyE8cFwxwuoaml4ssEqFWu
kTYLcmI/IJ2pKi684aVyWNRtgd/Tdt1i4ZZeDF4vP6buWAVmd0vo2V0juagO2Wur0twznkfLt26D
NcBLHqXKm9VhejD5Zt7N2n/LlFpNEkIWNb5IFPRswX1EybCa66CzVhLHQx+C3psMZV3kO8hGsNlF
O/Xfg1lyCPQOpyk6Ds4XR7/IgbiiFIN+eftIskBGJtwVCJnk57LXzD9gwRKA+SINcH/7XBHpRpD1
nqzLANIt5SIhnKBtWE4W75iLCXUI56Mpx1wgNVNzgHg9hT0Ya/YV/osyxmCAX9irEfufaUU0DscL
9RYm7CQ6W3NR91pV1M4SfQs5LLEVXqu58L6mQZZFmuaPeYpvvvNGTfM6wfSIjtym02p9Xt1BrduL
cX11GEg8R6AtCNpImxnfetDEher0U0JFF3DHen9QWjs9f/IJiTxAnb9UHtA3tkk1pZ1p3oBhItVN
EONLTtRlAi6dPiA9gQi17+Q/tWqUHRq/P3mrez/JL6zGa6vXx0Fgqr6a7qSSnK6EJaFvfLqu23nG
o2HTBPr69a9wkg0ifUe7lT2xZrfUvduKOXadWjTHNa3glNxcaq2AaAmDjmO0N8fUO+Sy/7yra+hW
GkZzymVX7L8ozzWHy4uy/0WXX/KeYv9WHemF1OZAdsETl5JgNsGtWgjUyS+M3iUUWTpECNAU8mRV
O4DS7UTC6NtPdZc0QOGYu1rIikawZnYp3W/HJI2n25eMYFRwkQqt0+j360mVk9Dos/ayJvbyirLr
nhZyAC5rSQ8YvQqFXN0K3nC1oMmGgP8jx9B/IpWv1lxeHcmrwgx2cgsjslICOBm6SkY8yGzxB3YN
z1agZwrKBxvsscwq2fP3vT6vJFie6lrCUPLkW/FMe6r8Wv7ykc6wvXwcXISWBnU+zZUaHMNj6Yfj
ASYAUdS0LZ08NHu+kUcBtC/c07wHMjgWG/NAlUnIQLz0zQS6rIu6xjNquXAJSzXDNlA00oSSjwDm
iAtvrUGj4KKxRrYX7oy/tF5kd6QioztBF1Z3cTe5UT2UG3MWfL18kwL7vfsZ75sqKnMpiOXAHaQJ
jrTSRNLl/JYW2i5PSyuh9V+OyamjKg2jHg9nafi8l012/dhESEj33rh/pBHBY5MUeSmOCYAyLMXW
bVcHqF/wRfzVUd5WQ1PrZpsWg9ZiXTBhIJXVMi9HGuhXh9YheKlZ53H2Gok3cSjGRN7QC/sfzzSt
0OrdCo+uoyvmBoANLbvuK3r1tRDJUkJCIQls5AtSz5I/CTdNe4XS7eBFdqizDWWQyy+xzZI1Pwgl
nueoZBRop100qC1FA120hS5BI6FdD+N0asTi+JQvGZRU9ZGCQThaYL0ckG+w/nw28OoRlI5u5RiJ
JKPCtee8R4Ff1XLk8NGobCFyheFqaYA57r1fplsXbOcWnvCxPHON8Nzd05puZ7P1rf7jD4Lm1gV1
CFlM32nxmOWTEES13eKb1wT0G65UZuiSsUjMohVCtCa+9+UpFE7WTN6JhIORekH3fba3hJgzEfYU
VVGt+nnksEzsf1devymYbQ6K1Wk7f7xACp68XVE2WkHGwkgoD9QDJJXw9hvt9Hcel0JMX/TJAOo5
Bw0vaUGNKk8exC4PZXfM1bfk3osNKVpQlPvsHDHXHbzSNLlayQHXlU/pNxCnfTMiRUO/IsxIiH8x
Gi2OKpQsjk7FH/BHWu02fdvd/4HetFAR70GlqKNibN8oTC0Toc0gky314pcCEhmorSHql0f9xIdE
0+XJ6QgAwobqrMCmXUC+ULtkFvcXqimoHEto1qA30PAJwQ6G9zzPy280jh73jnFUNHW+rq1EpczO
cMKsiK+r3BDGsndZRmercUuBjS9EI6Y+LUGrOo+ySYySYRGpG9ICHmr8/FU7AZBpjv0NFoAXGBnl
Tnx87mXElyO8oRY/sk3JPcQfdnLkJP1f3oO/CkckYE43AuI/+Gyu190S6Vse01hKFhBl9fSNPIbB
xs/F2z2NNcwhR1PTdgqs8bA2vq6bwvO73P7xyt/ozKDTIEYX/Laz0GVn7PpLPuySQvN2Lo3ewVah
4/eFGurvaNhoyjYIBYW5DCCHTqIN3VkIyEsQHN3hEhIH1SyRagnI8MjIcRgLBGzX/95H4nvlL68c
kl7zwiDBof2+1/m4lNuyd2mSmyKiFUoGP++ooZhV504Z88UuRkM/JeQhzdOwsv+vOFUc7wiAfMIa
UFULcz1wR3bREkI6zLVpnBcMpaopacP2Xp/AwtRdH6aqsuKwN26oPxnbSbhVUWlTwBWwVS/2r3a5
ct1RVHBmOwKWr6/HEPj1PaeuqlMFHynggs70jm+2uj22NcSWvenx7IwMDqag9IzHSjhKbvJfEEgm
lsBNzouMq6vJfJxASs988SbZ7w/bHICcR4QwnPTOk05+v+qma+5TDonu8IZwbuzfeH3agLt683kj
XnrEceXxjGzSIvQdRXSC4PIpTcPZxXoaO4ARPe/e5iykIUJm//SvSFEl53TCWJQ/fBlUjCCV8dML
Ju8orm8AvuxAtEjp80WJcUKdZEUbcTrGK8fs69560hDOt1PINEiFjKQmWO0TD9S9O/d54X4NaPa1
igcGGaVYVkTZueEtdgg+P3aZHhwWq6aXC9aUHg/gMyR9TkwlwgXD7HBwbCIGVq72l9Gx9/WDLJdV
n8tWDNarh78FWwMPtILB+nivd5WnyFTzyeX+qTrwhsNNozR4I3rlok9BX63HdekWm9067rQVekcE
tLXJJV74yTSy/qYFq+zayvTactGNSDXWCtxPBdWR69HNJkj7vUiQo8x0PZ2VNnKpC6tadYNOaiJJ
IvLOWI4fzS3C/uc1GHKDIBwhvX3+yuIGQxLNsI02Hd2rZKDhOHUQWRXmqQZoHOYDDoQ23chvjkQA
2YbbJ+qBRNTZEsxzkuWRjDwS+JYqff/VE4Ptanz4ahaQGUlqnMaSNFemkpX2yyZLOF4wqJG9hTbn
zij5RJ694n/RxumShWc5KOldNFsJwT/whhFVRVLiReROB/Q4FIxVqdlY2BUnk8Lp/rMZa/gCjqLA
o2maKUtq7A/4JOrojL+D8TeZ5n1afT/r1cqXMZHX6kFVMuRfVKY2MwB0V5hnkeNdZ4E6QL3wC/iH
KQ1y0cFzx24CLl1Y7ztKxGW2DyQBRt/o5s5+ahkU4lVDoUqRSQwRipmkYnOemzCYtFo196lMpcoC
SEsW+Dv9IoSEt4Gp6w1oEeAhMLBUhayiD9RNVAsWzDm56ILFhOOa40hL/gUvHABMDdKGClVLUHqC
ldUGERbwJSYgl7W76pjQf8dQko127R+avicPUaoDP46ftRP8bNSvT6CF7++elGaWVmRpXtFkscIu
s+BeftmwXTuadZ/8shheDpCzPuAD+tZkbS7IjF2ph9B+rSj7TzsuRHZyEq97jIbMJzBjO3gLAvmu
hVDDF4hnHkPvDjaaRFS0VQbmdHCVoenNUUNnE+G7ZarF8jqKByqVI6QmrKJ46cMh7grAf6XpZFaG
UbjweEQHysaHfFSXfBTJuyBsNQUhwcd0EpcveEO2t6npraRmdR1Zid9h1r75tjYZR3Pjoi58a92Y
7R/YNm3/UACehHJLxgExJj5q4iMpdOBZalvarFGOtEVcR5P27C3KaROXb0kfpcqEVs70dcPeojXi
x5JNcCMwPWNqwkrW+YOBeuCWpR/GXkO6bKnH0Oy0RMSbUGyYU5DTd1mR49QKBEEQDfTu8mFzR/is
FzDAnrlytPccbmXQ5kMC4KLfDQ9hyCexnVuB8VEM3ju26ASBMmGBrtuRo3V6QlzSYafegtF8WJWE
HQuq3Y8nyIEEn5C3afq7MeC1KiIf2XiORCBMgN6v0JKZrSDIOmeLUk7Bt+44znt3cQ8QhQIGnvqk
7HrupHqb0XEL3BQBLWW7WH9n3hHcamGYvqWxgLN5QpPaWF1vOxkTeTbvRmj+o6Uhe1WMRDgwpDau
EsLoy6nlCH+WFag5BqRz2zMubroNKvlLeORnjrBuwB+fUZuGQt9poZlV3j85v9WxzUtkgze5s3ta
pZZmaCXV74p2BZXMkZ+drGOWjghGOwij9DN+Vg14qZjWmYTEbtxljqQs63HjxEY8I36nqtpQon7W
G1JQVqVthn2lzdoNSDTcLxTaYSDvmo6YBRZbK2sDl5Inwf3s9geyHyEchffhvVqeJ8MjcsLREJNJ
Pea4BJWY7tneKqaU9uLV+8tOozzkFl4jkygKGLko27me+L916+KMxNPOKYxqFGxgjcZPItGa2wkA
res1lN/MQmeaqjnZLEPM5jxqqQ8o554wjb5+tY6AVu/8UekqwWD3sMGSKV92k3qBcpcYjc7M7wGA
PrCoYgg7p7O61+7pNHEy0xnn8uyxiRrEleW69isWXq3NrqnoKi/sYQ/LLgtngl8SsX5ud90yTFCJ
kMI6iS1+3Poi8x4Rqjth0jxCoWUv9Ei8TdfNk75ix0LPL15BU8Dp4xm1aLF/Luv1rPyLegcJzaRe
NflFfDohThqQVk0uAVbm2QLKO08AaVJPQaZ1crPQgKNXWdMqFzTVpFroLxfXcZXYvH0fSwVIIxjt
13Zdf07qrGlqX00aXw8T0PZ1zTF8j+IIzyx+d3b8JH5KiysJUgt9lzek+C6zvFQIdxeOZGDPGKXz
PdnnOItkjqpIBTrUbb37rdrG3b6M8kl4A1yGWY+PIiC0xdUXMdaJxyYPq7YDoq7bYr7rnrHh+PcO
8XQrC3rETst76DI28M/R22n1SxVn5u+hnuXAU1T3kKNwEVjx60lLDc6/6H5MFb0Ieex6IiOjma18
H00Ep5fIjxL8oPvwRyPgXzc/c20OoyfmB8lgDMMXqFmCGAt6HPbwE26JcFKMo+x/BHd9AKLJYqX1
5+Bmb3XyVVSpBOwwjhhd/4QIlvTutsVBkfwJn0otUMxQ5LcWibmt1LRikLVTajttwtqKQgogn5MQ
RlZGF5T/KzAJtiCMl6HldO05E9Isqn5m4c0aPfE6lfCiEep7852LUhEzTFId/muEB5yx1buc/NGk
+7BSy+OqceBoCDVFwgSFxzFUshpIUCSEMfVyBrFdn2zqPg8mZDAusR127n+GGUeYgu5ZvKGBpdqw
LHUHriJ8B+zOptV0msFXqyrLP4/CJa5WKFVu1Ao9m0H7683fyD98babqDp3X0M0mAJe1Ep3drnFK
nVAf/BjGk/sgnJVckoCLk6qEyH5C7/PNgEru53Bf/toX7NhD6ZoxscflNEWkVM3XXpp7w4KVf3Gk
Tze8XXSPLDjTWlFYAMvTVw5OB26+3t3ZTbPBRznU0+DwDXplgmsPAjei05uwxn0G/P0ZcUrGpTAl
jki4ofdprLnyiqfFNEbsYa/NDp5FR16N5tGv3lFM3y2CFCZWlmNZjPpxV5yZVR3/N7eJKHGwWlB5
l+zEbCFdprr+qybRBNL3yQjDw819wDdkBue98+XSQ2/8Qekvzh2A6m2f1rM8mk0lFYhyfYSRxica
Z4l/weZnEIC2q7nCkb+EUTrNceohXDWot+eDDa5DTicOfvlHyxkONFfsCO1r2TN5R40x3wiARn79
J5ucDMxaoenG2eccBIK+ljZ5ePCvK4+KXG17SKZ2S1NDY3yPYRWa2yuCOwbHyaHyH+/l3MLokbFx
xdmo3T7cMw4rWkqzUSoA9+9C+O0y6nxPCilXp81VcieN7WZ3iNKRNPTw4+xy3MhM8FhlAoH+r+kA
RDMlIUK5UOCYbPmb3aRrOXaFdlwnJ1BtBLDbaBixDz3s/6FD3owox8UHHn7r5V1muaoa899ZeJRv
OVMXhil24HD8l4NZafRYvCKbgd42L/mbI2rqGVjTmPu9bHbmoiZ3YzE0vfvPX+/BOFfvzDSfIuhb
GzydJP4eWQIeA8mpLskFM/y76R1oaT7b687ccUMNbBdFBDKW8WNhg3g54Y6VeYtwyr5LFR//stHH
hW5+RtlSoY/zvhms3TEjMabaFBHJvAIjcXF4tGDrHx7NWe5cq3oADnjdApyGcWULwBgK3r9nJ5cO
QB8F8zGDhM4uZJE8wGE1Ql5gjRc/m0bcKM4x27hVVok9OGfxwYZhbNNVR6OeBHgTac14Hpc21sXv
GPV0tQTCQtOxowZHZ5cvwTTUAa+ZklBSiLu+1JcdrIDnhfDBJOpJ6wu5pgoiba1itZmARxgvHpWH
twci2e7lJKggWhMGVhhQosUdrmG4ufV4hwEydFRWp+YJR+QIgZO+4EQL4b4g+PkI5Sb7qLpgDE9k
9Qw+PtaMFXvikMXaAIGk3syxXqGILMZoxmAA6Vu94LM6phkD9U+OcmP9ukaWLQzO9VoxsFkUNxoX
4dY+1P055TUZyatqiP0EdLLpxFfSGky000d4E9qmki2CbMdxuPwdCRDjVUw8rtsE04NULpQXibBm
hjZ3UsKvoCCoFMYZwg7u1AwTTSnAMa4KIqPcyGj3Fd4Wlji0i7FBI6+iZf+r6PNWQxTbK6IZUPxP
trUN5nbnyq8WSdLsLRr4nKqwfW9ggqJDzver82tK4PXsK1CjwOwi8CFCiJH4gRXXfWzBPLecy1o7
kiPcL9GsCuC7hdyLT4eRZ3R4MEWzKKmbaReG2ZPC2RSIHV50Ium8MHnr48vTtbHiGcmjy7A50eDb
i+LQ8xV3zQG4ffchNEPKw9dq1hYUDiHwd7FoF0wKGyW6iTS9jrTF8kvUgTd6o3yDETqTaiSM/9TT
xB5e3hLNBRshz9fBW7ADrZ3JUT6psE7OkGwMuup4EQdY2EAGOhnnsAAStDq/dGalGLprOwKtCXeb
hjwOM3jf0zpfjED7FcNJ0Um2WjO4HmcRgnve63tsI14qlWqQmgqjdPHJPW7fDc3XMeWO50jmCZsb
w/Ftvj/2AI0FcbaSXP0xJYX7DcT4ex+B1xbN6sqcYo6dM80dZ3L+L41xFARQ2gUjePAdwbo+CtM6
McT2h/W3LwcxmI6EFJ2CpseQrff95zP38xW+yo8hZVxy8/Xd5MXAE3te7YIEdJ6PGUKJXIH3Apz3
f2y4w1Hc2OfDIDbCjy4QXapJf2UBc5bhjSInPG6m0B6jQE6NROYUEQtJUgwMxuoeqXYcH7ePH+UT
S6Hs6LGsbdi1CiHyE6UU1V/FcvgXgJ9YeEtrkm3XZtN6YhLBENOgblnEhESkOdsYbuXU6SIS5Mac
R/Se3c7s8O6/MbRfEtXcD3eD9jmd3kt91I9coGUlYrup5fryN2C5riCd3oP/na1CCSlXc9n8k0GP
ADef7KTFDciHn3zzyDD3xWc3WXJ5gFtJau2e4BpfEOI+27Kk0/Dq/j0olSb2B6TYdv0HNL71lm0r
2VXp8kyb7cX3g8IvgDslvcssMHBKvfhjuU9mM8qJoqpx801btggnEKdTBhxzGfw1UgtrnawEYjcy
ItJ/pZkyZUXaJ/bVRS9jo/Ee9yXzwE5+izbk/EvT/G4eS1rH7KYIBF85yVujuL9GD4L4hubg86Uw
DMc5PQM06ry59nyWn/RYnvryGOeOiC2J9h+mLGC0848wwaTfaxR4kQ+NCj9wawq2w2o+XGIrBDFk
Q4Mcf0Qwpa/5CTU23nlnGrI8GwEYTBl+kMuia/5C+JNtPpZdV0buLRrbiFWjz7hhHljSSDJbMh0o
gkBD15XFj+MxbtNpl7jXIxZDHf5S8JxmlaxJWicvJ5oZ5odGKvVBaeNeAVYUzStWhZODXx4Wjcnp
spQaShUkuoPZsiTw3W6ZgvVb+J6lRLt5SXfFkGY1aCYQ2Vyi5CPGajdI7Ryp4VoiPKy3KsjxoLJA
GYp60i+D8l94uRlHysJj5M7u3ZgXkO20t0JNTJzKtoB7Sxa9qznV9Nt8sbMuj2U2uJMjcxaKNtRd
/RS/E2glfjJVhRXZ+SZIAJcHkXVQveBF0I++zk+qS4YzO3cb8Ta8gfBd0Thd4WuKs/hqMmCFIQV1
R50+AecObgdd+7s0AjfywhTbvaQPnmcNPVq/mUlnKP+BW2skbuK8HvjXwHS7cLn+2dNzyfD7Z/YY
RPx/jLBqPwABtLHoaD/iHIsrreiRCZuMqkjai5e/8MxEw1D+0UaIQO1EQwjt2MJXY3nKxe1/FFck
oztYdLSuUKEn8f7eQaGm6SwJpTNsm++RNoKaMzH1+XwvpQnr35S6WGDoYlgMBLlpw+ODtvf9E//R
hBVklnQkkIpIMKpXvt5rADRxjM3917lPVxGptoPpzmjPzCWpKXryEp3kM73cWtw0GmESln3KI6kY
hYfrq5qgNLd4frld0Hv6Kkrigo+4gm7pC/gJLX7JRHazsRCj02tPFjJ+OBFvR8G2JgrkTPyi5FPN
iu/konI2fiHMKHET15Z+ELg9TMn1IQm9xV72aHiRMxYc1QAPCPxpW1x+ZzQNh2jNjsPxPNBtTpb8
1KAmQHSUH2ZyIlvk08TlJuI3AoqrTtcPdMoGmGAOQIa2DMaxuUdzqsoGBGGQdwLXY7t7x5hk+dbu
ras9X+bGJ57kAocJoO0Mx6xqli0Kfy3FC4nwNfxQV1DmuW5+YmXAI+dgVprbmuIJhrfPYIurM7/2
gikIe2hvk0HrBqVPzi4lYLtLhTjp0CayelQlpQFF5VBHq/Aqrtf8TTQyxnIiwj1q2y0AyxOeKBit
AtL8y7EJqaixZkxI/jILgcUJVyayn+lfsx+DrY8qwYrkhqsSCYMSvWhWb3y2cKDrMVO56zo/UacS
s+RnnIuMlxP5+cbl1FliR7NmUcgCL5UnsJvKngjUvsXLQ3wp0jkQz7Jb/UZ5TW7Bi8FtLCX6sU+2
MKHw/ZQcJ57aoIiv/zGl2C7tkPjLxNjJOkfoHty3mQ/uU0J0aUEO7a6NaEogtuCl0jIO9R9bW445
abaWQeKkHWpN7G2oS0tYAB5kwH356opmhuEj8j9L6jgIVNMIZbfEJOvTCAyaityOZkhKmA7yUXvH
UFqFe9DDBtDLbZBdiu6xEWFHWZoHM3J7MmbiISj/hwhMaBcRcer5V3ZX1J2L6LrzqPKgXONruyup
95Ch375h4g2CZSShaOhkG6oplSPiRryFRtEyakV7YLhIfGy6u0XXp8A1saHHm4yky98FFIZVo0eb
PsNaPiaV7NsjN9BfekUASCRx1jUh2C7/4av4j2aaPoPdroXAMeiKTHYSBNtykF6kWw7nA65ga5gE
Gr4PvUVErk1dusL0gIiJuF/pxM9J5QAad8mA+mJT9LBzkapj5CQHWuyp+3hWh8xWsTelTNfj0sge
p2S681eo0Yvx6zNK+v7P3qPNsWteKae/s/degHzNGbEFa13KSCi8+9vfrJx0hr6O5MJhwrn5Jic0
Zbh0EUAApU9AhNdQ8UsIERQ/GLx2mk7ba7zGa0fC3Ni+Us0/GZ/65Qf1QOHq5xOh1S9TzVZ14aAg
T97aAYjSTA9rUq+IObWQ6DWXgb+zbGeUCyRPcY9W0UHWSg4efrPDA/c8FRpGO5aHMKiYv2Bme/mL
ElQeCbivFgaW4bAgG584kj3DPZyXWFbZgPSz+N7A4U5nq0QxLDv5ORz+GUXYKEtyxHLE0OmqOO7B
WDXcFjxxy2xEC1mtdYNj0atugDGkwtQdLI8xDkBJtAEV8LhGZrujzdf508oE76YFfw+MgZcrQhXx
qrDgM/P+/ciWQeBRhwe/wI1JCOzcRqpY4OdxXohr4WvxbFZo+bNZgTRyrUCRdru1JkbuegNX7dFL
tkwJDmQ+XcQFgbuPiQluzXz9yYkOzndQ4rOT5B38rAG59Or+EL1MN34zI35YRifqOu3tH3LecZK2
V7V2pqFrtlMqqylei8jgYrj42S0TDbp5XRPUscAgIWMW9erRo+sNqZwLZ4f9fJGHrUvqakuPgIrP
exNjDgwYDYJyW9tZCljDGD8dmLK3kAuF4Mt3cPnwIPf9FX+N9QY4aZmYLLyeTxURbqISEtYYL6q5
gkcexcVnYbcsQENEaDDsI7uQDRSOJNnTpYwdWBJUvyNBafonh1u+GPzYuWObN9aWA3PMjEQNtrfI
CL46IRjzbQky7+pt68Zlbmagw+uI2O+dSVG8ShWJ5f63VaOXCnA8w7Am2OwlSvtXOoNS4WnYcVa8
TOPmfrRrVDDFMbAOfEOfhBY9BhxL26GT956J7ZM8CpSzUp49nCWsdeuJv0LmRDwAyemRKtxnjRz+
7U17k7hEG8uEBY4k+vf+0mJJMirof9nJVhrLBaSZK7EjL/dNyDNBdDAcscdM5nTeVvrz1XDaNvuZ
YHYLz90aDCRobOAMxAtJtl9VO/SxnE+cy8eJ+t3M3wUuPCaJCGBUYuxxAQieqAjESdpKhX98FPxa
oY4r+amZl8PQxoZCAMy98tkG1vgPIkh76KPQv1DbovhXAIEQSzXVyYXcum6hXr7uVdTP9C/7gU+x
047/kb+atg0v70LAf9RH6PJPsxJ89w/4Gm9533jSoCnK/1f1No0yd4OrqAxu57yXW17dpQw6IDQh
u0OgY5h+Aqw9kIYgPw0Gs4co8WFTYSrfD4XNeGue7GBroaVt8kQVUYS+lHYHUibgrCQQ4K73iy00
VstjUC91ZoR3jySzlvydUO93K4ev5pWZMnTJX4IOT4svA8QJWKgXDNxZPI67SuqFIW4IA0MSIYma
Ts54rXMz7v/r+8gM8coGd36p8Y2xQ1NeW5HMCghyj6CKlGqJsEtTtvEoB7ZUPX8WkJV2SP6U4NEv
FqEGUILGFKJXimMV3jHIDRCir8hiNAyvyoIw1kkNXgjbM5i0dCJECwWwI9B0YUHAvri4KhL1GJL2
kwk5OAkbMxWqAoA1zIcgDepRCDYFt7ENRRdqh8l3F+HQhQ1XlZljbawj+QD40SaFqhX63dc17hdb
BHET62cnh9rsmYWTzvNfStDeSognkGeSAf9FrYePNiGN9+VH4+To8rVkIrnL4+QsbDbwoX4b0Tf/
FZVSRSkWnNudCRyJaTJ9kW1fRay0sIJIlmK6AHVMGzQnEFMLLGSkIDm5W91WSkY7eogcPfx4mK6u
Qnofpdjk2dvt/Xjpf8Fd0N8MuTmvTygZc1FUvpR0kHv1Nl5UO9qE1vs5u17d7OUTEJM54dOcgCmC
kfGClmiA+ENvPRGkJfNr1rC2S2XuJHidXfTlYo3ujAbOciG+70gOGV/46GTPXjJd4HKyGuRGdDUP
B/vnm53FGVEaFN12VaxvGbLv2p4z0zXLSn6hdmjuoMikBrTpaviz5Wby357n3HULiBmsXx+jyQ92
9B5k01qhCOtsfxvoN6Eb1VKaMbVpUXeHCFtOwM4RkpQFO8rSxlb8nHwcVSpZSjziygau9/D2W+5y
wKwWlXn2vpwO22hnIn6dgmIw8/yEOqLRmoIzjSVlDJ0XD2pp6k3Y0uf+I0eHGmodN6+uVyn0Ok2Z
5U6IWYrFjOzyLrRmvkfIg/HGAH6rsFj529e3XU7g9eBVQyTHdugtYVFezfIYypoE/osSDs63w5U0
Ii/58vZJZRNtUd0JW9pKzYc/5hKjKgSASZTp8uy9KtIrRC6RH2ro4QaIYkH7ofQA8K/yE48TAksw
IvDSwxl4P/ZZJjdzO6q61IztivXN2p5T/2ZPqHkqKtDlQqKLp+7KtFv6V7v0f1Lm/gfzXPqUWfPh
EIZgGCAiXIBiXFqkD1SFouPx+YVZymM5QaGowWPP1qrK2fQbITw/q68Oo9ivV6yPOYqVCGHRg+AR
DHva74WvEnYjrdx59Y8YpV+vhY/liciPIKOeK7oqHmBkl4X+YvvR4xAV3uOYAm4KTTd+8kj2ZWbe
JtwtEWHU3EAy/EAfg9Y1cAVe0bNdTQVL/RasygyK3fvItU+5Ewce3lznbTN7jZ3AE7xfVVUSZ1gO
oGvk0HcgTSidVHg+9n8RKXauEufwXB2i7rzJ/kzzqfVqnuIPh69o2TujbVu7s9EurnflaT7M2y5o
FSeK/Zzzu2xcGpxou/zRUlDUuNl1gdhwn9x9h/DGMaoMm7eKVdQrr+6P9Qm+oVeGIA2KI3sWb+76
6F8Ad23qW0NfxFJfLLCu5EP462xCkiyL/wBaBMExOuLU10FpPg1AufAqV/CRdlIGPop3Ng8qASa8
wW0ltqou5NxIZ5WCL86VwBjwc27IMBjQpgfqfMgxr5CfCSzfQwjSyt5zWBR0ZBzyNujY76uTbImb
sYiRTL7ni7uraa7dYOlgsYsO6EBgmhuFN684/C1/VC4sixh9b3TrshQLOdEorK1AwXmwe+JqSAzl
F2KdPw2K5n32jQI2AxURiS6l0xCXqBUWNAO//eAurasNWPJk0dWMVU0m0xJm6h93yhGTlF0C2qTr
FAJP2raiKTxGL2oFSfnSRP0tc0CrMbhd6TfA7onER3BYKOQnXpwFJ1Qg/y+yO0EFRyGAhHEfTi+4
B+bUIWBZfCKqoJqx5lYlw+g/MuQzk/NoWqrC6EYLb5p3STlmisxS9zTGjqMTlL6sfWJumE6FJyT5
tbIQ6kcly5vy6GQL8as5lC7I+yPDnVBkjxCgQ5+M5O2IXwA/tdI3CoKSAwglPFumdCGFjQeiFrD7
cvx8D/LAjmnUQJv51didCZ1XSuwdKZ0fsOSuulsGBVLi6XqqiG/nWh+wk+VXFsJnSIYZ2yyO7bHl
M/blDMTevBGZ3rViqZLw4tkb1fsgXR+nNyi79Dt1y+9rFwe4i4rKjLNgGJ612kZKwegw85N8Uj+t
KJPPyLQR3er97uW1MhzLYqlztcBozKP6ahD3gUyXxkXUuPjkU/QsKSVht6CSwjYu+k8Cr7Hq1I7U
2gy2Dn6RU/QH5rR76JfXwlrvl51APfQn7kz6JvOsMtO/uX8WTgiAViyPM9IObBIQP9CqG7O7Mrnr
hRBx8AukOP4Bc0cE5EbyrmzP27tu1w1Gh9s2zxKrWf0dbVGuo4AOlntYUu6F0BH8uLO7zzGGgluQ
kOg249PpSM85Z60TJ14H0h1BSRvEfYb7ZATcLAeyc2GgIBbWHLyd30IYN8utLLy9MlVz8bQw2OCZ
oVpsKAqEkagWOBgV4ofBKM+NxkcLEAOdnu77ulPPtfm4t/1CtqV9zaTSPzfl2upmP6LeBWsMdJop
8q/IbM4+R4LnsVX7gaWMVS6wgTSxGgo24c6D3UH14OsvzDvI8KDYVHBKHUCbSqZ1Rl2PDZ26XnQI
r2SArZ1GaDKSYYahFXeMksgVvSiWG0c3P58pUbAzGnHGCqpL0KSVmor1kXMly40zyzyExFMtgM3V
hrwiDaDlpgreihGnh7ceNMIIoG1hO1/jH6l7SC/B8rsea06shgsofZIqKHEokcK+DjVf1XFNfLcG
JS/LNu2hLU+CzacnoQeXR+zw8h7GG2pr/DhGG9Erzt1ngcMzQzBt/3uIxbniFWlMRnXhvL38P1Cu
itbYrjYu3EdVxn7HYncPMu/NVrZvdaz3B/RQgGXLOPY9R2giOu5PXrsqUM6TSgM81nCb5r9vHTMw
mo11vr90goPuH3PLaVf+lXZ7mLDa9L3i5K2bLXkRCRt937ViAMEtR7IiRQ9iamqzgg6XcWA6DmF5
U6Zci4sXmjjhlSDrDJehfyBLjiVWIScISWOGIZFQ/qjfY7g2MC9kgYvKTtRLGIiJvXkPeCLN7RLN
EX0gKEQ+ikP5vx0Es7ORbMS9jrerbfwt1qboAdtZBQ/zMZYcONGo+A01WKlmpI542Zj4IMXdtHBm
aQxV26Q+rUQBAVgrcSOFhWZOSxE3dGXIwl7MjOch39zmXfAnstJemRQujxUBqr3xSZRWsaTteoPV
Ap6TujQGuiQRnhGdNDrKd/iq8lsLcAQpFO+Lhb4xmLaGHzrxa7jOnjpA/mvNFwiP343O95Q6BQNd
YQJmkNBTRGcojugcAxP3rXz7DBSY21xDuDQEcQ92HiV6hajS37xwSu1TQN3RWvPNI2xkHgb8mc/4
j02o2ycOUC9f2ORrnqSLjbVFFa3iqTEDnJv6F2BiSEzzQdWVPSAQajnIcJ1DiYhm6tzf+3R7NdHn
19kDqWnhNuEWMhsoKHFhYotQ+0klKJok8P45jQhali36axygU4ladYOMv286nX2D77WN/b1GWAcD
4OR2cD+dLfFgdpZEw16lPdzqpp6PWXhXwgYZcPsSVYeZeB2KjoKp964ggglXjgIOQrY/ocn3J0ug
VE0HQ7xSIvxFzX09cXfMB08BAiYzFnRbdmhdKNZEJI+Fjrg2LhNu0fs6qNThgXD9/LUGc44laDA9
jlHBIWL5csAYfXulKdK6nPToObo8x1070DPYFcglCsV8P6XnJahy8C6GnktOe7d/9hN/0OpFGoi1
9hLN/M6z3uaZ5VQjl3aqpkIgfnCPhZh69LkIXs5l3A59gbrAZM9bUukFZCkdqJrZnsKuslJSdZXL
DviZ1fWkMOyeyRL2zm3LvZOShCv85sBV7jLH82UIKSVpuWiSndWmNOrCJCBzBW0FNRpfBdG3fkcb
rLs/Q4q5KWJSKjkQbJDUhFVGDU3mM+4+VEHzZEb8xvwBafvrGIbAKUqkBceEcf+/9QelOqp2KnQ2
ydeQF345K644/8MBr1wkx04zV0lDSsZvaSlI1idOaZaJgEAY3WPC8+LMweZs922vpb5qPlc+3N6g
vzNeRzU06jEmcolJxGKXLPrIfrcoDk3/7mPJF7D4wWNmh42NpAqIh+bawhmIzc4GDWja0PS3p4KV
7Iv5wDpseb1Nbgm5y6X8w/QERRY+n9haehqjl0OVl3fdKL208Hfl+DeN2bk0PoYF8SbivPkryqnQ
tqsRUtWkb1Ox6WIeSjRm9i8S2j3kOyCS2t3zazeQpZxkCKpailOABC1vMg+F+1vmAFElSpEosFKE
DkMb1lHGGUtPhYw7OC5dyU7+yVCoIk4ZlPqlwX5lfJ2jeRgyw9BiA/4GwMMk9JcTzw4rBIhcSeXh
yXh7+/9Slyms7iZu43QI5f9hQYOlSG09lnp5GK7/feHo1TewYq7YhbXF8+AHB8uLPrDbeJSjOfZo
P4JyV9K00X+LlPQmc86aNVlyVtlVDmb97DCl5oa33JfPUM2Aiv88NfgSLVpei0me1AS386iMWs/u
krM22ZlrE53X8YVDjaZFTNKIVrqNnsys4FN9uwfqOCCtLfZsI6J+fpdus+1NGL9d1Nk0gPy9t/dz
p44xWeUcwtpYjqH11Wz9WvMIvdL6I6PACqY/BjZMQ+un/zY1TsIoioYBY5PiB2D/cROAJw2xnF1x
9obuQMNEMHwGt+kifTx87I6fpCjoZx9grPR1M7Cg4Es6KWoAeWPZVjgKi5fEVWzrTVCtiti4RmWX
4B1yWGNYTwJ4y2dwxtQ4zkSLioXbRB5RzL1T5UTXrpe0zBUoqmK/sOsvFwRFSNwTyqiJ/5j/y7wz
JuUlVKdfkgd0KL7xelxEnHKuPoZ1p0t5yeL4hlH0fYph/vnyQyu0X4ysgTTkAyNqeQ0N6Xq3VtmF
w5Rcfpb/8OTQHrmP8xvPEIBiQrUpIdskYR76t0NvyrjDtv+Mx/AtY4roa/kKSf3oKxyP8uRXK0S/
A5nmIdugL8pD8+h5u1Q6Nzbx0WyamYyQG6MuFtTU9sg/S8wfXUTEorHrMHls4R1I/SXnAnKx1R4O
haq494Pv75SjCetIP3DYuU99kVQTvQM6wDj7Hxa79LgcGuW96eDUs2CPjzG0qhzlGvZ5eJ4UA2dq
liTRM10Q9w49egwz0Vbbw9Gq5VPyJk1DqxWpiPSKHlOQOP5qOIbdOj0XQorOHuBTo7Q77+aM1ufX
vau7bF/6ZgsWl/Vorv6ETuqA0u3G7DNGBnzUu/WB3HCHEbAl2bO+oeRKzuaUwXsNoujoY/VC3KtK
twJMz9j1UhON8+7slP6yXBgblribNxucLAaC6hMnfSVxNd+ibTJpPQ/COLq8qTbzrnk3k5LEp+qN
vKnsUXWIOWpAcVG5HUFehrEvzdBwlH0rCv/EHkdUdo0NNqMQ/Cy5opyLO4gaJubzheEufh8QtgcD
n4AEHSQDNDbZ6VnoP3ChRemGEvJABXSjzC2nnOmtbs8EYLVw5j9oYa5HFfppl/Nfk5X46uX4GrgD
79N7mCzRgPThBL44iRZrQGw1EauyeKGPjbgzQ4mbcrfW44kJWUa5cCJy1VQfYYRoK5y8Snr+sWph
QZY6be/mt8ahU4rlv/LfzMx6qABOHNw4U8b7INCYMztqsA0G9ppG/dsaR5gmbnQmmbAxEcgUStew
CsL3FrOVhjPmZd3ze8fDUfk4xSRWzNbt12Q/u29hO2tKWVMEnbz5kT1FBFXx+xksPiMEiseIi5Ed
JTbt6m/P6eWIbI11q+sgu5n7pEzlMib+XTy8qLmcMGW0wy9QjiuEdKSAH079B11hLEQmQx1nPm/1
m1VMrqs/2/Ikv+UQGJMHgozB93dnUUZYzONby7S1xisSPwmBmWx7QRTbaK0bh2aWJXCq/kbM7lg0
ZXxnCCeCznv7yJ5zfpA+6zk5mytINABhQcVkM69zTIL7REwk6r7ruMvgsTpgb4NMAZf5Lu5Qs538
Hbm7U6cSZXugcMihPOsOUGc5FpQsqduKAve63aUwbq2SP34RVK8Lc9WRiZqzedk1yt0+Lv8+qU/Z
QT7ddJVV52cf1i7uJWMemu5gwwYatgCfCd0b6M7y8lbLwt4hdiaoPp2XJoDOFBw7tpJY0oUY1hG6
DnEGQI9W9LoF3DmIR2NZXLYIZXlvgoHqsE7kzBp5Ln57UH1QT9e+Qi5uWP5hzemITLuDMi1ppIZp
BOwx8Tl7HSomwPosGEqcHCNuV/cSgHuP2mhM5MUzNR79jIKBipupZFrhnWmLyF/d7Jigu/2wRSwI
/ko5MIwUSWUycaqTJa8ED/yAKQtcV3y5Dm0/a/LsuVE3VbTPiYJySh0D3BuDb6wz0fUYXl2BGCHI
K0gseUl1MmiPz3Al9RbM8o2yPjJetDvksPGf6bbnPks4fedAe6QsbivOrJOOCeNtiDCp8qeFjPb6
dJqgOfiyAC2+y+MXcRL/aEZcrtZn1zWtl40VtPB5VcXp5v28KwdfguP4RApxx2T0zGvSKNBPzbmU
P8Jt6vnBNROJHkv50wVCWMjgdLMZATb0g9UwVjyekKutmqs169tlKfa4z6Q0jYjWnoOTTMxBWXIW
jIFzVBtYvzXNgpyGggUoR/bB8bTURIBIK3nxHvKQBbxdClyVo4reXmkv/Ybxb3RHqDzigVfHNY1a
Uk596utmbtfM4kPvdrfAXP4+e1xiuoSUWW8o/uusiTteyifcwvjQWjuLW2MNVADbV8C6mE1SLJRv
RjFkluf3EVXdIThStX5vlTwKVDlxfqDIaiCWAi02NdjNAUTuvnurkIhvtvJ842uMjW5oFcoGTc6j
sdnRQcng0SNRhMzDU8Vq2bdmfjXH1kRAev/MnxYqCfpaUigV87E5C9d7fB1QFf+4E33N+0iEHkAl
mmOwtO91T0SmUyDnuXuPfwktkWVpklXAd2C6keMMqXV9TGc5dAwv+B4vj43bJYMI499P+RA0Dwwx
VxP5aprLVJZwGXRI01LTg50ZZiMBFYqsEDHOs6JM0RCTo5eb5MCv6dN+ofOFf/u21UNEKa2Vq1Pb
8h8qafYSxthkr87VfzaVh4ElbM5rumEKITml4czcqHdVrOWWgQCazYA9B3r97ho8igoTf8HLBafU
M+f2UhJj94JJN8WNjvpuOUj6Cm1uJu1X73kmfHHTqB1U+6dPQA5YhQ4J7MuRVHPHTFe9UiScgC2o
yq2t8Tmqua5ZgTtkBpLNl6hBxekie232n8qdxkKQyiYl7/MSiN3Owm6FYPVyDBl5KcN7naj3ZihK
DV+KKVPDHzz5P0v64F+J9g2zS47ZbHsbMZOYqfafNwE9gAUHMgeUkLI0NxO3Se/CHE8GZmkIGekI
Xb8PwY6/jODjDkRPRQyBtKkk5niXKj4SMbWNkPHSvOaGIXcUBRfQrabRqEQzGfpRnsdEVQLxHNiX
qxKfNutb4qEcNxGsTOiOwOKPTE88eMethmA947bO9I7dEs9bHCYZorz8Ubax7wCanQfwV3YTrhDe
bXPOev+occwCW/t2RWof7nki0+R67/PAhkHm/8c1HVEIPQZ7eW+mXe8LbVJFFAvM0N1+N3CvM2dy
nrN70nfdHY/QhbjMC5UPeVlBiftaXZArVZqxSoThoP1d1vNMwtWg2wzP3ViyNmYyybmEvEVLAGLO
P3lebvEQy/Mq+IqdOne7Bs4PMCFtxajZnKSU186gk/fzcySEIOCzvVLOT8vKEnoJlVWs9i5xGmbk
bmngJBvLw9hzYOIUmbwlWfzecyIjtGKpO5DumlmJRWU5TqcUcKwZT/Abw6yX3wiwqqixUK43CCCf
r8acGWTQuHHV2AvqUydQQnXq/0hrjsBu+Y7MbpOAB+oHndsZEzRjpf71LzcSygBjrJmgi6dS6C1P
W/PXTUl+DMrEq8a/9bmNi29+yUu/ulzrLegx8cY1IcCiEJaRoAChGYd4e+Pz5O4VtI0VFB9PoDa/
GtFC7gN4kjTJsSq0tfG7XpL8OlpkuhxnACKkM5QbVHLX4WPdLsCPc+jzEVaNCEITfKd4XeE0e6sy
jkvqANm7fV7bj0XDARC5LGhcGGp+UoQfuXuStJqblVJiY1N7Z9CMb9LG6eGgi18jkAzKXlR+87QJ
Sb/6ZD0bJHMiE2nETBNEy5Dw2LjSv/dSG+DwRNH8IQtC8ZLimaOW3LscZlxdf1LdRIcux/tXP/3u
xOv21EiqvPpR+P3t5hurKLiGNCrYsZqmtcDjvvOqmloNgbZm3rHgHroUdxXWWLeBH1QRi05x9uMh
Xgos3rcbGjqhfPykB/gS04NPchbZkRF86yzWCMmmcaGmgk8vPl5NV9SedbMjRoST/neXTspqJq+2
AJP4roIh5/HmGyP2glbJRwyFsS/0pb7CvRBV3FFgAa+xBPB1LlXmBOAO7BA15Dhss2ky1g1mShcd
rJaQ7fZuj+WFvkFAUpnY3pTJkzwoxVHLXBUEaMl4IA437xFP9gFBi9vy4AOfMJOX7idBjEJ0jjp0
Bamakfil4OZH7ZveKmMb4sSo5DSxjLdjPlNa9bcWkUOPsp8YQ3WcCdBGCOtu7pS2RGoY9xc1Q3zx
049kfJ/jiFqNB14VC5wn6ZGQMNOitjug1/V+xJl9Do1eJK+PYlZfVzbbZ+/UivZHjr1DHvC+Wx8a
vKcifYcEGA4XlvZq2ujK/2/F2C0B0SUT5hDycXqvmnbRPY+0Xwt/L5FJ9d930/wkC/xnMn0ZsuxL
z0WoQGHt8Ys/TkEgKokU6bDah/L8zpJOjApFtpMQU8gHC5gaJ+JLY6BQocy2yYrgweujw6+VMr7+
yYvKpbJ9nirK6/RKu8+12x8S6aH1Jk8W0TNGOPty1wW2OF3VeUFlquzaiKtMz57rjpovtpDay/OS
Gl/syonDPlFbwOE8xE3ER1wwVOm2K7JpLiwtgQwzZ8pVOpDE3HIAZJt9DsLA3aRVpqjoTjFjlTPK
o9gyQ6mjjV3iQy17FqrQT3fdXU145y0Vp/rCx2c29GUtJYoSot/pGHyF1WILI46hCjC8cyvCrS7R
te5uzIXbf7XBTlIJTccePPYwgJGHxFRN6Ms0PsKkkEzDZDtTZTobidqS7WAKI1mHcJ98UdwfxOF6
i6+z5FYzV/+6au3EQEfNJXPhydSPfdJJEuagFbIVcGW/Z/64/K2rQoh5TwlSfJ8NcJDMbEGJK2HL
4Magl1MAEZ17iQV5yPx40QnFchcFThGV8XmSVH9RScliIu/W+ksBSRDFh7ROXC2WBVc+Xgrjw9Cf
xm/i121zulNeSnB/5rQ57YtBdqOuRGR2Q7ZnzOZswJCrNjQe7PvbqqUQnoabOrCbkTJmKdVA0EGH
m5hTpKzHjNNPnqze8qzlS0iJTihemYnSRMl+Ng4wigHI0du5PG/vkzpqyWEeLvv1163Y/lg77mQy
cXXalCPryun9qr5NHtOUXLuIfsbjZSoLDzlZE3d9J3hEeu7SOqtq8L+U8LVthUChE90clOWYi3tl
AGdirHyJt7LhMtZEZZBEmQqPAyXCBMqzfHm7Cnbvc0PvNUvz4xWQxLScoGysljG/ScYOuUcGN466
kkynBNhjBaR9n/cSfEgOlJdFA4u/Jzi5y5BepiHRhdMmd75ytTro8vB18LtTD3XZVrxpz5R8ijH+
BPHPOBlfrnqbow4cTmnuvcavCCtbiiIa3KFgELk5Jv8THnTa96h2dvSdQpB4leINl2GvgbVXo2k8
ephE22Mlwxa/HZ5gKW+uHSfmecb6fsc8wie2ep7fXxX+691mPn6s9xbAaePITcwIbEiZ6DZZBgjQ
jLjMmmlDQcwGLEf7bNcqWrkqDz1M799DY2YamIlVYwzlog4H8xSKdl6x7vQSDUFme5uIH/x8ku7W
ewgsrOCN9E1NPByPNP2tCVqvh9MPXj/BM65+UzEjroSjv9BpfbHH6LONM6hi7l3bVSCjxG+LPnnr
hXSYy8ahkgaoJXjnd2FtXxkSCMsigryWIaLdPN3hU5GAp2WY8EwY+93IotLen1PpJkws7g8nadls
d44FY9dCSGwNvC3TPW+EFf9uqFFMubzCdDeU/0uWVa7kyuZD69jf4nLK4sKchy1tvuC+SbGio7pD
HT/1dyCFrvBbY/NM2S33RM3Tg8LoDpzwLPxjKtKg2h7VpANjOYgatw9igwEkYSEtVs5t95LrK+ft
eNg4YUyGCeDsWp16RNhvVJ2A011OmBhs3WftWW+rJmeBziB/JOeG6NjreF6P78aq0cFELD4Byk3G
6v+VfO+SekLaR6ldtCW+hkVmmYEzZQoelsiwlRtgynJuSJH/nblR7q+tWSQRLb9EdR0Pb+NAtyNO
rdE4PexaZBGUp8mIvqshtBaCH4X948l4jaL2RDt/VIJwuFspVYwNQwZgFsJy1AzEZ/MLCrbu7bQd
zhE6NLOY7AP6XL28S6guUos3+tr9jkwukcZf4U3kaETmBaXcy4fW0ytdxrqDe+4ZTGRRCxPZeapu
bVEFrKyuDVs/9anwfVXDqEuYLmn9lp9gAGsDwb+Ee5YLXo+P54FAt1Llv+ZMNfx/xWK5GWCdTzu6
7da5ccvHjyJZ8IiZB9ADRLVo8OR9TWnMtg47dHXFiSWYpA5xqEaRV4GmV702SbU5paVxoBUSA+Cb
1jAynARg6wAFIpGW0HbGj/ZTYMjFjBhf7LgggBhH0buVTrlOAqYP+Jm+DbonebqrUnenJ1K86EG0
NGUmwC39vwKi+d2kJivx88/TNaQNf0nel1o137gfQE3uXk1g41CPqu4/d7iiGvKbBdV/LSgZNBPQ
mQkOrWLVZz8NaVQBL2LBoQ8a/8WFIxthZKfyvvUrZTMAkBNtxAjcevhPDNan/CWq+91u5aPWv9lG
tUEFHnVyA1DEKKoYQj9jSbCfZYt/cZNJ+7h5XJ+6YArWatrYcEiC40gX8ZUx3GwnWK9T5498XPxT
CLtMZFnQl8PTyR6Oa5v1YwFISblr8p+I3mUar4XOBn8xTSqllhxSMhExUh2TnVgTarkAs5m39BCp
ft/YVyhi+2L2LbhI9rLbwkeU4WwPUcyhYGSBfhRYudBnCFKAuA9MXLYeFDQp/NRapvUjOOKL07k4
ynmbzUvqCRPBZgtWufwuWK41UVzgwQWNd+igoWdh2XJpdnaFVvnrBsUFFLhTfBiVIZ3/XQwd+ulB
IWGntqz238i4Xy6QDlZb1myossO4H1tJpmh/4DDRxeDoKXymnEq6RRSavAlh2N0YjALEdeRpe8To
hyuEa1qB69aY0BhMPBC6dzd8gYoAl9lA4tsxpXqmdIwDUfY470hB8ndefGuy/AoZsDnmhTJdmPlg
j9p9EbnD3JVpyfhDqqd75kef8HkbnEWny8SZ21eLA7Am+0njWyunwZxYpkDJyGpmwfAVLd70AYwd
gLh8+Ur2FNHanmCxbA6RN6rYP6CShG+LjyJ0HK5eXry8JGsLl8JgUbs48s7LjIwWYRkJf1mrcd1n
ws0hQxH9t0VgXRnpwt5y4Yjh3WTb4faB8K0j7poj+UvR2iM8nVudaI75Cxa1NBJMS5QIZkE9xFO5
K9vlDetCOZ+tpq/rznqJQs2WpdWll3PI0w8HClBLFXuJKDE4K3FxM5irfhpyeRD4GgwVftvk1MPQ
V4MOlTY2dAjpwk4cAnrdRz7UsQfAcgLLapaWlFw8DI0obSbjwESBfO9rZwv5Yc7yYqmXj2pxvw4T
w5lxdVoA5b3UeacIPOw806hqlVDCHuTHfWWOxxaQxfoslkcepOuwoQ/GjCXjS8uKuEfEOzWGRxX1
7LfI6wmtviubMii6xelf58kucinryrzvFtWRPI76ZjKuI7aDLC2St78uygupirqWiP9LkM7/z//c
IjHuKA7wpUX6Zsj8WekCMXriUf6TPCLgSHUYNUWcQa9CD8y0eGj5Cybvt/BonDGqO2zjzHFDyzJy
6DU/gj4gFTi7koGBQkNH6act4kXRaLlDf5cJ71t2eSyvqjcL4zKb1xxaG4wt6SQHAJP24AMq5lTm
zAgIyleGb233Qst5rhc/anSCzXOlxJmMgx3qW2Nfq8gf+WE2MrAtwpbjeHKoZRO8pBcqqUUTl4ED
iZcnHMzgPGTkpwFHIE7Ms0maOfOFTTN1QbSka9ZtQ7yGu5M4GBmDqu4cgGViRrW8kJRuI1+xgaR2
8IgLi1vd1lER1PhSRtN6tFGyoGLJqw92y2VhUIlRrsZt1NJ1mDWWIazZ365Air498T349zYch9OG
FhJeIB9KkSgLCFZBsEUw1opQd3UFUoOwG8e2Mhas6gXPJmatwcK8rj5dgOhmZzOx+m0f/pAYkFv9
69Aai7NroXWITpf8nQV8d73NczOle2Fl+ZtnMqOEQULtT1Ep3RNVLRtjcuTF2xVJpNhb/ydLlVyD
I+EoGbNv09TkH/F+vH4yw18QebgKiMi86FvrfWLDeceV4Ug6/Uym1CXeGAWd/s8IqEUWOpdTrPTX
cj2iPy+pTyk8qsKghdMhgBMkdW1n9cp0Eu0ExpG2UeStMiDpsyV07z45m+knbquUCz44d545lDzV
VNeLCCDKiAdesh+bkGpOT8kKBfK0MBDgMXJ3vA4gzA564bKuMKkhsf0wIhEXpWe79gO6Q/mTpdLR
wDg1gMY03UIn8OrrhxLr9AvP4MLmcrCY9yVGbtHU8TtiXMoffCgYo0KxugorsH081UFmXuOwh1zL
hvb/bbf7SQMvgxxuHPNZmFvM+mukEmwogO9H6v8wIMDfd+m2+pCC6RVkvJ9+MMxzUw8NhXi1S2mR
SepE1mF4dMrxuPNrBr1fbTCeEmiHIxeu4lBqNRYl2vElPGc6B9AGtOEwseLnRpHxcowZVU3HFZOI
CWiRqOxKAL3t/BXI2xEMpO9C2/YIvG2g3oabCEaJdl/WOCe2vqLMSkj6O7DMhAAA9VmNm0pRVOfP
lIUlT5zEoHvU7zKRhtwAmq3PVyhQ0sSJv08RUrAqn6fglHRuQ2MWKGjmE0O637MqDXtaAOD5OkPW
985CtiKjmT8PEAC2kWEHRCNMjDaX2Q8Oly5WSpLMBRDuS4QwJnpSzDuybMwjQMzZmPTYM9Z41eXC
UzKH3OVTGp8t/+/Cbaq0PIXlFTyxdaXd3ELhJGOK6Z6pIe+VsxsRhtMwRHPhb+WLhxSUY93z7oJc
6LBYstZwA67XjTOlhysXYfMCHrbyOK/fuYYbsU5jNacXntD+EcLHJI1L3fY5Nbpm9U6PH5NTT+lo
YdsA+wlOy0p4zkIP9X8KBdzmI/3nNbH02pWgjoMTKWzC+uaEmQdlTIS2g0VTaOxfW2K29/U0ddEP
+WAjTz31Opab2lBCgsZ70qJJuf4GCHNCpWyY4k/ZPEqPMTZkyGdC7pMEBLe6+qAjpmDp9GvhhrwB
wrgnAcGuPiNk1abBvVPgp3aOFMOOtxY58V2fEJfFm41Jpdqr+1eu8CHBEIlJ+9//U+LxWoR9qc9G
DYNsAOLztRCB0fICEukoDivJBvR66NGwK3+WBO7y2Tdbj9ncf16XDZXk5Khuny5PubKAW/YGeQe2
mqFQ/n7+Qa8nMygmbmCEoX3TVYS8lf51Lyv2gFLOxkAezZQinfJ5nyymjSMlsCVqKNA0YFZdX6JJ
s3giifR+BhefNCHlNL7qzvPGVT9j0wy95JpAxaW3/Hgjrax09ZVwoVdbqqb3BexzcIyzIM939Byc
f7bIqg4pI6J/H29PNcuMmlt2p/iupXEFreHE83y8a/j7lDxG4GNljD5Gs1hBUzV2v8uID3Cz+oCz
pxA6r971HyuZKlitoFsjwRLNWXosfRbuTLTn1kbvSLaFdoZnmITcawroKa+9C5pTv4nLxqZcdo7G
LRysaAjt8zjKFCJ9SOGpcq2ESfWJkHJuY61uLpGgHjG7waS0XxiN9+nR3xOTnmHIazh+qI2WN/r1
kwuwjMrxNouDtb5BLADplFVx6DUt0dOFmTpxfDJY5bX604PNFcVH6ojXlh0aS4yoLrwvCSw8uNtR
cB50SW+7PYbHsz8EqjSKjZrMO/onPxTDVZDxhibVU+5KEaoL33XKm7uNNvYFeeboqplsVQ3DYcy+
fH4/pTlFI0+WBz8I5jo0u6A6bmN5k2MmQbI6bMynSGwJlFuIGVuaz1HL7I835QKmREq2lgn5wni/
lOUX6UKJicwDe3hgEfXuO2WBYB1SqbOB/EkDtZHbPk6Ebl0S6sDZjcjiurqOz5GIwO5RJOzN1DXK
XvLsoQiy4IdbK8zu8PS4j8tjRsSFCQsSxiSTBkcc5Bn/z8Ltdz9orv/ERvXfnfAxeeqsY9/BGLLk
2N5/xzWXv+gQMF+dy6ovVFCqmxaxy5NomN8txTs27L6nudUE4JAgvDmlF+q/kpfqtlzTnTC9Z6VL
6lMaUIckvu1oRbuur0MDpXVMrWbb2t7Mu78silciyhrio5e7fzEsTGN/1MPv298LZFCIhkQe8VOX
pATnDZNTx6XrNLLLf1FQmnq4oUMhcT3LeVaq//o2wrxsg+Xx8/ShJki9XHGPdq25+qzSb4QH2aB2
6VWCz44u0W/7lBmeZ9vPCfuzvyA9HlVEe5HMLHmSRytJCRameJIkqwyKe1qc0GzMTWKDnlFth/T8
raZLa9/huxLxP9ANx07ZutrpVyjts//gtGLmA6exwBEnTGrP+904kLsIRGnTtgTrLPBeqcWDz6/W
pGsPs8NoTDClXJp7Wd4xT2vBsInVQLOf7QBjd0TsJy1KMzwbKGrWyNzCIhjiNAcEFdWKh4woVStV
Yc9OFzLeEfwvqnniyXl90iwq4ktkCY3RuSG7GJ0/QlR8I9XliIohJsrH+a2yJywched7iMYzRQcB
JdOm4dlIhDfOAJK+B/AMjdEbZlE2lCNokzxxgd/k0xHZgsMkb0QTfFFWpdFstyQM6/WDSFlS/ZjU
scy3mS1HFn139bYBfsbI62V91zwSq7x13yMQQUVMlnStu1Kei/fxJXP/8wlJtxc9A588ePlDQXAe
6j0kKNam3Zu2xZwMeHm/Qp+wsFmWs4DtS879519iphphsjOXdFsNDb0OwRCkC+P81wYY4lGN5mnl
UzCFhdtVw+mNqQrtYguZ9Ln/041pvJ8eFV7MLGC9WlEYdbninjgdwHCaHatfNXA1pZrsaA5QLWCV
Z7WHLcFP3a9EbTlOWmjDtZOx44g2vrpP91JTDo59SLqsts0TL9QruFSjqD/rtVUvVgyGB4ORKlJa
Q5ceosq/vNTW5hTicI/wQB4WPKlUyvBrbjYKUANDh5nNOFjv41rXc/htI0K/1VoAKDDAkHkbniSm
zMQoohFxcVc76GsWj6GSIpqh2jOjY3cMcRxSXgw1sLlJ9TIjNHo3I+nyf1DEPXkPZIvtU2pH6Tvu
lhnNO/DVXIKEGEYGipuf1TyPtgi3h3AG/ohBWLXShgBLIgUyjg34O5eKV+JkOVF7bkqOO3sZ+9WG
LDNjwenUX60+du1S17KI8D8NDOXE3OEYWFaKvLMsTer/uirsDWWvvliw6tVPwbVKW/c5M1zal/rN
Yh1YAyOxTnA9d2vilPWIgVsd34N+Oz90s/Bkolr95OjKS5Z9pPUgi/UMgPNoPEfHge5lMtH41BAl
zWfnclxtyLoeLAYBvEvJN1cbrPsUvnBhvdhhSA0j/GSS9fzGTY26Ktagep1ISNIXWuXyx1diGhtK
hwyeNYcjvX9gGW1kuo4IgMa5ni+ON+5yrT1q7Qm5ZmMCpK+PhZ5v818Mw/mWzl2SxwN11f7t26Xz
8lpnoDriKHxnpP8dVuvyWCtTNs72IYOs3kB4NxXZXZR7U2KDhuGumRv6jjFwSoqSEfTx8CJbId+v
ZMPqc0En4XU0jERDeEnIRuE52fMqCF1FMRWCOi4QrhJUHrvSplmN3WsWlVidqIacusRwE4bJVk8+
fxurtHUB/G5+uCUd1X8cH7oheznBLXmt5sJXZPrLcq89xzFn/RxnwwUN5FJP5HRzdhcXz725UrFo
2KZNRj+ksPAvLU78RzLkKQ+BfSkvoNM231VgmQqsrvDPq4wFMVaQ0B+IF7Nh1t9jDv2/twuVetHX
7qtOdSyCxn8LXg8wzZO0YWjiLEIEJ00YgnYMw18Rd2XGhJDqaRtJwrCBkK2b5lPJUmDFiupOlPPN
Z7q6vF6PsUTR4OgOdG8SApUCm75puMBD7vvtfiXnue364jBMh7v7sq9aVUZC2v9xwpMTW109XoS3
WnlIunvpfK1WoNs6ez5DWkAdfAT2mz0A0cytGL5ykBW6gfiygrhl1Hgq4zVqE7wYRN/CLC1E/Tnl
APpIZlYkEh4J0BBA7QgiuBgmWxsPOxkZPs6QknmbaebM2n0+cGMB9kReOi4WF3EjhLZhxMewLZsm
AOctFsICWOGj2qwJlMJKkgyn2We54/75znGjux8w/Ge5UqOoLThNHQJc7l7bZxz4AKQo6TEJWpiM
dVXLTJEkcR4iYQA8e8liF6ysSXiQbJfLZciWWgX4yE01clCqeAweIgM/MZ6hhpE0tIgshKPuxKg2
VH4fV32oCsVyVmcBd0XligEQoBOHqeqp8YRNDuW2q/7y+ouCzyBxI26rU1gnYzjB36mHgBgnDN0g
5MGGrZxHP1m+G2YzwYFw6AH5IF3tnnJbPebu2jFdYxKP4x5lZfNpJmHcARuI9JKOUUy1ll4mB2/p
agzo8aL46DNZpLpa2hXGdUBHxWSy87L+QjptDP4oF61DPKRi+60E4qaGCfEDyy2FY1tvWyx8sWYw
GxofoAbqwNB9kFjATfrHy4YAy7DvipL2mjMuiqKjBb9SVnkTGpZAK2TE7SRCRxNVavJXLLxPSgi6
AZBB4fLFHE0+pt5q94y2rGtBbpyFTcg6WfG9Nl/7lTZV5+3ytnk/VQGEDUKwGxN2SWl76DODjk4X
im0yKvJ9Pxcd3P/sSpQpCHg+wmGhxNkkhCu4vfng1OLcL91CO4Hz4h97QarLy/l9g390GfqZVFr3
4ZM9y1tltqvNQUVsFhW1Dnyp2Z4/vDFSFXMEwfEz905rO+vk9F/oYB/x1eMHOkvneDInF+2IOIHQ
N2TkmreHGYqEiPp0Wv6CQReSL+dHTIhRMWR/iGReW0xTpzDA8ziBnKBn0A8evZxNjZbONWKiMD9k
5ezCc2Gr3Qi5a5YKSmpix/m7h++4hPnLNbvIHTkfpwT99Vf+L7S4K+QRJNqdkdMoA5SMmEC5fZMi
JhSro/pzcDGdO5vAvRn53MhI3YLvlqMrwce+fj5nekZt6FhPUcpKaFxfDue/GgguG6VJS37sRExI
rlqO3flhoBoo4nu2z06oBgZnDW0/p+OoeagtFvCFp+DcTYuITNKQCSEEC6dH88M8XQjQPosNJv5p
noY/XQsNleWLv3efw4OWvlHuPckQSjd6YGOjfBwTHw70Ol+y5BWu7qyu3ySQzvwMhHtkVDVUvfqw
vd9T5smKOG8v1GAo3fUgQOgt+enXWHQp0ALeA3eBgBeOmiTTE+rtCVauw/mwkQoKSd8VeIITKoQr
GssiG/36zUNBIIjgZfxlFKuEAbSPUsWtwhpJ3k7FmgHMAH7GMoP3ZrNKYeZP83CKwVJRBkLnF7sX
MgHNu8BjY9ILb9SB5qGa4YQac4MFkixURHlL/tq2cI7QZLGoxjMM0/tYOuydOKVQoesIOevj3Wev
mkqU/775qkzDXsWfNGra1YyJhHjUbpMkptpMOVkawg39DMkBHOKjgz9noq7DjdWwXIr2aA94IE3K
KzcYeQV4rRuyeg1LTawPCk0WEngh0DpyIyx1hl+aJLb+n9NtCTFYgUx+rzGdf5O+M/3MSjhxoyb/
lbkVV8a56Y7R+3q5UQGM1hWdYAjfflFXlAqkeFqnlxO2s53vCp4fyPXt5f0k9FpURJeFoaMtoVPl
QK+6ZmfbOPJxqjUcJUZAVplGvXWlmve4RNpZ78zUp2fAfkeWoXfdDXXCs9krzXqcbc5eEMKYoRP3
44THDXQhKfNF2wKVv3MRyvKjlPfWrP1G0JQocc4xUb2Hk8J08vPAj5DlefkoYNDtxCibedImzbd+
itkdTycpBhqZUoKERQNFSCzcFZxGat+q2HYe701H4gbaPSFvij0l7RcJ7RG5MV6hVwTNMshqNeJj
zIszwMELln8VtdSWOzYnP7MxfqjoztoxRrBhpe2rJkBzoknX+dshdYZuB4e6nuv1CwnkkS2HyrSU
uDOPZvIuWalnDx+0/SKeYi873kV94ujuWEi5SZ+z5rNu7zhma9IeouEj8X1gYsqmDNF/qL3ze6qB
kNSIOUlOZ3NjgmuSrO6fClbmuv81kQBwVe/rzSqCoC1whZHRQHv4XUAFUs0f2uGHmqNMa693asMn
k58qw27uq2LGOrWjPskwt7YuWYvq1B+IIC3nSLSOXm31r/e10RwCENp4NdBBbf/a9bx87YtXP6f8
+6WtB+trb02cZLuP3DEcqlNmfWyyIL7QmdPG8nJuKQ1cofs9w+TAerFkak/NmNrwF6y8DPcckIJv
T5byZmixJXxVWX+MUBoUd1InV9ZbHWgvU/wR+DGaUfJy+TZH/5B7VD74hdNAXcQpi6FskMdAziF1
dJGTpJ0Bzr20CbnbI7+erdrzPNoGp+DdKyH+tXKVB7bdc9e0X6AxoLPb/QGgHuQs7Xk6ATPijAOm
cLpNUOFhUYljrQCkAyTLDRKsBL3OZv7pVmwdteNcVD9fPfM4Sqobur41IZFm+mGfaedDdzGP8TRc
FI3BtctcA+UNXtDs+8bEOxrOSKL9W2p0s8HVM/ihXusxnKbpi9Jhuy42kmSv+1AuWhiZJ3q0wii3
0t9QnYGPu3D5NGt2grJXkQ5+pk9E/K33A8GAGpNHoOlySNzOOigoLAxQJlDmfUG9EaXRBqGcIiED
dcjbLQVPPyOuIIj8Znpx4zstEelyLIsOA78nCju/+HouoG7FWu5pBPFDHZFy/tEAtUI1QlNQ0gB+
s1uPSN54nGE+ts6xRncFnxvgO4e690ecl+nELArnyt+tpD5jk0n3qLgWQEeJdnlFEOb0g4qBkVcb
zF3Fr1xaLQ5PpUmWtR/yutUcOQ5UVXJEzOmH1a7cj90Zc4icj7qbXGDIMgqyo2OrceCKWVn99Ec7
t+rAXR68yOkzZW9AnHN7nMa/nhQH0jdsubgfVpisbIKXo7PI5IIv4syNjBHONkNQIesPpHCKn4Sb
Ze4fFtcOQ6Weo/et7Ie/06lmeOe//VMNfKev8xZGJIBhGRxMHFbfsw0trHr8EvNyEkZvgwBmJMbw
nvhLLeNPO5QwIZvTE1dtynQtEL2KioPfAiSKG5aU22ZnyB+j6D26JIFp/Gg0ofvuNiXiqOH7UfrC
sRdODvWxL6UiSzgoqAwjvzd3DL3qFm26e6ekSlFyqwVNsfyuxVEulyeOuR7Z0uXXhKTYy9WvqIy7
mqM3M+5OB5MFAaXG9CP3fbBRRxlC9p/gAbpcPbXQig13gz+iQnCeZ/Vs4A/pUBokJcOvkCOdyvCn
k/HwpCww6BbYgjDU7/Wa+9I4FT/HdxGJjsLkqrP9yqhNgjYG977V3aFRsRd4ET/G2CcgMYWBpNei
DdeSbgiomVUUv9dzeuXlyUZK5RRCT//Qg+37O2NehzDmL14DfdrVrjNtJAMlNugMEfL42Vv4hgX9
aqxGmGBFOzvcoDME9/1EIuC4m8ZET58oKdt4IufWfXuCk5jpSAPb0hFmfUz+DNdgBywzq9/S+sEW
8LjaiugaOkHn+aPF8vybZb2CVpRaffeuO1HZKUBltYSKx6/mp94QTE7WcW0cUz7sGLT5r6Sg/8ED
LmRM/GYVBVEIYToLinVfjcl4NmTs5rEa/djvul4dfO3/fIcxTyjK8JiNTM+5HP1q2OEZRHdzaVVC
UUV/02ZM3uKPZt2XrLCUQRsUGrzPdupDawM/m9HW1jq9q+BWc6nYXesuSKPaN+G1Ep2gZPc4BWJI
KmG0dX25PPfTJQy3/RPfm+AV4lBM5za+o0H6IKQzT6b47FVHP/T4+DIeWOCZSo98NL8m+uA3ax/Z
0ZGnJ+u/egLLqAYtuZ+H2U5HPB/BQf2wEXG1Mgzry3sffLP5iE7Q4n4B4U75/IyqyBzSP4lLrI27
uJ/Bj38Q6g3blQm34hXXdGxinmrNbUiY/VGEr7zg9pmd/Aq/+Ftk1h7ac4d5OAUWCKnXlrSshnBd
TO1NctGyjqI8zNoutDXoY4ogsvBSP9CGc/CXK+u6PaaC+yFzlxZ+uqe4h0blD2GYUP7UXvdhFLjF
0qCvn0eKlVqi9Qq6YTIfw1HELj75JQ58Uu07h1O1/9K2J+v+CnvkurIe1/a5sxYKsJeId7iJE8KQ
ohR9bBMySaVodBXdlqdltn62fycFlaKVylB0hMJjXgH/oRPnqcId2pxlgDQwc+vykZzRCTaDNu5v
HBE/kSy9+PF/FjLOwaEin/fqItMjBjTJmmCUkFhuYAxobmv7PnXxp8KrQkF7zZXdxnRUCY8GyR/d
JxeKhqXCYre7pLQXBhCPR4V+m+5zNU+99xT0AH9PMoA+NZH0W31ipen0Yk7N9hOsOK/2sBHj1CZK
0Ng743G8pNQJkrMWOb+alzJIqZIjwfMFo0xY4SJv9ak3/4/wTBAQLpwMKevQ/4KoMkKEhhtmTQJR
1yABOSWTxDtM7RiDzgUV0YZUY/RfswKrcI9C95iADTph3U9XDan6e4/YEvQ3XbFegUKlIt/mKbcQ
t24AharcdaIZsxbYHLiqExv+Xld25JcHZgOKA0eG59hGkNoZZYZKDCQuon8V6az8tmV1Z0KmZbfi
I7OFOkopRrm3o2WGQxQjSV9DiFkMFRZDptX1LSYzNvebH6z5q0ku4gRdIiZNPw7tR84MW6Xp9IAy
B3J1jdQDsUgxSFDMAecYYOG1A9Jeza22OGR9ciI79vCf+qCO8hJZdBtunmTkgaKL+B+SgZv18ow0
Tp/Qx+cQ874rJ9MqV0MMD0tO+uucUXu6IM5+VEU4gAyVyytu/0Usfw/lAgtH3BVVFBfhEFjZ0tEc
PlPSHvwh6BNShQ/LO09Xhfc328CrRHMRMQ3nhSksviqGakhkNn1ucJvJFPgeTNS7JneBAYBCNzzT
5WGBebF8Go1oKLzZ8Zbt1oJGfXcCUguAV1rVH+m2Rfd1/P6Hn7TE4nJZU2kuS2WEKaB5VHgu1Yf1
tVlp4Zw7rSw3mWL40mMbeQu9k/aKQQp1oxJNuFVq/pwp/5MJE6zTPtlw15IYjEn1QmvMxIvcuZGv
BuSVcApjQBSxiy3avGQcj7Uypg2Rmx8OjXb/KYDs8SxUBPZMdokiIKGPPiPWmbGkYnqnbLwXKHiK
2v1lZaP9wIxkofVFD4b01X3kUxL0GAncNEngzvidUfX6xtF+Baq58mXo1wdxJ7+lJeFKZU0ARuFW
8syLz5pjdeWgsJq7DeKHxJSqFSlxnJLOLorjfcWF/Cbs7J7NxENiinl/Qp9ffqimjOp/WS2yO0zw
Tz4kTebFLwelOj4taW4K4PwroJlz0M9n7lbhMqS/UdUpb05Nw7QYQehdKCIFkMZQWmFkhBT7uE/S
S+VJhCtLa226GA7fXfySlD8wXl0ua10axwQJA2EJSpZVEGIbUwH1nfwxke+4y9ynceIrvupssJ62
wAzjQJ//rabdkZz/tb09nIV4vIAHULSWY7yDIBd2+C4+hSjdU0Bl5nRTri+nQrmzFT0PlaBVD9f0
5k+fCpQq/KUZKhEJyHC41ielSsioSxW5hMHR1h1hKN6Z+u9Qn1qZzx0ufpadg38UnVt6YbQ5jWT0
3v19sEkJ27A7EK72tpr1kfmwDCAsk9ghbk/bkOD2vJmA5dqa5DZFJGUYQwdlxtIRA6GXlzwLGutM
X3fe0KlxEUpSRjbo5VzKpqaZ8yyvgul6nlarVc2icUku9af2fPeWLyYDfKR5+8av9LdRqlefCpsZ
C0J9wPznOqlL2YDaLJ/7cz6PmbD8R2H9lS7Fdqt4SvoOuus/tskCkqcqsfINFisKLOTib1lWPbO3
NWeapXASLofNxNLbb6CrJUCeS5Hf6i0Gdaz3hmZ6XLGaD4/UAZ/ig5HnjLvsXFIZQFIx/oB8LbeP
IxfG6DqI5stihPTLdX17JwnrRVAPHkNtM7b0tWGyYqoY7J0w+jwJBQLreGQqwNAluk5QYVH2WgoP
R2DzXc3cq3tmMwez1pnQZPRQXuD5ZS42/uY4B2UAMmx0h9FVMNO/cjngC1FMcbJyycxyHYxcEWRW
DcT7B4QJ6ro3+x36tjvKVKBfUMtW4jWMpm7uW0pcID1SLlvQlJl7vazoFEmEHpTv6n2NSWmXg0bJ
/Ox+QRfMpKT1KVq36zYa9B6bQ/j+cAvtwUjwP7dOTLOzvylBgoiR8YPqfDPhGt4INSH5ARtbQ+MP
EFbdr0E02QdRdIInEVDfxOKxKXy3KMIAKmwgs3d25iHrIzuQsly/G+eyzezSAIUQeiJMXxVwTOo0
57uyyWLbV1qAJh2SYn1QDQPQDjv6w8LRycdd7KO97Frnva1t3lhySMGiffX++Ls/EP/6siV7MEu9
RKzVcSuOrUDeHs2XWdNy4r3qT3SCKZGjA3qIWNruo8vf37e0W++SpTTqh126VxpF5GsJkC7bCOjh
7Z0rDTOT/HWZH/NEhD50cqA628F9/fhZT2mDdcYi5WkmdE402LOT9ptRpk8U3/oOXWzhzPu6ZZDV
l6eTCAy0p6JKcEiQjS7MSuSwP1E42DddpWComWMzGFbhtQrwCOeQu1L4l3QCTpzfJcqjtBkp1P9h
zh+BpmmeSEEBj7SX0gq4WYWac2OWh9KAS/j+sRScLxJAyN2exNL/tjT2Xef4cNbZc3Pyuq2EKJC+
5dNgU9teX7o8kW7+JOug3bsygjzkFhzJv+OuXd5ySSBllBpnQoAVdfgczB7s/IQ4vP7m7NxMN8ro
7DLepRp0ISx12PRcMaTcn6WQQ2HwcGuaoUUSt2nJ/HpHS3I1ZGgMriyVr+WVRZyK0dEUwWbisQD2
WXqO+m2WY6snDQ9J+j+sgoORHIK9r9v6k6emq5bhhFfY0nMS6vquAAjzJmJ7+iVX7FFkWhpNJpY/
SWLlOo0ElAihs9GDyyKr1DmA1S0RweZFa18HhzJzNXQ35kReYGGeP0Ra4eXQtgL2sQhZ0IwxnXMf
QpkhPB/I9J7D3A+vQFlJWvQieHhtGZVuLta9y5RAnzDgG39HzhQGRYPi4DOGQX/JNyYDcECrgEyw
TjNEPjYLSjKxZoit5W9TopDPysO91nqO5Rfy6pSPaRB2817RgHM1PgwrduKB+5MKNP/+U4+UJ30A
cHFDKAKM4k2t5nD24ZWxP/FtF9u/c1IbI3a1/1NGtXlqGOmiK5IckmS5/cGpooIOV2sLGlw12DqL
VV28kZL9cP4Agp2hRlb5ZBQjzI6ASOZmjIyfoLt+S8O2ZLXTW+fH+twtWgT4+A6TIfcJ3cShX7fS
7qZawFlEDV0kwVXOil1SbLW44E9D+09+0Ltodmhw+E6E2ccrTrH/jlxYW7/itkvp6BBC3s3T+9WV
WyjWy18ioSNdZYvsySLpxJ23Li4IbQqxSXu1NibvFgjLGUMu/OASRo3KyC/JEXKkzViHWC3wDT47
s7fF6dSQw4Fik2qXaiqP/7g1Ea4SCvc6pZx32xl8Jy+Q6dgNWN66Zt7WnAsn1rAmr5/S3EkfcsS2
W8UMOYj0Hxqk19CLpOYDsRHFQwm4G4zLY8ZewQ8nzJTaRsW0cJEWjb6JSclr9WlRQwJKgB7ONpwQ
EEgcymrHkdeHWVm4Wxj6nrYcotk+O2XRB0w0/PoxBtYfxBRj1fflfTsEU4dxWMfUY/pEaVIFrNpy
nbK4qlzbA+M3KfUnVO1E2HNBsXlD4nwUFgowSnnkVGU/ybuBvcPetmVdVs36MZnAfMbhWfRcOzth
+CAXWCsPyoT6aYhquqBYH/H5fuoi4Iuhv+lH2faeS614Oqen7ZC1MfxpGohE0+Vxui85vLo/qUYx
/96jzIwVMeerYrX2TUiXP5HB+Ur7BkRNtBfqkX/jhk3mtd2fMoKO7fEX86MkRdZ63PSbJx1xUqwd
7fqykJ8AFWQmeyaGAlE7x2aOuLYGRCz24Ll6bTks3G3mGom4g5DV12nQckv0r1uFyq3/GrtnPk5P
+dnxA4Zv7uEgw+JCsPH+R3QjcwcRFJzQzo9yXMVPM7yT6MyKf/tMkXpC8I2QACOL5Yk3sPs3JolZ
jIbc7Pv/C0W4qRLLSNsUfjUtYniWn4wvARjt9wH9bTYTeq7wgVcvkiQcwxAkS3bO0slq/QvDIjgr
2Bous8MW0eTaSLAotttUj51OxjzhdRKfJkXV9wpJwfQtJjkDJlsY+cmW7HTsXIwwzwmpFbz8FAu7
3P2CUJkrGYEIvf4x9jmvM7AjZZFoF4dXlm2J9flpu2oyT17dGaCUlaxF+3QEol/gFsejthJCV6LC
ANyevqk2u02v/42XV8pPgtYQjMtlnsjtspNrSXGcKRxulAtWLCmD2uMyq44Ocw9XahMUw77uRcei
V+isfpIJcky4f0HjElijGEhG1GhniNc/1l4Og8ra6gMtLBR4na8J/i7ZUj3rkMqLwsx525Tc91Ym
hO+uTl4Y6BDQlgjNL11A7CwkGuGGwIGoWlwBAcJlTbYBxfS/U0ZE3ffpVaXFD5jx4ACknbMYyMzR
CtHUqPYxaTVO31oXjM5KplaS3eOV8Bnx0Wn2HhP3xdgw7Ma5GJn/ljOqITNojWy+Hz938mRdjgXH
Xg3SUJufwPAbAaukYaDejBJ8NlgSQmyt55HsSQW+uBnSDELZhiz1DymcQjuv3VbZoLD3+9CmOfbO
OM0Rh5CWNTJ7x+pFLjwCvgJpiUOI95jegKTNP/8uPVKEYnCi+LWBnRk2Umzh6d55DO3lQ6VWXAIG
ubbPD1qBU5+aW7N8iAg1ccr7LAMayYVOABoamPJcAQkRxQ0PgJJZ69ke84rY52yH44f4fEVXEB/g
BRYkBR47ABcrcLY9uBhLY/IN+RQx2/V5c+LmiUq3gx1gvWGFQKgi0xPpb3Tl5tYWptuSgea/SBP0
3HFu7NjiISyCEmkgi6oz9h7/CbFtiZjegYAOhyvDfQjPLhWOkBiGU41P42uk4/jhJugzKJkePgzL
W+0f/dVo4sVnS4XeVTJhWq4TVPC9f+1q4OiIfnSe68O95VK0lrAey64Ti8xdUHhCa2raEKH3n7H1
cdhMOYn00c0ZPgkzpdkz90EnUZYOFh4hmQQbpHFEjLR5fE5ebxpi15XtZLYYqaUnNFt9mFJzZlaa
xj3fZLBQROUaTQs7kNv/QMJW4Me/wqHBXiAZ7kS+2PGlhDIWWUwSXL0tMaiwAFuBnVQjGT3Y6tXu
OjiCig5yPZ1sum+q2hsGE9HmdU9a4FsbKxMz6apxxxGXWiev4N2dGPwmrm0H6iL4Z1a4eTIlCC7x
1WRPtAWo2aaPJhmwTd6/Gz6yUPm9x8kaq6U1brlWT6HMhDunopSv0mLSc58tYF+fZK3E4mOoS29X
sRyLgDGgkh+GEQJsmbLuPJZSV8FGbdcv4icKsgzkuj3e0xCDsC0sI5wH0zAkMwdAW1WsF1eU4E7n
3FESFqzC0siouLTPPmngQm9fkyRaRb0PF6HYu+tUd5G2XJQVcnjNQz1IfqN2Z3jLkcGJfMdYmA46
D7d0dLMtp4i2UdwB0+SMqsJUUFOxXqn8PtxKfQsfQBBrx7DBZYpN8qk66CF8Sp8jOdA3YZRa5vck
vUg28s2dnomKDB8oVBQ7fVohiP+Wq9VvwMGiwyoNkDrVZan0mfUoNo0buRUhOeYlgiTk6zRLPhlX
cmYtE5+cUeTxL5HFBm8kfQntHJ0bLi1JnDbxWJRJ3k9ULosdQrn0hMYMlZB85/+Ql9+T0shupLX8
3ouAWlnCM1vWqB2xkqUJVId2qdzcy+O8g3uBbVfEv8/I73JsXFZc70KTXxRQDgL9a3e7FbPLJBvO
mAdkXx1dH86CEICHv2H36CuSnqjWPHpEZdIuK7a2RVLupwnMqev0/yMq/1QRTKDzeSYKG80Cg3Zc
iXGEZP+K9p479uUecbSKbCtHLQzP8ey7XzQHePFSTz4u1ZmRv5aYIWHWy6yZQF2UcouGHMc7Dx7z
D4uW52kQhj581ItU8Os7Wmvmxn11rFJm8FHFliUksa0l44JT+fkRJyPVEOWkEaSsbJniMLBwBaBn
HLUpP1/+TfhG4i2UKA0ci++OxKwWOQ+oOTqFb1Pe0Wt5T9PzEIoAMGV9UsXaHtu3C2NmAL9WEIOz
dlSQmL/bzHh0v0pt7eGtQkGi7FbSX2ySJ6riqX+WaqpwaiWhaMcjESjnH7aP0+xkKwkj5dPG3/Jv
g8HZJuewNwu/MLxOT4JMm10lpj5gGW54nxIpUzaU28Zv2kZd8BBlDKysSm/rRpUSl8tAob5V8nM/
9N3MGQVVNYLJaBh6ROlEeNBqN9CeEnYAaUiyA5BJkUW4tBsOZjXmkPI3aGsPpdrf2xGUKb9L9jXv
E7eEd7yMPzmMJx47LYraQ7WM3IY0qUf9bC+gibTK568TpwXj0RTqB3JMltqZin+NqSqOU4Fu2iAO
/HVelPVF4uapagvtOV3xUUVl+4Ov1ThGzWPmAq1cD4QGJaMGH8OIFG8esKzC/bh5XZMTR8+rZfOg
VzNH4WjWs+jcLLJSv4vtJr7fnmqbhSbrIhryc6XVtypUrBH3QAlDbT0UDtXE/GKha/L3hVT8msgF
fPDjsOrAFyGtSBPoGhbCLTgmMcmrH0VS8vTbkjcWIBCZUFWCNTle41pkO6i/4jxRfByCepn4OJ+i
+9o3OOnNPn+JzxOQcnFy9RJp9ipcygJDS1xSOyHVvv4G8wpn+SrGsyAGuo0j6lNVN1lDQdhWGjg5
rEAEQedHOqF8OHWE9K0AsGJfIk0iXRcfCwKH9/2pkpL4F1tyXt6E18COQU+BxthjViaVmxXMBBNv
joucyTOPP8MeXJcbLZxNMjzjw1xCOQJUaGlXkK3TpKHec9rRzJAnABuv1cFhAAdALJDgE3HrJscg
pxpTpxSBELRXWjxLjtlU7gE3+ONKKfgOo3XZRxJ3EJc+TSxM+NUPFpnrCeFRnl45iP0h3HRslqVD
eVvhylt1gAa4SWdqjnmdUD9TtIKGnN/KisCNq8J1ZTKuqSG2tBtPQ9pss26RDTSIS2uZh7GCqo99
D9ydidHZ181uh+VI0GeOTYnzRwCD7i0GD9I/xeSvlY05wpoSCrO+qXDlgVwWWkRlWdRfdEt8+yO/
tZnb7wm8L5RRDqf0FKE2r14EpKi7G1jeh8G65DLME2Fjxw63ZQEKRIjUFB/Rrmuazn97bPanOiZn
Oi1gQS6J2jZZKTnjn2c/SQkRuKTYZR2MVzSzXeI7Qd1xFal3DvgeCgUTXchI7F+RnYfUGT44aeTq
kymtjetme3dYcL5e/11lb+k/t3mYV4lP78OcfvknvPgoqxoG6RJvZ8Yly8FjFqqIuIQvuI4YIJvv
7BKuBdR0/j+mWFHJsL3Xafcx2DnvGZbYADvIgC1LUC7ssmLlr+xMd8y8p9x/4lOvwD4tQM/jUcmZ
rjfsPHSdNL5s4ugPuWkOUjFj16P9AmOj1xMeFXaJxq3p7yFSPS0quakK3/6SHH8VD6sDbvQ9CS+S
RFI5lhGTBXazOQjMWFO3lXgQVfjA/bos1MJK0CHADyTJViak4LKc7mOneBbyxADmHsLpyDG63TbY
AumimQVuDaWDRlmjYBj3rH+lyBlsVdsUpKJIfWw2wf2G213tlxzz2kCmkDf2F9cKF8rYxv4aqZfz
Nfw7xDJ6PWqEYYr3coQbR8skY0uWwgjvRic7J+CCCX67g+O0/f0nu9WKbjme8zcq7T26rttFKFU4
Yizc5bdlTHoDgLtAOQOJRs82d6pn0zznbh+hkA6YZ0K6sMS3R6NsfTiY8F3tRYtTguDBAu7I4FP6
UaqSo+aVI6RzRYtKvsTKefi2PauZTRNNNq3H7X1/fsybmLYg6PCNMgv1Op+y7uQ2wV47ChDZPVr9
b3P8ME2tkgZmAw4tj9XVMqzKZHnIgCXGlv1I2SfRNvV1LK3Pg0G/AiftwW89V7jatbzgv9IHgfh+
vfctef2P2xWjipQ87YQrFzvvxhsyrmZkxaqMp2L2SVWiIvxpt+Td/LP1i1OnU3GJe62QQysh86Ar
777s2Z0RDNiXgIfXk0Fpm1lHJp/nhRdfOOk9KdJh+z4VLcrU6yvhJodfVttLrF9m7QiZf5QKRVl4
DwM2YGTSQoQ5LbGKCzczWCjnOYz6YPBvCMCq4OAAxCdBRAgPBx72yUCmc+ku7Wpke4AWpCd4/qZ3
MylWP0qeVO1sTqdi0qfo6wdtR4zgi2nL3a0IQw2Wm/tx6Zb9sSecEMiRewZ6fA5sV1FkpEPIdI/q
goCuYTPltYPmBfIbfERhVqOUKSG6Z5meYu1E5WVdM7DN3JoqVvMUTfmZaaxZsJNWz6ByKWMk7c0Y
M+lPImCqVXbgHj8giBPKTcYE/ihtXgYy3jvccYOKOhYEqC8rbSxcCJfokoSE00lM//JMHLqYXTFi
LZBlFhGDzkJyB7jwktFNfLgKc9GjebTZhsO0HVV2pYaKq5XKy5ebMbUkPjScdZZrRkXCNrgh+pC6
bckf74HhsW+mPZ8qBV4qQoTDfYielhQQkEY3X9TLdtMr0JEFmoo25+vXRTj66i+JD6R1sNLj0hxi
h+TyXROKZf/PCTfGQs2nOCcfIBbJnVCIOYnhN32Y9NcOIKiL8Mtm1xWXr3x05tvfRjYequoogndt
qyrWBt43CeokZZT3bxdgh0v2nkvi0tPD2zxsPts4YMte4kwuYbdKXc0Sb63VdsBjlfLRFEMEIIn2
1jm1rVJ8beSzrxzjFe+8FlXpOesfLFR7JKi0XKug+8VIZAJ9ZB3Q3IJALvNjtd5Qni48nf9bbh7z
OkYRfDahOUNy1fQMv8VmxTBqxbCMUDixdf97DqV+C5Plh6xXtNOEwt08wdoNYSQKVjTMShLMSOBv
labyDA1B0b5HKZoNMhdFfJMIs1+kslnhe2KswIwoolRNvSAnyfeAkSbA06vSMu3unn+EDaD1UD2Y
14osAhQLTmgvzOM+keiNNzqrUAErH4NmHsXAkI+F74SfDLJRggHwfkF5dLY9RAThYcQjOwWIpL5y
BDCn5lFUUfxT0x8Jp1ZGhk4xtdPCYQaKP/6db+DpVmPxbKhwhC6+DRBnfy+6ErBWjzOLg1gFOzwv
K6gaUvadw56c6hqMegqCs7kaTTxhskTTfssH4YXbn64KaUykumufwewoHD9QN788DGfD5jxm4525
7mbpT4z5aANAhLzodxARJThNn6BzpAR2cduqPlgbIfiCthuRkOUr522XaFnTYtkHS4t9nOkMBN2r
gT3I6bB/Ki3Pr2fieA5snNNBJ6l68TQJdoNRw1sH6OA03kUyLm1YbNoI7+VbBH89fCg+QpyKOo4l
LTSim+t2PuPZenPZqTZbu7iityN8Q089HEQrSOhbGFmI5xFFfS4MqtBmP4kv8CW7MSY2g+CYqFbL
64+YB2zs11ri1GNfHOz3zHdKf4fLyKjDZq8HNPolKVfqBLUU0czIDMWjStElvQ+kK10ZrtspCWNI
/6ajlBr9vbZ51whQ0yNKOrfQpj5BNBLP1neBl2zERxBvfJJJIEnEuKrOJMJRteJJcX/2+m7iD08j
GAQcRt9nFgiRRwu9SLaKwqn2x1ZIX81/AVYzIyAZByjD1eYCXOf9Mi5/LXsezqtVyBT2oXVd2s7b
nMQTZYiS9ZS48HN4JsZtEnsH/sSHt8YX63V/mPTnVepVHvCtkYaqGtvFeH5ZPV0a+0Y6le0mk5uy
PuwmJlmipAoJBbpr1biZ0FX/M2UMZSWKKuMmHroBQ6jSqmYA75OpVuncKSH6jbvXZsc2lbHe8wvK
bY9t+tW4brkyrP0hMGK4L2FZQ2wu2GojWmwHjSf0cwS+IkSSLRuXo54hoob/yj8/AX8Hi31fViG1
PP0AFI1ueNsQznk+xo1OXvuMweYO89YVuap4bUgo0Hk+wnSdIZqrocYmpawwQc0COGiYbcjI3w1j
+ER9NvcRU55M2G5vn8r8cFfyL8LnKiGpLoEVZ+kRd5/YXwNEeFCQKU7hgkPScvwkuXpko04i1wdF
33q0t3hORwcvyjtQMep6cLdpFLKR4btOZ7DRwur6VB1XntWxZWHHpNBMmbsdBl33mvmnRfFO60s8
h+rOFogE7ETzM8j6Wr+Npv4y4aBaygooGrz7cDvQYvK3/0tb14cd9981ymcuJY0miNjjsECwbfkN
lQthexaOfj0P65Mvnq1xyIpPvoJ0n1I6P7PkQon1Ga2bF3hKiksceY0ujK3EVYa5SxGzgdKsV/Kn
U5umsD+EQ4+ShafcLQxqR9O35vaXtR5Pbl6LFAl0D+dbOC9DNuVYfpDloEIoFMEhxoYuOWJUc6M/
1ZZJM8YdQcWxpiciobaGooZSZSStcsZKeuPh8qAPFG0OqUS3m0cDTSvHw2JqmPIER6Iqa6/Dyfl/
+QFj568ip5VFf5dBsJMLIvbn45z/e1B1OHbzTehSBg7JcHFA2VA5ztT8e/kLgbWTJxheRWHeOYJU
ggocMww7VyIQBZXciaHgymfC+pA3odht5z/K4g8ORPkwggVd+ySPvFDGiuF7+1obDHoQhI5zNZxx
Rw2tlIWJgb5jXGlzhh38ea7l80V1nXkMDoLb/tfCOZbodrdz5ssXudBSYai36t3dlv/kt5wnj49s
+pctr7779wM5KqscOnPE8SFG99YmkzeYT6pqGwi2rnVO0C4HAplyl8up3hzR+rWSYm58RyytGVSR
H9K+LRfRZYq+A3rRXLM+CEEXVW5sWWitOXZJXcSFK15o6ar8c/qgXnZsaaINFZ8x4xciLgyj0j0k
qtPGg9fP9ghMzjDHt21uwXU3K3F0v73x3+mUTLJlGPycSWUR/yf6raWAUAvHvXaWTwNuSBKbTbtx
ADDOMvhT0s2aPWcaMOMVRlYSiwgmo2f/Td7hUUUhMlvP2EJXnzYTUhNWcpA3nIrYY2187fddSHTl
6wJOAF5N+jv4/r6qv7OWdrBX/CXcisQdRu5D7RV84Jop9PNUzEBCavkXmx++BuRoeATZbmlUcfAi
AC3mZU8LcMHaFrKdHerGBhZaD72vISQ+ARB42xBsZnBMC3U/r6JAdAaWxaGSL0K+V71Oezaj1End
t9vkk5qRReLCa82pV9yHXyIY8iV4z8n8slEAhSDxXOMR1/G5UBY+vhAq2MAFsZLtuPVwkUZhrqOI
ZeYKYCjpZ9ybPbbg5pGCghO6/4HqDhk5ugkcgmPs3w/xSVz7/wmQXDrCaqDtOZ1lNM+tOggRwozi
r1tVpojv8WrqDePBi5D8LfKmyEksuLRNhhyM5FlxEJU7e/nqMICrFdxo+hoa5X2xsBthsK8srQi9
yNk4RR2inN8SnWYWo6qcumf+HHp2PH2ZIb2uXurlHQGrQSCYgpGI0SJfKAuXyic+e6KRLIv4xaCF
V1qkMU3lj//vH/hKXmDcULrrCoLzQQWxYux3vnUS56qzM0/qoJ1NQEKa631dIDlGJX+c2mY6xUAS
Km5W+Cui+OHFzv0eaBEy+pPkujbfDdwXEs+PS0pei9Gc+v3mgbQli/JN0QG/nXKUxTy2n0iSSakv
HUTkMYpnBlN8JpaSF67DDc8Bh+BhEhOKiDHxHOrAVvJvyh2FNjGvUJnv30e7zENPWPNEiyCoknfn
7wx2X8z5Anq/JSgDpwh7eS2gNnNWWfZjFtpGV8BAd3njt8nV7u509RMI4sLXIj20QiqitSg2yvGU
yP6LAHa5e5Rg+4/oyuOaY+xJsCXyXmjxH6ZqnyQEx7oLCUQv0P4QGHeyhzUJhV3ZgzSQnAkRgWiu
PaQ5TkgXo0R8xRDYg3XlAUmCk10em6esFoOiwiroo1KVj4MlP/Pt8NMK/tDmVukYZKYF5oJ3RRAy
EmNLva799lhn6Bg4JltnoES4/lQMHIgpWI4ZWwSWzNPlfNc5fbcLwsKBeWPpVlTPZthJq9Mds3c1
dSZVwSzciTFw/YaYOtN4pmWnD3rf+JS9tDy3bBiU9hzqDdpf4iKwSdBSoWryapsSsIlqf6TFiPlt
jFr6yjAMQz7bbeiopIcpXCTXvKzGSg1bY+2K624hnMtyJFAm7PzxyTZESDkZO7nv2GFFMZV+o2gj
mRRmQBaUe1KxiJL5a0rvkz6WYr7wn9lumZKtKOtlo13roVTCQItthvpDlfOg7+VFzU//Yn2kQnAl
RgQrkq54hHsqF0e0S9VZpmzWo4Qv9cwjXSBhYU7FWzrRV/e42r7spUq9uJaU8N3xOrobK2kGwacJ
tKj+XcNE3wim0Y36gtSdYjquEzU45K3ZG6nKSpHJ30mKzAe25oI2TJcyUOZNbPwWMUF0WPOg8XmI
Bofqp+4aCcQ/t43SL8ejQxJEa7syKAIn1Phv+2kUfVoznwrfo9Fh1dm8hcrveZzO6BjImGutRF2T
t4gkdVIODG51vfU2DKmjs5do+JrUqdzuxa2GRj7oCryzqDtAepcitF6n+5Bf+4yGwr8ysKCDi1LF
NCJQ/OQaVCLrw3VFJYAHE5OXu0zfCB7pfmSwHUO8CreS7oOg/4WuvaaC96mcAj7DFGvmi7C6/BSB
KFTw751GF1TEoS4d4M2H08QxFnVFxJ7niGF5e+xoWu9MaStgR9Q4nKCV0W09yFwn4mzRu7Buxl/x
23wMDHXeITD4qGm54yhTM1MWVtHlmAUrWfWI6lMYOiFM7+X53lgRMwvGew5I/L4l1J6ezvQGv6bf
f1EFX7ogP487IqvTMbKzGRoeRppE+i2ifFXDRqeJ8g2X6WeTMah94Vu9f6MTAO0fDK2pW23TKEV2
MCNm/hYOe6Y16klN3yNOBaFhM969EII934lGaXGWqSYaOtqbGTUX9qrmnll45NOpRANfzsFoWbYs
mct3RR8bPGbWPQf+qpq2bRkCwGuZipzpMpuZ1rmjy8biwQQ99oxtLRcRP93FPGULsJJRaEZy4XxV
6fSC27e5W393pgkoltk6GDEhLBQIUGf9aIZYekf451VEqMxd9/TxXF2gTOvJ0gRGnKp60/Q+NkYI
OVNYMxxtseGhLHNO3QHbDvyi9KHl6uxB0Ov8S4H79Rf1Pk/F0he/8VfnFO0hATvmsuM1epi9eUhx
dQh8XIBdonYWF4YSr4kJ2fwqzi5uZOJ2t+NsR46mWQJvf8DTur9AyRjD0RGezsfCOABZGTvZBKYC
tgVA5d8QPA7gBEZiu3ouqmzPOWOKfEAXx3HdiWnyaOgP4gMyihJtTjlMNNdqtQ68PYCdSRGg/Ffj
dWXZ3idjVA9mL9ITuA311O5KipHwj1OwH2ZulIwvbGZrrYAs0VR99kuMyGUnY1iTvDDGk6dM68vm
Y2FF3ZnwmrzcFGmBzqLAUNbUed5pqqAl7mlmADchbRFcuubBQ1qZrT9bsOoPxpc6kcLLevLPJ4G4
wRBGhJZqCOxr/SjOr05E4CIaudEHpRc6bTXlUi1YQ7UIhsCjysg/9BcJmHY6BJMyhOJ6VIvwZ0pR
VQ0z/wNpGFqsTJ6evlkYRGx01TUnCkmnWukCRFmjxGXoJcjQbl8PYv8T6WULbkPHNDv90kGRF3l4
CvIOA/j7e3X/0OxhbVKNFZMcWpMwLZJb0727SqQlccleYqQPHGgDCxifRpJTTY4PYaPJyiYLMvIq
YlGvX9OOm/KV4Vzis4cTQeIKZ02pO3VAqbqDKpkm/13WLK9oBUaoXHkji1hzx+MtgFnAUcUfcLQ5
o/ZJiw03+/3UltJyFusQ9XA4OCD52mRbofbVphSILSMaf3XHE5aU10vfPnbCMiGRiuXxml+RjW0h
t2AkHyC/47gc8gQPgKQ12dN5R6SjrdDKFMztR1Qtz/aSb7Bq76y73oxWdDtZPKhIyCxRs1MOREZi
L1jeONoYi+wTb7JP6IibnaQrVkfsfIVNJcaOa02qqymHmhBfVPW0YVnQ0NdiEJBzxcexIzGYUdtK
Txtm+GWfqocZZxpKclWbvNijwCBPoR2jlzYvLgKXH5e0kWXS4/Vnq/4PeYoUCb4M6/asacC6lswO
yFac/Tmuyc2ldP2tIKjqJt3FiCWhT6GJirS3N7w+IwuiI0t8ozWr+W9BxwWUWNeD1BkXMWH/LpU/
NzNjGjNui5LpAFFjLPEXkJmVnHdxzYhB6UUypofd21Y3oavn0YZ/euIIjLhACBCrjsY7vfKb0Iqr
4WBhy+SBF5c7cqy18pMX/HZ9qzkEwVx7S25cxkWee7AJ41bq40cpMQrIxgTRozmYCNKOq1XuJj7y
9Cz5BD4lLmTjb3QrYRg4GvmSEXTdW/1652dUREU/6zCavbS6SUgp5hODCaCXlZyGFBTnLkuJ1aMs
14+2ggQSZjumvZoav3aJQZwdiOLgdYSA6z67uzxnT7376LEXAUwn1Ps8a3MS5Pv2UOKoT6Blyg2e
crk6fmDI94o08xXs+cVidJ1YybDgikwneQEtQ/947+hv9KKptCaa7/6q/3yWPSBWjzVauTOxG3us
/Zgkn3r4MzLaCRm9b4tV4v5r8KfZS2MQBN7Jt0g684sAkXI7NSejs8dbSsW9otIg4x37f3DSVQjY
LDL85wZsoD7Ip0ME1osqcbnDanPqyqNC/SdHjPdkRkMsWDvfQfuuU38s2hvJzcQG5uxGSv4u9UCL
Grri6lzhdco3oQKfjY2gSkMyfw5l2vmKGnKVnOl7+1FinrxY3rc7Xi2RsuC8rYe88zPQnozEoCkD
sHha4pdnc1EgfLl5lntI6TbS8p5pTlr3J8rChpAYK/gHn7ngwXdjlt2jtvIIun5s+j/yFjrk1Q0i
Uwd6+oApQo821EaM59Fp9ZCvU72+2hNpiuhGDTcPIr0LSgw16ubSjrdUXun6DGq+LBy8qhuIi0rw
RMiZIhXOiTpUnjjGiF2ettFuKEjwoTQJmWDY3fRajVJqS06li/+ymHfkd0FfiQ0IITr0qmbXAgla
RG5AO5AYBkRe/KfAzu1HmQ+Q4Z4oph9teole7as2kswYNMBXoKuTEGFRl4Ak6vZkHPi0Bp9ozuil
DRjfUDQigupV6KdbdyZNAQiB61lEvlH4MZyL28MF/rHocBS3ZVkJBD+AfITiPVIzgpAIdfuvUtlz
GzwiKf779Rif6IsU9PROeCWVlW5HxHNs8cwHk/dlDQhNhwnIoAsvtvbxKBezAPhThB47quKWKfk5
pV0wW3qIh6jYOM8ru8E+Nnn5Ed5T51qB3GnD4oQmi9TexkoJUc1BRHx78q2lWQNO5phosGiXjY2p
bdnf2gHgTLZ23PmHjmSt8oAMSiB3n345MBckvyRi88f4Ta2CFgA47W4slQ0DcW1fzbjxIhHHtNKx
nvBevQUk1QHtnCtKywe2EsDvgjaEgwRj27kvNWqQnll53Ky4AijdnxYHBgEZYcDExoXy5Ci9blre
gxQeHj6vQslA6Mwx3O8GysqEbHHpgCc+KI+12ZsWYm/9ilNqw50jS14lo3HKhNXslnmibCOCkSok
wgsRBLdb2xE/jfv/VWcoMV538Ggz+ZKVDuzittA5AWUTAYDn4ikQgsnhfwIrvbHhbs6ygsaC2we4
gWNEnSvxolWHbv9ucTkYRfq38MTM5hkaDFYQvj6QNbjp3s/FI0/1LHLgc/sFqYoNK1bVe+VLLAu7
xvfNCk1H0P1mIQ9KRaQL0EcOgOsDYV4O2r79MWGeirn6Z53IVRd+La+3XF2VIZiPSYpzsaqiD/xF
V763CkdsRzDR72GDQQVDNCvdBFGrBG2UFdvUf9np01rF7viE2Gnt8SlzLGSeeocbNb3FMZfQZqSm
vTgVnUcBvB+gvxEWIJuxtMYxwGYnx/SzO0Qtw5yYUzZUNjsioobJegWB2z8Bb2lSY0vUrKAxqB9i
0ndkFprWWHMmeRBLY4uoCPob5BXphAF7maimNYbQ0MnM6ObXhMLWzm5Gob0Qsek8Id2/XwS37mpm
Hoyj3njAds6pQ9uH3cwi9Af5kyUVJsAMjsonFzDYNCZIlMqJF7oI5siIYOuV6PmJl6itf9uZV3aT
51j2/6RDfl8EluaNPyirSY5UBzIFgholtCeg/S/ecxeRzQApOXIMFs9Ut7DUayD/F2ZWa7ibK6FA
AK7IIJQm/4m8u5o/YChsYXW+9aRBmFXxuHiPiVCl00UfqenR3Wm5Cnsl14NuGPCIQbtTK//+RcqK
EcbWPZsThjWLaNFGRnUw6oE35O3gubul5Ad81KtPd4ECxWzZptmGvrj3VqEpaf1idXgfcPkGcTjQ
b0gDZiXLt8YlE/LcZ7laIrrWocu1oNOCnkwM83mIGI6HxmBkm8hpnJOV/tAvBdFJDxFAkkcXLXvb
BYnBJZeEQNOFfFRUK4ay3BB1m6I8BTKNgi6d9b+tF8eT7q3NABfHMjToWyW4GT2sli8cTfTT20eV
eLQFE2lFxPwnTfCDGteY+u7yp87+UAqJ0rJnBU4o+bPYqY7enCmVj/cp+MyqEpbxMZCufUbH8pd0
o5LmCk+kN6usv+8ddEvMRDkFmCJqamTSvlXaEKeu7fXVvSk0I/qUIl7ypipzrmjr2HwPeraGeWKp
MO+9nXnUuxMTXuCz6g2IV2XoBsPSJMDnEgZSCXI3zCB0NHGx+uKFD+Ko9JXBPcULb/d4LsQSvFgC
iTkttg2Mn/ldfr0fRrx+AbRF3eQQPn0btbtUj3hizQmZKipmtYEzfEzOBiUIU5NAXR3t0JbY+rjN
pVrELXiaxPK8YJwIcMjbq2/mZ1ioVAfgUObTss1I8qKbscvkeZFDcbeNkN1tHkhlWLT5IljKkSCT
lGtawn8FkTb3gjy37UmRuvJk6brdSkzmo7onReFixTdn77/nhYajllSjKKq1NinUph5Q7ZsXjfmj
I/V4KeCgnshAaR/BZqM5mEqqTYKWmE3YlcqwF2nbHwh02Wek/gO3V/GJZN7QzSUHAnCMSfTf/yif
Re4QaqD+QbDNAry3KgxtnBtAKTQjB6x6t1L+grTAhraFGnhbykRIHzINx+wzUot4qyLjP4yYzKYU
LsOtl83MHHvYv/tlNEmxMoGRzOynandIRofiGfkXLwDd0+L7kgUofEZNEjIcOVIPO16I7fSYAcMY
UpPfNgKkKFSk76vshfjQDsGgMcU53UiK07oxlq0eTK6brYC9gW4xIeOeQuvdhi8DIzFm+OCXwUef
17tovlKgOzKYVMfKu4Hb06AyO8z32er94vvwyfoFElXQlaB/TH5uhHKaFB43arR/eaA6DqBOWocC
gglcmBNcjhmOGiO2MPVKC8/effG8sSJ/NiXLEyKQFRQ0Pc2r+nOgxeDVNwvHu1B/jUCgBcKePrJt
hRfrW2av1Xo621AU7LgMzRBBInIxvipoteL3V+yeWmA4A7dd9fjBYvwz6xb8jWe4foL6b2lKOIqK
u2Agj2Gz93pnnwoothcoVvg4ihhtNpfUkA8+ngbolIWgVKx3XgPzwyolbs1/2HXSUB9TthrlMqFf
3+9cP7xOSt8/lUfHPkEydms1+BnFFQEyFeUS0e/gd66fuXTWQebkOvmZNZeTHKnOpeWS3C8cDG8X
Di/DjYdgmvtUlxhoUqVHwfNp2IEv6vAxS07dHc9aUezXn4ADpCZRo2Jq3GkRUKWHfhPN3W3drp+0
I9bOLCVhdnTZ6fo1JXToOrfH2NokSVvVhmhyLZPRAidQZT+FYxTsxWc21opmLH3eJPSDJg+1UCSS
GE0hW2+OtkaZTQVz8wHHKZZsOHJ/Vdsgscek81LoXzSiAQO2qgzoczqsBlH6ms316/FG5ylgxHm9
6aWPE/If05idhB3ayLTqhJVAWI9XBngUM8RDJOO0QbjprS892RRi/K3j0T3y0i8PL8AJYyX06GDu
fwB2fg9foOK8iybH9rGFItLwxrdgAsgA2rG2BxbbD6bODX4MgPoBnvm3FP9qWdRWL5gXuiIgW8TM
jFDx71ci9nVmyUHpOKZKgAFdqhNlkTJpu/82Z3oAeT/uftZ56nh/d0R70oBLkCVhUNs/9lg9I0wX
xlVvWz4DaqKPZaE4MPzUvYCGnGMwnFW9k11lSe60Eyt55f+cin8MhWYKjs+KUxybZOFOiVjry3FM
oSjgn3emAE/KbJv23QTSj/Euc+PZ8FRLzNefFO7m1KQoznaIS2lxFSfDgmxmLuIoAxcZL7V9gOdv
Ue3WQQ69LHPY3ZGoQhLC3AiFRmuddj2xAO8W3TaHDaJ0TwVrLlSDgtKfGYCFexCo/7z9vta453q7
4EtiL3EHnentFTvDU6+D5UcEvSE+NuuxYAijPhAmSzubRqsEK7ZTnP97tnYOdOgg8lkzdtWNW29B
IGkzd6ocF6B+qD0iFjY9weEuWedY+p0D4ncKt2MZyEsEvnWu5paV20pTQlbLMtmzhaqM/09CilT4
yBWI9cvlqzINA0pIIc8cG01MjALUcmiQuI99hTPLQaMvOiKaWs5rJ5NCkTyb238+naztZWOb4uW9
fxtzRNU+VmH9djdLFJsFOEywIxXFin4rf7NJA/vWfX3nf2x2NqbbNEgaCSvdL/LeounfNYTYFG6a
qObnCAbNtoPhPVcFFo8WX87pYZ6VcGcqLTK8/Wlp4XcAitzbwR2NJG4/PdBEBBWMxqH9awMc86Uq
flmtYFgLpJ8EZee1ugX8SDePxevxUHBkIybUHfqJGtxMxQxopgT6whvfyRA/UJkBi+qc9QTBJ8ud
YdjY9XhV1vxCRCH62XaYiMk1m+APVKjpBiVj7/96IkG0Gv2IYdjO1aZX5TNPdbKbEaj85fDKFEgL
RL/BK3/EYkDJIXHhdULmrTMDT5wP2irth9Yt2VOWJ5naIrwposwNyO4H95gspDWl/WRKwLurOl35
llDs0Apaq+qovVZnV3ekR2bm+4eyutvtOAVP/1+ozsKLYd9Dr2P1+/5mYRv58IXjiNcA26AcSLcV
x8aTpkL5CbTq4Mxq8L8BoCQn0BEZypLpcY4RZ4XjeqPDAMl0xxjcsHuBH6v11FshOKs7CufCHIlM
2dPObzl2z8ySBCXzTH4uOgFT1NVHoEU6LKI+5ZDN55HKkQk8dz4Rveys0y5vhgwIHL1aihyxmsrH
NZYBNHJRxGksgMwckljh/itbu3iBpQlbc/VaFFh3wawE0x1iwqGAbAcf2CpSYScpkeOH+kxg0kji
gE8kUKdjy045zCUk1ndrzCiV6u8JL7WVLbP5DwsBCJPGxIjtf9K1/Lip7YwSwZTF8XnmC+ajawJN
c45etHtJQdbNwwWLgGMNRPCJjnm3KYieagoNzhc8h/Xm5TZRkkyjsIQWX+YrUdLuXk5l68wzoCT9
vHkRmgyR9P7Bi/IrNKRMlceS2hX0MUpG+xk3mPXuKCCuAxvi//9bD2WHDCxXmR2NWyfj/SpSYO5+
S3f/DuIwQ7uSLG3Pqyy/RZtHDQEOnLZC9EzKEK0mHVcSxQnqwQB7uv2ydDe3T4o7NM95o96uhQAo
ld/G7Y4rmX6XcqC3gRBU3btLY4LgG025axwsBfi+VXWFrViGPMNEXScuCwOzRLwkqY1VsaEKW7Pp
dwceQPbTqoBbMXrK9V/KIJFobNvvbQa6EgXA51z9IB+9gb1rV1uYynCVVjD1wQjLZ2ldagKfEIaL
Y5Kf9o+AR6J+U6lGEKGVrBu3ZsV9CS2iHWlrhBcBi2EQVqeZGh+IyDvKIyLzzvaaO3EtynzD2C9P
nAIjJG34N6ZFiN4Rxeug8prYCgSGuYUk2LmR6VSw7x6pyRhfpXFG7BBaC3ETkLxxsAgVaECl210C
Gz5p2wZ2FGOS0uNPIUBpFOX+mMyYGvzuZ0wurrJMcDBHdMEaQeChOlMwz7197ts9X88j5+BJtVcd
kIRgXG292gUb+M/KRI2mkyIxNO+HNEV2NPXMWo6edUxU2D6ElT2QMPKTjbSyw1hQU9bfYFtLHBeu
r0cf4sKL8sTdQyqjNKA3T9u4LdeoIf+Tn6mIWgCc4t9Mkxt62JGntl6k/quFXvBeCYf3tTrpoRNN
7ouEE5HQuMGQYgzuHXUTBOiZkJU+7znOSBHB+GCCSxwmZp7pD4cYbk2Qw+rZ2BJR3R5I0EoMzfgI
WN06fSfXkBXTE59v3JwhnvvbyGD9AZENdf7BXMhgaglT5a6mTwdg0TBkiOtIbi9ct9wMiaSajd94
QQw+CaSyaEiQia0PzsVWa219jNoEmbXzvJwWA5VmpXNLcvvp00izTN8ei/Z9Aukr7fVgIta9ETd5
DKz7YohNlaOqPi8VNyqcqw8UM8qreilw/UEzJwHrq3zrZ17hKVR/C9TYsiBOHchqsVXRQF0SMzG/
EKwlvzRfi38PUXpSYB2P9uhlEwnCiEFTC86xxVD7bFOtbYtzaLHgbIHwp7LlXoDHJG22Lbc8X8Bh
klvhI4q99j4A1iELFvM8oInCVZ26XFyqE54L9IODF4j2Md25Ohz3J1eNa+mWlDEaUg8Tv8Z9Jxbd
XITC5NmQwbsj03WSsv07N5BGiOS/Ckmvm+/t0lXeU8POoGCG3OaCTpv74CmcugKaOVbkq/0MRNio
zMq8gfVeE2A5VCf76t+nooRn+N5ewXmZ7i/TqGEJ+MFjs5WvFZoMpmqnPUxAk+KEuCrQHEr639jW
BTkTPfw+N6GWJxRf1QzyX0hVgYjIqGYw5QHaqQ7zAQApbG/kLoip2H4DUTLu6W5vPr60ReNfGNRE
kOOuzcIC0hh1F1ID7+XjZ/A3pGv3qQSjfXO1mSdnlQhijuB81T0Qy8JGLjBKcqW9xdbF+iaLUkSY
wLGqsPJMGEoiMwA3IC83XietySOCkelTamtbio18oL5kW0wZXiFVcfU25yuWq7SYchmsVd7LAy5v
Z+OWYziMEopS/fyjyI7RRIk4yox4smbemRu6tHj2sUaE379JeVpZw65MPMWBa4pXU8+Ir78rOsDu
as7rxsIAoMh+7Xk4AmUOItcvkN1NIkYJKaJ2t4CoamRHg0EeRFtnQmGnI6oeBL+au5P8rk0n+KE+
I22niYqzDHCaWfEn+K8L2z5Lf7BCJVAKjJWIiAsD9AQuu35edF7g8aJn6dUeqCeGUCYmULa7vJpD
EyBlPIoj8F1LEN/Ym8YpFr0IAbsfq6x6uR6aBZaC3KqJyACuxpyDkN4BQ8YXjz3UbzztlLf+YP5J
FQXJNQQYMCx73TFgoSTkN3ww4Im0xmp94SDK/eGjw6IOQdKOrVkL56V+1TlPWNLgx6H2fGn1bscx
b8NObBqRD98EJ3UkAYBBrgddqNGD1ym2xfjPcFvixF5xcRH8jD+q6Iz/AWpd+dtJ2Mnw8Ndn8Qxg
h9xd3+XkExgpVwVHDwiTvRgpaVAdQcMVQZq2m4wMnRXLAxM3o7ODZbaCfZfnibNlg5KvsU4e1YMp
umtop5Lc9RvhK7PZxfh+C+vX+NNasyhPt1xbJuP2jhwvv4y1blhoVttUoqZAD0FOjGaue9MDXGZP
RoULPDydiZQ+kH3O9KnJe27oL3+2K0eYtarmIZTfknTHUrJ+zxv1QL3sjc1aohyyAgYMSqijv7fe
bFHsltRplj3Wiptw/cjdiLNlL/xKD0eyrFdaIpgyP1eRU9dgNtG8v7q4S0xg+cSUzoGl79aTsmgG
Xby8lKd5/iCtaLmY4MX5wBVDhqUtZF/bmtBmUcomEK8V06B3KpGaYSBpKNt+OP713huNCnzuIYG6
oxzVqPxYk9o5ZZX+dW7rqx+xm0N/J00ghX6B7Wdp2KJNgBUgD3PFdVnAbhpmkD6nXB6YpiQ+Qi09
NYbZ1Ji8hn7BAL7FUZqNyhzxZFbkZ3Ukh3WvYN3pFMUfv263I640by/QOn3eeGI/N+X0yITu3M7r
G5DejemKcOqzfNpci2mS09HbvDhXVtZIe9VN1zCdDPl7dJGsb0tNUiYBCMsdx8W8m672QxlZs6IB
DQnOYpokvH8/wcty/F4FUCfnyhf9ZK8D+rL93bpQV+tCtArT7RJV8maYJabxiURpCLsGEKLFslTa
ryfzs52KHuOQcyTFXK7KdszylyfPr5QE+JSRd4LaQnjBmk5oukxz+nmWtegk2pgeQkh+vSjmL+/3
Xl3aU6FnRBVhdIPq+r6+nuWoQsf0z+q+PVhWiAUo+oXm6zUF4INVOPOPNjMsobJKwO7VaQ4I/Xux
mhBPGZEFRYRHRxt6HB2hGB26zIgFjFxYNRBy/SxcSrsRJGqexH9fY47AoHTa3K768NGqS7BSNFWc
q6nMqE1IakLosG2C6YbttMM2ASBIoPaGKj3KBYMBwm7YpkCL3Z/6Tt36th9h+pqAh+H+TYEjqG2A
YWiNWUyLGzDFHgAhP+Zhz77g6WaPl62nib1k/rXdmIVi+JdOzZMIXEBWMCTTBT6++c9wMK53T90R
86IDmpGnUnIU40CwGmCJwINfqDQ8oYHu3uGfnp7A3lgcYb9xBPOyTd1ckI/G/bQODxuScq+VFKDI
mxCnAHnVnijm6YGO6gdr3jUrOZTxTSoSRV+znsuuKHYhfDjIeARAWF34tfzfsVrDZTefo3qon3jx
G5QJLDzyBDOV6RtNEe+rDAagdkkrb/Bvy2zvjsRR+gjcNyQWsd79CGId9VaHL1faA/PT8RGPDtYp
1DwG2fG10/Q73qNnbvMJxCstnnZehRkk474ymHbBzmtBrOtBQZE7AEwGcyt9Hn8JJNI1zeQQFae3
dwW2+mbAl9nsJFDSutlpgnyLrsLyodo6IZwmMw03TZx3Xm1VkaZuCXbruAuaIguPhZsPnwponKpE
4c1Zmwxr+dnL1b3VqNJxP2R3uZwHVngIkOtj9NTZrmpvz/1vRXezlrLCDYgFzomwXUs4se3X0mfI
NeEsjVA6vONxxKM6EmkIwl/RD9sKOfoWoA1HSxRLsO/fu5f+QGj+qKqdz89IJALyBmMnpeiGTtMj
C/IpIRo3UAADHe//FbkjgCTD3574/49ysaq+Yrbr0Nrxh3mTrXSCcrpOBvZBdwBBylr/K1QqN/5B
Z7MCwa3/J9MFyP5H3gWFtDI0d9Lwl/UiwuUgGeJBg6aV3WSMCJApNMEN+AdmGEZwu9crBOJa03D+
leRoRApqtqNJUXlJKTMdqwVyG8L4YXqG4XI7SF48zhgCvoCluze/FAFvWJsbiV2op3h0ceYtHgMP
DLpifowJmawaWVCZGyb/Al6v3dchx/bzmcLzN107CQQax2s7LtEyHWFdDBbkPJ2nY1cc6rDKCrMN
kVJEdUCO094YiCGCJeEwonCx+8mSoG21s7toFeyZXEL4n9RiLomvrbzXWlyM1zcnyvGyub+YkjGs
e1UxPp8zrPQDQjuYPMrlerbjtgzUgDqsNRQbVSyaL122HHnFbMjCEvjVBostTvJrQ0lXhaFDBexs
EsgLAwyLfaG2+RLZ7ncHMd9DlwKwQYED7jMVJLbkIMBhibMxIjGgc4KlSeg2nQrAs/j8lfh3vPRk
rqQ1a6XVUnkOEvhHLhDUS50jHK0NysU8Vi4eaLzZj2ojg9aLSHeQ1YUR0HU9WPMoynQP0vB4A2vr
PEx2gzFa4G2wr/Fs00RDWYetw7TNrFbive4fGOro5vlTiDhATPqydgjbaXPRgNrfFp/CdmLDZz3R
axL7Av5Oit+b+X4+C3FittURhQilffHN9Lk3WevtoanhX3c1se3TsfanjU9GXAGoTBoNkGUOU/a+
s3rSkx+u5c1CVNlbl0I0b+V4S6k2lxg3jc5M+DmdaKouw0Wcx4sl+wAQoAh73tINOD6iteMGCWYl
tW2W+ml/bsh4y7sGvfyLPcxzzCyStLYAiDGOQyw/kSINLGQrsyKDRAC+G3j0UsBOq0moax3liTYX
OLs6krfQlgYZYgACNy8e3xTHeIBKSEAjWhRmCXiGqg2HAOT7LCl/AFp2MqB+J+LMtpIVcdfHAbP1
QwtL1xw/DA/j2NSH01wSTnEeUDu1GInSZ1FHOxwO9NRYOugNRSceAlfE/BSrh3tclyxJqAC4WJIr
wHbN/YjMa7H4HAiTCoDFW5tVizEL1WoxlWeREQwFuLqOUQ2/L0AUXCADRqbBzNFKaUSVM5UJwD6L
5H4P2i8F92wJnC0n0/m3bp7ouBN/rbPADAq7xxKiOJxwzvzJ/sHZHK0HXck+ai5K2Nvnn2wTfmxP
6S01ZW3GYLnuzqTgMezUAwxnfK0lEVoa3x9bN0jS24n6pUX4/gRwOYinAtAG4kdbVfCHGSc25GMc
xxw5d30i1OZeSqJsnKeyuL9aHCyOIHGPQZ0ekrlHXvBPxjdN+OvFwhct8OWl+ZLPEo9CzUCNKg8b
g1a6udOnWAJdgCq5ASiDJnlY7O3YeV7WxHDeWfSZOb0kTmbph6IHz36Ahp91UXbbFqTv7x5JZPGn
+fMtpBA2RNp0sHjDDmc2xyhBX8HM/4FcQwAOfarw7oUwUXOmv7OlALktBJA3FrP13hwvHH1fizjs
11BUzCUm9MhMpFqhGdnsotgbRF/aArWUW7+ycoQUkgXOlc4evf93iVWcd0yRdmPWG8EBo/6dZOch
1WnqtcnikCrkdZ5kFT8qBm9/laBVuk6OcHO7sWaK2t4U2Ax2oN+/TFAKas1Zhy2zFgbn8sG7HyAv
TcLtpLRSLRhTYn+tjvYg30Y68a3WsupbLQqmR5LhcyxyhxZrbPjXC4Ge+7LKL68ayRahDhMtQg5V
A8HxFcOd4v73+hwIbkCrHNU2kiJnRL/YyXoc4+CAnwEO/OTVNeaPSccedfRj1XUCm6/OStFeMBN7
pfYocQysO339xHctm9EQnJKEzIt4GwVjQ2+c/dJWFcd/dczpP5yrWAXDiv9uqlCmL9Zh8YjMwuTX
++lH19Ie9o97n2UlvlRNDl5RUXubbNCk33DtNKXc4lRLIbUJP1tRB5nf4yC786bmHq9T67ykMj0Q
2m5LKPSJlTL1vQZj0mZHKJU6D6+CTAV59755zDVxlaMjNNncL1acb8Zb/sdVHnC5jl+QO+dQj9iy
v9G08Af1LclVdc7q8aKdNjWvBB+bRq7znxAs9gEYn5GCbQrcC2/UXNx1IaxCopJQ+pAUmIj6/5N4
FTYuWHAOVrYeAQPnyusowKa6Z2g9f3w9hVU2bNQZgecIMBcw24X/zNj4571cJE6uNY2ZVaeA3Qty
yUQXOjyNPPuHv1Viz0kDeE+XtaH48523trr1Dh12+CmiHcsDrpE2GeXw1y1TYPKojprMZjV2/Hpz
TtfcIM1T3jAUjIADM4zq6KzODq+HnAxAULma+g3SAavROoY6XxgpFtoynUg1WHt6qBp61oLSjK6c
7tLe/yUIB1PpdJXKYUQYqeCpo8yriI7hPbYIpzNiY4mIWkwEQyqlUDxuoYghjhQwxRsnuda7W8dw
JkyGKXe1Qx37AmalXnfztXJxO/0QyQ3GXY0MnLg5HMD2qaKq9DYJ9beEqzWwAwfL98biGuwJSP9E
aemzQgT+c0z5S2qB7VVJxZ++1GVaKWC7RVC4CRYx+5x//LJns+liGuPhme0BXLziWxan6yLuTCUe
NW2b2WT8q01kEhF0bTIb/dR6sQuZTi63WCkWrvIQN9Mo9PsUxf9Q9mYfIlnI+YVymiD7JmY+mgD2
FuCQ4QX9QbH9/q5tO6hQsxBFotvR80J5Lt3gyhveXWU8/QS8tb+riIAu3/VIqjhEHduVTIdRSkKL
zjF+M8Ne77o+XhVvOrYxpiwI4z55MrVeCk6n2Q7g+YEcahdpqfsPb6i81gJEWPfMjfzUJ3jW24vC
QhWDXNFcBF1vKV0Kz/urdhaXkzHH7ToJ3V8dty61U4hg7L5viBSciDVLgEnc0+UeJ+SXTVWEaNv4
1I/dD1NC1kgfpsvZ/oegS5nzyusUW01bocyN6AWWTVo4ONkWqN1L2Q/VTezaElAq1Y3dvebRFWX7
GWNW4kpjWJ2YJr32vezCMdm3FFaO+VSS9JmxKdLrS2LMTc+q5RE2ExyQ29dd7fxz3ASIP8Jlg2wh
DNVVTAUhT9tJqEJbxq+FqWn8dHMWfMy8rSbsKJfRKEB3X8aIXX2SN2b0d6BbkAGfi47FUvHDzHAD
LTrooyQVItKXaObkWuaQ8lFYkTysmkAr+4X2XbqLdHazNCwpFksqqAhnndiMILASO7j+OWVrS1Gw
vY7bnvW+b/qiqu7MR/k/1CzgLQ7cl9Bz/Xfe/cZ+be1xdeBlgEmaJhAdL0I4Uiigfq0yZsO4wIWK
hCm/hsis468PkHcURYEYd02YsDdH+W0fGDQTAlUv14lclFhOiDZSvkQ64wjZpW6+YdWqZuZcyC75
EAnDi3yRPs2NcBQ0K6EaCODAcSYjtGDICJIBCsQAA4uGqH9zTb7JiNjE7xSNi4T2Bh20fVrFYEAi
icrYfRRUyw3Lc48sSxaT5Qhq3VZ0FwS3vi879qG/fVJnQY0hBSH4g4bRKPpsnLBsljlxBzv9iiRs
k0S6+opU9ZYtxjWgBKjOS3p420vAm9wqEPSFGkSqDzFEYBN51VKjVXTE08UOyzi1mzm/ItyGmMZV
Dg/NfOf4GdJVfWgfgvUFBIWRutM/pLSexgkfbk5SM3T4oWh/ow241XKNiFDM+cy00nTTGjdu1/tW
GezDACXQ/+9PIt8pu0SBXjhWZz3IgLpQznTebvR5z49sJAfSk5U9agd/DTKcptbbXJ2mgoZVUV1A
MIIrK0JCXfF57pOdCvw4uz4oj+O0kdO6IDjGt9LUfOUdRjU985i6vfc1/2VenTBFoviWcGzhpfEf
0MxD34k36hfaj6aZVUoMrwTIDHac59dBXbs5xHZ4gaHIZyv+4lDk08juDeLEJhCodBvISAlFjQ/E
pamnWGbc4MMlwLqDpg7vKEvCL7WFTUX9v9Z22zM4Vxpq1maI4LdECrMFsLHrtSeK/v/ec9n5dIWg
b+z/22h55Z47al8WrSK8uDrDB5gZYVCN39CNgP+QDiDJJb264hIUCV5Yh8c4GounoHzZe8bWkdE5
nJGypGItQ9aVt/5yXHmE9WgegEkcvhbTYbX1LJ38bRgGU9yh7v+f6XElg7ftnlIhbOh6K+cs+gS4
CIWzRJogGK5UG+WUV79vwyB3+6pWpAK6LjJBlEGRfLZe9ffm7eiI4vVkKNuKNl6KV9gesa5TJ0Wz
iGWiwQ2XbsQtuHZLDiiL+bDMFg9giS2Gz8eyFQgGI+iqxlE98VOMHFVKuxYQ5qxEHk/yfwiSGwWC
HeZuIp9h71SJ8vRExHNP88ZYYpcE5N6npZb6qechOX+94kbqu6n4zOwBL0pufSVFUsjop3tqufqq
+IrttElZnVNtCjAGDzfmsr3q9AQVtB5yKZ62bwSTQjwaEqDFq/itqJRrsqBzZPpaVkehlmJOA5ne
Jo+TZojeFYwKVkeFFgxqzUZ3A6QFVywxMXed9VUxVwTVkH+aLy74Z5m6ubz6kQvXMVFmns/ti98D
ws+WmVNza6BOPbl7nRCko6lmhnzZH5GdvqeUQncGblowGwc2lXZ3dSPkUPw9kOqqHOdOuZ3FPbeR
9utWvNT6FmH3Nkt7gxbdh1BSwlYFvsjW7MNcW0DIht6oKGQOi4L5iAWKcz0PRLp4/aZVRlZOc1FQ
UoM2bCKHaj9SfW3fGy3UM2dO8N7bf0p2mMltNNT3HiSSWLdItw+Cp6gTxD8pDaLQuvfgWkS5e8L4
FchEdanx1pYIYP4N9+tRMRo6TSmssM5IyuIQPnzPBLntWP/LaneniX5ZW+pBLWzUSmKoxpegyUDY
L1dw7nszzalFS8TcxpbmaQDWjVlTN/anXEh+2+gxMshNbFuSQ+1DsiWrKn6WpAgSeMTMDSjHjcU1
jPsuAGgIM4YojnSB/g8VjnjJLvNFlC5Aa/jpMMJjT5QN1jXycTGgSavG3MT053XnIOzLjK1ofT8Y
Cn8unohdTjOJwaDCuXCQwcnRthhaByka2eCtEEjZRmYhIGZGrLAeTam/RPv3ekc61rcmlBl7/Lek
Xz6+GJgrQ061jixGtyxFEyY5hPrgSHKNADbcHDgWo9qEqpZCswm/bMtAhKOve0SnpQf0MGNpJRzj
xrNlxIEq6TQJxtBkfvpnYo+s23xSPUUJMLpixBpsAid1ooaK0SQTfUJ3FZEFD2eeVX2435W5/rv5
FpPvh2LJRjAsb0rT1e3itGDHABW2CVyan4gHb4p4aSzVwUl+YA4Sv2IwBIh4jHQZ3PlwnMm5gIUM
mLR11nOeZMvhO2Ye59UVsaxEU3M9glYySupaX0KXEKumo2LMl8UOvBoS3Gll0XDt25xcFynvcD1T
UqR2Vyqm0IQgQ57efJ9SqDL/CNFby6iVRYm8Vvcp2+DF57XyqKjjjLNzFWm4ptK6r+/42kYJHPjQ
SflAGXfEVmiUbBwQHILQTxxvlR2Nm6/CzWtptG8KOBk2XSat9QxZAbyczgGRbWTiVn77sWc+9MJ3
qugIKbz6xai7O3yNS+2dWjS+ViBGXP5Ug/hxj091j6NBaDmQOTbEp2OGoItImYDlGecHbyK9+SwN
eywjbRa5LPgpjGWda6b8GInjc22NzArxOYQCZqYMU8R6LptUOvQRNVKaE2s4w4rGSgJgiQ1jBUjX
0NYoLg6mhvMg7i6j4nLcZ0JUUF/ZOSJs+SS8dCDLKPUgxUXBZjyFZi2k50Rrskho/iVOS20ETaLu
2Moy1w4DcGd+Gmuk/l4A3fvfbvafTZ8Wm8TM8m9IyJvuOJzjj2kRBc+ALbF6WFKHm7XhxsqCiOsh
M4P1njoRULrQOK4UT2DBs9U3ntyUsY7aUzBTgcDORvDkoOXNzkfmscHQkx7V4UF3WIuY5f6gZ5YL
SavnkDuXUfwlcWJmaY2nZ2yzEOUeroKKgQfYsGI1TY1wdx5pbh7cDDLLIT4idXrZkKtH5o54bVqW
XiCibO+Ts12eFZu0mParzyhKtg8E2z0sgLeP6NgHnmGA9GZwxkiDrhSSBnVRYaFBJCTBS8KzCpmS
RvbDMNQE+Psc20K0ScAKImF3r+phWjFmv6yN03kgKGLlAdf9aIh8RFYvL5NeHqCyYeCuaOSaXLNP
YLsdVVhdmjVjZUWgg4Vpk+u2gocC4s42SAIV1rkWmd1BUXWMMWjCGcXck+tPGwT/IFThJNAvDRkf
ZRGKX9zi9EYiXQnBjqaV/9C79yADiltteR/EaNSIJJZwzjOlasop5DH4ag/spUL6OEEQbfH0gC2B
2R0ALW7EsFCDGUz0KpVZC0xTSQZFsMFtyHyDOSo5wLj8O7LG0A59A51/Pv3H53zSpXL7HIY0/+8R
cmz3Ainxb4nVC70yjKaZIIie4kZQhAXZRR4RLwTcWRsKB7XqdLse876w5r8WmFtkxQhObb7/ZA6T
7N+51h98JYH5L0exyEoO2+N6ll1cEPEnGCJ0j2L/oWw9AWqm9THvayVyYtybMrZdHjaFZ1Hczyue
bBHC4JUXNrRSRQHRfKAFfZVhvtapOQ97ISCL0sVuJrNK5puWP+9TtgTPzUFXIc6tZyZHR/sQEart
DRebD81Bj5qC1+UqHH6VwC5AzHgrhxiS2WkjQeWJ7HX9I5D6tiw4t0BMT+nBV1Jjwk1fey82V4hr
OHlkEQe5ojbZjcOiGmb4dKnEQvF0eMBq79fJL9YFWvnG8YXT4RuW0As/Ra4tnjujvuowuFv6fnhx
IsuaYpRw5Hqt4U2AU4x2hkkKLO21DBMgu72NFq4be9e4S99Yd9GuGCVOFsn9JhEb3kuZd+CP4wJ3
CbPmUfqiDKKTMKJFOXLlpHM8TkI7WLyLWWvOt6RPauQmc14YkSG53zfl8YVOC9t/gkxqRLm4r17/
iepiH0ulExdiepZRfzXcZBe3CaQ8SV5PGIbDGZys2s3OFUwJJJWIvoTepOzi0i4QjO6gja79L/qn
Rm7ZBXp/pPLVqUuRQXNau9gR2e0wn5/UYb1WusvWwGEqy5ieux9LHk60Ybfd7m5abWksu86nBxja
jdLQ2nWJGXwwWM52gw9vi5jqTBcz4d16FvkBJlEz+M6ELC9jAy5Kp2NhBeOSuoprW+096lS9OZqT
eFDB3+kQgTeQjEL0ttyNKENSgq+0I1MEsAvdC/yp0pMZNpyW4GVSEIhBw9mDqmjWqwvzrtb88v3p
QXkkn4dGibfoGeP3JWuHNtyaTBHWuVimy8Z1RpucUSf3gEaIiJ6++tdUac8A17jcuKUAL1E9bWLe
BNyet5bN7o0JMqzF9ChDT6ezy8AjHN3dzL7bgRUpmCQlcqV3yQQQtwOSw/LQyLziyOHHTNtD/hTv
1wzTMYTBpYgT2qRbsc6Dq12EoNdqdaflAw1edAXsC2jGDCFRLRxXNhmzAwiw/XMm4wmNqiAyu+Af
gF03LyRCBTCaTc42/Jn3Q9Lc0Jesunve5xybMOFtx9mYZr4IH+aG4cuPjHjfP4/MefNqoSWZew2I
tUh9GSBZOh9GWOeBvLPc5NP5RX+Q+gCuKchkt+1Ik/ebfEAkF/BHp2hawMxsvZbLsIU3NUMVwiwZ
BojTBZDY3fSvMMYIRLEPHVRGRR1JmVXLXljNhIh1+CoZw0krzpXqRoesGDqAn1dyMgd7XaO8YPKA
09pQTR/Zny0UWASkt6PuDPfWjrKEBntEQATYxVGowwHftQFZuSoBUJK1vK7LSv2TQ8Unmqnyfmub
vyLZJK+xEoLjUjP3Y5NNDWqO6NjCy/sIbCBqX9J0pthA65eisM5X4svNS1ZLmxa8RGlw/Z02D5Ug
RplkchomYxkGQFn8Xju+F6kbJm0MVJ7EWMvaqgaY36u2bSu3Hi5obFafYYl0Enep6CHtBAS61//9
nLO5wv4I6Rn+eVPEKTapL1qOpX+Oxzfsotj7WaFcguNoW6L83BT6mDHUu4ILuFVtQXfB+q5EE/EG
lBgQZIEgewVBiRX7N1HJd7s5S1F53j1m8EHYPATiph3l/He7ud4J1OeSvK9qZWuv9sMr84d2dQha
ekhZdXWqA84gr7fv6Oyifv/kze1EnA2HgRPiFRvIJRlfPqQLKa99gQfyr+Abb8Ponveje/3Icc5b
y5nhb/u58CDR63u3u6L6b+poyDKeWMsWRB9D2L4bkaQZGbQKhWs4+oIqzzRLs5Hpodq9/9jOkTVj
uFGMnBI5DYHg+rBYDtV34wyd1ua9G0pU13dzukOS9OUut+oG+ZYFjX9w+4qdJOYd4/nJZ4ZzkszW
zO5ZAoDuRhkWegnd9t6TON/ECWlrha3GRNe875fhWJkTQ6y5+Abu4ijHNMcX+ARD/iwz5bcnI6jI
RShFPfpa6VLl5hj6LMDiCyOGl1Kt6WgfR2ERMblfVAFZX+N5YSaObhZuLsJCMuX07UmxvoZDvabi
GUWRyji5zxsYYNdr+/44crCTqIzp9cxTqtfTfw3GiGP7LfYsyOsm1mRYJjGdo0qgrwf18czRpHI4
s65R9ZK+/qLEHXgS96tTCOwXgJlLzUJbE1/dvdkB2wxigc9E2XFyJeGkKfCHK0humskdTmKxgKkz
XSNle6D0UwKUrykr22ISejIohAnAJL4nza8pSBZOU/hozDTkejyRkH7r8UCa+oPXQnr53dkwz2SD
O4OdHu2rf8QCOSSvSvmhi4buujJDWNDewVjhuWdTMq8YajkaRsnGe1xeS0/F4R5cA7e95pIziwTY
kvK061dY/u2ykK7tB8hgmXx4Bbm1Uyik/XhO2HY5Rv6yJkQkiHz1VKT2DZbCJqlSxlOqVQtndeK5
46Tq4rmAOprhDyyCf8gXKWlw7163m1e28q1RiZsaMdn97bjDecz/mDU7hcu+e1arKfb5hK7QJGuS
Mgh2VucW1Ezkr2YfmNq2lYubp1tXyWuwVNiuZHwUWAYbGsCsT/ObNWT9j2lTGPFNk7p+TUnAETIo
3E4joYoXx5MK/Rz4Y9IWR8rPiba7ngdcZQ9OWEVAhDrYE3vntVj92dC44ka7z79gJ4b4HTZvcLGR
QDRIgqwQflKvp3nqObrAZkTofpvKGP/GWE2twwYSKhcztdjkv8dw7BJNLnvnpNlCNoMYMKmgO8u5
6ueor7NW7AbEspO7D8wNMWgOVxMzAVBukBEEpCPoEJSia6VMfzFk1iU95Tb/gU7jO2dzLV0uy3BY
JDWvgz6/cJ1ePCFigYdshw30dlHdv52RYjBqsu4oUE9dZ/5PgrXLYWlu4SGYzfXcmpQV+HJJ6LRt
iegIouy/b0TMz3sSJKx2mJTNtCuqDsoBiLc+2feJZunq9dB0txazD3HZ+gtivaMU1UgCPIzqd3Og
fZm6j5xZcrubGSCqbA5BLxfE/K27wFmddNzGdanevoREKpp5chqjgoFDNqGBSmbLCRg3jExHOmgG
tfsSuFryJ2mriCuI2GViEaXem3aAtMabr33JmeiEjpczFpXslC3mu131OYadHTd8zW2oZakkQzmp
FTNfP5YS3PmImxjDHVniL56C4/64i97786rW2+3A3eh5csGdpIhsmcZ5C/nsxO3AjYaINLSvcrlO
x9Ded2aLVXdUulclUirt8F8lTJV7NqUBu9mhM0eDhmxun0SucR/lIDm7oQ3wyQvOMJ0T45qSs9z+
Mte+9kmWklAtZAjgD6w9NZRTZCNJ/5EoKyvl5WGQjMblgW0DCbXnzPLa6pH2rk6QbVq3ogVQlGCv
YFacx9Auu407lsk0C538f5OVf7GyXvZcpfg3MrArSgj0966UPJ6FVaFHzRk1h5MgrRHK9Y8UOWMP
st5x5VsXC0hmZSCKXajZYYQauz6S7FQLHdA185zHRW6fLL2+lkZjW+WV5lNxbjJluY9cLgBVq9w0
/7xq8YtuYQnXJLBqE1SX5/PGODiUR0oRqqDIxFO/+H/pLm+lNS1Wm0ul/qzll2/SNbF7KlqdTUIt
6Xv1NhfsK5MUlyQRI0+rwrIJsS7VGU8AH1x6OFYV+MB8OtWwuQge9cGCT4XBHHPgsB+88vbvhQpF
kxUZmQATsmKYxdEio7Z/kVPgaZIQPYMFtI14TVi21tj12MR78SrE8/hTwbdjOxga1/+EMoLViyBb
W0Qd56byi1CoFKNB01sux8vlfnMER9bMiFPziTXAWmcd3ntwo/inaJ+UvXKJBXuNMf5HakApv0Z2
sUf+IJ2jbXUgEffeiTPSdY839htZrxAB37+QMx+akHANdVcBhmXwUAwKFGdHsdo19neCAB2njbRi
CSeFTFdJznTSGfXH6yuhyCds9XeeVmPk50nbuHHhxLSZimm+wmHrxlhNBR+PdfPKft4noc8YHKZT
Sxp1cc2JJhqp4qp/Jhan3C6khnNDrFq9dKpdHrJwvNfsQKxNORjUcKoh3A1cGkUiXigiTzVeVOkq
XjchD4p440NxfEA60fU+S5WvaIho42rvluNqh+h5yfMLrdJVY44X30tiLrjAcyaYltYOdfPHveWW
EIZF9QVTe0HY3bp6ldb1NmVAY40hpdZxfmpYYXI/cl5SugxxV2wJ9neHolQJkk1z2ALnFrpFlY7V
n0pVK0y87fHu+3/6K3ZY3KQ3LkeREpctD8NloaH7oP8ef5nGWSUF4dcvnfXv+mQCDSLwXFa+95bc
tUO/9XE23jt1k0mG86aiSmiUnG/dxUWERqT8oeBDa448zpj5L+69V1Z2NEEyqlWWpJbI2Pz3+qib
Xl5C74ovmtPxbTzFNrWjMrNJTbdAbMWQdvyxeNoKkQSLPUKquWliMIG6JT2MXDTeANQTpodTd3HG
vKsUbX0/pkQT0JxYBxgEKoA558s3IXf3EYdDfTb5yCy7gp+WIeHmj4c5+rm12tCdN2Mys+ljM0Ua
aQfrkWSD7F6fJFgHfliQnWzJD+e4n8iE0cnjA4LgTA/WDRQFdQ+URcyuoAFHJnq/9loUyfNIS5zg
xEURb2DQYQ3iRvwjAACMSd9bbs2RtIkQ9sa+NjD0L3kkkP5Lie9HbpergFkP+cxMsKg7iTxVHdYJ
oB31rP5yQA7tI2ax3P6nlax+mXGvAmSHzoO/urWh8YZ6iWPzWgPu2HWMBVK6bOfz9fzGQGbcEj9M
tToVpNVzEG7rOnpgPDTPabYkPcL/RMU5ZHFNLEk5LmvPAp73ahd2PmV6C0X17Lr8YkUcddwem205
gBiCkzfWBDhRKs8JwnKUlu6EZNgrLBB6XIClZDKoLQWRIRv5TYfYZ7BqRDg9Nf1srzo7H6cwfMfW
mepcJLu5Z3RgNqF+id9bkEEG/Olu7qHzR50p7wO1ZXn8/4K4t5K3FtRQA/8zfCnYY9w0zFBqolTY
T6MjUCKE26VDfYcMSoHThQcczLWu6M+D60OPqdS0r0cu5tLLdYaPBBxhPTFUu6KLN7tHFNI9Hry1
jZ9NpnZKKyDClbnoQX+K2RILnRe4dOl0Vhi4iauv1zWltqVH5u9s6iO5L0FQ3A1rwx8T2ctlO3LW
4PPXHYnxHhVZUZusdoI0Ctki7w8KOE63Me7pHf9O/su7nlAtOR3V/SMlNYSlh12wpSnpAlToMIKf
W8Vakzsrx1NUg+Bro8s10uKGO6AxH3CcrkCqiXQ7Ly69MDcqe9Nv1xttRifKBlcuyIyiJLEE34uL
E6E1Bd6COPgN+0lByySC2cahMRI/bNYEXa1SMryRsQzN40XHNmGXE7oaXHMtvAJm3aHr3iJ/8wEj
gQ51LGbFBYuks1KpVrrMtBt2p34mujay7oIM3jEm0yDFpoMMEgikljxfDM6Gm+sebMFrOQz3e6ak
P+c/o77sSkTLC9UrIvmwkmKEcfn4dg9EtxVlOXcsaOhzY04Cfne4WK4njISocLCBUg30gQ3kTewc
GyN5LcixMkA3jaGrW81YDS64dN5XWt9dmbBOlGfOVjrTTDXUFkayY147rFXjN54XlaNJsFlQu20K
3yfbUDXEq56wdBMGYscwOZxvOsA8of3Q91+590BTcro+VhM7IqpV52Ip2Z2qxjx3fdAlNF1TA/eK
mSYyH1MFLeSkdgePDAHWHso5Ym2ekjeeTYoEqKc0hbj8DT4olLqgww9fwY0B4e8h6jHcg1TN24cj
LUE3fiXZmX+UbpeLva62HL9fUbuH+uRShG39n9jlK9/VetMTx1g8bqTWQr6oJU22xbwHqITzO/5O
S/yfktLu5CAVtQ4EOlOp9hl86Af316STy+e5lTpKfRuoSbKhKnGp90inzygBUY7fclh1tff7ncja
HtHEQWQWOpSOhZflieFCQ0cHTbZmF4dgkAvE13DRqKQWvHvGrrt/EIscp9GYmJJDdwmSrOHHoZLi
zKVgWmPRHpRVvhbNAARc7PUzuNDb0Rxt9MTCIeXoR4mW2sC3vwTzRb+jboM7Ha80yaj0phRYCiIo
96sZxQbQ1UFMTe9S115BYeZXzlKX3pHL1Tkn3x4JG85nbQy1gyTQEQbzp7WNkT/V82RQJ/KolFeO
HPgvwhaxavrlDad7kxz7pt5xcaK8PgO0ZEO+QdlKysk66u9x5COguePi9DjXyDpTO6UJlXZSSApE
5QiSCn8R5elDEgJ0n0sU5QXlxYXDe3YRvdoo3yq9HYA4+Wqx3nyG3DMwR5r8o1TSipUmWTvQIH1X
PIA1LWKmMe3VuVz+MPlrMUqNeV0UPSjBO8aY/v+SdI44TsUNf1d6krV2VeFUi+lQDVN/rOwlySD8
EwGoQibtAF5t9/CtnFhq++o16t1KKtKkVoyJ8HMjVuILzlq3nglOTjsQUTen+2bHXi7+mrIQb5EB
9noWUIjanohkH/8HqsAWuRmcuvr/BR9KNQtbM0uXhXATgDFSCV5cJQzxuHsh7JHuv4mlOdQ+BBdm
nAhS4Sqgv37djxOrRf5bi0aTWod96UggE/xXksSHvETSlPn30G49KgFYYPs6FlBj+QOjyVJIHT7C
WB2oT9wR2tUPWlQeIR/dGLdEAsmAuun1Fi5X+NLPC1qKjJJN6bYg0fbyt4j5oz9I1frO4V556zTz
P3JcsifePnj4CUQXwWg5HbglE6MDoo/PnSKno/FHrzeY06nZQMvyiLTbvMdxaiv/jo+ZR3BQq+r8
rONUOrSzvnrPzJdryhtTP4qDXmycY4dDQrdUutbL8SY738epQLrHwLLDgKhLESioD4chSTK68zXA
MnJz02x34GSwo0wLQkRil2/Bmko/+rPIWCKWn9F0RnQ/ubC96qKjOxKlZtOYvIVBkreddY/Kxh9y
kRLgW2wQ4rBEd9AR3iDDPL32I4p54tcHnJRlP9Y3vHlpu2oNrltke+Uod9st38KQ6Y/A+9WXnhgH
+dzlWf3v3mIERxBNKWX//YrjvgfzTCAmatqjBkq/bW+FZ+Atqpp1bo4Wk8gTobL5CZDN+FsCu0vL
oJgDpZz9qAc2tdNJAUxI0QvpzVqfiomE3W7dxGF/zivcQytNml49rRR4dJGIcGO/uG6PisG2c3vp
D7A4x7IvXSm4ZEA2iDLGjjeh+4JG1gisEWjqE/q7tLLLwuwEP5BkTqYixpM96Ef7sMKAn72458jS
ZIQJf5W0hiRTFBqHkqt3A5upmrKUo/UuY1kLjQ5k8R9OgPROASY0rRcuQK5MeKmq33EahXneQJ95
a9jq4RiJoLmHMthtIa1wurLoerfVcWkDhYQDV4MNsVJUe6CL2/fHjBZjMIBf7zihR+CwRnAb5k1G
MCS//dPQ9Yr2M5lFoFN2BdYoUTCOfADYFXncozyX82HqYgN/CQ/N0sOla0Cq9yCU2GmQILnRVt+g
LvDMVEhBVUyYCvRDJIg5D4+M6Lny2dQGQ8IuVnqewh/RBwt3foX4JCUYeh230xKHQSrxSpgtIZdR
BAfNR+aiLFWnEITftOH02oXD93XRUIm0/ayggOWnXJJjcM+MBm9f9RJh70KK1tB0XoFUJ0uxFa8X
3bKgzHIPtoOUK9T2qKuUspB13p9bhwCR4NUwWEWzpqX4ONoe8ZlvEQWX5UieG1TsfE4vKeNpIYls
OgqrHyCuiat/P4/vHqlKZHRHL0VMRWj400EFYz+/FzAAUpL30MJ6oSFblA6Kq3LyX+WFzDzMCyZf
1Hr6tJy71a1Q/GBDmpfUCrb8wswm6L1lmTdVUs0XeWgepvXgGARjeFEL61zv1yZm+BIeMra4ttkn
fdASa+oRPJrRZqUTu3UxoaV1SUZr4zvNyoSuAZHWXnzEQU7Wa7t3prgNpwLkyahmDXQh5jgwzCag
BusHmqa6Y/haMQunWbhovUnRyCp4uCMT3czwT5JP/R9KeRL8+0hiuMw9qnMeDbfC8YHU8uWHIeKF
Ek1sEmFFUq+O53esqBCcQLHzfyXjp8J43NpuVSVM80bDZoulP+ar3Y4z5yLVSaKfJltgWaWGg+Nm
T0E+uxCfXtQzfO+tVBr1QF32ixBh0QYbKEbaMcuRJyXn7Cru8v4hHU/+xgjAs4Efc0TDZ1OptQil
pkbeLZd4Jttb2u/m/VUcn6nqQXb9olLH9QE50yqTK3ts4JeXyrjBhyalKlJ0rEhOPMuXV7Oljgfp
K3ndL/YnViajIvavkALrvF+9XoLkoVPL+Sn3GEStu3vFZRKGDZ7tncQv0dsp3oK6oggwYP/gXE1g
5eMJwMYsNuniW/7oaqkwjZw4jK/Gy7BMwxnqfu2qP6S24HUrp3lRGdw8h6/iEdhZLmSOlgBJPcT5
adiA8t43y5I/2HotzFDt7IrrggzAr74gHq5PDSiFTUYh9VJRYQm4XZAebPEYXZk5Fbu4zChDj6rn
y+MlY9ptqzu3XOtNPmMSkXpy4BQjk2ZFinLt+AU8yRcKpJxyjkxx4zzuEnG2F3y6tYRlWU09eKzB
DUEgbMG0jinMA5h2gcVCw8cQrVpkp7m4/q+Jw8IT7N2SDSDdvrWZEhI5oH/f20YWmSLVz0NEpxgt
M9pwiaYjXChbWgq3WwN3BTWzAZWu7UQO6IfAFbM6Ebkh3a8Cvbo1DCWLGLLGKTUf778SyUvsAwE2
0NcVVpCs1F+xW2vB3wOVb21JwNdcA+5enjRB2K2IsLqdSf+i0kOsxCr+kcP/tgmX2Pg4guutrpI2
2rCMsYgVNK28eP+Go1MJ+xGPX3cZWeNabmC6nKbXloHjithS1sQ58C0bAaHgwDSieFpQaLqOl16D
I8qrvwq0g1K1Ajd3tiSbgE6CO//dP7ooKMadpupZp5PfsDkFqTS0lgzN6uhIEIG6h6QCc2lieNFA
3iK1noOmvt+uDajFuG7YmLQtW+NCne4mcj8A0EPvRB51nmktd0NNPvV4PCLLSM/PE+nbbwludbin
iBECfdeR1knhQyPVG3AYVQmTBZ5dTrsWeN5GhdL60RG/KgyEe2aJSgYQp4YgeK88CBDeWym1fpdb
P7JSLRXPcJ6wtwq7uUgPI4s/EWqwsnus9Tp6mH+DVRNTzQAKbZXG8KrJKltjLc5pNuO1k20jO0Ri
oGZgkqKquL2thE0HaJG0Dgru2ya1KQ+gHLJRIdBtbm+2uPoHPJkqGqwGqwcyw8C9qlI6stPMbTFs
mgih3AxlDOijdSDTCSpC4loIMBSTZ+jRx1eIAct/Pf8ndESSebCBgCmNoV7colwBe17nvDe07+ki
np7si//IWKo/cyj1RZKkt+hIp4uN/9uekibYWcftRnl+TJdJybTDZSYJV0WwykmF1dGgBH19/879
EZpDwu4nK9cuehnZRlWS86E7XJF/f7eIisEKoyOQPB/CECFSzO6EZEqqDzXxjO2aK2jos+PicoaV
PVUMv7szqWGpkjaxiY5xKmytBrIyOdFsngN+qGamLIcUhKVOUX2BIL8INBoUODcxQhBYJxTX8XUH
bKGCB6kTC4/Sf4pfNiyUvZV10iF9KOuWuT5htnCJHFOFVyVB4DSAgdss3jL9dA/DMflPJcvukvIf
JDyNX1TXJrjnQm+3YvD0as+gZJQ5ZHOOKSzIzoCGNOJP0kJ15N6vsA2zqPmLlOmsapewCY6kzXmw
1YrbVSys4hWJRfO5yo1hCA8KdG/krd3K5qOjvnKyowDCk2z3y65xK5SCLkzvmdBcDj6smZat6mCN
1fhCuW+T82JsKHJJmDrw21i1A0GSrcNS7k6tfz07D1k07Vye9BOsqcZxYF3nuGtCewcJslD+Rbho
X735BQeDdkngxwSbL/sjFsVmkPdTYsAHlBwmm+rlSNM0qC7vqgZyixgok8hQplGpuDqwcRYwDzV9
6XUQdp4kgcwGpHoBKHSRUTspYMXyPSn7A/DhigQB8qsPWNr/tEdkpLkLDbIxlWy/KGFuJViKpv4e
G1WyYLKjee1kWVQmrz/G6nEy05yNlX8ZsgYhWp7sqsOfKI8BF31pVVTJQ1S8/9pfPInTgB1saeVv
9QUUL59mFqrFYSXeWWhpEqlvEGeXAZHQpMcyOsfVNQoZKkpPrWJ+BQa8mLx9giPsFIyoC+bUqnEd
CvmhW7Nc6Nfpld+rBb2wK7XUqES45eyskGn/ETlE+N36iJ6Wo6WkzSyqoSPkHE8H9miJMkBz0pXs
mKl43+WxHDTh1b7GMuDjmdw7hn9A9pDQNjA24sxafI085FqkbAb6RcvTg3EkJ69YffovG9reVkBY
AAu2rmdPsDHZh8eBKYeywgGRB7sW8Gf2GyUFop2iyiDUpTnG9VSWOfem6nu0Yxrfez84dn9nDUw1
s5v6GBpLKRXEDYOlM0/RAwQtiCsUGpJLKUHfjN0QA2pl+3itJ/OwhAW77R2YMOsoNAOMwKowQzVj
SbgwJ++vLWJj2T1hEnxpd3lCcHlSftepK3L7xufwt9X+nE2TtCPtpsGJ1iWE0oKWpz0jrNRlRZXO
hQHlHjdHWcTtjyju1nLFpei9w1Ypgfq7zDAHhKZsH/pm6pDBbwmaDGkn8VBmHOTvA7OCge7o+j8d
gNgqwux4a79nUmd+AyZo28pRDmnea2oz8rxe58l63j5N47cIH6fUW6U58AfwQkoxLAWjrMRCWD59
MQnMzVY1twuyRKg9Jb1CecEFx2vz7/fY9+4cB+2WCLrOibchloa5WT7Lp0CbLEcXGW18/vymq5bL
aKx+e6VquEqaGweIkjwfkrt3UUKSU1NypyV7ENvUjWp6aYeIdqSIumAvFBvm/rGJoQldKJDZgCdt
No9jPZLWkXqYgPdjXJe9C97uSEc5QpzmFJaVDDpW2wVfF2xMuoHpaLrLZzgkHAC78S/Vq3r2L9UH
Cp4uGyCHoqJx+zTjWksWBD6mfEfJSkN897WBM1DwTnWaVCC34VYQ9qF+Ds6OJpj/T6EOv3HKsZSz
xd1bDgqqZS9RVEWtDJudXkkptsLitnUJa4AZ+Q6jWO2vzzUKgGuIqhLAvcM2RL4dENGVwvpXo3pK
rbSNWhHdEUk9rcmyGLkhumCMozcFOU9DWveaSUoSOwBC1OodfxLFZ43DM4x0w9tlaSShjXJlY83F
TITo6W+GEOkWg8HMRw6ayDvSGGUSLBtlLykvhde/6SI42U7oGV2ozSZy3j6/APJ8iiJPA0YAdgEO
rWRArZp/mmVaMj8IIizqaK74P2yQMl4vRhgUcRcyy4MnEUV0yUeVb0Pzw+2PIUFIynAQTt0WYhsd
k7K2K3wGNXAuuoWmp1yg//AOBGsokLZwIDEpX0SO5SIzJS9ploaJq+3U5uOLvVNj8S6WaNTlja4p
W0YMliN1626AgHT9z6jWjj8W5hi1uEOLtzZNHwGh0/VzGyXFPuCXPw4UpzXCiR0ZliZo5Y4g8noC
oD/ITLS8FzO0Lgn2g7RQ+jJY1P7VzDHBHlIEYe1n+WYL7YysU2m2PJT4eTFPzNm9wSKMe7seeVK7
4ZkN4KSUy8T7GAYvex0tVeqngu9JWA30u/SqowxulwH2PLlRFVE4WmpsARKnqSPKPn47efRA0d2J
eDIy0MF5W1uQFEOBzULhQ7r+ulGVLBjPGQ0EINujSJAD9AyCe0ek6lsZ8Aaf3dP2ezvpOSUnQOGi
OZ8xapjkvhdfnMxJuFCdSwHwOsAYl3v3fkphXQI1x2vMR/UMnkGgDPW2Jntn07Ceqy246fOfuiKw
Pb6Q5H0v/BdzlOPbMThadUcXhgxvJYfAZowfFMtw6gMUdHvxLcgYn0OFyNpheoQnjTFrutXbWgJY
2MR8OyDZWT1d06TUWm7W77wEL/Fy1WiWa7sQLbOulBMeKYEtk+JQUHhkVynX3U6MVNkzLAyEZFJu
HKrRjZ2X1omLAJ/hB8fHs6k44bn/ZA57edyVmJtylh6FTcYZt8atlcZS0KP86ppiQeOP0XSUqFwv
OjEOMr737895haP9oidhrTNRgcTLd1MmpxIpOMAmF6wmdhkXbd9xqT/ZNxf85BnKeh5PBPGVaxha
gaexKYRSy/BV7mu536mRhaDg/m18RIU8HJEHo7BLk+cixyDbBcIcSfMJ9l5DUwws/70eUNczhoPJ
+lWZIMlIJi5IEL0QlgjiOi+HNrnie76ssGql5+RPXAQ0vjU4sUpucOnAV2hG0WwSbE/eK8qSpCpR
0KLLCbpasFCcObqI/vI9o98w+PodH2anH/mZEa9HUtsIL91RgOIABKfX6ZNqw9HFkwZVtGUcobWc
6V4g1WgdydWznRABgY/ww6KaoMmyLyIg24P0jrhO00x07qPCt5JrJXtDelmwsfCyeDSSH9ER+O0M
N3n4jTTqPqUmIc3+BDPvjfWvbackbGT3HYQ/vT837Fx1KRGoCSiQRb1CpzA35pf+O8tFujQCShMQ
5/FIlgiD2jaP1HPD9RFk7pAiMuR0VLK+hq3pBCb18y7KpX/+HP5wI22ruWfbTTg5lD8xQukP4ajU
TWDwTMgzKcDDjp9AsD5P87BeOxTXqVhzCFvwfg5dqCtWRdjyXsmpWWFYJOKADTfbvraoe152CNh/
7KbcDbtkKEAemERhYi3WjVltqdoeBewATsIYOjr0KGpY9i/Ylz18fovd6xjrJNjzM6FSsJHoHW4I
fTR2foGbp9pSO7x3DwNizjFeBrzOpxNKZDjLFks3kbK6sfMnvKpbzwYYsyiVttMbUoOPs4nMXT+A
kAwc0SSPp+5dPG51EMrZZuL5VXdMSsInEvL7aMzwjtlcs3zkMUPpcs3QvaJxkwgom1Z5Tn9p5M/z
gQp5XnkaZEe0T6xtyXENmtuZRW7+jwf5lZJvGKx+jqcVg90kaIH8E/0A4EdDa00BFqijncd0jLgu
Xq/g6N+1SSsAJ4yPv/ADP+89JJjKe3V9g3iSGWPV/ggSDuSvOnOS6+iLrUaWICeBavhcvdvgOzHQ
iAoyRA9M/ErXuLMLKUu1H9puFlNi5FM7JPhsrHJXXf7iuyv01k3olINlu4pOkjqxaSA6gKtjDBta
xNa/weW7CbQkZjS9KoE7wCqGnNz7LyET61hrbpStIMpAlmkak/O+eRUWsfDrJEjxeKGRn8Va56it
NbtUbGcpwKCw2/5u5EbY8yMf7L2LkDF7USfJhAHdhFmrW335X95uWmvGSvxW79hRs/k+kHUg4XtR
iVO8TsPr4HrFlb6Y3hfOGJw0gwdRqFvUq0slvo/LI3z2u2R1DyXItyB0n07SzIqL5s3p74DavqW3
htdu21RXhNN2Le1dj19/rBhjzvfrjfVDQXWwVuP63I1+vWKLM12/s2I3sUGHTFbXOe4iMGIth1vn
WIkxTcLyoC6FWfA2hZteVIKUrZUckJJ5Oz1/+c4zA+sp3png3x+FtMTr/yxpzTfMrba9FOpRN3t5
Mj4OQjDgkYPPkFG1xQ6ODVc9SHCfiu2BFAjb/LfWQcxYOX3ozEU+Wbx3c57tLB/nFHhoyNvDzq1r
yO4efcYGd3Oc1A8Xto7Scx19BFbmJ4DRBIB9p0H9JEvaehRrRZSoZbDrsGJZ0K9viHLa7Xh4A1Qt
FfFtHTOR4sqUONJKUOnnKI40+6w8eGpPiaAIkB9AwzQyZC4ADYOf5RuKiQbNJXT9O5Rh03/9EyG3
O73M/oGSEqru91VSG98fB/lYm5C4JPlFtonaWrmmhVyOERYvf6i0A1bgz+ve5fGlFpDUCruLyY2+
UjRdVmQFBAiDaKrNoDLdc6J0sMv5dIbdvMKPWOnOFdXKpxKigA3NAzDue0WA02tMpGpz7vSO2q0z
C9lgKl9LThF5YroR77N/lGlnygxZ5DD1ESucWRKrp8lzaOhd903yVmuCYHJ7XM6M0W3ni/toscqi
eq0+JsctOzMcVKww0/0IcfcSXt+SgZxoT6Jf6lA3U761r3LEdN2NQNVQTgqwUFtzLOSTErVb6cRx
ihOS804AsyAFDRBk+LhP1B8FkQ7kVDUkifF+ooLPDEsZ3sB/bvvrNfJgIrp4CvDEUP841yNC0apS
AX1KVZzDej3mi4wzCSQ08j/qS+iZ31QlgeviGp/9CdmoDsF7f6NgydRi/OryqCoo3jhjAptr5BmX
nsd8MgErCHdJxcTkwN1589GRg4ZgFPfFvD3itHjj33Nh9W86s0Q/cekSfoLdB338N2omrHxdSJt+
PFmw5/eIwWoSnrZRIBXmCEP+zDRpTrH9vbrKdootzkM33+ue48SBvDPBj99XhR5CutXD+hfEUena
aWNtfVWHa7K5aJoC+6j6+O30QZFJbiDtEnOZfkz8zHLoYYrd3CqDJgoxY39jgv26RZ0DgDEoRSIh
vZYCG4HqLrNi+YBeEMmCKA2tGR3tS2UBXXMT5+/eX0BVN1XuNg2MTXUOMmTorZBv1KqLn5+ZBZAo
ybXcbyhMGXf/bPaQGANJnGRWz9IrXIQHxa9/OCUiyUL7/FROZcNquPvljAbbq9xuVPndblki4nrs
AVII/iEHp8pSCtXiN4gMy2Rt8QX0X65O7jf4KJ2L5ECiFPtAMRLrNL37Nbd4zLx37nBlUK5iMDr1
MBZVe638TA0Bx9WkTlQGBeeRHGRWBQtBGkbFgHTTWcLlEZPk1PQT29CW6ccGRzyXrw/O1juByQcg
+WZnLVC40M2OS44ihwB/pud76ru1rEToaVn9hjJw1mpBNnoi6hok7FWfzdfXa1oBogCXt22SWvVz
gJoknCIqsaXHVNDdCDza/F3wgt0uiqz81kH+DHSdsj8gNiYQQQAwSPIK7GVNyY0XogT0iU7C6DYc
XsZs7Lkd4Vq6eFgHg1Rgo2XM64I5rLplayutHKFVqISPdZFKo09E217+cntAXhNsxgWgEP3beIod
jqCcEUBgV7t65Y1Jc0d93n29hA0uHEyPFYX0wzM2seqnxPOoEPAnQyvuGnWlJ/TlnPeW9JZaoIcM
6gp4rDPm5B2wsZ057cjh1mZ6jYG0r/0OOdlcjnk7aWHsoVL+MUpvo1KBS+LMbipWvVOZ6IirVAl0
MaqgOt4NXfDZN5oF8hCiENiQ5X5X6CfHoHAXf6qBnbEJTUxkJ4MK5lISV3Rv10OAnXmNaV0tEp5A
i63VX6USEbqcyHspxsOcbgWaRzeaRtVAO45nUYmlGXpIsM1YT7myPdVNOF6E0gzOZK6YAdtGMrVK
UPt+PNHWIkH6CP1yuTQWpNwplmSYcDFMtUGC4V8zJ9NEBAqJ/V36j5VUo7vCwzfDP7wOJkMIwQPl
iAyNetkwGTbXvy6qk8FPIoaK4EvfFv2j5EeVO2a0eHvTyPLIYgXvqjc9O4HZKzS9MgWoyn4xxKdh
wy1P6yho+ruUXEFJ9ju/JuZoFkimiJCKJsEsUav/D+970ti2EwG3ARuLsrTlAG1N4VdG53IjsCt4
CYoyrUfe9+2IWzDejM7AxRCKH0PV3RXsM6keZhI0aU3loYlJWFEerW++nJLyJSnrCzwXTepq/U5R
ml3ws9BcqmAia0ul0jSMhmTMtkvddKXMqWl22Kojj4wQ4yFMArEq18DS/5qK+6wLBPNJum8Ynwj6
HQkahbyCSai9pUGY5WM9w0P5oStHqJADeMlRysYyII9UWhP1dGgxE/384oh5nVE9M4BTe57jsz0Y
3r8wKw8f8316WuligWADvODo0X1WVFUPr2NbyC6A86pEwQQ8VDa9WKG84ZfOGYCRsp/oJQYWWFoZ
UVg3jK1YhRTJ5+RztlpSvupc6hSBovotxmmG/pXDwKFYkmRMpEhYwqTn1inMlPXcCewF9bWwpX9p
WG7SFP4HaR0JpTY//wTEQ63yX05bDtgS82EXCSr1j3cYvjwAY9HUzuUqe7vjteMrlKc+ITlH1Gac
06acTeqy0ZR0AWrUL5s6Ig/74xG1tTMmBAoUpPYhtpfnVztuJehqU5a5D0M35Fmi0i8gxuevwc8m
GESIY4k0QcwzF2I9b5EBZREAHGuLtVBHy29xeKAzNTDLZwNvUr/Nohe/d/APyzW2TQaV+452i7pg
1rQhZIWYPJmw2DcqRCuRDf9AqhtIHz8OMsRNBpty6pLA6yF8dfEiCdpq3qkyo3rIL3Iv0lheCVYP
t920HAmKHnigLPbnLjcVj4e7dY9ht/1wn/rLqFbOrD29QWtVnE+GUGV8HjVHWmwTpqeebYKNUS2x
O98I5QIc6AemshIi2XrjelnsxhFupF6ZCZfSqiIYrurUFvH3t10n/4om/qR7HsT4ftc5nsC/h5Z8
y596WS3Q4lxjpYmPnbsbkfr4mM/69rB1cYbxtfpQUQq4VWPDCJOhGqXtEACTtyIe2iMk/km+X6+a
i6/cBzZytrdbroz24ff12TGuxxWQk5WPXDthDG2ATH7jvUAZiA7DrZh3+4AnAjHKrRFjnPwMMgBl
9ZCVIJpVLrmvbPytgC5sN7Hrg0syo+hdp5dmxRDU5t86HJt1OSJGNxFP9fKNsibtqzsr4VbQcys9
IPg5xbfRN4Rdgdhs37aI6BsqWHnOYBoMEloUpQCwT0p5CByT6i3zIJB9y/NHP0acsekVEgFaY5lA
tvfSejMoQ69sNSvoluLACrdgmhxia8XvhZHpbxwLqmGdqr9z9ipPiGCU96ebZUiYLt9INf2SPWOX
IGbO3fJuJFr2e8ISWq41bcqQXnjlsvRUTTNyWRMwLyNRvxa61LTLs/7BQEgXSecYYZKkpuOwOdDM
3ivu1fODjTUJGN2dZZrhlOOa+pUJDtEPLK67z8qwGrHnKyZ7Aw0cZdvZPYgrKMouzOzvs0UsGJb7
cAKG+4nIjn8JKdW5L+nSkymFuBWSwtvZ+ZZWPFUwPsYRK95dAfP7vyux8fT2ZrLEKXweb2P+zzWt
hZQ/mlm1xnTBbATKYv7Ve4LFzewnM/og3yt9g0glVGm1fUdzOsoDdbfB/oWrIwf/pN1kJCcze8Q+
UXo3D0qWHCYQJxYUv07W3w8yl4D6kfwdpRi+PDgzJGK1/Pvzbf/JvIU3Ewn00qIVGz95gQPRzieR
5HSQbRYXILxvVlAoSKCkoEBb1HCqfeDKYyr7+EFflUhsb8f1CZGT2fFdsyn0oNR3sQYM33mcryFD
zRwkz4/OEcAVBAJq/Pbb5lIk/08WwLIURmUg5ur9lEoc+NXGliKsJq6Y/rSSgVGcPse2EWHtaSX7
/K3GlZGPbkiYTXrVcaGq35uw9v1VbtJwyjJcGxUbf5L2bNbZxOm3kefrWWJartHr3zPav9qf8aJg
eUZHLwyAfL7caql5u+cqcujA1il7YnLBB5WpCYAmq18I0vhyFuCXa5xoa3KXA0DdoPLDfiCGFGRR
qlbRKXjkCesuihF7OcDdd18zMklSjN18WvBPstzU2Py9M06C60Y+Pc66x2VyDxluvrVRCffrK3LG
cuQp86qlR3Ch8uAqfd962a2PYl/pBLc+PAXKFWBIfcmLFbISfCcJ6MbFMZs0YLmhkiCcZa+mM6yV
WRF8tCKRS/EUgUCIdfdrxXx1ybbC2hnUIfv8J0RhyRulvdyUlFGCZR13uaZabJfNQl9g89ZJfgZq
4+IEUj+N7DRupL7jiKc+ysSPASPO1NmbWvOoHm3/8PlpJzsCcePh7WtZHvjvveEQTtGqg+axzpoQ
BGE12crzKZdLmfGTiuIJPv6eKnMXFah93vOpPBdNwtbQc9XahwnAeztQtsEmqhDBQt6VhM5/R9GL
ZAzHB+S3D8DR9Kz5L5KefpOafL3vyP9RmvECi3QN/psSk5PYpmun63PKHCqLTTTK9lz9V1IzY/nH
vul1wojjQfaABBbngtQjKlqWYL3OskJyq7LSMbeHROX4ckaqCzDL8XRNIthf1AVVzHYoSSsaDQsX
VEsF/X5MMTx01wYkkUfjYGbK9qwJXipDB93FF/FuABb1D8aCFhrR9emYw8TNXBQdrqoS6MRyYBn1
qHTN8G0LnNeD5SrBNV5+pCjX3AziuN/lTFqydfvUzysWWUwwWtWGe26xUq+XgsqSxZEpkK4wjmB7
1cPFuFhNrcA46YKQJIC3Lk4AVGAFpiekburuhqZS3RTz0JBqIWXXb97koWZ4pJcb6doc2fOwR9tW
RLuzpBS4ifQsrmR1YSLi1+ztc0tHU1vdoTg0EWXy97cCKR8jNXpycZAzzddEZqOZcRFL0PNLVl8J
skZkuP4V/iL86FA6hFKj+67LK4eGjpp5uUJoOGsN3TRhCC24saGddMqWL0oOj6FTAZevMGhRj8RD
fwoIxIVB9fyth1NX7QH3qSCTzBx5p+4Q8ReMeawLzHjbc3yoqRuaU4qd2CqFD4r+OMM1m1Rk7rnb
YM84a+ceAgrolBcANSNjb42loI1b4+xkBw5IpN2+N22tJdbPK0nk4B6Jriql+R8QON1id7/Wno7P
EZ1Su2IhymQBoyyGIe/Wg1JTFYXAn6EubSQtQjKRweYAcKaOAeWBrdAtYO93Xrm7aa2+gfBh9ruZ
Qmo83oZr/1X7GOdMULauZ4REQZnyaQe0lYMrfB/24Ex2aFsKxTjeT3jcv69Gs2e/1W8M/6sjDsDa
jDPA61njuUVdqWR6LOd4pmJ/sqhJA5u4jeVoq/ExiXKIKrRgbex56LLti5I1Qf6ZxUC6amtg5f9x
jGigeeIO/FgPw+dKuC3ZU3FuciTfc9f/dTq5DO4Xn1PTlf8WquhE4xA0xOE+K1xkSL5iWOlfWBST
9LwcrX5PxXswwF29DJj4v9R9uKmTSVOGyDJTtUV6Mcvp1S9/SG6KFlhejU66KXDKqLNtlK22syxX
bOcXb3cc589HQn4AZ91rCvtidIpIFlgM7ugyaf/IZN1+IiIihMeZwsg0uvbtSE2KlxFmv6iBwcoT
o7HzP9N8XufDUZHEchOgjkjz0lODUZtlMjyMCvPnvvT4I6WbE42T3Bg+Zff9tjFr5Yt5o1v9PJWL
ko4OPkhKX1qX9raZ3NtHrEt0MkVyR/HGcKnJHPXX4c1BdQVhrfa3hNRqxWrOD125X6s9XTGBqJ5z
Z81v8i0nHPdUf1yXiYAHpCkz+RhJBPKeIXPhDKcZ1gp0FWZklS1s1TrAdCO6LSDV/yBG7cUbtJhf
zDaB/AtNPAXH3sCxNO9++IUcHiKZJRg3RJkamuRmnKkoK6dnd5nyy83fzfrrQbGEE1zW4VIYdm3K
VtKQ8V/DEfF2BbUWs/ZyGCYtHmZcJchPhsk85o8xkYyt25NRYIgRS0WD0Zqikj+8JS2TGYwVH508
UXtSZtTatwtEHyfKUeDD4E1K/qRvQbzL1QJCnRyBeTA3wpgy1osvQXpu62n+/nKUptETBUhJ3NoX
XqsgBpml///y9nQfcLrJdtD6tgVhJDTmZBpc2jfFD5U0r313fM6zC/8QrWl8i29IdYa2g3djsg4Y
NV5zCue9rOeYzoTBNWI/5HXgvx6k/n+sClVSFBzmJ+2sEgOkAmjA01FswgJ1jzNOda7lQXnMHZDU
UABPEySiIU3Xf2yPR5pwBP9coXy8ICx0ACIvPBlA4U0StsWEfTp7591rtaaifVzYd6mQhmNbLhG0
O7+DjpPq5/L2w5Tr8/6wZJgLJqtPCplzXE6vkzuIm0qLc5tYO1I+VeTmqUlOh83EO3rD0nThvfEp
U1R5L27CfS3WQk1528vMU0M+3+ZiwYdWgXWCMARbNUubSdj03kOfpl4O/V7KUpIMTtfrrYUH2xz7
BGXCb/oUsPDX6MsX/Yq6A4rEDAuTAxLwLxp8icMiL4Uw7RHdJtZVGCooEuSxfFTrUqLTKlL2gPrr
YYUHqwXB0dpNoFiOUfsuOiAVCCiI1xtq9+8CKunif1faGZ9tSpGfyO+e/rQEufityb4sSNa3sB59
PfvXUZPqvrQzkm/TqROpLgbwWfTQXxbtzNIgswZQFRdC3H0R+P65SMpWmumko4Ue0TuVIlOL4/0B
h+x94I3TurVdw9jz68mDWrO8pyIT0E09z7VdMVpb1DS3SP2WNkJ8+9G6QQwYS1CbYye4gP/kvJCa
e+K1GpvpfB93Svg1H9fZulGBG1sFcmjakhM1WRnheF4LGn7GeUCK4uRhS03Ba3sbpC2V8W324n5l
SwndL+McAeNC9830EbL7Oh/0k9slKJI4q9OlG+LVPt/8Ouar3srhOK1t9mOUHZHNbRmpY0HmScA+
y+I34zs1qnPvy/YZsxk7qLNsB+i/oq6kA7LXwRhHeIGejtwJahybAKDFVxn+Oli7Sqp7FfYaj6OV
BoqjygPwudMCR0m6qD03P0mPbinlvkMArS0LFnqQ5GXhX0N0w+IoAmxY10n2U/5KXSXyYnEvF/Ks
WLazo1/cyZvDOYfrmvd9q0Wsro5wv4GTN+o81HaC9OJmeyDLlXpbVmbwdw2l34kDlAFEJuqszwlW
mHZHSVGoK8wPqql0KFzfHcHoolS+qctL99ZTSeVDgpX5EwULePniD7LYNYUEmow8TKGAXrOLsvQB
E3lkA60tb62wZOui4OeiS24S6OIUqAdeXJmH/N8Ql2n25Q5g+L0wwPy/W7BV37KlmJap0nMUNStq
5nDl3rIarx8CDcsLXU6Nq+o5MHoTcUUR7ExbWVwNBzAyQEjVkPmpWUIAW5AsdCThiU9orETyvKWC
5a5ASXIl8IWLcy53dRMW+VWEouklWdSLiMEGlpYOQSPooZQk2Z8yCnmTv3F0REgztDOUKozglkD/
OltFYzlebcrI5cjJ/S01J1OS3LLGUiHfegVb1m4JcLp1xow4ceZ/NxsAIGmrHKs6s8gjUdtuZR38
76kj0DTC06iPU1sWEFmAP/U37VNpbajtX1Nckt735XbER5qvQ9i5wQFn4so2AX5J8Wg3jg0gT1uD
bIGICv1OPHIHnCkFFzyd4sLlTMolgev+V3cK6Bo0j7NUXMhpcWw4px6p0fDrWPvZy4JRg5CIediP
PovjEO7cSYYDyLysIiW4dRri1wNr5AaYS84Lki2sGW2xB9LBtfsa65iUgK3K1vp3GonMkkeGx8yX
erUZEY6n/in9b3RcW/LRG4tc4IxqURAByC//2jyifenSZ4qBfjB6XhPZXDBcadAtYR1Xr2FBbXyJ
kXUlNwRLMgHXQSuYEwmMGb1FbfcyJ3ZxvO0yOs1nZxMiVqlx/f0n+uzamE66NI7p3jWEKeFJGcyo
2lU5cbP+aSF0lV7MxOVHj01dv66bkGNNQtoG124eA4afwaGQH3wdWNgG47APsNQxNRm7FG2j4088
mUQQc2B1PYZ/0u2b21vufqhX0bWxcrL4ixf/M/DbY0PmvieISVhBELb/7i53s9cawLnNE8+JdIG8
6HPZCSVNu6OElK0z9wR8HvheooPgvvTQAFSznclsLXU9pHq518jrwzQule3smKptLcInLzUrNw2/
0COLCvlo1JtycRFzvzRs5SnWnVBzyHAwvjD8Iu8p4JruwfYvWRL/+t6YA7OsqWKLCWBOb/g+nK4P
pwCQRlN0egQqgjt70d7EqLg6SMEWYhkVy05tl5khq+4ANEG+kRp60/qe6HXSR2PWr3Qwj08JNTz/
qBNWeVUUrOnujhnU9q5Powpj8yw7q0y+EsEa+55c9AT+oAuiflRglq4BSo1hWB/Cpw2FBY8Tf4ig
Jq3Or8jOTBGEivhKHuedPbuOa3OOSOZ/pBmtjpWYk/PbcicojMOiFXjQ+Fn+ztVu9z9OsTLS0mN1
hRKgsgj2rYx6rcHmcs42tDYgDoY2/i6MR0hzfj+xUjG/a81ljJcv2rteYsOR2cA8qaxnAVVPkseO
fBaFhwsy8Fpu0ySF2LmNEz6hDfIS9oJTUXKrcI+MOC9J8a+x9Eb2grC4AK8JLG0RAkV5awL3pDRP
n2R/R2WmPU6nO/1RsP3ctIcMFNzkBIZcEY6t8mxk+QOjQzETTu+SJZYBHI3EWxhyIdHFQoPxLT5v
gZ7ib8AIFChIq8rP0KWF695fbEuMETuX0a/7YpOww+AxQL4Of5zeAA28/g55Cc014LUc6wRQhRrh
x8IcX+s8UJKJeg2qWUvPrkicILbqqLk9Ukjso/lC3LVNM1GkwolYdetOAUXz04J56t6j4LbajhFN
9KRnPzG06V/hQwlJc2NdYrXoEVWJ1n9RBr+7PhTI+9JarMVhlw1htqYBPiOx7U+Sxy0Tdbay1mOe
JfB1qetpQBOaXeMfleslf200PgKA3/L0cRuEoMr9Dz93XOy1kDhtYKz529s0wgpm7osCf6wBIVy2
pnEkfmUNHFH1dzlJAmNFnvWtrsrTVW/xm/fME85c78Isd8+XCcqlPOiHy+pkd7rYQGWuBcmGnoJ4
iLg0uKGbZOaAbOvRUvHcbxkS5Yg/DsqlJJnv7D9EJWDKfgRYno2vfS++QIY3lw0cvRUMHzAoAAmP
raIVNtP0jN8V4gw6QJhtnQpU4HNB99IcghgKcsP+oMi/90XJKnoQ30AYLDJIIddhGROP3Mb3RWWM
tMKqgpgHiEKrSPFb+kaAsY3HcXvOImPhhunVRQExPoDW9bM0EaPNhETx8dniitGPqhAZQ7WibVNJ
gnDFnP6IsZpCp3wMra1N2PecbzIIyh9Eec+MhImq6Twf3H+A/hWbzryHXDclRyRZ/VPC2hK2Txsl
psILqr0kQMQSRfCF+zvgUV8tm/wV0q9PbTAadY8GUFGS+phIgVooyKfjnGmIsgWJqLoVYLtyw+4K
y1N45Ex4cSqOCf9ENLzpqkEYbH4sYLxQdQ6lf3JD/vyKUz3FfDe+UV9obiWKg7pTZh9b712zUKEu
GSeuXpCNhxt6HAHXqRPzfkGXSR+AdrrV/uL570ml1d05xZcAFYCGiIg9OxRjkVEfe2taJ+V2JiN6
cvvSvlihN+EJCNyPuXtMSVhr7CgKcZZGxN1CIh/2M2V0DKVMnmz330qLJvu0vFUhuj0nSTMpY+VT
BPAb4IRTDFqQ9S5RllFju2QjMyULU/8gPo0RGgE61Qj6pGms43L4WJT6hQsJIFxKorIezLkycaZ/
Q4qW8wMwX3QCnEZ2HoqW7xBhPBPtB0rZXrKSLkmxdxDhMZPKLQ4PDUhhEPhKE7MUqGpJ2xf8G9Uj
+HcgTtUicQy+SJL7TLBYDOoGYKET0fUPUIhHO4zk9qUhXh91FuQH9YirOS4qWgDwCBId5bSaMoKE
n0REumbmcmFe/0kaUbXqVIjfqa8GYhM/7h9Nk2+f3eWSD0PdT01D624WjDTAdM3+lSMKgjL6jipy
6ken3wSnLfGLB2IRUEpsREN6j6cio8gSHlkX54x0kmTBVmG0Vi0XRYNimCkFkCgwsdkvjUywQRD+
Jx+PDWOrvS0B1fGynYsYVPYhhthTWnocG4F1cvWWE/2h3WWHmEpQp6rkHPi8kyXHsH4ZGU/YKt7f
fR7vA5jgdakrYtau983LglqP7mcWSFyUoFydO9e0w0fXN+eBuHIheuaLD8NdwSc8b+W1OUt1qCua
Ecuyq5nv7UVa7H1ZcIAuDSTS9N+eprdr2LvFig39hSuU1XJrdxUbMKwVYdHI9lGqjNsPPCaQFEkA
VVP40gCcKDpravoHQJ/iJwguvi9Lg9k1wx1P8FDOCkCKyaSl4L+jGD9i5tjK+RQmYEqdAfpzLQbv
QSY4FayAR4f0kfCLew0IUZRqgsB2uqF05kAA9QZZM8DIkl3MfvU+/o4L6sgaRCLYKDsML0SSYJ6e
/qVrHSRtSRBjHj/C3ompEeIFYSEkHGNzmeK6Y9CKrQh6/ZCRjuBd41RT8rgGFIRKHmAicJEDRtk0
y6ovnCBmSApX2OK9mE1gCI1RirINLPoj6vLNrv6V7PNjfCYgqQNoJ05gtJSviV1CoL3Kv58pwPjE
FfejVlxH0wW9ykvDH25HECuwBvlgcpjiKW7MJsVYdWMG0YdqIm09Hu3oIUILAhfg/JwYu3STpl88
K3EjyQv7lDV4RTIaaAuK8eVMNO3q0LeEuU6Eb2DYS2ENnkpd8ZQS+GSqv4Onhj/PNb/k7hI6QTKh
bRjzDutGb43Bgbq/rqOhLCPXfvHS3CBKweOrUoYT6nqegqnYqwFFgj1njouAf1hwMTG0LHuLn0rx
LENdpgiBPaqAFkr9B7Y6jxTz4XwyckYxiUH47WIH0mZPirK8/9WM+piv+mZ37p3etkTPaW6tQxO7
bMgXsuVWW7G5irt+21XmiXRtkI0+rM6yplPhSwTYq+2+2frgv75QacpG2EcxsmRJTsTTu/fHvJoY
fJtKlWY1jUNrdC+3OopXp4WtCGP4ptLKK5xr6mI5hvXgOpupt9Fsz1Y9/TjZkeKoOXy2qccK4wFF
p/wVEuRVv+5QCCb4YsUEaiiGeokhI1quyJJSQ6ydDfwfLgQ9kv4MXhN8jovyU2cFmTEsTus78cB9
bPhaE2eiTvkzU7kX54M8WsedZH1ieSGIw8T4aTMEteRmIddkEZpB06YU9/DitI1Jmka5gI53I+AH
v+y8qo8hR5DP1sljpLxL29ciMboqDXl6+xpUrt11tqGf0jTrjC8w2J7FFldqIt8f0qzfNRW5tf/y
hjB6B4KHWHGMX5UdW+3K4LHGMWM7g+dJ4Z9dByEgwwyh8whaHq4Xs986tlI+ydaA9yIiVDnszHSj
kwGCKtHXjhSYZf1L3T549yc0k+YKn4SuLmcj9/z21wd8ivlETatBBkPgBNFmjqqYLal03OO0g6AJ
FCaz6XpuYMKgvnpll+Ib3iUUJmOb/eyQdDvyZXKxuFbWtlwdsa+R5V7NBgATODeyjQeBQiwTY7JG
HY/t/90yVmHVfW9TLIOZunwYtnH/EtaGPmtjO/00MjJIm4S/bUYnvIcFtACgTInz1psuYeyTAxP/
S6D0WyQPOsQzKNxeUoG3PgkS2oP+LMlMwrRnnaLWcLeszJiJ8/5Z5Pu1MGencsMjT9YKIitSLpjI
bEVwCdEZlXr6Jh0mfX+trdSq2GIDS6AyhqMntR1ztjIMpZhK+dGaEHT9wuQxJ3PcSeLnjrYAosnm
IUnuaErkRCjAPnD24+Ko7AmuwFqbF84O3i49lAsnsuu5LD0bs5cJYXIomWUO/FbN+3DFI2MLokab
GwgCxsv/81I5xRXMYw7Id0QDPWEIhPaUDgnV4ngP5Uub5K0/k8iojvTW/+AaK5VyOVduENgGxKa7
+7LuJNpDFYvJyhACi2KzUIJKHpjUPHgJ0Q7swuB1ca7/nF6DlUcclQwcQHy5ikUa60C6jGv2vSwA
J4x0Pf2bUTbCHov9V8QmHY5eQypNsPxuHLWo8Hrttm+PPemdV/MF7pSAmr0Dx0f7vNCUdt2l/xOk
wwsQHyF1DEGI2mZGqDNfLpj22DANl/839rR0dKzZ+GsP8T1gKkwL1hwSzpw+UFL60ekA1uhRFOxd
i8fmxZtY9uzlnsqMI73i5tNMN2AMP6MdCrNxTXeWJu7XVM8kKyhPf9VL/NdElQ8K+ROA8F100zTO
1BG9AMkAyTw/GJYRngPg5yIdLtPu3ew7UB+O5uhgp77knCq+Qa6oEK2ihHQziXx69wh07yI04rSx
gPhvXqMU6OZCDqdla8lvgzJWcmmkhvlpNeaP2HUlBXlfSi6aBq+EYYssqg2/PvQ+CzIsZuZhCuKW
CXpwozHI0wYkl0v1sW5X8VyCZPxBcDKey/MT3jnAyqOSUk/l7dz8W7LLkQc3EYylUf1W2ym/rAjF
t7pKZVleEf7eShxeyX6HkcIndDVjdHTjoNQ7ofSxtmiHSMEzTeXFKYrqiNJSaWeGK7Xk2DGJD6DL
IQDHszHPYDEexl5Kl6gClUUUYQ5rrbmbltyapeKT61vw/+ticyCED1LtbN1RdBFGu+9cOEfolfI9
4sP/sNXR6frRFljz3uikZIUPVCoGXJGxLxwzQA97/NnCMTaxhPBBgC09bsNtSYwMJ1hsiT6CaUrO
KWYUyodLrWTRh4lnbhjLW7KiVMQMrdhE5i+4GfeI+Ai6HzxCVWwJYUgpv/9WK9t8ZYlHX621i7tY
/crZlDWtb6QcUTAhgNB3/IVGITfD3JJ+FgYViM8cUO4UqPRfk43bCHfvUOon9QdlBuMfod9KbjuM
lbLBmWcLmGs92uTMxMScf+/fr6OrPPZSM0k7kPmiroTTBHUYl6DSsFMRZMyrd1EgXs8HJORlDaII
89rwIuF/fjNf/jf/0JScVRyZIm3d7j0nlNEQtmmCLSoHv9CUPoF9SZZ3kPi30q4WxYukO1HE6n3f
wDrcVMJ6Y4RC8ei68D+l/c8WSzcbuEuFEvh6bs7RUQ/V50oUXhg8frIhQ91FZUBXx/zb7UQIwklf
jNSVuGa6wuM714C1G+CUudXpdPIKop3OKOxM+X7thtmttBrFw/2/d+Ar4vOXD50Ibuz8rHk6Urfa
BTZt+R4wnwoaKjBbRV91fVvbyQO2bGsTZLJnWBJK5+Eu4txC14Qshsl8UenXHZVsn5uLqHnCBt+h
F7wCyhP/yitQUlEGLirvBzs528d3rIIJVHEKmik8KqeVIq1D1oSld/h+pxyn7MpvlQcBA/fHvZCr
H/tyuFjCsQDC9DMHkuoaNbNizzMvQeT/hMwgWU3EKa/wbtdtx2ioTBT3yCkNntujxx53vQJbngou
KDqpOX4W/oP9UtnAa8wnBwWD0DHGWbsVRU2IAQKRVNhftDrP01xTwxOTCARb9FyBUiyAk22d6cOY
juFp/DnNet+3O0oaX3KwM4y39UhE2aGXfoGcNOnw2+yNtlfG9DyC+apnS0YSDsnj2rklLyEIzpk+
l6zN1EYze94ZMuNth4CGtiAFZ6oo6CAw5VtYiP8AtJB4Z7bxdB9b3j9i/1vCvrdTpmLSRh1ZTQ2f
/O1w3+pWVv9L2RyjTlqQLvaHgWEropbRB2kTHz17qKXSiWGDvr97rM0QS/kTuPEaNYnh5mSmQy/H
os5/h5IsyRZzT4r8m1kItYbGNbZK1HmH7H5bQLCtqBLKsyGKEJyF6SN97tJDLHMHnLig57rb/GtI
vtqOEBMh8KnCRk9zzTZ+zgA1CvpFyoqTQIWO7LOANa502k77d1xuO1lZlVunp3KF2wU8w7RTjhyv
Pi8N3OlvPGbBVCvQfMeVycJSBe3gzhuWOB7vKCTnHwB1m9jFw/lp1Hk9PsZ1mb7L5IAiXaA89Ylk
K/Ogqy82/gSNnhsO1IexGMYenoE8hsRzEi8RpO1LpPbBwbgskLmLgFA+/4UTqJvrqIKjnsWsbApp
9uz+kfo6SdOublDoNA2w0j1SbKA4ZfynUcEW4WbT9sUwuEOIev8eN9O1CzngQd5Y+t0JoyJ2efU1
qaaCzVHiUzTvQoVhMkE9cJcwJvvnxhXgOfz7r9ImDuMu6qpYcMxEaTvjX9F7fr34RGYl29V1e8P7
UIpmA+G8yd5At/xSr4kK7s4od33qwHeOp3IdyfG/ZfQmzh7UqkNVsHUEJM5Kzq4I7W2RDWkwmjiy
wHDkTGUpDLGmE4SoIe7AeW7lY1YKqm1/Un2cwesF4Xj3nt5aMLdN5wqiKQhCdfs3d0Rzd4ZDChM2
IM8puoWGDLkt+RjCYoG6dAl8pve+Yfj9kKx6QDTSMHAXqHgQ8esqchiMV0q4QKRzBTAvL0RjaEVq
traNzfQn7F4WWLdylr7v6tfR4T00gx+eqZ/+qFI16iO0jfe0Ss6B0EaYF0yE6OcwhVvWkP48K8aF
9NAbHp2Buq+Vfdyq/klnp70UUT9MhB0SI7ekrTKBDKZQ5pN0Ar0yPxK0ihS/Lqm257Teh8Me5p4u
g8SHX264Nq2xCIaRDlMLutVROh4+K6/IjNBIRSK0CWD9jKBdGBTIF5+/6cW/EW07NvzKmyJI3sZE
7JJHFehRlhAOh9EO/zQjpFzjw/YPyeSHjOjX9idm41waS5+NhGDCSLfc22HI1XEdu+Cjj7Q80TgZ
d9rjC/tHBi4tdrwF0+svXT46PKPzJEThMJluZAz/X4zMqrWVkzSob5NEhhztL8Cv3v5Dm31Wdaxb
3IP+p8JLVy5UwjtJvG3bqpjvFwr1F6Q/LVLQVGQxm6D84BxQ7PQPmSKEiqqJRNasfkWtwna00I8P
atJY1Pa1H7Tm+08/49xaTAJaWFKbHplUooq2CQA7SVN6ORsReBI5BGwjfqNNvr0MaL1uhaDxLJ81
QeHrurttfjkIvA7oOVD7byK+QfSheipNxh7xSl8DZoyaCU5+9WlifbePkxdky7j4OnNg3EfGCmra
kypRb6vR6JAZpt3AD/q44YBIfUpwEcQ/qrP2RlZoghgsG+4USUQw/OiWKkoBOQLwt/cvOIBpCAiP
/nBxcS65TUCSojJkQtbFA/uTJEKLGfvllpamqx7N1qJgLTYl9BTmLldKkVbCaQPjGIHC9HX4BzzB
odGbnwErZ9/i0RpG5ixMAlIiFuEBJkksQsXObV14ZnbAhw8DRyXEwTXIrquf1pqxgnNqQGBH5NJz
4hp2JJwNvuxdBZgY9C9gZjGhloeRytreEehieWL6H1TA/BJDkCpWjjTVRAEz4B4uc88diC6++8I/
MeyOSsHpOORePjXoCkqqEJjvHSOCCWH11N3YkVOIqsNy5YSt44nblU1+s2tF/sQfvDA0K+8mW4VU
4Orq3zcFeJtjs3hmnY37rtUL6uDx2FZ5c9LgfN0bLJejtvvywwVBbYsycGQ40Y4GPeHRYOP5BHMU
0jcayAAI9E5HP9+7OtjUZb99J2SinPgQvy8SHTvuHGqjRLMD8na32dgLsh9BWBv6hwZoXO+suqmR
QJt95XDeZ3c1AT9EUdJLYlDI3ip8RCO07aHBmHOtsHmpBHdcnjM0/F9tkW8hctgJMvTEcGIqeXf2
op+ZXIhwV2F+yJZODLSXWFTgjEKuPFB1UPW2YeHb02HXGbu09UJNsLeBdg4r/0UVadZ11RrnQVck
7ZsjYunbP1DqpGlu+ssQpf3BKP+d7DSnR5Y/608ntklWIgTU/dr09u+sFMQem6cK/E+xi+KSCxtv
eQ1C8dRR+9tfVTDs9+V1ThPTzitoAEdUleLcYnuxSB8Kt9pfaw9p2H7KzosEUT1XQjSK3YnWh3yR
mJkZ/Y9bMzLsNktm4XUbbqbfUoI4Yk/e8zPi8bx9dTYZl1C6oS2wjqQGmens2eObBd7fqX1zB7Nk
kF6vUBgrCmguBBhTnLmJhTrD4/U2deV3udu731rSSCXCbGsQsrY314dOciU+EPf7lNsENZwL9rD5
SOQQE1R5ngdsMXWPg+3TqP61TOII7lIsTlLHSclhPmeQ9wnJdbT06yOdP+2UOaSjO2DN4DULwf5u
miXKQQB0Lgf66x3ieIw5sAEUq4sTQPEL7ldJvBnJ+6USuE13d7bdKK7j6QAz6x7dPc05K+hbw3N7
S8pO39LEt81KIvX4AYBrAPyrU3QW1xsCy0IgM4p6oJaFbUTFGTWsxcY5CUIWMDZwu8hvJP1j7miH
v55DYE6Mlz6OwiaVo7vU/h2jXT5SuSwCs14ntekyj+QUSBg9eRtHyyfz2r/ntrqHIQjXKCONz8ph
4AqHMloTcCR04Eoiua0PshByel/kKBPrvIlGj7kAuDQZyc2kedfun22CrmrVSf2wgSBi+47X/scU
/vhMcvbhlW66sVqyQB+mMwskNlJPrX2A+I+Wi4oE8t1WP2jJXsT0bpWQz67dP/Pbf1bCysQglvb4
Ee7UvuPtalWL7Rn8Tbjr+i4m+0yPkykSC9gNSPYaMgiJ9XqPii8GCkwbRXDuQSqrLF0xsAYnz62u
eceQLPrn5st3D89ywYW7OYGzxxPcBXs/7JkQbfkKPemwu8GnTOSdklIh8ah1JSiLY5o6G2LDlccJ
APR7MT0mP34lSHhKjT6HUHuWxdNBfJlXNVmsdEJV9GqhAOJkzkr066kLp3WvLewkwKU47efctbyK
reEiy9v47NdfFD5RdEOS8dgfgnAocw2Dv4QDunwOnn/YdD9IKASUmI47DXSNSs/Bi8Ks/TN0U5SD
4CmeqQ1DqBUQzy+HmybX9e6Vq+2KWuJYtRimfeD3Xtc6qL2gzV3DXmZMLXHIZz7uQxnuntvZqR8R
RviSb5uDbU/JkzPrO6WKkLsGgM8U6zzJjQxQq89ehSuHcJSvTebqKOB7kbOolGH04I8dBKmreH6t
k97bYRrS/2ne42KSMqR+lSWswLh4tacsMVaz9qsevuVMAlzO7ExrNc3Lxtj2w5fU3x14xrQS6Wuh
4VXE5/qr3T6ceEMODTlAOqAmH22I4T/EIt36tGvIC1PVHnQTfsF2IDz1bDP8mvs5qQsgtx7DQkcO
cZ4CY+rkqBSSs4PygI3euHRyBT5VhqLw8/7clKcdTdd8h1WGd9v2O4lM78QNbJgNYHZ0LHOQ2gLO
1T8VY3ZkujkVP4+p0okN4aUrvHsMmC7kj7lEgFwjWPm7IAw0F/SVLwBe9agKGPZouJpjYsVeqag3
aXpDWGMTCWeqC2UyHuVhjNWxviG+C48AzIEDbDlqujW4WcHpkzRgvyS2w0GaXKP3UBlHtGXh7fcU
cCXAM3vNwaxBInPHbdN6LccFwstJmuZZwaEDHHAWLqsbPn2InOsnct9Qo+Oy44zTLPaW6CONaER5
rmeOvC2s41NK3OVS09jwzE6AkGcDYUT0l5gfLpZw+x1/wegJ4+nGU2QROwISzm+0bM/odUDk1a/b
5kp6kbC+r7G9NdnITRXenIBMakwuMpwudXwB8nbQIgxzizvMYAfU+UNwLMPtR9pv9HTXu0yqJYC7
RS29rEKGmYzkny4avfrAU0ibibS5vvyiIvAcQ5FcROEHrois/Qwu00FvPTq7EbHxNG0pM8UbXwAV
NcQeMmDakd4SAr45UJvdQr83CN3JBZPO4zvUc73WdAAlfX7aHh6iNQDDAkb3JP1IPUr89qzG6PQR
HRGdxMQmRBm+5IBEvOJXcM6GcI+8lZD17JiNuXn3zfBa2V6Vi6pc2K8aIilwZPAgwgFGUL0x4dFr
c2iUWbwFxWfYW0v1sBJlnWMXJ7d3tnqmqdbQZkjPkmmjZQ7+BVCLDnTCp3cVWq28m+/XmCnI1WKC
GWtxrOnCtreMSKjSQNozFi446d02uQQzYj5AFbKnvdSIxw45H3NK61myLZy91XTILFLbn2f5wJFV
2dR46iwF/92rkRa9mG424VWUfCD/hxJd3LQP1R66XlTk50cW9lAV3G2Mgl6jjaw/7nK4Stjq0NET
pXPEXvvsXbqHM7n7zyX5/pJtQ1uQdOwC8FPQf7vOBLSg4BgdbDEwgn4sGUyJ+nTvlWiJVSLVRspx
/SzrF8mGKa8E/eil0NR062fhfuVqTES00nwUFeOciHyxQvoR03SH7RPhkyOe0VUx4IC+wBDYuYsW
R61yzqcPAWafnfT3QEO8ar+Fq34kcRbOzNfAffeeNbPx5Uu98+3iF8ZwuW8U6BRgtEEtpx54QooZ
uidJBJ0I7Tpbbs5HOxkeczgNHrWMriXatun+W9ddTV1o6qAw+3TfAocil4tg/FMrLY6cQ3DzV0+E
OBndLwusPXNf7JNS6mF+vso1lY6gEIEZkxo6Rc2jl1e2GHSCarbt41cn3U5xNVIThTwOMPDlZUbI
NcS2ckqEbf3LjPadr/9b9KPTa0MGGc8Dfy1cD51a+5f+W//PtK4Ag3HATfAVPOgJ3gx7Si9ldyAZ
uCLfgjcGglSrlmq9hwRcbziQMUtdtHnl6F3DZ4QK0VZlOfFta4acADFJtV2AfkT6M7m4BPJ9bbNC
VYsJ0enzBwirV6PaOb957cQSQGlNgaviNX6beQzUXkzkDmqhL5GGPBJpNRHmZvR/Iolqa6AcK6vq
erZoB8Ce7v+7dzg9wBNYsUYjyzTv35yvTxDKfHldSqf12sfaqI15d7bdHxRhwCbUFSAvY2dO/pkh
CCNtNtcaSbfv0ECylcAHzQxMCpp7uukhyCuEfAJf9Hu6dp9o7V2yzSrr2gVlVo/1FQR1Mzgmu27w
7LTGQJCCzPyjm6HbvX5nbE5CRw+uOb4zfE7cqkwJtbQa9oK6q8n6SeUNoZM/BJCfPe9TiEZ2s69f
q7A87kKLtgrdpz1fjRQei+h0volYqFmbVrF/i1L7k+uh0TdGmkWAZ4Rs5h9LcTKBsmnFyiXPOppz
D4dj8+SzsLqrXIrRSsg57OCVN5K7H4nuAAu3tYzqH9Z0htRE/V7bl544SQRK386uNNqDLuv97ffU
8IxjwHowBeXxuaK/E0JX6oSaJDm2qQHcR3pibQMEFc9iR2bGsqrROvAxb1hg7xhoSAnhdTcgCV+p
eqoB98ujnzycFEpEPGFvYJYLA59V0Yh5RoAdWSB+YJRxLCmb+cmlkF3fTpILlkSs5tzI2DoIvp2t
1q2fNRgf1oFGlwARoEi1kexrEmAP9ukPBhowl2zgW1GJ99qvP02dAoftvku/P1anGMgghObpsJnQ
2uMIPpB0IRFR/C7AYR276v7WYDNN9uDJpkACQrJ3F6LsKH4Nx/QWglpBGZVoQLvJGV/gPjEHjk6H
gd6s1OiKduih29UTQHDcNOzx3VgusZ8eCcau6pg15c20kK1yUc8H9he5xC1IAXg+vfpLAEFdCelp
/7yBwoRTRJecK2Mk1iuMirPxO+FVUKvALLe4w3ti1oHSmnMD17RRRSNowiMIxv4ty2Fblsc8O5Sw
N4qG5CLeZDZ7m5UvTqBaXLw9YEghFQPStIEdldS50uiLcKCBHhB+bczGSUIYLbpFS6/BzyaTuScl
WX2O5RZm4Js08bfmTNvi21ySHKTeWJVnLTMzVo+YEa7TXq/YGR22I4kP5/mrKLIDDahPigI0/014
woeuonllKaL2cPSpJkSr43ak7TSnaUX9ZeiXf7q0DgbXEMMNdKXySOCU8qCg0dj3BGc5ZKtpREPk
sUtLU8fw5RqaCoE6VI80IJKEsSua9oiskbB7/8Kz7yrmJqdnZoe60DmHE3fldk6R29u/+9fOCCha
A+3B+h1LM2ddAaI5JTiZdbSwYjWdoQvwdI+nAvgTB/Lgp5tyCy1cxawbpZ6gfdW7pEWi9FqxsCt6
/D5JMNVrx8/ickHX/KkdJixOA2N/VS1SgstsqfNJ2TKpsx6vKN9duKZ5QpxVo0RCCeUolisYvOMn
kd7bRXiEr++X+TcJZkwUYEfTifQcCvQuhpqtQkvddH3mjTrHoQzHtyIi1nbhk+vEUOyjy75E7/IR
6/7Ashf+1/pC4ogaQAE8A+NEJ22zA3X7Il4yZ+4ZAMFNR7rhvPnsX5XJTi3gNbvVC8H/mw0QG+RX
/mOXHq5HZMEb2Sthl9MCsoyx+VHFCXvcowAO59dEn+6Z210w+yhJ41ePTvVsmTElJ1PzOzG/OJ5b
KNwT/B+BJdUXlDaaWCwnJ3vUrY46FJaOLwFCbGe3H62yIRkuDKGWxFqQdCtQDhdryJOJVyHsUKb+
88kdrXSnaJRqZ2cibJpd+JX+XO5TuKLxXxnRbXjcjcpjZxnsKjTRsqzlQmyvriotDoKH68KE7DIW
VH/G9LtQumbuKWtNQ9y5rS6K5ADNWHhYAtApTMNrkiq/hU+nHCrZo6yG5+i58KL+jZiZb3j5HyGB
5M5PhktXE+4JAAmx8nuznyE0RdiIpjItFmfbSibWtO+F4l+9vO3dfVlYxX8S4HT9n7ZqxS06O87h
nm7L32CZ0zA2wezSPVmGwKJM0mwlEogxxLYR8Q6PLiUcjepMyY0DnYH/VHOVJX8XYNLnH/2jsdYd
/lqEfHtILb8WLz+qQ6vZwbKgK1QkualhjJfXY9X5mkPO+R0iV+T1oV5pOtIzPXmPugn6PEnPXu5a
qqKW7QpjsengfhpTy0qqtjJkimzkGO2/7OjfeJjZ+nTBkTMdmQW51mS2t0N6T+NNwXwB0hl3iWi3
WqZD32guC5h0bLWxI/QONqcBwmI1XGRMAgfRtQ6UF9p92wWhQkPJKYLUZFn6AvVwvDRmk/KJfgOR
+DBYbGkfdmAXZ7l8TX75o92Vgqwgwpf+7HjWRnn3yYhbHopg8hgasstoO1E8mOOoz//nlXuxDNjK
dKxmme20wKGhr7L+dPjc36jEvmlBY674vtcFV4Jk/U+44MyO+pbh7XOtui/voFSemVEoJW10XSJu
rfMIfOn5XLWOeK0WpkHOLw3/cGl8HYHk02c9IkWOK+8sLwA96Ch0wTlNc/sV5u6ZdcurF/Yb3Jfl
XPEXwaBrUg0WrveHAo7zNDNWpRk/IuzRAE6F47kvZ+nZZ853fEwOvCwCjdW54Dcxa8zwmKsF8iF/
qfY5gG5K2DBERJXsakkTFE2aNdnxc23IxZ6oBKVnjlIrzGC8Rly0+ViRuyJBNkNSv5mB1R+/hT2l
eIm4U0T/Svcs7FHEEK5MaOnM/QsPRbat6DDRw5vphCBHL3aOKTYhAfjAoAdIcgBQKkhOGk4rW06Q
kJkzQr6Un9MdoDrOoEMGYTkzzf9iGClQlYZZlrGuuFT0mhO1UPcd7/MnjOWTssTgJDSoWM1tiGbq
AIba5Z3zfkb1IkwyM972Y5KzwTp5jIr9kPw4veJwNQpYTOkpjoK7tUK4bXO5OFlLXxbkN1of4zXq
UQnACoNPa41f1goMNcqZXQeOx4YuVCRNw4bep3HwX1EAkIgCNOMUyVSe1UT96einhvE2FS46CgYB
MMu9GwUsIHjL8GJAi6C+2WGkoymiOm54QwbEEN5+8xmsHNGRC1z31ravI4BWyFIB6ihm9BzGUtn6
kmXyN5ET6pl795x4bMkjkwHJpBVmmKVmfmhmuAZ2ytlMVjG9vknaM5/F/GZzYmbGDi4mn4CmZU/f
Z/r7CKN6oIeFD3ngfLGFDfChBC45qLbAY4YW4kLscZBVH2KP2TgAOXGoCGbPKbEM1CVR4duuVEA5
qAMeWt1LWWS8ofpGCPfVq8IUSYaBxE/l7qOSfMyVvc2SK38GPEOKHRqf1GSwGUhFMUxFyZu6QVjh
g3QN9TKYHsIg9e8vc0YQxee6ZybOOXBXcVgUov3FBi5LyM55AaSzG+wHtAjLrqiu77IiBcYbn5/T
5OoE+rAxetJ2QukG89Iu9Jf0QVyqJJIM4+UkTxVnpcx4jBHI4GbQlWAoOS5eWxdd1hudE6yfdQdO
YSTLu+VbuinhvhIKM4aHSvV0orLO79e+S26EoDVSVcI7Fjjhm+nYVKBhFxTRgsQm18f00SUk7jX5
nuCreLnrmP4DZ3VimePeRmfreCSOEy7brmaGMTKB3DB4otf9ZuoulIlhgsBOs2SUyVWEKsKdmCNv
iWCPEspRF09hHJJyd9X7oSTCzNeuMCpuk+KnZMmVStyL7lWzLUO2z44A7GIw/n1csfuk/A9Mo7OI
JD8XDOwytt+7SZK5JDedag7U0RcKUkYk8DQvOD+U0BitMesQWnHIYP+74Sh6ykkz/HT47iwTqLlc
aRuhAEYRioKwbUDKnCWrciuJBI/pw1uuFAQfx8s66d6x6fpdoLQ85BfSob3EmWvhxK2If1XIufTB
EekAxMaQQ3iFOH5u+MYjlvP3oH6GPAwRACAsI+VR0xtpLrQBc/beDeeKd+gxcDXbQJ4ObcliZiKY
6KU+7MwCbhSLs2GdMoU/ibykZb+IDL+6RqtcWaoVul+AXhgdeNmAUibuVIwfdEz3fAZUKzvzI6J7
b/ADUVNugsx9dbGjXi0LuDbKrZQIWVZ5bOZJQfLCeKZlnDkxi+YmyqmIKR2ANSHT/aZvoMsFeoc2
UFRUGPn+65SDtQddTg6D721Im5VWymqBNFKdwSYaWp6PtFPw/oi8NySFRHi8XL+O0NM5EtYszCcG
KWo1KLtwN3Umv6vIox71muiiDS5vFUi0X+MWw0Fd1NDCzFODs+30YXcKY9SsBDKuhehMgSGL4cim
wxqZ5j/r3So+2YI9e87uomIq7JduvhP1Qglh5VcWWDpL/kLcXanjDFb/LiH7dOz7Pb41nGPsaB+1
RoaVZ1lDFfIAgiymUh6N/IeHOqRoSBGkL1QQdb14Hr2iraPDCLIxw0xufUgHN9H116WPMKM9MYLl
3M8zb6EQb0nPcHEkdIq6yAvz4utdR/s4pTRTnPW/6Mvd2epRog9CH7k7DUStl5IsesbOvBM4E2Oa
4GHyYh+XhpOMqYMXyMGMUnkmFye4TndZQzRI+Jkn5H+GXN+MblxpHPNIr/DpwHiyqmmn3SvoGGTy
Araw9RyYCe7drZ4Pg7HgzquxALBRXTy0JOD02mNFjLqoDu7VkJED+RHyGPMY5pB+V6Bp1+tOdYxM
LKFf8gZDxlYlN4fkD1SUMF6LTzIQ+Sde//DYqN1c+keDUFzC4x+8EbAECRw6xqjNaGTDMjjrr6RF
FaS6e2XhZEI5n7pa+A26BYZ+4//QsdY+0cKingLYnLNyuUZA9UVsFEHCICOl9ogtrITMj0174A7S
AbRrWpYuDVJKPeqaVrunM0LDG8x2oCQ6/edtyncB1Heu+u61ctC3Y+Yz/JfB7DodXEVobCiCx3Gv
LojDlJCnxXMhDCZa5Sf/wArWl/nSvr7jUHBtqLdLjTjVIYLfPW/lGXvMJX6NZ97d4OzUVmPZmpJ3
YYskjoBeV3ERX4bVn/9x+yWjZDFtEJGoc09XanpyXAfKdbfxU+ocDIwWV0d9mXSsPUSJdEtXAR+V
808/L5W9T5h/7Z+MMG5xyS9ecRfIIg42K2KMFCRpquknEpZnNNux5V/jx1fisOiguYFaZcJYFxQL
WU7n6EXwAyA3/4sQgrVpEIuCXyz0mcFKf1IA4AelXAfmBKZIx+9ujA+gA3Apssqa68ugg0pGCdbe
bcAG2mGX2F2UU+gp76VheaDqFFJW3by5KVEve6m5p/NuX1mwf5bgWDPsjfxiOokiGs6w2hqE2jro
+hbKG8fpT33lSyuk8CPdn0vDa5qt+uwnDBa276HQ1ZUNMvfOnEnq4jQ+MEaN9c/vHWFXz3kXP26V
IqRIOSQ4wfurzqIhqFT2csStrSopKZiQdJq+IP7dUEsEQDG3riuGcmhF4p8+u/OkFtt3QFozHz3j
5k47klBD3Etzw9/YzQZDlQJg/A89gE1uc/1W9e3JKE4R+RCEq/kPCoiOaG4yc/QO8nzdKr6xy4ZG
l7etZqb9fONDLgLiUa5oXn0Vd8TrxtNRuoXCjzqKzLFgj+JarvEVhzILKcpznCAEEZmwuKuAEx3a
fKGndCsbodLzYm/9o58CWgYXvvBH3Pre8ZRAE5QBKeg8Z7HP/H8CEg2iaZ89sU4dmic7qAar0n0q
Bpq0WSRsMYYtrxrsn7BiIBosuU3mOk871nFXIqoOZtbuAfUGbPt9DjhjaKmOhGuYHSS4KNs/npWF
SYQ830Dfb4U532bI+oxmS0rROeQWHXCgp7IY8F5j55niXbtI06W7oP9CZ0/daursvMtBGV4g2tWx
KNUFd/BkDNhTLgL7vWiuvgETTGfqeLziyzEGArEXGPxxc18aL1QRPZXJwa7dKYQYGBIvpYZqXuYJ
0K2QcLrSrT1r4Q8qtEuq24/KS4I1zM7iWNJnMtOeq+Z3W/yq9N96QCB3QxOuuBA78H5P8mIlyLy/
Cirqu3kBeuLvnRdOMN1mXwRZqPQEdRZNhcFBdCwe5uwVyjwoYbflcLjwB+Vx48Et5en2MtumheUd
EUnkf40BLwakUpqwFpeWLcxzx9YOEuKi5TRgkwGt8IZdR6QtnIEnZf/SYsiNT4SRtquVOedN+GeM
BvqaKNMrNV/6ymL2m+KKaQYBzJ/bJkWmI1n+/lO7j50B/UrnCECMpD3IPCcwp+sBYDYLTO9Hbqkr
otfG+ECDIal80nOsaKikm/DkYlfhwwNDPrz91m7F1nFVWO6OKvaF1XUzjX3KwgA2+qiVO4T9KYjx
zn1ObNVIpNdg+joGbr5ICAe4oIcXNJNgTLhbO42wnrincXHBtApeOF2aHF7buIe8H0IEMnJWfyXz
Pjhd9LgjyK0ULDy2SUGk55wEGuIbHoVG85lLnJz4Yyg1osbgUFcHfZjrpKN58tbRZbvwKWMpv/ct
FIalmzN8qsZ7/YsTOyfLx0oV51xDGj4H5bm5vmZ3egiX05hAKaqD9hdJ3FPDinrLpiwEljlxZXYe
nnkIr4aDJXfIZy86GJfQ0Nos5cRmdgKEPuftx0XB3zRV+24MkclgZnyDg66wLSakNrzd2CStl4D5
i0cSZwsEtuG6d6wRBGqvr0kvsHHJBNWV2UVCs8r4R7PDEN7TcOzJxxGEN80Lp++uzq7NNtLACC0P
ZsEmkbClPZJB8QZO4a/8lEtKmr0nlNqaApUaYF5xe0IMELX0F8subXHFiV5fyC3Svqyb0Z1X6Jal
ObPhgYt/dgxU83H+mJH8j4zKrPYezWSuNzI34BRskv3ea14zRrVAhfowDc4sVxEIy7NdvnMfJ2NA
+Vc2KIKE6WWVLWTbWohuTaeM+DcCbF/5eHeWai83YsCSqdieUxI6W+0+H7HfM25bWYf3PKaE9sZ7
6Q5gvcLkJ7znXRTYW6kgTgBIQxSEUI8SSLo5TB98tguGkORsy41zMpmxnGpJcD69087NQg8kRNkL
TXuGNEreveJ+Z2uSlSp0XwlXAcBtEOn5kZdDKi5+Zg4MgFTywYNsIUVlVLMALgVl+J1+OiR63nDR
oHdJBi/KSMX1r/cN4+E/3AL0hE9Hq3HrxfswVj2cTeUfQU9F9mW9spgXGZMfZTjhGMHlhxqEi5K7
br4HvwhQZY3bOHMhHTu5hj1kocTEllwh/IOWQjL56nKOGGa8ZJMY7alOsfbnWmlaHHdLftH+5glA
cg16q6dY/Y/wDg4ZEutBnV+2GlGA/nAniqKgmhWuTWsdRJ8zi+nUwq3KNgWaF0/GsH2wCpzjt1YW
l9ZzPhcX3wi+TrMr0q1pcwRPiQREla6k6lfFQ6fHTuU92luWAAOwIrorpL++xXR+k51muSrh2L17
3vdV64jZPRO0DqCfywEBtbDm7A6UqYGZYrS/1dP24e8ztAbWJJjUx6FK+LfJ2xKUZB+PCg3T5TBR
lV2YFgOCtYtaRsrfsrBjV2oqEYUWS8U+uW8p8b8X/6T9JuGU7a4xaEaZ4phBDDWi41J568gBml1C
irtKP02VUpoNhI7YxvLtqo4uHzi/ynGfDLLzexxX2zkUUGurIFiTasg6nW+LELK+wRBEpioxTAMf
c6f2cmSQ0jrXl8BldsYmqoFU7FxcW1DCXYgOyuslCX/ae2PiTsO87lfijZJv5ZG9Mc1R7iiOi4xh
j5CndLikj5Uxj5j5glOtgPjOrDGYi7gbJhkbo6mLn1MIDOklDZ7QJYh/t16TErtwmirNbIlKmDCY
XhfEnjrPK4NT6YwJg0KdutFEgatI8Xuy5CEsxrD/Yomwl9RDXprzarlg4/hexVFrv434KpwUVI47
I2xHLaze/80Q8zmTuwht+IbFFscxHvjLvPx6bE4E0kzGcNbDb1yB3qPA8ZZrmFmxeVlrmaD8KSwl
hl2VJDCwf5yx6q5Rrsq6v5fKCuVj3xyclCJ9dWTxWy9s6a0U/Ujy57FHioqTJq3l/Ui+RXSXwJaH
254xraV9A5zq0ee21ciUJ5xGDmdkrHSbZhiMfTzAo+W2EQL4YssJtdB6vVYV9I6ik8k4t+VZgHH4
eksHaKxebhBwdfAuu4qoiah0HLYf1ekucc9ZoPWGr/hAQD3cmxuwMxFv3gaZaaOkPedCMFZfVywH
o08CyUyB68/8APSxDiwh2f0zdL/N5c4V+cXo/XCUTp3P+HlBggJnFq1SJfYcngimjwvfVVn7M7TP
RUhh7TN3DrhO4pgLv17WG8RejdcsxfClGPFe9n1k7o8LO8Os0Y7VpyGgESTYyB73J1WGxEZB4dWH
2TxG5OAacJ/uzt6kFY15VcD4H9/dX7tWgQlFAvgXXjfnRLF2K0SXm/w2dKIrkAQ/ovTw5YAOVsSL
IxOFrNPX+stRsZjDWPlBaWwIpUUHzpnGGIGmpmXfK6rrvwkrhP2SL462D39/+URCV9mf7i4A36sV
IrirkVsht/vR8M0jCrHdbaNFqsEYhkqqlzI+7PnpnCJlJXAIw/qECNEHEzL/bpx810EVEGiAD3yj
3Sf2E2vICOfeUAybpn/zsG6Yj202DS6XffjcKEn4Cb8gVjt2ZQs2scPuK5sFqbgoQQVM3HN/cpXP
8jr02kDRRy9aofygMW0yi7TA/pF7P0hDsIeCxURe9vYQ2bVgeCRlDHli9XV94KUT7YfSQPPgT2un
dpcY2OKxmJs8Peg4+gxEfjzpFYjr/jz9e5sb6jZpTPjqTMro84CVfjUAzfbyjQ9IcuAQbeQuBOB+
f1PGv8aQbFbqmCIvGgq1UFp+3h4C0dgIWaO1ZtAwwaBQIprhnF7bsXs8M0EggGiVQA7HpZSHnu0J
JO3ggUmV4G6xiCdVj+q9IElzNqLkDP87orLdwVuKY7yNBrM+Te2Cl1+QMWn5igoxxHE+zD01Zwg0
0l10FQ/MN+0XJ87NCEfFSZSeprsn7JZJDmv+vnLxMWLQrDwwhT7QcjQOy3dXKYRdOfDSDlPRTROP
XXONDuYdfB2G8pJzoxnzBjVfDYSDu5inPTf+JmT7b5DnPnWKbeCTvtgfxeVUFHbHAgnIYqmMCknr
lZtgBsi27LWZ2Eyx6hYJGpS1WleJWivl51A8CNVfB0AZL18aFN9AgORbU5t4Rs9mykKdRQ98LN0u
bsyojak8PrxU++VPXsEZ6g3GZCbYhOLt44mUKvkQs0q295VJKjrJH9s+l7Tu+LZYqsi131HxgFRX
4mPQSWrlhrwr+VU1EuI7U9YcNwl+avPm6s6WmY1juygTYciUsoJOZmvwR0glY32EcwgQ0eIz+by1
LnVVw5Qs/ekC4fidnTcHmboYVTVsU4OCqw+8CPvhOj0I2D0yF+qjAX4zWJDtAIcO78ShreE+Xg+e
9ra7O9SAhSrCAptitotp4d7oe5j4LUwyip7fgIkVuxS+RNqF1Ez4AvEKNmFXyuPtoqHY4JXVfqyg
SjI6IOXBBNsqtIx9ROUOKV6hWVCs8Cn8r/UTN2HZis9Oe2bpF8tfO4zMblcrfFAp77LJRkplZYhX
Y0Mp9Ak03KhsbK5lXoo4qfkwr2pMMB7uxwahmrQfwCDD+wjQfICMZUH4ridsitqrKC/PDf07F5t3
ZRE8btsRR+GZ2sByy4V3x/+qV16FyjscSLlbrY8kg4IhWLMZREscwMOzhinYuHPHHGtHEwwEDtgW
/Yg6BIq0HIgg8nEz34CgHqP8DhEg47M7k45sQuk34XrvkOkGL7dk5yx9m92mbwlN2elJx8E8E1dW
SqsOlcVrWQbbxS4uBbgoK1fiEJzB0kjfANwT8NTxTrGnXWIttc7D0olhrd4dvrOJ/g1jymsGJa/0
uvS6Q0dFJJ5ShlvJ8TtiIbI8CyZzv06cq9VL5TZWs5mejBSHGBcLO5VbsmTZU8auVnhuiAUb+wdr
Al+KZjGZHG0DQxACZc04TgyBftRByFWmCbUaziDvXRDyQ/DJZxVdV+56vHw16AuocVcEaIrNxivf
bozUZXrpeBHRG/79WQa38HYlQ0egylX7x7OMaqVkFswQtB061fEwC+DZdddFB/WmquN1e7W7V+gd
4cEKZ5SvFYD1A9kWzo9ltaBscoPBprEbCWBcFnm71usqVQCQfgtQEt/P4K5ZlP6hOVB6emct0RE2
3oWDztA2FTZwGYDgxKqXPdMPP8WwIywzdYyH0VJ8GF/3t4d2PqFJ+R+PMxC+s18AjsxATd0RUVkI
HW1QYq1b04y++c57rD7UUU+hWj/UxIasGDmjJlf95vIQcflNPzXMDVmh41ihe+D9xGEqb5uP2hwX
pHYJPF0zwdNmjX9VqhBm5DsUly4j2fKhxCrWMiRT3OuFiNYq6ayWQWHIUmXnWo5f/J/cy6i/1ESG
THsJmrEPzAsPkz4xShGEJZ3n3oGBmfx5VNPph9K9yIveE1DiNI2DuVMuDSWZuXbbwcGT8i5xNA0W
SQlWkyyZjThXNfcDiLeu+LCNKXNvkxqdSL82dpyU/aZ8S0dwqX4Pk7hdHC/nN3UWQwX+qRV0chvS
b2EbUzL/XZDTtPlyNTDjTHj4U5arRkn9u0iX0dJO/oHAhhDMgj1ugiwnd+GVR7V6nmMwyWwTDTvl
mrmE/LmrUEetT9p5IBuvCN79NUiJ0/vG3MzFc30j+1+R29zQ/zx8Wo8HEq+oCQlVYJgh09/OH8oX
wrEERxMWP02kZHCra8Gr0S8vfE1reEaHve1VfoDW0jvT/iMre7Pd/ACNpHj45y2RQ7u3tAsocCNl
Lk6GlbrgWUbe1M//wrMG44x2SDrOVquoWRzniMG5MrJZgryZ7ns0JG3r7/8SAvaj2XgINhmU0ygU
5zBtwKPdlIxVyYNt0tB7XRVjkM94OgfCwW+j0JUIUNrXQwMPbqOCISBqDyyUcj+W1L33Mzt5Zt7d
9cK3ID8puEjXDize53nFYJPCNpeWzxw61Qrsejg8sY2yg8dJ0XJGYjfEtX67Rax9nSul8e+D7Lim
gaU1EZB5+5YJhS7Qez6b6CHK94UilJsbQX8Qh49K5eGTRr/hm8vf1LFFFaC9INInuGX39+InMgWs
6tnA9FA2JqurhorbMyWd+ISQr3Ruy415voRe85Is7GLk40SYB1x1qPLi9qJpcOCeXhjMQkisF2Ej
gXmnbZcupiesdxFutj4bmTeX6HQS4emsCdIFG5G0Oa1w35JIA6ytLGQfzVS1XngTmKh6qzh0lx0a
V1auanBByf9MKc66NYi6AkU8Ji8ive4ldsEnjbxtMA2zvO2+AcAF4xu+daI//sWgKeEjX3smDQqr
wW0cvZH80SveP122KYvG8AISxytUrhc8Zt8x+A2sDOchZsCQtU0WhF/z4QVT5p+e8bn2MHeTP8jB
PLclqT2iYdcAjWcDr1lAD6LjX94F6U28KwC0R7MKu7vfUuOdenX5xIS5v5kumV4YTHqInauWEqyv
bjeDonvhMzi5uxNxynidFQvSr6HxxUBuvUwwmoqoqgEswPQGZ+lp+HXXFTUfPh/bmqbaaFBJwUCP
X/262QpQg7jMY0bleAS7ph3wRy8HJk+kNe9rkXTviYpKkEIMIm2SYvv8XYrWavJ8zvG94A8/wLE9
8Ey0XsgAVDJ267xT2f6R4QIRSmKtCryizdyPjMyDMXEuX1AXbMqT0M1PDqJQdOjJVEsQK9+Zx4K7
2N24L4cGnIvxuvEaNjtFR6RmGSHfdMUaQAO9mkdJkUWvThchjsRpxcyhK8ykpe3Wy94/KD0MI5V/
cek84rbCL0plny/PAJZTb5MKoO4DcZMtPnsV58KqH+5CQHn3MveS4CiKG1oRrh47pDonAgfzZvnu
XEbOoPFKlXEOdAL+c806TGRJmWSu6BJx3m/I75zV4AVquie4JdmGy5Qw0p3CwBhqvOKTKTV6jzma
6nDwo4kg4WU65+LpK1QLBEzPZgw6+c5yFaxDjY7y4+chYZJEMmgNh192tpxdf436QPoBb1fEPCBK
laBLc1tUGY3qSYOz6UC6Y0C3UEFVIJrGWwxCteV1n2dJ9Arq4bVzoNZjmphrVcPHa+6509c6iorI
pzlS2CnaQK2qKywuTPfQPu10UGTPxM0/4jfjQgV1QdqsdWW32TON0druxoQp1eyk94kFgBQH75qG
rrTy7QO+LbHHLQefVQsT1lZOc51ykSPSZO3rkuacjdD3GqRYgamp3yj7LD0NNI0kVv4ptPDwmVwk
QTTrR4YQxLe1I+oSg75QLgJ5NEx3KFNoqdPBaKFlKM5sSxR+d2Xy4uoo4B/8wK89hGUOIPs5DGDM
0DPboR36NWu6OfJWzfg/r8uFbxpnyTmdoIGGzsJYDDR1qlCBWvRJuKvarVuK9rwX+NT/sDj2+Eum
mMMoA3ocJAkxwfUGgWFC8KS7+IilPhzNodiBT7/iPW7B9OjlFaiPqyJ/7HsJ6gb3xmUNVaxwvDqV
qCaKOrE4tqIn1ti3JtxWN4pRH15sp0z70TzmD8NiWy8ffiWKUY/h3QpjLYOzKu3BS+W+ccAY2Lf3
fP4X4G9moTH1aDmdSfh2GZPGkJfvvAqTei34G4Zx3sAUI81/wFhpZUblBdSLo36KasZkBcRceGZY
oyD93YVDebwqMpQ8vcXeCMQoAqZvF/6ntY+1y0bNm9XEZXd4azmZ2ZWjybHrsByC4EQzBVyzx4xy
masoUd1VoLeIq7RfVSTf3F8EOEEqYEpRdLDDKQtQOcIULIpn5Rg5+eftjyRxJgDvxTdd1fn/ISyV
Eabp9q7rCV63wRIhREQo7l+WD6PZ4XxFz7ph4YGLeCOAOLRBjbk3hND3VmV7sxpYGRReqmUOts1/
VCGMMyUZMW2mn9S/vfz4R5VWA7d0VUzc1d29/WUMCCyN4ndnHWFVmVJfBmMFFNUi9wcS00KGQ3VR
IaIKHTIHqWzeBGWfaWAhmX4XnkP3NvGBezZ9XUFPZAf9dS6Acua42rB8u3fEQVtTsfaT/hwAKeeO
lvnUT0slZGfWJjfuIeps/uiF1hDDpKuULl5vy/lAEx2Q5XOuxeLUopY2jjH3SBP7fML22K/PP5BU
yEt82Ng2cUVEVRaIC0Kv1gc4LcJWkWIl2nGm/PXyMm0IoALwsgr+Uc5OuWIG54gnXae6jQ/7Q4mB
0+KYiQ77+7BeRcdNSV+oJg3ZFlKWhczxr+ScPy081kkZORFXbv8BvUmVbSJsfviR/z5929E7kQJf
cLZ5H+UbJebt+hHF/hx2FOGFtAtaU6HpkrFEBKrHgHZ1UJ3o51HMg6LcFMf+i/0+uE2hv9YDJ1f6
ZpEg4wOuasnTOfBWaSbnc4ONtMJCTVVCytT5gmqwbIpFkTetzlRJRdUUAGiME758rX0aTkKFF7n+
IHQEvqLx8AyvsUPiAO16aOHVSRM2prDOy9KKLMyL8V9MsLw0iUU4xBwfQC4uuxifGDpO8KtFSA5y
1o3RQ6gixc0lOHwBA9a702H7zTj8YA09po6z35ds4QrcKbuhAhOS8bHNK+yE1sXmUrNQ5pdvLEoN
ERxAjxpld3i70ppw851U6io5claBWYwhFy2M6EuUi6U0ewdFUkZDLPKpgWzdc5alPtre97A6kY2Z
T5xZlLxBfTxXJj3qO14mU/fm2zpW7wPu7eBfp0EUuKYdQaJBpoY+awD56KiQPCPoaLrt1FBcvGNP
ezrZyK4Ope8EhVdN/EDHryAkVxNU7nJckUyfi6QObqafwUpic7Dg+NiO91mYp+kbAqIxyS4E0JQu
5ZyLx4gKGMtoZxAALGRh35u/45XPUCAi/ABMxiNOWkVl6fcrcHMEbtPz6w/jZAKxbyPLo9XPM8xY
8+FSrbpeV3aRJGTw9F4qOXzlMWoBiCEBjmLBdPx72PENAFfFZOr8ms1Z5g9zzH7en9cEh+Y0accO
PxO7JTkio5qIa9ZjJF7oYnLoBM+25fDY81GZxQPr1p+6w7kI8VeI7bEUvWMInhuT04POVhJdV656
H+gUn/ePnye8/RChwzJ2GNvPFbBfAv8ccC6QNKxPPrN9mMGg77D9kwJIwcGTbaQXWkF1IXBa/8wC
lZrqzF2IfofgjfjaC6eGueSeZsQjOX9RwVoDoPGR2Ub49L3DQGvwnFk0/ddC6MVFlW1UoW5ZcGqe
6yljEm130LS0k6gnT5SgXmiprYwDZqZ0MA4ptuyzbOkudzJX6RokUniiOkfBjUQRZDTprh6GxSY9
/NbTTNl3wx8C177Fk8MiBew+zcO8RjejrhAjH57VVbM6i+WZjGfKts+uxJ2A+evhiLok+8JtLws+
uW1dzRYcyrpYUp7MU23l8uOZ2ihEyKKqI8auesVZSaOcR9y3g6LXbuSLfMzAt8S+BcsjALfRrPhf
CYJPp5xL15/xJji/ZPs2KWty7R8WGeiI8JloxmPUrQX5lNpbBWWxliwPFEO51P2xpzII394LeYt8
Z/B0dKyQ1c8JosUoRtNYnael7E4pBAux5GzT9CfS4s8EufRYjfoRexf6FOqipDn/asOTC7hZppcZ
MxZFQ+nnxDFaX1PhD1aosQhHyewqeSlGcZhuqM+IoAzzemTI01KMCMHGN8a5YEUkHrH1mdde6Rwg
Mm5YSitdMuJixIpO3L/BZeqBg24s2+N93wUZO5bmwdAKFdu29ZBtqEoDKjQNus6fq1X1a4rYehfT
bZtpuZwnKfMCxTIhNjUs2BpNDnzeZFi7ERZDPjkLgdGtQpkMIi/sDaoS/T9c3ho1yZ9eeu+aDF/K
nnFDV4TCNnXN1rlFUpxr6j/8/wFvrYysksTq9F1pX+PZQGhIgGd2V3UbAA3w8WlArrtG9Dzh6Qmq
AJE40Py/HDXVz17TZIqcjFEKsweB618yiPcQTfaAi9H9XN9I40Uh0VKmj3QHBCPROXgmR+bzUhU2
I8NaQ4FM5HkRXx6C45IRXw2ALip+Wb1nlbJxSBr3eyzS4I5kw0KLe50Q2Lzi+4wsi8lUoNDokjQo
G2PGcDAe4e9LEqxQcemzi1c5YCyfB6VGz43/HuTU3vJc80By5svWszFmC/dRjKjNHbe5kGSaSuxX
Q3bktaWLrHzPi6WNLk3uomIL1siWcO06q0rtYFdtllfJlMn/5UaarkU7Bv3cHhJejq1OejoSWaBI
fz6Keyv34RY5TO61POWP2oZtYcPsIafEv54NDcRbyq7ztgJF/kmaY1Jal32Zc5fpEh6mkSae5A4c
7zLWgy2Y3IR7QBtvgttwl7gvyJCGstyBd/D/c4SbD65JJObEu48E4CH4UeJMeu3Z+DbcaJd1OrT/
C1tCXVGrOI9N4WtUAEF8+ShXv2ghyufqOiRY9wRs20iTd8bgO3OZeZjggweTwMt7MvtXy5UUPtOu
7EmXUUTn35Hi9gaOYVBWEgunJaJQFYTSIUZJuW/gdLS/QJSMNne3PkL2zMKqnCyZ1Cnzk08z6/A/
NcdYpefWXUVlS1D9IK0OEfupLCftHzIv1I5V1DdSSFz/basNRtxbl8bmJPN5vSniOokd2NGFsD9A
GTBx4ll2vsbdZ8YQNTacV0z1Gtr8K/aHOQ5QqjNIJK/bHF8weMCAz0ur3DRW/Kyqv3HNNSgbqMl4
LybFDRwVPxvxh/O7/3trfUsqIP/0QajRBWOnbmYbUAX5ydSP+7U/nwpt7AUdVHJm6yrnmwhGyIw4
yWLc6yXOTi3s7zhcZParJFUEhgzf5EgWkfRn8zdPjY/okxCz+y/lUyGWQIfHhJUcsHtTLpTr4BLR
wS8KFi3QQqM6lSjesr19luceTramz28L8VFpcQ21MnqKHoiQD+78krIgHB9f4D9TbcOvhAbnhY28
DrN9QEUFYQsVUaBRMGbStVK+s6zaMMdXhmO9IclPh+z2PDAgTR484U6c5/mkHEdRXNzXiL36EEfl
izZvxjzoAcBrR0bS0BuKS3BApkU3lWVfgvsaHX3hHX3d/3BPz9eKkB2CWr43R1UVLkFygyE7z8j5
j6t+tnv/YR9X0wDbA+B8AqJyNvoo2/4UddqViSxXJpo6zc/9nRFzqS8u1RudLlNlSQ01Blqbqcfm
/t2vtkKfBJ/WCWysb4LA4zypuQZ7jTRuBaX3jW7JU30qgmiDoucXRqYySrFqaBC6vYnNYv0A0MOC
j9CqEWD+uo4DQVbNvn5IcqOxCeOnqTmNdxadnGaXqW1ljSugswOSGXguC4Riw2taHR0Y/Y9pvs1W
YMlO/aPf8sOwYpyetFGroVQk9RchvCK2SeaJ+KALQysTanzkMNXYkU80hgARds4MJhDNqsbAsTW8
SsHaTiyQAlxlA7+fyip9fcsTazmJRHJAmR+lFGtfyPOzpfrxkdopqQNoBty6DvuaZIOkpFQjsh7S
iSsz5Hy8/RSFqx/jiQHxh4GYTKjVPyNYeaKFkOd6Yjjr4m0vwrwqoQbqn+dgwm1VIQgDsH10NMxU
luehqeyn4VxgU4AGBzJohkQE9EYAdnku/gw2gbNDjBOeYFJ/OFC0a09j3vvPxkzWm3ojWzJeS7PN
M7Brl0YiTCtj29YqPt/4pE4uxDW6TSHgyujz81kvt29Ee+hzupR3unowuthOCCbA885IvlPKfeOR
tniR4oeaD/TXrcBAtpTUrbNpDJN5b3eIkrv6zBbGaP48K9xB0NFOW4uPLAAhY4qZK6T6xKtg3R+a
mmFmO2Hvd3uHNnuvx4fSxHRSbmbw1ffbktXMiOUlHt2CJ0aa05RZauE/FOwFKF5VoBOJtZRj3O3U
LfrOIPMLEXylNEuzX2FK9Gq3cpyMjRrWZjqq3uBGIPHo8NKq9Xpr/zvhDC+V1cTPKJoGDb5osH14
Ys24AdEm0rWd3SI2DJAnSB14HHVjT8sZqHjggxjAisft7Gb5lb8EvLFsgkHnuEESFPCJY6gqH4nf
x7Too5UR0/QV9cTfOsX8uj1Cl19XOAKK0ZQCIszO0/FI4BI5rcHMgD/I4NIf/QM/w/1WVEp2etBA
wIyEry69WZSkeu2pjHNhIexLY3fwMfa/a9WK/uOUXrqekB/Gyd5VGwNAhjBZC2vZoTIfy7dpocYq
Ftsyg+x3RSKdOlsbXWz4BBAC9CW37ENxwxae7JOBpT220jg29Cd9OZXmqBVUfEBpr3wDwfEUekVx
miBJxOFaBjI0+4YlPlxQmZ0lbIOjG5UrcREGLY+maoI0Hpi8RIv7otCeSUXn5/hc3e4btUoaClvw
eVLNfcY1ukm7cW2eUt7quepiBbMiB5jtbwHkajR7hdTHvEElnD88Ei1dOOUaazWgTKF18ktCrpgS
fDtBuP+0mBl1Kkxu4YSlpMi8iQvMKSrdNgwmHZ+0DJUKTlvlvAe7fKd5R2nBvMCc4yvoc8UEyeK/
9DpTIUkX52lfaMAiKpG9mtAcwTlQLwRZP1ZqYuCewEI/B0QxgElAuGtnsc4A8syW2yaJl85Iu+Ze
PUFauYLsXcqpmPYjKCO3OG0PoPjRTmP7t34H3gDWlY0tszJFAw7LN3tGGfZqAG0ZseBxK7T5LFTJ
FzFHgxcwpL2DcTP3aFdq54OhLOlxXwB8gW+5bRytDQAh7LaZYp2gufK5USJ52CAiMyYPwQ2LkF9E
Ba2/Me+pkCmaj2+TXqbuRXN2dUrE9BT7EDakiFjr8bu7AqJUwZ+WZioewBI2pnNLTyMxTeii8H+r
TeRZ91qIXmQfCusYcx88XDcMjwkChbswx265eKSCo4/l0jT8a6RTlKGzBaqtE3SYcL5XDSBwnBYw
xvuNYqlCAWeur1BLdHJ16ux0HwDYB5MJn/dLs13oMQRZsfyS3k0HWvmhQz20bvoDWnOGGFtUGolj
wqetP2nd/JJWvRymXSqFj82sgiQ8RBiOKr6O8fbm+/izc8GFzJ/ncH3XQrcEf29KuOGj60iqBYp8
k4FfYhBQdW98uKNZaUYronruNoza7tm83fWbBEDP0yJlg6jDy+UJWP+jVZHfKT8ABSEMpTbJIgcF
zqfbtmjSaUE2exJOosPrg9mK1CzrDeyMmvK/33SfYkWgcUmIRqHXTdcPKMpv22r4PFxe8WyYcdaS
wfPLltGMMj6KmLdaAFoZsDp8FsmmOsAukraf6lzcE9Oz9QfgQBCFuGsc+mkGEwjhtdQ/fjCtv9ON
q2PhUqk49MznjFvhjX2IEs31cKx7kr9NPeRZQ6yH73ev6jOhIIvWGgg5R0BYW0FsxvJ06IyD0/AZ
dFHMoCy5iBf8dpK4StNpd34EVGtAmOw1zi0gaJhWc+SGMu1JyGIB4ZzwkrrI0vlQvEQ/+W9xhakG
g93ktlDB/pLnpkderp5z5/GAj2ZcLgQr2rbfS3qhtXVpv92TV89E7ZZ58L/oFlzXTHrBb2TyYZCf
hE9So1hadpraxbq5jK7ty2m2SQDT1yIK+RzWwo5H85LLbtS+zbtUBJ1JX6PbLNrjvTru1GPbD8kQ
ILaD9eEfZ3fo/0ib7b5ExjRpGUXisie+DFbO6AIZgTkBHMTpxZSMQQg6hMvTtIN6alJddaZK47Wi
6yiCZc+VIPiC9MDEYQJI3ULwrZ4kcE7rDEcyY6BwAalMpdxTV/iEpUuF+F+jHr0y6VwuhgiNk9wO
sJ1/HK0rCvr0sU2DcjTnQTy5KflzKVUXzoeBIjvcqg7x+x9G+wL0SnBZbAMgD2Z0PZCqib27Law5
cE3pjrA8j82sCP86ZbwGL6uvPf7oOn7H6/hvum3VNK36u9UUwJWc50k3h+9Bj6LdPNcgaQS4cb11
fX1fuSJZbakOhu8juG8Vkr2+uKpuZlWe+YCYxUxvjiLi68ec1c8yhCjIXSlZKW4tZFcwdEa1BXr5
UDngfCpTxNiywW99U2N+cMqRWYoDv8azbhhqFuvpmdj1iE2bUQYtwvvIlc1H8756Qma5wBcYdEJb
rFT3HLZViHkMIVqnYR50ZFaojTtsTYIW/nercHLM9vjPhOtFv7TJBDt3epMnt74giIOXp0j6rySK
XMOyLjVeQCfVkpwyDbTps4NJhjZMF6vIQjA8uuhUXkfTPvK7/GEK/wOpT494WlnTxsJMMf3owdzM
3jQ1w9zZ4Wid4Jhp42PxEEdCbM4STWR+AEj2xCYbt0EZCjL+gJbqzSjUo3IW+4S1jF909DC0Ggu7
c436hqqc6Q3sgX4jps2k8SfeQ5ptVocDKCAm3e/PtipOOOQMmuaaj5lOugKIXreZPoqfLw4NpXnu
Zcfr052sWcuM3b2eo9DJ+3dBx31mxm1PvZv19higfh9njioVBj8rqV4kwZ+N4KOdE2YxrVlaDWEp
u8JWCUOwv+eeySuHuxomGFZHGffFV45PcJsrr9IhWlZrwUJbVrVlqaZbr604uXVyA8f5hgg9v4/d
v2t3okv6HDD77gejfeycpK4P7W9FeSdWPAFCWh3Xb7uSFdlnGYRWtEou5DmD+zIJ/r8MntgEGhUb
SreraYsd/S4W9u3gPletync34hzceI9XRgL/a3tjfL/MQCVP99XX7+aVpX3R8n3kFmYrDA6z6ia5
EK7PeHa/8gg4j85b2ytuBmKerSpgAvKvlZyQVkyAZI+rAdOtEjTocLg58TT67A+c2hojaPUsfrEQ
CRgTDf/fjg8ukoS/sd7xgqunL+GIRoMdnRFDgHHDs74x1FQ7RZXYkSOF5QKcRIoIvzowMUQ5oXHp
EiN4el+E/YdudfpNywhDe7IpKT+ALLX8qjZYpsi/93Uj4+K00l9xXcTbhUUDS4Gy+pIu/mvsIqi1
4czy/n/W1Q19ajijBuLCAdCqNEa1O7D9AQMfdL6bKTBR2Jp+72nWeMdaouTclmOMw8fb3ZaTyBBe
S8UmN0ZVKyM659910HHBb0IsP1wUMx9XY1bPh7tbnX2ibKO7UKOnuOmlz0Q/sfwlX/7K6WzfOxqj
QHlzBKYiffZlyzb0yXGyZqi5cXCM9CQL7WZSXsZ4ddd2hGnx6ypeUuOKq5+Xt6RtASCbJ5lZPAOT
FZUaR3OHR6IGmvFQZR5lH15VtS8cXCyLbuB/AYb7hdjbt/YOXwkVMoaudui75aYQ1j041hnOStqN
dVhRWAiuUKOvOI0UXVptaQPJHGH3FF90YmNyLorZxECGcDVkpqtPSSPMJITJBxpDJZ5UoPwQXP5e
mpMYZm1dUMrHYut9GLwMJIVVaqI/WZnMrw5tWF13DV9XTv5Y4+TruckchAfNb+3rXl8lbW6RRh1v
OAy9a4vVmX5S0pHkzEGKoHJ2RXt9ocn5t9M8QTrTJHipKrfjoNeJ0r3ycPyPT18n/EqpTg9ITtU/
SteLDlc75aElu8tInbpERCNBo7xL7Urk79dXaSHJwXPGF4tYcbBTaOuh/tzRSDBhx+Evqf4pZDNi
jj13VLeiVr/84QVHaLnH+ce+YBA1i9p/Q8Xx+l9cg3TnHnreGSM5CpRahqmjV1FZZDTFJBhB++2b
JSdeJgxkjmhq9Rpao1wRWWnBDl2D9E9GB1t+p+cYsK8ZqRy460bKCBu5tsw4eNkihbyVnsSlEfgF
AqNKMOqvrFosfiWwuTqUXxIMmCpGjvcHHJJ6a+S6AWBx2byVIY+x7lrRt/e+FpLjNuVe8aDENrKH
z0HeCgal4AQitIuCcVdQCA4slz6/9+iEXk/ZmbsDI1KUREdh/zdG50hhlhTqSabvNgaoVas7gpf0
e+BjXbvG5kfXSwCe6y33JKW32f/PWAbwcLCQOab3hKJG0za2m4qe3pWTuAmRCJLAyULZYmy2IzjP
FZUR+h9mKhRsnokWeAq2swYa60gT5JcHynX6CqujClrEvWxv8A6J8YWEvcNeGqnTukaBGaM2fkta
AKIaN+PpJcnXxfV5e0DoyLY92V5lQseolUTfhpZy9lAoGA40Lt5JNOoe5EmF1tgpKFLiAdX8uavL
QmiauN2XjdGydptA0IptifhWooJklP4UPc5z5Rq8tW8rq1SLqpiZOu9eHNodKwdJbJn8L3v/nTtw
Xq71ZqsjNfEfP/2lbDsWAU5PAxsWXcFNJRjaJ4YpbdbZn4JAaAu58SfUfGVrIX60hJwmQx+DoFYj
dLaj3RgvIIK9pYjok6i+48r7HX4rZcLUh3V7I1cNcOxJJTI6gLlGtz3tnX9D5saDYEm2mOlau3bc
nyLTwpwk72MunJwlTJOpHXwCo8dT0YpDUw+k+PNM2VNLUtIQN4aYItP6BPdR4wMVA4krnwydR0xi
i0+UkywV5dCRtwqGwckcP7tLMfj0xn2sjNttlIWmSw/iVp8rzjAyPBOjEalZMnYLj8xGKGPPgexn
Xk9dL5d4TmLeRLhHQXjvjXh3xkK+wPfnYQgRFDAX4lefOjkmFq9YZCQ94ZkIVw9MKkAyN63Vkvqt
8rXMP27e20zsQhjiMM798JrwfpOFM6OrpiLHVRNPVCMlYEilW6EOyMfZ2R0A+M+Ujasmr9Flmd9G
Pi+9Bk3Of50VgCEPRD6ZzZoQ4WjTT0HfEb7zUnkfeyF928WlWyMKH4OEjmM6o5KbWDnvX5vXfv03
4/ysXAh/qaA+OMZSAGTEfZJ1MKqEK91IdRAq2maVNKSKwAO4Vf5FPtqYkXqmvfRGEqUe26zAMKjB
G079eWctManAUbOJ88G6BCzVxrWR/UsPMwJVZn57L47IGOEUwlDFC1opNSm7g4mxVDSAGJ6Et4cq
Nh0uVtPrRAAoLdXxLoDxrYat36Mq5CMpKcMsNvrMBXEN0GjImlWp/NHUsKBkyWNh9XQDC8o4A4CL
9YVNp9LrYwh1ncDx+CMlPir7vg8obsD1BaAE+E20+fPzutRImCEo5qTwxwQdWgLSIbSpBYsWH3rI
p37tUmftaCoBmdanuvlNALlmDwFwZNBAM2BHYfWNmEFAvIIm3tnbAEg0yUDqWp/W7LApBW4VVr9p
Omkpig4rzdUPwzJc9B3eaWRwj17caasFC+ApJGtvcZmmfwXHg+YtHdYrRFkWXBmtnoV/vlgabqcS
0+yrD6S/Qj+Ex81hc+IWok+D+0gH8+hCcH24Q9WAOMRNY6bD+FBFrzF8QrqzevKdX2rnJxj6g/p5
+GAo0qHpH4k0wmuk/TESE3UeolTta1UJhnfSgOXlz3UeDBjB/UijrdtzKzJ4MTEc1JQ0W/X/GUl9
RQSUQwSueYEg9Kuus6fPcLCuXrgPjn6UHv7Xk+coWgUC/6Bpzti3OTvF8mmP/6in7XDhNUDHde+E
YaykJkk4WjhNn4WGCx/KNdSk4lUXCNIPDs+VYcKPOfr2PYKcoe3TzvzOYujwzvX1TYbUuE7mIgs7
wUs8qXlXWtEo/YLXRguq0VpKDN7EZuXGmMOvVYyp+KYRh9rYEGWT9KCzquqa63CAjenFL2rUfrA2
7qfFadQYAggQIqU3p/uyx3lClFxNwrirt8Q2/v6ISwMtlwIwM3KB0qXFvK3VO21L9FLlS9EA5bwZ
G9uw6GXgIsq1iL+AWdEff3NQjjeGWXHsCUnqfE8wvmExtFeg8z3phx/Y7I2gYGkswv3ZlebDOiNE
lTZe5QAq9flyWr7d7do/ktKP1dGcuc6T7qLeTp0qJxn5mptfsEqm2x/lQQMoAENwPjDaLgKImAbL
9cjQpC5sNYcGLVaJP4dTBvsyzgZpAw2fKTlEmRQk4943T/KZi0kdgG3Yl4X5Ne0bqVZarqS3LLa9
1NktVM9ETWzfErKtgzDYjz/z+JIA4Vfw81Tz4XU25KHF5iY3+Lx2PWtkvMeO2g4E/13cO77t+/OR
Kqe3Os5DFIfcO4Q3PPq4TkLPqilfX579uFczSIQtnbZnzOSyGo5Z1PqdIYggjU6hVBa9IS73qF2x
owg4oJctaANASUnUMZKvbPzDa4g/ndol3oXFOVNDr0ULitFySEzzFwoY7sslO0cIXgxLMATVsWfj
182vW4Fd2pfQ5+SDkEmYq4t5GpG3jSjiRWhs5LWTuqiZxrLVxUfFGxkLUuWasEiV7bSLO1CYTaFv
b+fM+23e/EQSBFpKIKvUQMuKab7rwSOqjrT9r14ZrJbCcwlttDp09jcAao6t7bUIcLPNPlxgPJdp
5BS15rYKVv99jQ85uZfwvw3sFy8KC0nM62wp3b4WCZppfX4oMc57XkOZZ1JVtj3+DLiiF/uQQO/3
pjpOsdU89VaMq2fd2Dil+YnM+hJPiV5UXmDFK5W/uwFqSCsfgjvMsDLK0THxGnM1N1NFRcV71AiU
qAzDfH7QUzn8qYm3hapl0ZfQyJksgaaF8q+hE7hKrj9y4ULtQkOTN/9vLhezXp/8zeo3FyZt9VCs
G8pdM+trdjeluSg/6AW7YEWqMuTTf84wKFFkFUD25xkZvAQBDfpns2UcZ+patMEF63jWiHqajWsK
2oNTBiBjm+tWWR/+X+oR8H212SDyzwB+4Xwzch1GruhK3u9T53PrsYOtCDrcqxbKVg6aRC5ODQVj
sZeid5tuWuozFTG8W+fOSieD0gDeEEJmB1ooxmyC5DrBtof451Hk3wLWpoVI9b8f6VueKakW4Azs
uTajIjGVgZOCd9kRJ9H+jFOwFgbbsdnKBZ/2XjzFTL8jIG4tTVliRK6TDW7IP9WmZj22Qh4l5876
Zrop5zv76dU+WxYW+J76uI64dbu34yJl6TfWP1X6pSuq+ifPW1+yQcDRMlA8zgNhLZtU2YcnvgYJ
14fBYT2djK3U4RG6bmMMM4uN/0xj+URN9RTrhRbXmvxpBfxU8jSVMkbCLYnC41w4Ty+z0W02Z6gO
Zy2Lh6sr8gSJR9ysK3KNbpNpwtkwR2RHPuhXWRwMjifbSOtDGYhqRfop7JNJsoirf9HcLU3U6wkQ
L5uZdDSAKCWS/2iD7GpNnyDp5Gi4fIV4Uy1Qf8avGh0LjBfKaPldynKVpFn0tAUUg9qhEgW+tIi1
VX4voAPtr9G0IAhC8oHSz3GK96K4bFLFXDhRjVKFODYAqPSQlhOrFiE/YlcTL6QPAbRspUVCBYNl
Jl0TAfrflwQZVSLAQGS27mJmVmk5FTsYOi3OIKaIpNTQvM7E6+0E6l1Xo89WRryQjA9Cz/py+ZMp
QCDYbgLXkGx9JFh8ouERZ2gZ6L66J8OLdyQ/TTPrYu7378lCRLOL7+mEK/85QePQMinuUnjJyXTG
nSyiH5p043hnpPmrIcElZ0eZd9dIx1RfFLIfigEiBOAXf9DScD/lp8nT7epmdgKRmawZD67wFSl/
5jiVwz/xyhDo9a2Z1zUbZqGgT3WAxkfIY4o7srX8XiUxDLRSeqd8xTfyg8/YkLF1E4e2vAIXb3Ap
0BL43SI2gTBA558GaS7zzqVUOeTQ6o9ykHn8CdBE7QvD87Ef7o5TNTqcCHgsqtqfLrU/WqyGJH96
jqH2RQ2YSRaz7Nc789FBzp62gfSOJJ8nTDYUotCUlivsTrnFm21w7a5PVZceL9ji63MyP4IRWVow
EuMcMSgpef9EVn41hVvkU4NvdH/z7POQGqlNm39mxA3yXUHX9FQuIRFhVwHU69mzFl/EZrwDAcMM
q9lNyyIJ7wwmP5kyjsz1k+2znyPx+qZFlWAPsXpyle+busx6TP+/jDJ8EmKmttkTBI/rxtAy7fIY
aOs0/JudbrnWP9aLimP4MD4oBMCJE61ecQu8sxWAme4mOtvA+BWMiNPjjVtWba035uSafzodqq4M
WPee8JFkbW7j5P70FJZfVrJxcp7R9BTjWSUR4O1mbz3o1qJtaOhZnkVBxXFpEPiLFd0bwpJXbXt6
7OkDwfF5gWqrAlW6/Hp5fecEz9HI62OZ44jKliZ18rGDo5y+hgNGEpg8IhyeReKcs50K7rAQ45aa
mOvOfjOP6t6IejTIrAYJHxZ0ELc8fwre9FaTjchJ5T5HWJGJKn76aCMd9DnlYEx5p8sLMPfAH6XW
EGHCRY6rZd7mqi8gp7zWeQ0qoXiw1+uPt6HIoLBsAzLOTWm06r0qVMkkA266vFLtFdbMEAR367Uy
tUCIriKNCUmGGCCY5iP6nqDF3eegfkghLZALQl/PAN7ZLmhtCJvnkzm44NB75luzzzoASFXkz7BW
WyLEaZ/b8D+JwAeQ5s0JGaCzARhbeB8dV7IAurfTk5OtVa5nBJ81PZpxqnd1GX0Xy3b+oZS/gRPR
YzJ/KVWBxz1TtCrnFx6DJnql3TIyionlF0uYlxmEB2xBtpBTcbcaCC9k7Y/nCAihjRwi6KC47QXE
OyYtBVyoDa6VtJ4cuGdqOT9r/DXdd/l3ylG9QjMzBO10pfWjo9HmG7gjZojTBI2elJk9U2BBG9+F
h2QwgfWwmUaxJM/7BbAgLRf/EX+Te7tnEK+IuJa/HaeNlD6CSJMXIZJrGM+HT+WBYogTnt5UmnLR
69rDB50bmNtaoD5Np38yKuEEL7dkQihB9DVjoO2DIWglullmnAVPJhWmsHYKaYzaVO8+CxmT6HUP
rhyoH7BrN8e1+n1Y8Rj075Nr7CYR2KyBrWYY0wzxvdtOWNuCiDVvcnhLJQezh5kTSQHCbV+ZQHyU
i0+DnzltelGBABzVX0PzekcqAYOPE0q8pGtFvZdUiNrYo1pueJ2CWkPL+hULF4u2IsOShhswojDX
WDgGvYPGWFzB3xjv4TigmLnO7yMqfpdtH6XaKoUUEdtKabDzV0fsww7t2n2M4dwPYZyXlUUk5VVI
fFnEKDq5ffzslezUWDwad4bXEH4LdBeVYVJg4L8/cRWevTMcsOk08iLX1UqIJsdoCV2oh4tQq+WJ
zLNApl/BZomWGXZqRqqdPlxayg4wkb3L+Cf7QyzErFBmPL0Dpt3BUncBWeRi/ohebdSpRqC+B7zz
ixAQ4tagr4Dm7GhYt4EjlMSj3PmBAbTOnpH59xb/WJHuYbqn9k+PJWWoK/np6aHHO1Z6JvVlhtqh
t2bG+g0viLIloFTERWayfmYHpR9a0gaRm2rxqSO13t3Q/G6+XGjoVMYBxKl8wJAWPQzo5pHlY+ey
KFpw9w81FQM6I3MWQ7QMneIGINPghcjg9itwnq33jmBEKqSRarOYCzOFwqRNMqgivNtMdj9J0bza
0ZdEyepfogjihEa3/lpzNyi2VJqosD9Lx61oTZs2mMMc45txOeqnRHcf5VczksfkrKAQ5hjGflpM
9h5XUN/v9VTjapjw5+tP4JJTptGezszGyA+0KTmb269u0kmRp0tBxKVXRVCilEqeCZrJBtilGQOU
O+14T7heAmJAwwpAZvPVEaAgb1E0J4Qq28D1nRriqJ5jQF1t3p1MuJ4270zaSDSPF0vuc7bdge8M
cY3sIIzx46yTFdNwX8U64r+Fmy0xYIXTYqIRcIaCjIWv9x+wmDA5Hm1JFxfNaNyZtF8lh5BrpvxD
zRIxH8RPrtCN5Xdz9zWA9XVQTjraJrhluN6GkKDR3e4gvY4qeqtV+ivANaWa0AOraD0qL5P6qKCG
TeAkfKcZFWvmOtAnWMh+1lu+gyT6EDhtgw49TTyZV8miTAtoCvU8RJ3FArSGlC/Yb50RTaOAuoXx
Yp7u/PjKb7LMHa78YmpbE8dk0DUKo5bgsb5lYMJJpjKDsVZX9sJplAC7t3WWboUaiuBQMhfww8+D
buIs5uzbi5/qogABfzuuoxAhOvfu9XyEeJ4AtmxqcqKhhD2pf7oLLtnfL8OiVpxe+AsIabLDryxf
KF+gYAV8q6wZkxNRNCAfun4pCm6ga4D8r1vaxxn28idb7DZabXEGRQGuDMstKtD4wfzy/KPXg8I+
XIbZ1uVa934o7VL7qelTehBQkFrPa7DT6ZxMM2E/LRG5FnxhSG49W/P/nA4iDqFtvvGmHnS3N7IZ
csQpVUedEHJmiR8U6adYj22ysLGbfnb12i8qS39iyD8ADi+wQkh2FJfPhgSftgFYhdYiSYXAVLJS
QfrvUTvuQBAHEiU7VcgVFt6p9hFDux2aGdKuSpGJblagm69vsOaX0L5tNvFRlHBt2P1J/0ZjEruw
5ZbmtQLj/3C8lKYd9c5p9FO6KvTAcgP96o6899hTM0Rr9Sl3ZhDBYqG0tsG+S+7si8yAc3OcysJf
Ot9bqcUNGc4kpnQ9OoXjLNt8TwdQwUzeoRuPFahLdHWnMCsr5lW8j4PlazkUY0Wm1IU2jS3USiDa
Rb9uGTCl/VAmVTdE41qrX36tYu9xj4Ht59YN/81b4cwdENLlRhqSC6U4aeLc5ua5wcfjPcvMjU3v
kX7gKcWA/Fa7nVo75rsQLLyLBItgnRceWNWgbJAZ9ZkCipv7MkhANyyDl93AX7kixFGwkmmM5f4B
LTfVnKMqZtaqxheGh3dnAg+Px7pS9xtXdopcyBVFNb0R9aeJXoD2Nr5njVQ6gbqO5JxcsmQYdseJ
5/qwx41jhOqk+zfgKh55aPieZJbCDG22llgWxb1EIWz4r9gaJ3pPSmiy9lygbMV2uXLFOqvwYof0
Kz218wx97G0sqsr74VcPaZdK90MUf8Hpk74QHyUjy5inkHyfXw+FYxLkNbiSrfTGxIxRjz/A3FDg
v1jk3oAYSisvvmqifrzAF1Mi8u5U7QKUH6RjBXBQ+ffymJMQ/ES0S4CdSQtSKrRxQY+entgdq+hB
4Vpme6Kw3140caR+PBwY/pB9M/xWmXbN0CVFn9da63vnSTmLZjzqseqaOPswGrc4v0fzh/DGAooi
bFn/+7DApZGJI9jN/NGJS0hEzIhtkVmTyIYRTZglAO1ov2h3f+QgR++JGb129ooZFGucnDjQbD+p
c8yf9gr7mf2gjPON3OLXECkgWG6Wyx0U0FsbmyWB4ES2827i1C2jWsbd0arUhHQ5c5agd2OGT3Vz
6btmDMFVZe6sZlFQtDCOQMnVzx5OwLV7hI8a9OF5ZZRaFOD2jfVMVVruij+GnmjPli5uLDOFAx3k
ZW1yXn6S8jSEgJSFIprKZqU1wyg+GI2zaBfNMWstLAr69z3BGMpkUedVvqAxxpt1Zysk3QsCnils
oUmZWkr5sNGhY5y4RqjK1ZhoizuVTsbiP+T1p6A5Y1uQPYrF5CwWaRY4XrPCPgsy6r+gk3gK7g8g
FayIqSROxan8y/FkSO/jxk5sol6m9wbmuuBlYLPLAsMZPmgbfTCjm4tazQa2jb4DeHHcReieaVUT
QTNG44oEIoaV40X869ZY+76SsrjuSwzBU0O5URUKMa9NN0CnXZV4bAet4oP01IEKeUGnYoPAzwVq
6gZeUMHrDEpCrCusws9WWg7JMc+twqpXcecJgvDNDHi8R4Npv9B4L7j2RLI8+f5yT2MOCNMXl6Qd
zYjWGw6KIA4/YX57IwN7RgH2D2MxcmtehhJJIJro4TJcvzOLOnTEXoGD63K4twlEvydyvADAyi84
jKYu8jnteCjgtU965BY2dskm+DS2GRMxhJWlP+/zmKbeefeDEs2MVBV5Tt6QjtGfuZJEsUPHGlPS
BUofRYx1VezVeBLVQXUkSQ2ZIUyo2yOTMnYndlCa/OqziLgc64H8nvq1OHASETvKVtJX7utVQu1M
vxE07tV+wUEv3tMIicMrUQc1YxAxf7o8/uz665RHTWhlK7dspU9XwMQUzrc/yHz6r2s7Vkc7Z46O
1PtTtQgtQXxMsu8+QpXVSRlqzUb8cMZB5ndz0Y5eHZGwMNF9WT2ZPgwyCTQAaCVpyNaRAzrXaJo7
R8YwodkHQrxQIqTLekw0SoniF7f09rGH6oyNIohcG3Pm517U2o2Q0tIycmJPJlE0enJCw7WDJAKR
tohroNU1W9nZFJee4XCu3TTWDItfsEL2TzzAtCl+8Tp0JHyQepgF+fSfEKmUJ1w/NHTtLJ2Sup5U
MLxAtZ3t0PXmmeGUE/b2ZxgwKW7DjaW3ICsyaTzbz9FYGjD0tBxTJqyJE7Ce7Igw3lW6XdC3P/ht
HXrYLvqx6PCYce92UU56G9I7pNX0IbU2QxlUzcoMnz8LBFZFG08x2PAn4fEObmJir/aQLWOmiJ5J
w5cVxjQQnGyMvSUGj/wEopPGJvLd8NX39EEgT1I3f3ImexPGvYyHVid3ZrQ/NWIeL7xmlWHo2pMG
1jDPFxGQ8IxlCU/0yYXexNXmyOORoPaqo7udspH4B9wDrIwGJw8BWodLl7lGNJAS5OAM8c72UYZm
zhm5E/EWfwelR5eVbqwaKXM9Rr/y44z32SBj6jjv23qI+Aq+bevKd3RcILqQcgINPEAwZaEgbfuc
HTIz7bjfupCbMSVfPkxZfETU8h00n5yOa0YX0snQcRD6yeNDFZF34rC3Y/qrjgowOF2VCHiNpwOE
eFUHCEtG+DnsSg9zdPZ7DNNge/IayrcMxPEphbhgrcQaPGnaLIDxfhInbZgjSSFkszDWHt8W3sAE
28gESo1I2IgN5qSww9pCanffW9k36z5+fCWXVz+E7YfRT04fO9PeKgfWvosLnxiXOzt8myWR3Cl3
cnUaa+XKfduozd1sLBzcfHIgPV91HQikgnGcommd51AfeqfQTAvXi56jY/yWQNZ2pUMKcXLExXXM
JGcZJaYXx5oCFEwrluHTaTdjGmCDjuthTkMflUJZtcZc2Mlhkze1ZgxNrQhSKjTh8GY8azxTWF3X
T+Vqnvoi56Hfhvo/XNZ2dmx7VKcTA0miay4f5pQQXtBQAJPRoM0GMb6z12ZTrzbLW/RGIberkDHk
kfhv/hQvnCIVVwEC7/PvP/IoKqTZFOnhIFn/48P+rvd5ORszKlfBixHRJ7+Rav7AuFena+pmsLgW
5W6U1W800D+fdaDnVzXdHs4RQz9CUHuzAi5z/xaG/PYJNbo5i3lQhmb34xm1/siO94xcqzqAcAFw
gmgNypF1+3CWaWopu7aIKk52xyIcMRrjU8EswxY5TOYDZ+GTDcG90eyKvcDCK3Q6hyYF0OMo9oz6
GM1+KhFTRjFqNS1+2i5kuyapnD8dwbQzC8aDSjgccLEJiOd6DWfeGWNAqS+kPXaKcElJR87JcTMa
Kes4YNsleQxfOKH9YPW1DuhUIigmhfl3ue0wWYLQxypWOMPsWZvGaccdMW1pJB1lJlyGD1Wo+pE/
eg9zhjFy9HlxX94MjKf+OVXf4lbNT284VLdxg5zNCqU6cLkHqWzl+ySo/+7U5QXUdPmBNGBymsXv
n41LHPkSy2ePK4UEtdgFHKVc88u5gitd7z94Jkk3R353HTDosVQB2ox2vhrmrPMqY+xwXeA+0l79
o7ojV1aJ3eGgtvYxqWxmDMkmXnOgJUUv0TjUjZlVJE9qaqVadj19xrzfTzuW8x07wqno7Ep239ib
HbyE8tCUy0vmLYpvmG5vsjeKUYLwPa5lbwjXWLObiHw9weF0vdQ51OZvFFsPSPtHnqqDg+xSenlr
RePuP4Dh8+0RbQSjhvEcrSMrhEu7jh7ujFfczHMhljolGha5g/ESwS3qdSvevZDiaAFN6kRKwxYt
N5CfsC/yAGilKKd5B9VCxPIq8x74Fh2+wTOxIqSCbErTcrzqtwFk0sGr8cKYSaGKe7nK7xaI0GXa
3CvXCfNtvcSZh831xdk2k/BPedpVCcaycxd+8KwGhbXhO0us2FGGS8/0xRQwYRzACd4uhHNsyhXt
gq+AhSXgxylgk5WGCO4wTrech+eqSRlm6uo3Us5hIrLjwZ+sQ5j0XqssteBJHDTkpiFIaNKrC0k2
1u+Ya9Xn8F8oFr5aXB1gfJ8aSX8160jLoRtaZHdQASOU5sL8BrKWo1jjjHpUzDK3iGuF3KaKT7+b
lasJy3z4qe7f3C4tUzzTZyV3v/24TjZzrubJJ0s02CsjjLe2XBvLzKXwjKiyohjv4dxBmi4heRhs
qYAY2KHSsos9aTlXfmwlF9OYkSqF2O6nOd0TCo/9HATXoiM0lIfxkFZInuGOtEu8Gx6qpDMJe/ZM
BJzkMWlgkuy3Jzane6V7tPelgr30c3Gkfl3YvnKRlj5ebZcWnxgb8ptmQY4MgxxBZUiT3DfK/AeU
p8mDU3H7IB9TYUnO+46tFT4BQ7MjaWjn7h1ygRlsLV1otg2OnBuHXuDe+no4Op6qkxJqacWBgIWz
T81wGgGbae0SUhAFB+jfY+vXtornm6KqC9gjjIfEr74eh6t3V6l6fzZAR5K6wNnMLy7ez/NhLj8h
vnhvZwv5g1MqpV0Pt5XJdZCWZwVwfz6p5FLn3tfneqxuzLc4HLiKtyFZbmDqaU0TMvcVz8Z9KapG
/2JwkoP+VHIhvUCnu0n12yehY3LmKfX/zCCPdNeNZdWriIVPdTXxlUUA63u5f0X5AyNB0Sm1dqJx
jq9YLXrGZt9K9PXVXD97KAYy0DV8SfT/aTcuItsrXFZ+nr3/PzbADuaLl631GKdPO81EfbMFwKrS
/1drl8yBlx7z6zUTLi4GYkKMxBqQySmtcXNN4cOlL78oWnCesfwhZbuAYMKq31BxMnTEbTYGvuGV
Mg4u31/Xcdv+G0xFUQHFmAWBfTbcmvzS82H6D9B/JfCSf2GxRtUV2NX/pfEyaKpXkH/pNrFm6Wvz
U3biLt2ccTc8X2ouexKKr43JRVjh/+yFu5AqaCQLNtzdkBnyK1S73Qc14/IFaozV7QZoC7jPpOtL
1/xIhSU3ybxttyoVtshxQv4CLaZqPxbqWNLrd/bnlzVuzVYocttGNdMaVuA9dngCCIQvq00RNRyQ
0IY+Ck4aG1QkTnCbNIF47tYeeb1KJEGRi+ARJ+Vs4mXygErx4O4MG+LjapvQcIhLGwdJoDUJd+Gp
WIfTGhJLVaJx66mlKCvCgKPW1H7zwIMv/7vmQ3ZhCuQx/bp0GF8QfaXMvKcRxFE2pa51uRyF/a9G
CbiMO5qP593h+A9xDaopOcw4ZxQl7xpW5xgcKvFb+RPm0ovrE36Oy01cDSP9sxugxHL4WKmsPwqD
7HzoCpyqvzDsD7SfxFw5L0h6tnodGzHlrrc3lSRlAFMJQ3vkkahhIg4NpmEcyICdttaa6CJ9tFMK
v+dPFZ66CbI6lK0VyOHgFugfRW/9pQ/ezWPm+BygPoqpgpzQpIcvw+GHklO/uiOhO2sYssjXRK57
x02nKTUYX1kQx2ehaba4pIwMCkMIiED6dwumHuXMoKRYX5PTzh8oPeJxZZs6ag1l05yXdbBQXTJG
xuPui53eJVgs59dPBVDIf9Wvm2A4cbd6N8PRdOsHEjuTMt9YPC9XO4yB8EV9qvbE6ut8ktC143Mn
a7aLgUJsKJz04TkX7sO+c/GAdAKtbWgwRzkbEX0Z0yela3YBIlut7foigsrQ9rwtG4EF17ah28Wa
qDto8yHKOzyOoSXakz7aDvZIWgZO08/5LDQt8OHxCzSG5VWBOKjpepTwyevqunFrelrB+umvKdw9
8YGAxUeJ1LueSz6xoUSz0o6fkgjA3iexAxKvCXPxBCeiyo2k6PhbxNJvhtgC4oFb6RCSCABYpfLf
fayqKAvd036BMIF0EyN1Xaq18aqHK1azj3nyBkEgEHqBOZTcp8uH4Nb/ij97YCHUuyt7dNOtH0So
aMoyhZdxEjulPEJLqym+YMcrrPyBQbbx1SzftUCrtm7hhjsqkT/cdt0ArX1VZTEySzaAkjq8wBUc
vyYmDlgFfbSGo0Ku33Z+Hpz/0VoVKcX99woMLmxzXEbEZPy90CvHNbJ5CfKl/O6sGdhLge/UH5cT
Ip7nSDdsWf2mLytp1SkFFs4vRrh7jfp2CJGxAgzHXojhU6A8/EOpWCf1M/1GxRd7CQ6Zc2xN9DnK
R1VlPWBgApK8Fex5oiUr1rC3/ByUYhYppQlNVmQlh1ZOpUbdnvMngxblWzfv73j+9ePay8DBQ1YR
Fh8mocQ45ifZX3m9DPQzN7v94kETnjArT2qOFfy0Iv5AoN4yQ7MQEdw5L/MYbQAIa0xJimPadvL/
TuBQF9PQznd8DkIcbKZQVws0cciZFVcn6Y8CWkGEgY4KgHRDpfm40IdBYA2C4qFsjT6ltrh/Gtks
G7wain/jTIXkpuvvHv0idlpOCjXC5VctRh7GzTLb+t7mdbbUIJNNYhXwOwcliDCgwswEIMrQPk7x
jH3W/XP8RDGOUNWo1sON9pJWDUW/Ote3Z/5CHIbq+8v2jI+092aKC+W4GSNGmgtdlvo8APMMrcQH
uQ0ibaesFSyXS22xczZBq3B9KaeEb4IBZlV2iFXVMZrjtTnVkYZb3yQIFEKcU2jWECAfnO50xRp1
tPlppc17woUoGEnozQmChAa4kctMTpkVvkbbUxxAPqxEdo8KmTATExg2BKiFRKinpOFo/Dd+qukL
u7JVA1Hr98heLSdLCb5nSCedN9dMpl9i/C3P+wRYMe6abRfQa4+E+cHcXLECU92qS1nwDYoxzaj/
05mnZgs61x1DpEm1kguMy+6BRDzPJ4WPNO2KhVkNsrjvgCfnIQNL92yP6zn1I0LjuAoXQ+tXnNut
GFFms0GeLbGFFSWSP/3TwAKr7EIMKIKfBOsDQITTyzhFG9MPeMzAAeH6Nn5WvtxdAC+ig5KoPqak
oAvkhNYrGHnulKhODH6U2DvJtpkPTY8GLsfQ0Vbx6wTl3y+lldezVwoXalgCBrBJY/mVTJuXFjVB
y89O9s5k26NhfQoVCXgYziwHf29TY8CTC8Bjlji0sZQgJUBI7LRzQ+mc1mitDXcX+BUVQBswsUsQ
sozsUOfoKLpYCcCpekuqUugprmmFudaKcfgEQhvQ9iFnMe1mYoBj2WDTo8ALTN6tlF+oDFQsGHM/
6k8UeKnrcZgCxSVsz1uJIHt0N4IMFcSOIyDUW6NDd2KD7rh3OIe5hvQDykSY7QBdJjGHP7Yk0xcZ
yw/tHNp/tdrPZ4pXfrUeMJgt8qUpvfi84bq7htrz+vYlD+6W01GGX2UhRmBu+CdFmJKHTrD97Qrp
VeZ/YDuSSTSsFICKMRuVPYbmi7qF9qNTNnht4TLU0JW4L2a/Rv+d4gsFmcBF7ntNxv+F8Hhs3b2w
DmpU4L3/1vAyOe3ON+m4zE3KZMDsweaf7gZlyRJjnTup8MqHtX6AH5dpqMKdsVpd7CSXCN0KBuBy
ZvBMfAbYmsSnXfp50CaL9XkpBVRvgZPtuiyEgUxEdV3zFSr4dS5+jJRRXZe4OHavZTmOa+Kd8qb8
uYFCad+rt7qZIFMowbYWuakg+zmR41y7vUgXM28FO8XgyVBV8U7LzgDXx1AferoJq3dS+Y6N6vx/
aywzPaKPsCuXaBsk9uLhJ+3scLMxZ9Kfw173Or+101SyxHVrT7g7/p4czIqoeEEUB91X03SvD9/f
Jr2Pu9DFmpBLo9hrl6J15nrCWyGSirYWdECZdYuDb2dRs0vvQgb9uspkJidXBcDGPYup0BRliUJl
yzv0Nc0C7mPJf4nCwbEAbbfnPRytrecuzEPP7RAHShB2dky5wP9cMXLJBAaUPba3KkhT+mEz/V9i
lnohhXCRUWPRg843vywYWvFazqaxmZZjUUGJdoiffd/blKnp4yhWxPWxGmABExG1qPa1hBpzYoSY
6Zvl5lCOnmGF9Rwde8dHgvRhcu/LEBoJTx8dNVg6vSAMubOwcrzsn4HLyqNcRcr5IwOuOzYrXVd3
QTIDDiBnY3aNaDNRMAY7KFSn1gpu97cDABaExzbxvRbq0gZZvT6ktcDfmxoI6Q8yNRsidP2/5Q1m
kIeidZR5bGIMgUs3qUCVW7dErcUPPnTdgfQK/S1sjbXcbrIV5d+wIBQ1rU3qTUnKbbLuZG5I8xKK
IrM3nK+Kx7gnLT6Od2oumWmC+aHhhGZD1rNlKVYbrhWvV6v4FFqipTYm54tuFdmHDLqK0AY9Ujy0
FbSkhN0d1/vc/9sSWLlncDDW0Vu93cgdBQFf0M9tNF8xcr9FACmmeCRdMH8SZL9C/STC47LKeBzQ
zRh4G2ODIYRcfLLDP6J0cCylYpWZydpk6Bew/gZgP3jmOmr4/4YF9bVqpqkW5XsC9m5yNta8n7Xa
grjpqGyX5kA6gp6WyMyrYWyFTQSp96c8jclGLWEyFGuccmbTM0G7S3tWq88RPI5C5ASX8Rz8Umze
o0+BsCYgJMC3bqwOJ+i1mKP5fvopF+GZ2kQSnTwzLwrQ5ObI2uV2dOgwmEdtRkcOfs1+Xd6h5N2W
LpghlOyczX02W5ZJ8OVANLicRrwWnBApJBZG12xSMKsONeB/t/bahzNaHhPDoKCs9x8dcC4RYLNr
QO5iwKbRz2cTNRnfU4NuZIhTW7nm7RRBbjVMh3ICP8WG01D/yTJ5eA8LYyPP2o+E7GvBLv6cg522
pr9iONNSZ9s+sBxCg2bEgF1f7H3e0X0YyXSvrLXfCJfJDTCxU5MPh4dM6FbDhKZnJhLMONtZleA+
U00Y1iUU5J8wGrF+/teyXlNpmQ9VY736PPDz/w9g0rVvYwi2xoxnsz7DV2iVZmcWb6k59EkjW11n
NtvAdpxfeXDiV73Eao6XCo9PA7g4o3drzO8ClkyBjvhH+1Al+Jt1v7f8uZFKN94K/3sGtra2GoTP
w+fGbincbI7Qrqdb7c2jg2QuRGHbkVvLGRv4PKks1Kv6VBWAxtWU/JUHZxz+85iFbncMh1gTrvPd
Hoy0lWSkH3frhqua/2xmQbbvzJ9ln4rdJVCdCBZQ+eBrr3Oh5umEgkvRNbtL9LAf/aQBdSaEoSoW
gtDu1L2BYea5QYZofoJ4sYre2O6CRxSt6ANmf11okbMIsMHvyfpdyGGma1k2YFPUIPctrcBaCp33
Mtvz73qI1SmvNEeUEj+tXQkPq6ZiQtzkPIL+uuS6W44LN/VEnCzBvVrgDpFmzMRcQf69MyMsb76c
nuqO15WwOvRqBAIpopeMyRrGSXYMHk3siUFvgTt4uNSb+qL3GdwEJX/cdoX4H7a05lAWbjNU2qPG
nN9A1TrXJKGGwIq1kYpMU5XvKf4fD8dAYE/PW8a1g6dC4Bx22Vu6AATqsfj9qaojVeiArkRSVei6
Zkio9HN17z0gYLHq5vh5FoYUawnaEdFZIqhYniFWQfVmIV6kzVF3xvV9Cx+Mufu29GsIaXJz7uzY
JFoPATO66nPJESDA5O0yXpBsbIlfOxG77xLNI6mj/GXauyHVHz1GYDIP8KlbItocDOVHIHKdd/aI
P0nQ2ex6nk/ey6WJQGZzEtC5Mw0ADm1ThRWqxZtwk+PBFX7KxyRxn3IZ7pnwb2YDi8F37sWijpT0
vXrelNLewJhfefit+QZm/L4seMeNvihcHFuB7pNwomxx28kZ6qtrujL17W2f+yuh4KXvIsHmeq54
+1wIrjTjDmlAy+nty9p7BBM/YZtKoayZwYv5ot2oKUXn87IveWhyyxuq794o1W+T5+R3kXcJqrG5
xu0FjMlnRQ0pfXpLtekjxLIAfV6fTzsLYd/EkOUMLF3MEFweXhFtBVh5F3fEqNPykRJOSUwhQ7ff
6QykX3nRkV2xDkNKjX6y87sbis+xtkQYgILjw46Hv+HZVYcu0xGnFAPeHgK8ek+imy/chG6Wz9cb
likZ/Z/Im19ei/u1HGaqMK5D6LO+LUPB68qvK8usTwYe5nsUXozV96y5Yy8Ky8qdNJS5Idm71Wz4
XTU5rrg4fsJjxNZKGQSLq4TCqb6/MogFZykN5CJ/xfsIQlLLU2Rfe+03V20ybQzcOpPwMuYaErTe
efAcrpbCaySzy32YCaPKlCiPYaV2Q6JjD0bJZWa5/1u98ML7uzu73JcKmdBbnEuIY/QrJ0X4rdja
ysulqlKD7srua8q0oKRQ/QrodvO4AdKZPxmRAoUQYek/ze3QWIml9iNdVd9SrZ4yOJMJuZqZpile
D+B4kcebH1rgOpnYTAadXSeyTtFbk/bnZ9YXq8kaI0A1FD0DQi5Y6wndztMz65Qcs25UUgzktQCp
3z32pUo5iSBkVhngaRIXSpcbfMYokUf1lK1kT0HlSFrXQm62Ohx4FBOpiy0UWBmnNS8pFGirmf5e
+ASJP8ErEy7tnzCNlRLyJWwtxA1JKG4u9SOPgA6/ErIu3FMOHmxMfT6GteptRIrQiLn9s/IcUvTr
AIN9dgrLWP4qAxbE5yVymH5Umt0s51aeaFRQCGVnJYVe3mCuYA5blIHJ1X/QAUu7iSEdCEmgjypc
x8BPB3/lnPiVecXlbetCXqfvkN0a81oOuVVS/CWOOqEFt/EYN0+5+AKmTV35TR5KEGywkQYXT7DO
pjgHSDGITEI4At4nLnRJRSrzVc4VyOlg5faQOQgsHp1LoMROE8zt/kW4W6EbE5TOqwWFjqAdtlaA
NpBsPbXhhynTSEXciNcUlKfQquI0YAzcMsERgdrILLaXpW/i+PxUk12yfyJPf75SvAKOsz1BeQHl
pFeGbaHs0xtMB4q0YOZKHXgv7t9mThB26cOPnvTNk5YL3zdmr0+Iuf/4OxIw8lEG4Od6a0NhnmEX
E9lOcKt902kIupQKEh68DuK3juAkotg53VPfoU1Y4I+gJOiyTx9gtlvTkKq2bkJ55YriasLWqtDh
k2B5RKFbqHt+bMK63AN+OIWUwosw1CHa8W8D4urEipipW0lubTk9//Ntae8NFDzFgTz1j7A0uFgc
RS+ifXqjjB7B4s+VIOouIiRdqOwP+EbzYMU4KqLZmaogan6/7GWGHlsvQnxxVo0WauCNefrkL6Gz
W+SJLHCkkV2NdocUkj8nCJnHlFktr4m+fBXiPFc+lXmKb4rht1wikMDnFBF4/iOPs9icbj5PUQ05
BHKv21go+CzbzGrpo7edIK7njGMx/M7UkyBUXc32dxpSxufuq1TAke2pq1+2l4gOys018kVaAtcl
YsC0+sKpBTlXsLAt18e6oUm7OctFXjRqOR5oPrR44Ol97TmHDPDwFdpr4BnNlaf6+gc969X7jjA9
92Ym1WdgaBMJVMFvkUk9gPTQTxv6qumKQDXlRyvWbuql90VW94dCxAz8OiOg2RJfMPmUQQjGiXPo
8VemcsXjKJeuSZcSyndsKfk8stbEzzo0XM3i5D4Cs12G5OETS2pNNk2/S5KB4HQ/oMRzKDbSoVsL
QWhHPp6e1l94YPbCktQw3zoVgb74ezJtJEk5KEHWGnV9i5nxHqqVID4vRJybiLUDIOS3lrNWAhAs
K3cjQPJ5tu7dKQwLcDIi/SfjnSwpQFRqAIhH82a4cLNk1PAds3XqUIn5SYNtHMFwMkOcDtn7Mvdy
UBu1LwRdojOHlIDn5KjNY/hOu8MmEhHl7mXu4stDpl2QkMSh4gMsG5wASQTs3qWU0TIVpZqbaplg
YOt3yJkQATEzTXH8qUwQSVsSi1qNoSVpVCs792jGzO8jmgCwMe3TEtPprsq3hoqb/BQBDIkpI1pL
WcfiIXu8GRB4nPvGyS8xkjX/jxoXRPRs7d2IBgy/AgGK+kwuPMrFwaiV9091jH+OyEALkYSRzI2H
beF00iqSbUJQYAH34OGhCdF3q55bYfut6hfJJU881El7bNgbgDj1ennIfOlov8uKYk3GTRH1P582
bbnPQpPRRrrf3MBqsjhLJW2eaG21OdBLAK6+h+t7G1umlWCLxxeM93AuITO658ojP87+wtb9U4cN
wgj6Xgkd5p0pzk6Jf+Hm0dT1f95Vhcas1LmjHA3cIawQopp7LJFbLb1xL5FdPZjkbfKARmUk6EmZ
24GT63LsElvE0k6K56MvXr3nNDM3yBpRtdPfe9HKqRf4+qpqcSaDfdMgtvZNpUP9mT3ufwqoWurK
jZx8wMzhmzbRHAx/WvkI8o7AcU8CPpxM0licq17YBSzLMD8VU0SOl0vWlJB5Q099pL8dpkgURUU7
cdk+mBK/BnaL7ktmCsCSJNC6MKxiAh44ndsakGFUc1xhufNS9m+/W6966t4V3/ch3ULSGq7smUqJ
HVU1bck411f/W2308/h7EwNeNXPHpFWdaFw0ZAyU7H2VZZcYXDKIfVWxxkviFJX6vLJEW9+8sUzo
jMXULHnWyQWBqTxKDknpyaZplO3SgNlv+gKX82JiPGmVe+Daqr/2ABENB+G837NjcKkCJG3LwuOh
mP41F4XQpxW4oZ+WuktLrqQKTZzBDQaihz8RIy3BHYJQ/Sb3zrlc/IYyFrg+Rh325I5iLTKuVcpe
msOp3lVXUh18+9sPYEHIuqa1Bb1amZ1k+1cCSp+PE0qvOmbZohkxPqP6mMQG9iQmAizFIN1Ae+Sf
QNESimngpdskhJLQoQpNAnMR8sW3N1CDDPS8T1Sua9x5xHtWeJDgTExxxfdIuNgUtS5b0WxNZ2ye
O0V5teohkfb6PdzuuZnrCNWSUYHmpbF7dWVxv2qMlRhnSwTr/OAlOxFwK/KPOskp8fmXLLDL3W1w
YJG1buVNWLIpErNk+8ntgYPBo0U2bWYluz3xYVybn9wb+WtrZiSLTcBukj9r4RBxjLtOrtHThdN5
BfY1c9po4iGk/hqrra+jcCj9B2T8ZzNvi1gOfZ94c0Q/08w9Wz27fNTd7aORIJBp1diYdaOBNV5n
iyJEBrxFvemVLaWMhkIZlcChdgSHLWqOaNeiuKMkNJr5KVudhI52XlvraobX3LxvD3d1F2xSiFUc
bFHhSpE6bHo5bR17JE1jy1K/hXXuztuT/laPW/TXaQ+DaFllidnU7mcZTsnnM3KZfSIFTTcpikLM
TDfQ0zy4qb9+9wKMLG/IfYyL0iGTB4KFFBl6cM7WLjN5kjdDLQ6P/H13DPmEWEy0k3QdivhLzl7q
QeX8ka0y2saXkIPoMc01XWv1ep2CMVhCLAmO0pGCyjPNlDd0sSUH1sAx0Wk9b5YgF5qAnt3eOyaB
65PVAdWLw6JRZoSRCt8kbllrGjn15U32hDlMATtiYffrVHDOO+V06eOkT49RsYsoeuNR87n7plcY
ydhGm+tEZrxruybHRIhBs7lPIhMR9tuehmU7CjiHEOSMDnaaX5mie2EYlIj38xTz1guc6k0fg0hb
MaPko1o7sgawXjGlF4XklrChFLNWLRGHP6DIElQKrsK7OkjjYRnazKhq6tIrgoESoPPL1fkUYue0
z2D0rXG/q6YBKY9SjKozD9DgQVw4gRuV2grL45t8Ifw3jA+nerG2tW+cel7Be3BN+wb2T/4+8fLr
ovR/xFYUGydgcD2QexpkmiBM9L2Xj0pkrIpPQEH5yNV3QhV/2TT7hxzrLxWaf5KFAPvwpJ+PKBqr
R3WSTw5wGJfM2bc/gytc4Ed8XBXGSMXktWEUY6VlmJZZ2Z1VQEb37dyfU+S46kLncLtgTWLeK8MA
DadlBXgrq8zIVce1BjWCc/UIlqoPKjZRDPo6jvJT0MIxclj0p7bH3rXeNjKyJhDFNXnBjg/7iHcH
zEKBsiu325HZ4T8+kFES7sW2u2hHvWCBlVjH7TF+kAdXJcTCkEAFNvT9WXx4nOrgBwrVYpqBgHfL
d7OvaH5ukWqLN5qJsyf7r6wsBIYmAB5mZotqACsCHcQYuD43XF7Mh/pTBR5S/FjETg7NRMoY9NhV
dTgYDvQQZAIXF1Cqm1YXbrqZnnDoEBbEXd54xBsQfuAfuFbLIr0HgHooMrsislZPAY+BIoGBBAWc
Bc+BBKeJSYLxMrT20FBhcVyvNXIGyhoEFyyE7RK1vlffmBy/1lkkRpCgk4bEXEiJE16u6W8J0WFF
XeZStlWCOedgsZLNe5m8poM0kxEouqnZ4ep31ovBst5ZWdsNzL7oFDBOMnhL+bFhUnWYWPOZfp+Z
N0L8YbyvlT/ijgybwBmr35+BijKXXW2kcFcRQN/y7qCaSHWqe+C85EZg1ZOjTk8X6DKq8EzdmHBx
jKhxPaAPmF/esRFohSWJ5sXllVZ4rdzjvxGdSDpjREso1Ex3oKwcZXSpFYuvIe/zgv4QJ4Oy/jUh
6bPUMNOgJYxQ1MCt1vgZu0JQ8eDCbjgVd6ZdirDBtGTdlA83TdHu5NAInox78jZbfTc8u42RMNx2
aQMuIARzuw90M1MHwIPYqRS/qx67MqrYqm+RBHXAw4fatSb+2dkH2c7CUPsQaxTD4n88ln+GQrsg
P1i9kywDGWOs+SRFHNtRHkYXwKGKEQUITJBgsI0JZcydEIvuJ7tbLnvksTFm99HEwHcy9avH1/Dz
5+qMYWVVic6E72IPEUrm//olhZcQjo8ic+rTEkDAj4P2nDMc/DbNTwX7jVhfabVE8ifPwwQ/KWLf
ItKiUnLszH6PZZlZ/X8pO/rGyV2bE+EHjFL7T3ZXLB+hLvS0CMyyomi3KPdczXK4LBm0Leu/Y7n0
yk9qPC2DxInRWTiIuDiVbudysUOk5KDlTKjqKzCnhqOzWoUyx9LiqCiviEb62aiKj8/zQs5N3uj0
lUuJOc6H7NWyJlfJw3sRBZTL3P057tH3Pg01gFGNe0e0WJFe9pJQBxk0eynpW1d00BlyBAOKMTsY
adY6EE2mne5ttMvJia40EwPZDPnDXZp2he7vWkHYO5r5lZCEt8vRtCBkOk48dEv6FhIpM2BquVRB
QhRnjjABk5HiESC755f8bD+bzdEorBGUuCxCM2zgx26iEPpRkeD2vXc7WbqvxVU2VYM77iAjnvBp
/p0pvt4cHPmH6flKxoGJw2ggWEWPnbgBMkXosxM8S5w3aVFHzNXsc9BEoTxwQn6I0s8lrg6Dter0
pVysAW6EcSoGnK9H3qEo49EjNGm03X1tmfH+u5hrEq+Ajq2DdQTFjxrKj0cu16R0wZ5o5AFvmcAH
uGud5VS/puqbl9wILiPsZht18ry8V34Jqvu+CJ0RM75JAXNGKSco0rWN4DgJYSgE9h7EDGdJSJoG
ZsyvZ6Jy29CQD1XnjjIRgFrS+YoDQxy0SnNELd2UjVOuMvGN/TaEKSH8JC6ptYJ5CZvn4oP3ZOEF
mjDPoAygL//ecKV3eO0h4GNtwkCpdnl5sFjXYSfkBavlO+dOZxVxJTWZoF142wPXjH9DAmh+4kla
zPaa797PEnDurIelchpwK1cERKDjPMsO57dblZSTUJT3JBuSM/g+/1eGno0jdog9DfWMNRRLAlW3
ASB6Mnpu35ha5+tRpREgE3xAJoTVhELAVDf1zBKROAmBM4HqDscJpmqzx0ekGO/NSd/wH+gaVyi2
TlLWY9juDwTyDIu7z3SrQ0F6zQCoZmjgQzedjuqgIdfG7XhMRGeYyJ8Az3HoZBQSh/XAADXj1qW7
VecVvk2V0Uw4EIBFqVPXb32qfj0z4Ox30cmg/EeHdFwC7LIIJ0RZu0f3DLU/NVud2L5kUbNSWmtS
4Kg+CFuiFcp3P3AdLf7OtLcP4JzoX1PZCp/fPhgAgMm8x0h23s857jfCZAI7eb51t+fjjuQGVXVm
GaDjhYbDHORPPd47oe4zlxwBEaJhSOh70NF1azZS+2+Ty2+0Gm9ywLAediz/xXTkN/7Idq4s2fo7
KwLP/Nl+wMMnPCUcgq3DDoycswu+IwOWRQNfpydZIK8hPOozn+qVTBfWlHMcsMFVYR8YN2JALPMY
zY6ANsdNA+hrHnUPOBYkYr9+5iiGs/oXW8zmTOBH9jVpHtc4AyrcpplyoD8iFej6a1N470Qpc3pg
m8RP2McO+NHFhKrNBK8Ldpv33HVHLMQz74a+QkYCpo+GajQKfT4XOV7EeQUjOh6UAPSIL3OBv8FJ
TtAdSJJLZ4i2lU/PVkPMxd8e8TjlUb/Hb8h0jqplHXoUl4SMRuacOluzSULXNpEaLW/Xq0uXa7Th
pc/fB/eGCxSaxjBVxszJwP6vSsulUFxNFIFW5faMEFnLO8QKjIL9QPG/PRnT9VosX/MHaXDQNYGO
LqE0ul9xBkwHlCqGxXFrEXCDpQQQPfpv5PT+sLq+u0lCcfIo/ekPklWwLy4hEcqIHUlh+6HjNVGi
M/qzVWNaWPhoC/MXqxr3RpOo+uxy/RAZhUx234ycos1lT1qutBhtgHbSDt4gJKd6lSqkEHQ3iIFr
ej7kCe39i9L0K+u2ioSIhCPl0IRvEsdHycm8ynKgfRixJyCqk4NNRSA9T1AzdtdcB/MLnvmVCUI2
MsmqTuiIRLDZFrpCa/vHTmlPVqRw2tp3VEEiAHYVXeHIQmCHUIX7MafIdn9AgZZPEXZmOpqPo0Vr
SNv9yIpy+8Ntk6Lo2I2y8f1Fkq77H40V7LNt9XlVGkY8K7PcjBCw6hSQORy1Dm7u7sJa+skHrsD3
c53Z+5VrEo3bWrVhDhcfIdCYfmdWmrpVapWp8YUN/y6ma+R3dWWnmzhX0iaAWmnBH2O7cbafrk+l
9owQoBgi2v1kZynZvKM9+30Wj3P6XsEymC0j3um/bPe6ql2cFqx0I7q0WINQ+/HqCvH1qT7CjApm
8nnU3iPE4U5zzi+qB3ygAymO6VgErD42UGVPEEGU+D88JTYLCIrWgAjLyYFeNAE4c6hsTCndI6p0
24iXGuAdjs1ohgoImlEIUuroF6aYWlOgCWnj4BCMvcVVCVT0KvXJHF8k/7uPMgdS9SS03yv2AGAT
lBTYrZl7oDpYuCnLuo/EqPUjpczylB1+aDIHVeh/Us+lBKgliFPy4QofenHlnSfwodHqRtdAiIX1
mx+HOmESOvNZ9n/r4DLH1r5tk1SvV+zkDWTkmfTb3rNHK3HtnhCOQkx33sjnMB6ZgsZEiY1R+IMX
fG2l/EY7ia4Nkaofm5bW01bNFp8hkCtilxVQLDZZjOAaBnF86KcmloC/Ech+expp7ntHLg6ORorW
gGyiXO3I3m1giX3Bmg8WE2yQxxGi5VYn15TYS8GPWNDKxQP9NrmE9m1v9VSSF3CAAqrbxiNpcB9y
65cCr8LuCase0yCVd0qE2LiN/PpLnxHzaXNhl3JlJoIoiXIghMSwst/Z3BRr/wX2zZjqFGSPrUfr
4v3sIXzanqYhZvzKBIdja7PTzkZDI/YsaipDRgvuN5aMOatpeZip2EKdTzEEY0LrKkBiETO8NAja
2jIS+PtNgBgYuhBLvoWuau8E4WTz1INUl1nGoZ5ZyIKj1Cqa/b7i/NNmwEIigxoxcdqBvRRTcYav
F1WBn4TbzwlMF17aD36r269167ZtSlIysBFejYjLzSkwtP6LNpMU8vgQ6hibhwZN9920dhUyVBAo
ueEFyQXQ94x7YR4C8Ouohi7y5kA3vzAVsHvupWr84NIXUKFZwZDvvRZ0T8b+xhRag7NaSxsBoUip
KrScNjvauA2zR9U/DY2yG8bhG8cjL5YfcFaGbBCu5ByVSUuphgGCyz/9rUg9FwSWTL3gxHVhZ2ab
3ghMHRHJZTPcJhRecPDYnwIEcZIi3E2tNgAtpPeZXJfo7Bi04tqUV+3PLyto5qtGs7an6KvM7n4Q
DYNyUVB5PGPY7C57vcmF1DTv8RpBntiPp1L6ZOJAXUAlbMd77mY6pc2AzACpqC/FgHkCjcBCnJ67
ux7XCUEfNiAiXzWbnhuPE1X9emCVC/JKCk6ud9rboItufE3s/jngoQsIfH2TTLzcNefqDKQoAXJB
z8AGLzvTq6Hb+7XbsN+kFqbzE/QERS2Yf+aHOedsoZVmwJh0wiR665Zh20PRtns1S9PmUDWPhXe+
lrFd9HFxe4oyYYVeC9UXgGp6O2vq0YyZ3DMgeVEoZZb3n6dU5BhiMS7uTnQuw65P2tgBinHAKJsO
FAsJGXGvuDtzROm8F8hHrPahvLj17psO33NZgqPp8SlGQpgFRBrFdMn9UkCh0eT1Cl0PxhbWIiIj
a3+69L5bDZKOUJP8yQXPIUQLtL4wj0YdPiIbaTqkC+aaJRAw8b7AJXfeTVnS2b71bzLmskTkWP0e
mqkfCFzpxUOYOxCfHjyCmbr3ozEg50UPCgUDxo6R7gvSvj/iHH95RLQqWAWftfb0h5vQ2YM9opL+
+REiBf0Oby6xUOBkBSm7kLyqe3Xq3JaOHZJr7CVtwF2G8v2vgZPB7rXRPiwKXTGKmIsIti66e2Be
ERUy6wlUFUBoVhbJbA806Hp+ghBYqZS/+p1dtJYlbbPk85+pYWESKMvUdUJEqZ79fAbOOHQ7BO4t
At483RDulRdNlQVKil7+H8+6W3vSS4e7GDVkJLz8jpn8OIBZS2LOMj4NMbUEmFwMzpU42sbcV6MP
SYJ6OfkpBc27UzaBgptZ4M6f09d8u7OBSR7cAysy80E5Da3mF0m+2q3jrSIR294EZ7YoYpa5IXyr
4AzVOtwCIASv1CgjH1xqH+GutV7mr3MCs1lhrW5HLQmU75TzivfoLuXQ9prMjN7nnKA9Z09z4Ctd
aAulVnPrbTtVMR7+yBZdgpxoTAxJ6l7Hy/lyXOkFAWjQA3iuUMVc8ZeC9P8cf4qpoRn5oUAZZ8d8
/9wT/nb/swYRjRia+spTdwoAwMvW9bEcVyoFdKahYBUtjRLUjmULDwuHiE3Wdh9L7Y65AK1YaFUJ
8BcgfC+8baK3aaWFoaU1DZVR92U9hj4iObJlSVDlYuev2JWLgigZmmIZbJrN/elc/Z82wJ9tfFS8
QT3vG0ZAYShagLvT86i5m1OTM+BSqEN5sh3A2TpP9Trvw7U/RW98aNuEv7A6R4YWBb79oo1OcHB9
guyiYOrbE0hxb5RbjeEHPupldG7f0rK5qkSZtlHNPTdddx+D1ZzDasaRKk5zs1vjqHFxoVD1ovDJ
91QQbX3afG7viqJ2Cxo83CP0KUglskg7d75ZC0gHn9LLSUMi963njberaYW749hntFypbW64QLZR
n6cn0NwoKWIbY9lu/EMu5Uf9T2yskHYUil+ZYw1KRwivQ2Lq0cKAd3BWa8TSKXNhDsO82U0EXyKd
15rkpakB8YCfpJoKQa7fwJQyKsBlWyE3Ba9GvZw59pc5NMMF4u/K9A6Iulm1/nKvrBmeVqw043OQ
yhtAsR3JNVLAsfIeAi9dfxfSSPUROA9OP6dEiGJ05l8yd2NuZiS/8DWN21AYeTyMAwkqY9929GfQ
eWS4dzH+/TUBoBzTtT/IOJYaNeIn7zWsn5ejzX3I00U7DwnOlzSaKeZeNbbUxgjFc5n6g5/x7cDj
CNrx5JbC8D4p2AzRV5B4cKh68VdKUTw5nx350zo4Bxi/7it4Z9R9ktGgqpka84Ke5pSdQS6WavOj
PfqNvGjDELt2KmTL7XeKrkZVtfAULWD+u9y4xr4C3290x9TQzr6sgPlfScMlWgBc4ONxg4JfwRHl
7UBf2AMOFj0wfiHcQILsVeFzaffeSaAmRbXx4/9EDSmr2tS0cqHSsPz89mR8bWT1WTNUh7uhBcAQ
4dIR370CI2aIMEnhmkabzKfo0u8f18tTS8ymt2ECgL9VvxTf5iOhXAdTA+HChdo5AqroCfycLDyf
lV2zkSjBWJqVh7EkHiL8nZAUOX/R5kKeXIpH6QBCfIs2VnmHeUb5jSCqqdShIwVIGFLrikFsni1g
mmom1/GA7hRaRncd1ZDrL3FBApsgIJF3G67OQn410vGEORulXi21bO9SaLUAcV2AsJRCNTmFC0wU
sA9CJgekIKYDNLHIDzvHSPJsXnYqgTRsbKyL2LHQADcFGhnL5/3C9bqxnHYAL3MlARvvF4Wnvbi/
O/VLjA58d+tt13iwceYWZ/AzcgKsvz9XuVQm5zucSeZaMBrclwPEiwNdCLGk4K3QtNgAIaFUaf8A
K8PdLvGoD8Jf9XilgNfIMT9BMhnfAhQ7mRoWLFG7EggtJWt1mspsJwW2Udb2MKIOhRrpISPILmkH
qtIxfKWk0v4lOmJEsN7YugIyrveNSl4bMaHn1Pi4ySW9RlKDAO8Ip5z414aRu8iXs1EOSfcwdzKV
tk1UIRa5zZEbhMjMCxE0cV3ypWQJLLxeob3Qx7qhyQe0kl4vhBwxVGgkZNFZA9wo+fVpJKyMiS0W
EN61bpxAIm19h+2sAYynZ+oESJHD50X1HbvpjFNZC7elkQV8DSUOQdyUdvjhWrupR58br/3oYBEd
gAHJFX7WblBAlRSuSfUVCBsJLRpeig60R/nTzNpaYwYufaG6rdSDXClNBhcrXPHaJkqJbSkaNI6a
5KOLA/Gbl7/ppAc+PI9kgc1mvmH54PlYV2AZBRLJCo45tgiezrnrS78ZDADefdd/nGkZH0jkNThE
hCM4ONGJeG9YWmK2FkrHat7SL6e8XQQ5nbGKWV5C5VYK9p5XM7ouIeeJ3ied3C8RmLZ2SX7Sg9zE
tWn8oETTqTzLGBt+C9SzsrU0AU+I5xsUl7VQPcyRA3mPNjhpf+WkFKnw7XXIMyI7lQaWFpK0xxqK
rgijDX3D5+SuUHTp+M8ZpxYFnJcSsXxBBdeMGAbmSPmoOJ/z63AuqZ2NBdIVC+1i3teSP3EOw+BA
ND0OLFwiSfUR59rJXxrYo3/lYySd3tMPgDlioaGBiaD8QEe0l2JkoCSk8FqtP5KR8pxGQ8zZqjbl
JfToO2QCHicp6LiPXQrxHQH6QywjujpUx2xvszFUuFz/885I3Fec5Y7OMsfhaQQ8M8GtitIET37W
fOTmxe+QeSRlM1hkMblkgAxrJ/tjzp72EzWKYxogAXdpzWXtKJ38/y6rMwRHqf/+i+rQiCOU1nJ7
CrGxXhvhWJze8PXlTdKWdlWh7AZBkFuiGO/nCGab7WLI3rYdzcsEoxl4/TBPJcvyLC+bbrgF8gby
tSrlFdvrE8m+FPbEUbXQI6pssNHJZsWQwwrQsytwiWBdhy467ZiaAgBWd9c9kQ0T5gWRxj1Vztzi
aq+Ns0KgO4gtKKPekoE4ZKZRGTGiwy+DZ7wBpq37Q3NnqPccvw3TdmISPBI8QUd4G/7Y7s8LPUtA
rrhlqNA30ClvjlDyyJQpdqoyMN222hU5nfVcXD/XFrSSuqyQvVECKBLFpaDrW6I3djBSvFJrWUE7
hmkYrv6r3VHA62Rc63DmODrDuyjgi2P7XSvm2qIr6K5UewzQ6TbqgfkR2gxeXp99FN61gbxa9qZG
416Ch1jKuCbE1t93sO2YGCv/Ir925qfWB1K1S2+SM7ICChkikZDO/eKHRuge8bVI3KGqZfQvWth8
eBbS/yeoT03CYS1hLtdE7LanbxU6QoRfV1qQpWag4zqgEdTVxh64tcjsMcnz+JeACVw0Yiq0dTM+
xiAkG8arTm4lU2hNpSkaw+HN/xPnXeaqxoyN/elVTKrJoBDcO9nvZ/HsCy9ru+LbqeJ8shPXhJC3
4Pv2JKJb5ElVr/7CsXL0nE2llWO48nILPbs0gLQOVZuWsDnkZKTaEZpS6oJCi2AZqSSm+HcHzFPs
5ZozyfKIDNql9qIRNZqDxnOXn5/2aduroIhSUE16iMe9xBAiW19x0OxvEkX4A3Sp78je3l507Aqe
QL4sjpVQMsVoKjlNZbg0yU9hXlb5LIy+nSUy1ze3x0Akl0PbsTMuJSh6+xjmu5KgPAR7urRCXBnE
iSP3011qp8WRRN7vGnRH/TqajJWVD5xIr1FmZQqSjOEFPfMp5NoH+wDNXZP21FMBImKffl6EienO
XmrSYZpmnyIb8AKSxX+Nq62GWYb6vTraJio9jzBNqL17UD2RdqzCQ80D3u4wsIRH4RLdnan1GMcx
Nx4/hFey+53x2Qs9ReRkOySQ1m20J5Q+RgZfxOWa32AiBt9/KcHA1gPSSJNCKk29zFnDvly1vBc/
rirLAPytNw1jrYYZDloIUv01dG5k5BKIBb5l3nYhRCwMBximKVWG9W+tgLbFfdD2Ffudq9306FD/
AiG6c7kH6YtflO0tdHJO1HBoE4EbzfDAHomUG2DVxoRjDggiAkmdx+uCGRzpWSqNqdbOm2ozqA6Q
UecGHI6psbOtxxgjUJG8EWQFBIY1ElZmlTdEPyFTpY/KhtMnDEwjXNar7762sVv+uqYKPu46WXgm
sl6D8lXHsGE1kC7/kdRmjUvQ06rtbUveWsUQX4+DQl7n81vWNj/LVzpg8svMetJbukfHHqN9btMx
iNqVPknOcviOs51NHFG4t3ooW1EXKau4cSDcQX0DfezsFhFp39RVixaOEeU4maxlUiARwI/FcKr0
Elux1cPRUW0tX09nIAXdgaR4uDLQDEFUged+5EKI/LZEzooupZRhIs74TFlnUTa3Qng9uFpafFpD
BNoH3tOYzrhqogs1UhJmwBpITnQ4urY9vJeOqcS3uwI9l4VIcYlqFUQVyl7IuYyveTsGLscaXzRd
fQ6g4tQIxaNXsagdeLlIeRw9ZlWcx64QVkbTDOdmvh9YkfNzI19io3Unwk2SxYeMJL6rrRONwPZo
cVORBkYOHjfzePuyR/veUNExqBU9y6Oh8csZUUvFIOtu9FgaVwWskB16y8tUb0z+DWYLo5K1O/IV
GXes2JCNvR3NAiFnLEl1bXIbFSaI3VEYNigqvTohdz3DSI8BADSBOmp9duyicymc1Egok5OPoCTW
zDLgjBq2jmi1Pg3CT9ZW3ZQ+waDbE8OlzoCDosV0x691NeCwu1sst2llJHrUZNwInsTBPxnVZi24
vLpl/YVTnwQBwhGRqaKpM1zk3c3yeB2DgfX3t88yFSfQe6Yl7L19vkF1zYm9t1KZs27VJfQtGMty
gaxrLQF7dHBKMmmM27ocaNCdQ7dNkjGRZdxYZeIs/0Brc4N3v+ESimGBATwMW++vmlPJDFztVK5V
7KfuKPLgjB5TTJ/e5xkPD5T6poRPklVFoE670x03/kyFHXvoKMPvMjyzWEonAdciGPe5l8yXAz2M
nycHolnHpiTOJh7PgtKymDH3ic/d0HoyBzM33wr7neX2lGBoElOTzcN3xIfsl3fgaBKsHso3rl5M
AKvkkbDhGQKrrIZOlG9Cw4EuHzYQ2zeitKmTbwC21LLiX8wdF8ZI9JOb4ERjThqTgtNrPHn7lifz
3JvKyRH9FPZrIhVbWVk1gvUknJhmC79SnCV6cTwnLqV0E4o+FFDePP81PC6gDdq5SQZVkPKfUBTE
axMzS7LuKl5ZxyBnpnlO93YwliFtTNtp388fN+fjLYzphyb+hHQJ83HJxdVxShXkiHOL1MkZYcOF
uLUwcFvT+W4qqnDUu0eG+HBcyIs2xzIhbnElSqMjrZmcNu/IT3YxbT9qV2GJT8pmMOsi8yCUhBu5
bVeGR3wBCSCNT3yYYjhj0EH+98xWBR1K46RsF16ie+S1T3b6K3oCAkwmCyxqU41qe8AuuNsC2mYW
hvHyeQRJM85z6wiymu2FjdXiE//VfL9cat86x3y0NsLsCbeuD2DSRS1M7NY4IZiY9mFnWSRIcc/C
2sewWV9FSHAynZOeAyogdGgG4/pzriURM/74WqUGgwJGNoM106xM6jyGOzKH6g/CFisW1KmKOWwy
XB+hJpw5g/5hBuD2/Jf/N70p/QOpvshH5xMxBkCGloeoi92XzPUOXHJXBRlSrojF5ARy54uScjx6
uueKULHXrwkj2jgUTjAehiH6vhkoKSYOuFdd7qxb2T5r3/ujcbERV2wXco1lLB33y9l34/lqP0mH
n/LElQLryfOuuSDErSFGMMwtkCJeNkUubjx91UDjkm8hwflBGnb4/k3XbqHxfCVTjRxyy+vMjDkY
896gQ/mEIq/mPqbSsPyePSk45Jt11CIQIaKKhjfCjKoM8QqcBrcfGT6kh4grzEURsS0baHFtUBL0
sbKVHYhzEkelFYUe7id3rhTg0SNDAjS1taL8vAIaMtFAaVVd1ifMjD+fxx9T88Bp1178rU3JIdZM
e6Q1LVh/rX7QPrYYQ6PNCwCsTl9YWK0KVxaOT5ftTMDFhVnpLUWjMwBpiZTOk7ddWlkTYNS9zjzS
mDMyMVWFpU2cS2s+DSiqMqMWhUa4PPBMj91lnVlwkrJOeLOqI5V4PT5pTui/4uGlHUhSJuELkkUd
reTF7Poql8owCRnWfj7qHejblBK1SHgAFyzP+7hSTM7rhEFpLvV2a66PNj6mUFh+8BKFiEt7KOwV
o0bQHjj7OWbtfGjwp7Z81KL4yhxncYdJn+h0rXktMBl8eFIJmyDmKQQbsN1/GWQMkEFWTJ264JFJ
xCoQVqZvm0CtDIVQ5TiASeg51NlkdcijG2wREWAauAzE5r4nb7IgKmzbNniFd0uaKesJYerzfTem
d8ODxx6mNhMOG+u3EbS9ylOZSgu24Vj6Ewx+JPCHkC4wrwWFaaReZ9hMX9kDEtw1hn1npICiB65E
5muhh4fVVsftTmXGnchDkfNVLxkaPX4WEIl2DkfhY9D8d+cWdu0EUTIQ65mRagLuPdUWvy0Tt7nI
f60ahd38+Tt4fUkfBIljwpI+e2WaM7oPnaGK58Dz4kJBZs5uSkEaOmg/DrwblPKnGK32FtC4u5Pg
NxrlmG12uDasLqR4AAAqe9J5e97ITeorXRPUr7gN06d43pyTZzUqTGCooiuEafLrVzPkLSw+9bg+
GoTtmOfUKPmuXVy206orlIdPb/6fvs4Fv2/Uw/SVcy0NlG9acT6YVESQ84qN1/THH4YfmimLPK81
B62pHbAd4+LndzAa1Ob2ZSIHeUf+UwNaqmn/RRYEPU9TW3RJ7Z6BIXV91rGKYzhbG99KE0UNsauZ
Y3y2eNjHN7/d8d2pKa4NTj3eD+7mua8PepV4AqKNCTBaDThp9/UqixMxsByOHNwNyT83wCk50Q5c
JSjfiA3g/IHleC1VJURbGULvJjscIOTaSSxJ3Q+6CBrBpRiErQOX0hrCvFgzxjJY748WHu1cot0R
CxQSHxTF3HKoOE9zosSlzrcAc93KgMEmn8Bz/AswmJF94exbwaa/wiPKx7+J9Zjobj+xp5iANHCT
5CWUs+dAzli5Mkx/q7zLcAh0CY+s66F/CeLf/WhjGutV/3RaIxqvYeYw73I8m4p1RSB5ZuZB9lAc
dk2gZLXXKNotDMk3f1avXkntPFssnNKCBTcnR/tB8h4j9vwCuScYHiut/c/E9dW6TqC5bz9QQDV7
1cPuU6zQLvgiLwiPKsS9R15gP2kbPRLP+yUYShFqJRsCnIPuFtUSN9a7bIPGMA5EwagRUNjUQCV7
gBeq9/0ySzWv7hpBr4mgh7gR/eZVgt0jrrBSa5p6ywIk2ezATin6pNZivIxwz5EY0y9dZp/NAA84
ni6roCD9BwQ1muoKsE4xqpghLy8CrtHlx4plyRPGY/X+CvrWAyna9yBdJOStYW4oPcwgkJP2zkmD
8KggMBJ1aAYettcJl/wAd7dkLlo4HBP/OEYYGo4j9Uw84vTCIpGJqxi/JrsWv8kQCUbUN0PcMHRu
o9bdguzEgssJ4BktDxdOL5Jl6qauPOooU8MFHCi5mogaizsN+YsB7OsNQq3uGdRQ5X/mHtXVtqfn
J1trwhX/6VLybJerQQSEEl/Y22/cIijL6m7O66QQtMvWM9PkmLzESft4wfZIUps4RtkaynyiME4O
TKIQTleZe5+igDevXK5/yd7IiGGeDHy1nBJiJtSBrWfl5wskyeHPs/OoKdw2Xsq5WQtl7sDC+PRx
drfARUsLwyNwzBJXsjihVXMQ2xbobA8xLerkBsMALl6NcfBO8VxdUqoUF87pbIYIerAhExV8ebhW
+2kpB/mCPOEFCh4JV++HOb36cPzCFbJK4IbxlIQHJi0ZZXUIwxWJPDOuG90jtLx1dMWyJCLbeS8A
QWhtTvVOCMh49RledXeMXKRM6C4sSTX3PpOECS13JVU5MnZasLJYuhjs0TzJPr/qbQHB3FiUdcsX
HlnPMIaCUt8CqdAuLscA/cpOzvV5egRCQ4NtgUDGPQeva4fb++/llPuDDk4gKbLYoRZs/TrHyf7p
17j0ds83Q4MzqcpUjS5LM0nITIRS6EkbHvFm6tB3tIYKW6lTe9oRxMfw/3zv8e3TLWIrZf/dXbQp
UKkoZdb0AG307U2+AKGna0G+VuqqHIEOVfWJ+rzOF2nHAyHvJax3VD7czHWc/RCREmz3bQW+lFZ9
l2k9bnxRHuK51/BfZEciEObnLAcHDI2+E2USQ0j+oMRXCajrpF84Wwh9qEshnkODGMnkTLJlS/h7
DFG4NgbvcNSKehv3f9pV/gl1h2lBQ2mc1klWoD9eGg8Y1iCV/+dnz5xQmRpOVTE7Ps0tHbU3lbLn
6uvFWepLaCUzJHXHJyAMEoHgk31AqmadsjY17RIAwLouo2F6JuGrnITWw7W37nxGnc2oSmiLFcXf
AKDcKBagUy+IxMUJTBnbdagLhcxIjyxwHaoH0vzBLoNBccyhV28bnxPUxzKxOxqYWoZZnUFpq2KA
jUmBy1ogEZPSvnXEvrSLe9NDIvjn7TrRGldA9gfvIxglH7jdStxF4JpTXijRP5jQQ9MbxTUQjxg8
kG7SmAIgcYHXu6wOf9A0wSQ+JECZBaFe+AMLBRT6zoCz4rPuYij0uxjFwghYMM6eeyhngjMdFIq9
vgu/i36FIucwS+GtdN22RutGVGfyU/ZxQqNgFjGxo9gUawj1zJ50Ipr8ZMRYHRdAOPmWwVvJ98dK
X6Ll97W64hl/psWeljjl7wpL5CA+p5YQDJX+s2+LzEUmiOp/nmm++2RrIjohJtLL/QlNpcEkzkbm
709UhQJjUnMHVuyvsWfMetB8fAgG0S1zXXwgwHmNdAsZhyYGsky1i7LYMB8RlTrjOr5dk1CeCJcY
EEohE0NgfTsMrR1DcR4RAgdfnLCqdzG/mrV74qnx3Ewx0qXMnL+/t8U89ZLYWcfKJrIO3NkUn6hw
U+S+xoneOu5iQi9SLxNqgcmEo7gMTmQ9I1WIhsio4ocv90AjhUi01er0hE22VpCgR1HAWlyNlxzL
MyxDuyM8XOkof3ChSYE5HL+mhzzc1Ma4Ie6Rye633I1Av9KKYA99mCF346kkREMM0+SaHKKpqyed
n8oo9Zmnq3/NFYNxW2T9EuDgNNK9wph3dTfeqdFuzQ2inp6KZk4DH7SEwwdplFOR6vzUSElTM2hd
buapoPqx+kDrLpezX9yDz/RIJmO2o5LPX9im+JgxGMIEXxCYMGZvRjQmkuzOojcdWKyjcqcvUMvJ
OuZDPCYTQw9Zty18erBon9IqH/XMdBJ+c/PkN1JWw0hxPQre10MpJ8w7ioexODUik5AMNdn88Mof
xQfQ9L5pP2GXd5rdbg2sJrlDTIJPyqN4Xmyy4qHTA7QpQQq0FU4kda8CIVdH8AETkdo2Y4XfbUsH
V1EjhQnMgMu+dJyXYU8mcRmiegUfqddjBL1a7lJhu+I+1kuJQgq0z+D8yxOX+pOhYIltaybAFQfy
Dhoxx+CCcJlck7UoY4pIVJyWHAz89RNM3g+35SGNk3S7tSOYmnsX0fCeGHDD4aIiSsmNbQ3eGxF5
Sm9rmInN3AwgFe7IDV+ReH4cvc1w9ZgoeO+tMLUJxC8wNuTSQQ50x8DxWlBC396wbDZnel+UkfO+
yeUO6lu0wKlsH7KuMuWE3UO66SKyM55OLdBERNy1asrqBZXA+ZALfxRIwil16MOnoZTWolrbj85s
lYj2vYALcyjTHzh/T0r8PiVc4HEGUc3lRPBrCIizdG7Cqt7JukDYUP15kAW3NMdJHwzaA0vPHiVX
MPvEFWJ8xKgeF909zj3hgStzG6k4pzlh63tAHOCAgXwIQ2ykloRYE0C3vnYs5qyMDkcWKNBK21aI
HjTM7/MduYBXhE/7lovkkI2wT9E0hAvYxXvVRQdfVocdk5krgT3I/DwCksQV8TB4d8IBKMeHLUf2
cxlzciOlv3ww5v+0arGlUASkpD3xMERiNW98vzcnXwMtLVCdOqJF2v+voJQhk36ayTYKQlhB9nii
VLyUPb5q984ptAQS/OsNF2eRWAiUjzidWcYAY5UrER40PPemcQXCQBylqGmN0JTIDgMO+sZ/6Pbt
R1DQt8UrK4z+4pDnIZAcHhD8ZTiBIjglIso17Iy5NdigWIwyPD8pbx7vWjX7TYtZAERsrx1cJvYp
7xtPF4HyNpdmd9rg/lzqbS2/xzCJvCQ18ztjIYxPOmqH6S3oNSE8dq9mNDf5z4xhV4f2ajoskDrR
mzDlyd1TXPSqK6gF26nmcjOC8yANCrmstWc0fOC9xnba+FNTUK0kt7YFxYv3Xxsme0t0QI3exDV9
C/2ocegKvRVyKqNznsWfb8KLX+wK2o3p2jaxnycNBS6s/hFDkJntpb544DwHriRaYqm5diqT5M6v
222mzkTtaDHqIGvg/essCQJ9doG0FzwTGJxo3dth4FAJ/jghxL1Nzdo0oECKimxx7JKT4HA3tPPZ
8N2RQbZzbHQTqeBUmau8/uXgGaPfxNVv/7nfQRGRCTMDrVdd7a+mjMjgst9tXJ054qbM76V+kccX
CtZKBK0mG30CmSE/ktBDiIqIpmLDKzXGfHfGyp+dyvTku7i4kpxzqq+WhnmDjOPjXp7OXilELbrL
H4l/971Y2iCYTosNM54XYOQn5Pb4a66CEjABTqD0PnncE5wQEemXO4DEojPxvPYkVM7TMud9hBsJ
vkYiIi8nowTZmjNhlbV7fqYKewTCB8znv/zH2OQv4z9H/RgpCdKex5XfPWWOAuGDZs5fIqQ/enA7
tRels7j1cB21e3gFrBBGzRQZC+yktUaK+8jCQl0aW8vRK1uw3DZCGPMyGHXLsQx0QEa9U2LYbCrw
uJ2Mf8pZPWTp9TSepahT5vZe8khvhbBtUgjf04RSwZPZ+mLQYrBUAbrPv0CDO75kWLbC61fmqaWm
MxW6w6oXjfob7Qyc6RSPooa5WgVIzutTDYOMCDM2B2vYxL2p0WOnnY7YAFBMmSdpNe3zfjjkiMuP
83sXcJBwgz1Fsmb9Aij0UD0VDInTrjyQnYUadDcHzLYwhsTsqgkc+pH817B7GVScL9bQwBWHLr0A
+U/3NcfL3traHZMGbWx97x8Wj8/aMzv2GmXenXG0Hhe4sGGHAG+o548vB4F80FyuZ7F12bahdbyG
dR2FmL5sLePtH788xz+bvdluD16Q/nkdJBydalUrMOC1y3QO3DqdmnL52rsqha0v1j049PGIaeKh
/JmGmOzRiTZW+IIEcN+M//yzPgS2QvUyZR6SeBFG0V93UcI5WfZc/v687tQ3yJ1X6EtYCimTP8qn
Pnl6oxKOxNQ0tfdwm2P5zEHXk9ExHHjO0iuoB7dHp5adKmilh6bga7GxkAxmFjXgz2lf+DtPE0LA
/co31p+1wnGwdAM8TDOCKulbLhCJJMmrQqTKe9qgQ7mdwKZjISMlgEXPVQiou0C2/KEMxT69tJ+3
/Xi6PPrfFNahflu5Jpnr7mtgJMfOIEHqcxPxZFSsXROYk2m4Bit1w9LxLhgWO7ba9s9O9czSfjyw
KIWIu42Tl2CU9H55T6LbZEa2NiT7FrgIftxj8HeRL4emzcineeZkIUxz2ABe4t8fmJlmw1n7tyFs
fiKTROIeOspEmsdvjUco+cRNJh2WwLUWmEDq17YhfcEx0Pg5bUkFm9FEV0iC8mrGJDC/d3pr+X7r
eEVEJVCTSRMQXuPG6Fx3KEC+R4QBImd0DFCe96ZLMVKH/Cs+NzTC0Nnqsg4dT8HxLI/pQtb12awg
1uIthMtlPbs2yvX+I8Dbe6W33cOE/FiWkfma/HgQBDdkj7lqGdqe78VP1b7cUzlm8BEqIJDtDKqP
aFFDeUCc+0MM7/86jNbXnHvwn2iXdVoDfZWpYd4NGp/KXJV670vWYVx6ZhWlP+iQkTjx4BUMwxFo
ehDhWcQ38mLa3LMhcH6qIDLsGJheu/15r4y0ABDfGP9N6vpXi/n+/vsPmraH+IcPGuSjrIIfnVK9
LJw2kiIl7i9q/vlshMUNDEGKZ1RaO6TxhrupPI00pipXqLmDRssAR79UYOAsGUOB9+6tlMHNOFB0
jO9anocs5era+7gXjOmla54t47vnJGV+tBElL6aG9DS91NgEuTH/vjXN8oHDOKEhVDSnZypT7iBi
UEfsnjHKfL5K2dMtI+pGsDNb6Ygj9Df15riIGFg/KbG/gpkFGBNyMM/+SD5Zfkm3tUcKITo9WFT7
S1nC5FVz2eF7fDTEu98mGIpzsd9X3YoDzPrafzPJyD5IZq1/NQSLlo60y7K1Q4yTfgLtxindHvYz
9okPiYiiyMSqiWVG9MwEliKtAIfrI5S+2p0U8PJsBEXMPUP7DLo7J0l873p1YZk3ms/0DRbUjO9/
+tdmZvtCjVt+Zh1bWkbJYakuv2pIV0eUYWnj2CwL4Q1g3xpG6O6fb6OPsLOQIRuXbbjNtL2kErd9
3xgcQhKPY+alz4pNasDns5pLwfmAJDvdY6XTXnoYhti5OQAmgNAYn3wa5VcqjDGpRlBHllQXkXbR
BmjLvTLYUIEtXe9zGYT2ehhg/YJVpFXnYXhFn/vbKDeOjbeFtMqM3PaOIvehmqBogTC86wuU1UEE
GG+QepxqkQ9UbATF9zyb8zL0ba3YpeMMJePS04rGQsfUl1l0ZCb6S+Lu51Yphhe5HGiqcdx1bYjE
mgSurYofJYa2+Oh08eQRvcNMIlEz9IWrxldtrmY2+3dnMqqalcEu+ivY37yML71vWIkck6IsYYEA
Oo4CPBgBEaK+BOreKdw4Jt8tsvlUbW7F6lKpS+Vxu34TWzPSFmq3Fl5XvC1QNhaeDGcr06XFfkpF
YT6zQ7Yp51BRhyToCoAXEwtoQJ5cchdLnD954sg2BysILYZhiDQ9zsbF3vYLzdnSk+dTwBXc+nO/
1v5lieqnH5Qjq/bkeHGCk1TcoPB3/XN1I9oe1erRM7xXSv4ZtY7G07x1OY96hYLf7Iasm+4JxJzL
NBIh/m65M+KbZhifm/MYrUXRCgQR7lrCZBaaq9o7sJTI7L1f4WSsfzbKbkzmEpzJ5veiJ+0b3dQY
/utrfA/3AGtVxKCzFch9nrq3sbLv1BalsHYbM0fjI+z5cnvGj9wuyWWTb2JxfpfQmgqpXG/o8+B0
tztsfos+JChLmEVems9wHwg4+1dQ+VZ+kxR+okVZym60yB/CAO+3a1pb+tB2+Ad0zHkc3Nm6E4cu
ysJIeh7Jur03Z5Q9Wz6r6DIFeVgsLAhjXg2p6FZBWk6Oi4g475zIvy4GYE5qVgFBaWguj/FqLvWa
Df/gyvuEVXJ9BvwrAc9SzhFq8Vczdd4k4EB99jMBZU7UtzTG7uUj8KBXae5HIKo6bf6NMQmiuN6T
grE3qq4WONuj16415k0txVgslCk1flQIRdOAMDZQPXpNcapsZ+O4whITBXWngvUCL4CVi3GOp2J0
vq00xlTLOZbWEqrNHPcJNtfimL/XD9Z6WHp4EmZLe/rd0zszj8DjQrq9PbofDAPvgtFxMrhTd4pc
6ql15Z/j1o1iAS5xdK/TTRqjHvHE/g2wO+L2rhLzuPiSOjMp+UnSys6da5vKCN+yMMLHiKdpDjPg
GojmGkMO6sv/RfAPboEi7t32L5+y5OYSRE4VXk/kGShlYwosIn3t1VIwKlBj6tovNL7fdEBvQsr8
F7b/CUBvBI0doYbyn88EDF7IwVu09El8I3PK3PFek+OkUnnjIejAYvbJrzzuKV/UVgpc5gvsCQSe
odbUYT7aVAh6GufIQdRpSoh5AJpa0vvJSCx4oxV4x7xUzs7AjiUGmutfqVvbVNpjLjhxkjyhBNex
HqaRQCTz9wDLhuoRlYruerDYIVgiY3llxYfSDXs37hKRmz6S/if2uPxf31XDQaXFlfthvbrICAaf
cIDzuSlsGAKKp7Xctx7VIj7I7ZOqFFpaK7XL866eG8ZtJrg8vaKfoGevwkZSSbca0BqThaoBk1/j
208MxgQmB83q95A/Shxxv0+mqAYFuvCbSZn6E/fGAwkTj6O6pFXmceFNcMH5Lu0UDeR0GW8qxsYL
6wi71N4MAeQPsBkDopQ48S9UUCWVvNUDWfIjVzftBux6yjQVYngNGA3y3RjHvt2Dkrb8yxhYVN1Y
hmUwJilc1oZe+RXEcaTdSJeVYwA8fDRuTzKA9tEV7O7myz0x5PvS2atS2YceKGT9cqsbNn5WAL2e
CPEunTe5jmB6MZt0gIZSuWOf6E/axiy8RpFWMNbm/h2taFfHLqf2807xm0QWAJsYlDIUgnsPGbiL
L+D450AED1TZVh8biy7kfLVVcg/xVcEy4SFk4AYyXMklAqZ4R67Ia/fll+EiiKMArORvbD6EvO6q
+HxL+EWrQELaRACEP+OLY6vdN+blmmgO5AeFWlnKzdUEIAxoS2zrsAKW4bdHe2znEbylklpLT/hY
ozrIJa3atcYEN5q7SwSC7OQ7t6elqd683qRrDM43Pds+TXjf4PBL1GzVO+caLFtIFHWJwS3wOiHi
QjxWWhr0AjsMPSxbLskbBq0ybrynYapkfy2J4NJpcTTLgDtiJie0gW836Oy6sR4WL47mgbiFab+y
8jJh4lvODMxC4XtECrufpa81+UDKWp3aMgHUYx9M5dEf5vDIL0LKV3gshXVOmlrqzo9OJ34m0J8F
o6M5qreC1bZKonOM2oi8NrfQU2xEgdbaL2rht9qQGNYLmnJVSqVKP8ypVKYRqJj/FArOT/Z667D7
baV1mbOsDiUQndDzFavqlpVFFsGN3H34MDIwcOsN2f48ZNIa0qG4iUu29e4qvwgnYSGl6GRC3zAm
x41OEuC7byNdb+tqHvm/e2CeTGnQ0jA0LsQ35xEIQKrPSYhs7EsEZ6+r4lulniRs7fAcjRcXYMMF
f3VUewwzMOyaPgbFgY8mPtql3x9xmye0Z7IR023U0sGrFHlKbAX/cYnkgUGVYtRtngYr4VhfwXud
Khdgksmz8dAOZaeNypwUrq2mcaTykp8ssloXvKiyPuk27hqnpLHlEvDjm+wuiRn+mALG/Ssi0+ia
U4SuDdRo5fa9ERBkY3evbEypDzPHgSIN2vUwPgeniDpcDgMTHfzPPAKZ1BRJX7ehQAhFAZVZBxzL
TmL9Mnkx220GuNSMpFvCsSuZ8rh+ogylpsTw/TRsda1Ka6QkiehV4eIFsioF4VlkxPQQ+2ysCHA/
aylxZsLPqWGzS6YO87w8wsAEXh9G9/ZiG5ynFZFk6zIGof02KY6spclFEv78AH5DtZMm1n2TnBWk
Ng4YIVv5OmYmrinQkdFEBQbBcQbi3gOZWNZy4aJKTXgxyjBXdqFHTXXFswTpoVjtRGP4HOY90wk2
9hytUjQS0LCJEj6akaYgzUC150KIbe9rYmT7uVj22zN5dmSY6o+NkMvuKHyFKeApmLm0ZRvIJns9
CfTEJ8EA6MB1XFwg61xNTV3ed2AaNj/pbYVEIL7YGz5by6mnfndGxHfKqsZ89yT1ZKy0WCHX/cHI
AASDA2HgvBWCfPfJH8gFMConTqCtonZp44fqCxYo0OPgpTzcBNtva61jgO9g+aMcz2yvPdB4XK07
ruCXUMbCGBqPvMmcYOB1caS8fNwg3ySKH5UWcgdcioXQtmMCIepUYJSfTSTi3NSc5QZa+tDrRx9x
2Z45K/GPfGyynMi5939sIOJIqknGcgou6PQ+G5kx9ZzHuisTLlVCNbhmxJit6b6UzRmi3TmdxUIp
mufPk5nMdj+hGIph472RRBd5sGVE8jO1Eh8Eirr8P0qYTuYrqYzcxcG/xGV7OiusR7MIGx/gVXzg
+vo0ibBxIks3Zc35F2h1WkhEb88n/+STCd4BQNY1NNp51quY37YhgsQ/jlJhTBQAbAyx8V1NYUUB
guQypJPiMPdqObhYPYv8r5ixJ4+Em3QMsIB23I8HEJdGSc6LletW5qhB1RZq1x8CRs2GeYLIg1lM
oCQ5kmzzQnR3mAE2JBq99k4IS3NDcDNho/ZoaHe4ilWm9R06bP0Ua0Iz3UVyzfnFrOfIbNIPoDTE
h9lzVxzYX2mTfYldnfAmE6IEmh6uHV19Qg8dmt5isJlEhMI7YmAtBG5XAWqJwiAmcg36C6hKqJL4
JLQGam00qRmYJaV+yZ1eVogqzj6n3nu+7WSWydXpF9zlWz9z8w84ga3umsrky2e8JeabrXb1M5uo
lEpwo8QwHKk/wWFvqOOb/BEye5HRg7rJScoJx8jw4N7FNKMbq+b/1WHm2PS9thR9orn3Cx3pDC8M
E+2xf8nyrhIYLm43er+jS/5I+pqwUjRk90VGXOdVs8PU7xZ4RzdFdTf2XllSUOSKVBLBMLs9Etz5
DKtK3c060boTqlZQld/sNYN0Yqrl9oFWhOfKz/qfUucb6YlaxDbVDYMjjTU58tfxPH1hkqtxGy7V
yt0Vy6RU8QEFINjd1DssF0/o0/ORa7s2d0PzJ3euqz1reMn+yVe3HAADT++J/McQWwrgHegOFyXc
uQ2DY00FAif3U2Q7QQ2JD4tbrML6h8apK8eLHss7xK8TXwZ0TnRIGo7jilrCUNmbK2f6HRU/Q+Fp
dEc+8satogrE5BC6v1h85JPEcnFvJoE+jGccJNJxQ3nmGRVQ8MYQ4HzHC2gIQEtwN1wvDtVyW7h6
urxKgcvuO2+ZWnastJXc+qDsErwTE8PD6VrY0kOjyMImh7O7IRiPWhUEbIQkNc7fCWbhsR6bm48I
l7u0OW6AGozAXnX7phITUXpClXC1NzXu8GQVruecnpfcvYBYXxsdM2Bkth1MbIL3ErFQqcQJpMMs
UK6YKNxiM4BCXlBwWFIh21XCeB35CFZQPUkQJzbM3rX+uFRr/jurm30aIEM6xKqluWNU04WKiQNF
Ua6Cu0CjjchYSxvHJgwCgBepWQLSZH3xthvXqhX+QN8Oie4YOcG/tLJSNETa4JTYCK9Ou1twY5bX
3sB2ic6h/3WcdS0pUmnt2mMMtFDUpHCuS94xc6ltMvk2GGIxiO56buTzmr43eA8T3Z0g578ZKOYX
P7puUqIh++y/jG+rkY9/A4PHRA4PW/DjKswmC+W+DqwFv5+KihMfYBjst+zzHoFGv4pkW1rkk7RO
LI8qX1Kesas5OXNjwKXuYhnL8jCpfn70c0i/BGXnKL1fOvevn/+POMSyy0jPZS3VzJizoWwCP/N0
e+wo6Y7GitY/hFj84uRPDOJwbedZuHWwXxD5RdPhcLi7LUNBh5lJJi7hx/UDRk5hmOnPMt6KNalP
HJ0gKB8gaOc9sSZlhhZjip9cgR83BhZB9r8qYPr+RbYp7Mm1Dkg19eK9AYZZl89kfFIBESCwON/w
qVY5RXU2rm5SzyjhXiv7+/+CNNcGYAJVBg1FVyFYuNrlXM5SWb+tVXx0qBBC66SMdmmmQbSO2fHm
hO3acLRj8+fw/Ijl3Alxopq5R1g6qO5QJiggzV4kakoMXFvBlW2l9TkHmzaV5/HXkiB0M7Wyktly
GFgRWVUCwI3aoW+6/f25G4JSkhdyidhtA9stLVbN7z/7qCgV7+8SCnLwi0Y6dn2oNhYFIhwTR+d/
oGaF1Lh4uV2NSDb6aZuNuYvkfKA2Y13aZusqceCKqhUJAJuStR/UQ7y4heyL7hQdUmJfNyPTToID
YqdKRKU0ukww0y/JUnnK4EX0sy9Npzp9JLacKQl6Ih+38jxph3zLQ3MNQOnhvBjdpCPUf1sfuh46
k9G1hiF9RQw+ZEhvMlGU3KhrHOU7MgjxprQsT2y676osbR5ImjTi1naLPK/XGpSbq2I8t+oSrRUm
ZErYShOpHqiU5/DxNQ/sLzqpnwbXVaDVqVtdAg4B1634YxRArcdleRmR1pnqlvWxL+nxL5JaiQmd
VV33TEeRWCPl8q5Dmmt6TyoCgmzuqYVvMbZUrnBcDVK+flaqDN8uzOqyxe7YfjDQMDbsBRTxhwoE
0oJrlqqwQmw0/9eX7KSuRdojsYIyefOoE7gCHPkrtTIORPst6VCKSdTodmxzSKMEchPea/8CbEH4
KZUaSjrAYs9aA1CFaswkCSD/jDhBCtCNJ17dfbaS6RCRakFYs4O4zDcwLFulXf+z+5zYWnsh50Mi
wDrQKSVS85FezJHSyXuA1JMQJSoX8L6LXfJkhUrE73zeReFHG5LroA90Pc1NA4eBrhmr8ZCTX+Xn
37UGD16udanJyG9SR+4easjiX5hx//x0ABX9gtgVnJP7mbTP5M+MXT8GKvo2qbgWFdAdB4bBZyyl
Lz1WwwHaEF4r+rd7JT63jEldd+AsDzIcihBuDuUB88dkKOlvlTFDIJf30ZDK0w6ZCOwzV/72fs8P
IBdH9MYVzVwAya31mGNtZLwp6BZ+bs775tC4SeBMzWWEWyjZnV9TqYKMAN9zVFLZqmK99GByhtBF
hVoN4zE++YLxkdN1ZZilk6gBOfS4Z/7RMAWIUf1IzMo+RX1fo5Gl9iwljkXaeVtCZE5sWX4DNeft
oFeGKoq3SIy7s+DxsU/8Cg5n9CQR09LQQMzhZeYBPV0vZscHu0TYaBYCTR7HM3E/E6wegqV0P8ze
otnr4hKAME7U3JXhN4Xbr4rM7EPOouBlo2wi0CmyHnl6tQhRz1jMjZSPhYlHIJtl6O6qk6GtvcJE
MkVSYxDSg8GTzTlfsaYV5d6f7rgLJg7w8wBKHBLmTUzDfBDvYXmCGI4pzciipOx9yMK2MfY1t5Pj
IGDyuaTrMrTnD8aLs9xbNEZpr2NLjW/Bh3gNJzv1px4k/J7/zVwAIPOlzete0JJVZIzBPGMsrIMJ
my1PR5DlNwIuVzJ5gaBjJam6CDI0rsKX5HTZ6M2VcSrS9pEugJsR+2j+gBCcNo6UQj0dycL0GjHl
phpzpWZ8YgybkphEqCJEgHc+qp9h0xvyL1g2LEM7K68A42/rv3/S+RK14X5IWuP31P0rSp2dXA1E
ka9f38imxivaERzXZ/bxTEgkqG4WfoKMELPgXuywG4d/4mHAdp5UecM8oq/TTAXnxb6q22nVt5GN
ryhSrmBbF/5B22eukjD1c6Aj83DIV8wSC7yxoy9aYKkBn6a1FqKJwLCEjsxgerEbMH1dSjwY+ZOK
NHikc/OVjPIPhn6zGFTUhET53c7E+GQrcCxoI7FltnvsSE7DrT3YYFy8Ho6p8W2LUjHVqWrwNit5
5KQociz07o2gXasNjj8v8AuebJ09VO4eEXvnSn8L2U1jTcnHYclxXopY1qHnQfGEcMIZuPiHYCCa
FwsquK8zbHvuI5XKiYDJEfKhA/L98e4KLk69uZ7n45bchYSyQgw6YQnZEkY2XQ1QNEehreB90hyA
8J39C69xwDMABrnq2CrStjZ+AmImzB4GWo4ZYZZ/ZWlEVXMt7hynH+Y3MJbvOVER2lldsklK321m
/IIbwTn5VM+aJQottw5cyiXukGVqhnAepk4iBD8x6YunP7fzbgi2rv4ZAtyUoEToGaN1PCXNrswp
Jzr3Y/QnjwWF5yLKtxmuUZlsTsYyvHp4k8RAIiqHIoTarJ0sEV99I/kaDZ0huLFe4hFMjQ9ZIy6h
KlO0lP5uf/dmG1gh2LRC1UrVkamJzzo9esomkP/k45Z6ABUTGWuwQcGw2ghnQdvAW29o6CZdnXpX
Fto5Biolr8xU+Y+Nrgy7E3yDa+VD4NMpkS7kElb/ISiAIGJQ73MeYUqLRR4qvfTGNon2/8hO3XHD
zy5MwhefDrO5yD8s7AGVgguDPZ0VJnie4/kvuRUU/+CQWleC7s7oxzCKETd87X3uJtqxW2g6vray
ZYB/OYdNJhG4FQ+05w7+Ar/SVyHIxdl7B0c+C9XPuEbML8QsyE3x6BD9PYz12fen+/celKzystKA
eTHuLTwYV6SHBDe5BTyC6kByyFYbP0VSQ9npby9HNZRqMYzDqQLJl13xjEU/bqyTChlU4NFGPtKa
+EsjB8hgA8GS8zuudn+AgNNHo/n9Rl51tFoLstqI2/4L3Z0UFdH2hcvNvTS+E10FPJIO5KSyIS+h
IyKvRjPCHLFugGOlxwUESRQyFKlQEuQWCBKlYeRKiS1hVVgNfpjKk8IOb6NNGPSPJoix5c2UpK6x
PunIpW50f3WOaar5fLL20/4a44cXfoFqL0XPt3SQyP6qFMOrFdTvk/7WpjmiixBmgG/Q++ufljBH
lbV/9U+SzqX7PhH2aBqRW9ATGOFDKjoypXxMgt9H7AyLatmv5jaSrhjAEttIDVzWpWaWokLwh2/6
SC4XQ0x3YyqxWc4gB1v4HiED3zG9ttgSHv8E5+Dn69MaCjKhPNMVkmiLcsYfUso2VlAxqtR6azJV
WWDHziEzWLAL8RLk0sGTOk6opDorW8UmgtZ4jI5E1uAfP+EiXA1DP4qKA0J5clhyC7f3btNxYXk3
3ihF3rONKCOQd9268QACziQJLYa/mPBei5Zp0lfblP4JVVAQ8Q0NLwOIUR4NFXQIZzN8QxrrhV+W
hneacqU6qdHRQWSQAxpoOfA1KQW73QMC41xyUewEIKyAw8GfsdKC92qNvs1d2V2qb/E6TKXUSciF
svtaLrWZUlEex0Cn7mgfaGdyEJMyvAsqe4BQiFTcTKn2gwSCvo+ZOPl4GcyiwVmak2gC5DLI3HwN
IPLqgRreWyglm3hVHBTZgiEvXeOvW8sDOYmpx0IpYOzKxIUfusRODoslM+DgLYrwOsBUm0Sq95gB
4ZW8RX62zuYVC7JDHgYZcpm1ue2klcI0vbYIp5Kwe9Sb9UPQE0aVhsV9lIql+EMJ4KCiCHnPW5H5
JzdxG1W7echnwkgLLNuaUYv2zvbS0YAoiG9ss/X01W0xx3rDlyXop6WIv9b60r4KDJLxyP3H09o1
vRkbKS+D+4bPBmNtIt6Z7XlegVWYD3S+SvLo6k9KSUPn5ysN9gndOZs1L14lNoeUsvHN5OcfZm4s
LF6MF1wvi2YcXARtA2l1mhJo0T2zXhRv8jiEEqIZRPbZ6mC6hPKkmISRTBtRCwpE+5rGxPwTabQ7
a0gE4TioPprhjKoILrHj+qnMrxtt/6Z5bhecZ3ZP57zf36FC5Z3syah+fsxdxD/TY9cLVRKYwVLT
NalDrIW915uM3qF4PaGGb7r0x8qKkp1dHauBAuBVlTvrkvydF/fRrX/lAtk/SPffecVZhvyBZ5Hz
0qkAzlr6zByFyeuAXtbd5y/W3xe4w0yuZYg/jB6ikyfKtocmiDbuOjXjtmCyBmHcC5DLENolBHEQ
+O7Bu14yn2oHyVD4NsD5KHBGns5I2b0Ey6fXu7VYRjv06MW6kLIVk+d2FE1jPduTYGPIWDs52Dtp
cxYtQwIPiS1zPfH5r/vxwUEPJzkhWYGNZtv6MfueDeoRxb03kjlkA2ZrPrdPlr9ULQTs5KHR52Ms
ht32Rmy+kf9RixGKBZ3adV/FrmNVKMKw8DfqTliAXPZJ0o0Tn0Y4NMFdqcbVQj9bnzTK4f/ULIOt
atdRnIpbPnzayt659lUkmBeg4n7+pTkt55G1qfiqhvUBgqY+DH/OdDfa5oBIvd1aoFaqEppau88p
BC0Wo/tZWouk3mIhzEkQLkeCMnlQ6cLaaSYxfXfHjxjWPTuAJZ0/u8Zx9w0oLfEGWNdqmlWN7QiH
Ap9H2xGGJ5kUYIPJqjj5gkLKyYK8gUDzYloXY7B1O649+sfvYwONbOto3T8IBIwpvflQSE4ge2CZ
IWzw2NFUjO7Qom+5nbcxBoOvCC9sKEQgNTc1hZxr6GjhOJSA97s2RZRzdGFzMtfc0UljcJ9b5Q92
wHA/qHLldHR23Camdxt5/RLWcZ30caIY7Q/kD2xIV9lqJwuoGg8Oe0Rux82VwcuYF8xCAzKjUPDP
2mEQJhChWZwGgJtjPGI+7vStp1lzlemYkLAV43hdRd4849wIK9L4ATY949Fh6IeuvZAGmqDkTkCL
ENcz7RbSLSvm5Tw6kM87NgXg3pKDd9IT8s5u9DZZUMEyLYV8y4EW4pWnu0RHbMDQGswh6lXJ3i1Z
5V6qWk4iiXYlbGpzwuV+rgKDUsQboz09cHaomXO00PLBYjJRme70KiZhTmgTYjW9dZObDIH+n/Wk
6amSU4AaA6gsXknyjjt/2H3z3rzf1Cj96EtP7AwHiy6E8bajXI5BVw0GY/0+9attiBsNOPSQq7so
gWazckcw8xIxdwiK4KNnB0JOQla8IRX2rO0JlwrYO+VzxYTyrxuYq/RV/+s1XlTdAEHul/LCbOBR
TUSszsCFzNA7L2vVJvfxKr3+gvopgN6HUgXaq7BvWBnIQgWDFuH36giiFVp1SvdMmfk7Bst1warX
hLVX0exuTYSmD9MZ1pLx4UM4ArrBWSPNZ2LSU4NtSGL2xdqh+ayLwkFmGF7nMd5wY3zhEdgWFJC/
y+JYr1BvwEx2wSsH7M+caNkgH/v5sglzjJOS4bv+nOAJqcoc2gAxWpUcCXK1+YkIDXNrMyP5OwQL
sp1PLLTuqlEoOp+bJLG1W6RaT44370N9SspHFxif7CX4DQ1F7c+dheTWEoxjqcJs78IOCKSxlmLP
dH8o/GSKORpNtJ7LvJumGI99N5zPPlryug2ucfv9aGvKa/HCTKOoPTh58qqwov3NPF7c752LJfMj
IxQxFx18oA/cScC7HU6gfoQLuSswJJia+lm8m4wQjpdYj7aLVB97WD0FP9lWirDRiBz73mLIpYd5
PV9wiAAii7YdXmY5yG9k82nRovrUQJb1bE/U3Hl0YFiY1LggMiiH482j1pbWxXpnXbzugFu80fKc
2FRsPWzQuYWyoBrPI52N9RKAl+CXLiNoksaKOkuFOiKAR87VKIWnPkxt+VqPDrtk32z5a7Guklmp
PmUqlQLRa5Yrrt/VugXLtzwg/KYFBKXqA3OhVBPSWluuAYJONLELFMs1r2YyLUSobBvdKmTnI45l
VvsdfNfDqCWQVwOV7vFXwpiGh+eq7kyqOeeUfIFY7Gi1ZUZC4oZsch3M7aaowa+YUezZ6GXtaqiP
zKvfAOmQqr3QPQ4Tu4y3XpIMsPIEabpWTlw0koSwP6DOc5lW6h+tUx52/ysYksex61zCQhCoG1Cp
IfBQVTe1DINWUhXmDQerYSOqwnPpM8FHKTJUtFJHjKlBnSLXO5w0zG0vl3bAZYDhsY0NbQf7v/kM
hyWPgFp6QCLYS+wUM8uMXOOT+AUlrRw0zfRYIfj9WWuLOSnuijigntAIy5m9TcX2wWK9FawDa+3v
rsFPZmrpK5INqHQDcvbusJr+4NPRjQMBIpgJt+9XQ1sGgu/fvhVkCVnsikefBC/4t4hZWReirtnV
l07TmG5v1uzGjL9VtSEcZBR0JwD0WAtdxkQgpvjQVd3l+B3/7DCyW43PRcwCEiUn3NKMr38a+IvZ
2ocouQGED04aeiC7ug/rGyL+7v1QjpDYosfOH0//yWmdQE8D4FNuV8d+bCBZ04LFHxM8rTCojQ6z
+N0cbdlOJCuwwPtv89FbfpMoPbtQ1RvGbrqn6wVbuAfomv41qd/jcRzT2tG2B6+Wl6sDEO/s3AeG
MwFMGGvfN+I9ybaNSDE0WhsqzSzddb/wdb1dtt4klp/CpwwvFkVrfjY5xAsRXqNedGdYseLZTyOZ
RsPs1eh96891QnnyqgFMPyaGJUtfKiRLG2J0veVKqVLbVHCc2JalixC1+1dn12oUaeq3cE7HVNtV
/Sk23aEbpsp1K4OHr5WYGZHCcgsf0wcwiRn02kvylLfuQt7K0Ye9FBtBExJqNhyhXlQw7fVum6FS
/MenglujbWn13TgWNA1l87+rH8lK/Stt4DdPMFMZetZIyFIyc13Y5fmxt3tdXQA0EH7Ox0NGKvIL
BSRk181iKy0NIuGMvrmnf2tEIvSR8aqC60oBHFLM6wsxYmkdBKzD7f74jl3B9PWBJpyV8MhHobE5
RsuHQfHhCP/cOWb4RWbEcUX2MGiCj9Ebmp8dFb7EZI/8uohjZ2d9K7ktYK8TXNXrvzgqSTE2Saje
r8TWi08Dsa4wx39FePpeT6eL5Tk5vTSyFUzv8lVg5r8PRJvLG9zP8lIvQgcJ13rposYJQyHHRDOO
Lu1cMov9Z1wygZ4ldCzkWSYyTKSvufc7VLq7UogxX3VVJHao0Kn6anpA40lPrZVJR7VeQtveIjrz
7jKzP6bKCz9h7gHiacKpZObElU+H7jDOLFnyAe6MfU/JMlL+FYO7IElhi8DgJh1RX0z/yTKsLc7w
wwPEBHfYeJtg/0UtFz8HLuS0hWaJW+CA3VQ/kQbHHFVkMR8qxfwXHtXpY9WQFWWfQDvgebnLUUII
FWhUao36UEy4tkis/Pgd1cx1yYz+qTwYurWAzFOi45lLojnJ2Se9GuscfqY9mB8ogWTNXf4lvlyM
R9xQB2GJ2aDOjzVW+isfh4bO9qwB6vSh9Tj9eMgCpoAZLYU2Gqd4+dkamTGUyq3jN3FPa0q+1wrn
pqeD7/QQ27lZmBXgZXaoLPjdS540ZVPaRQU4kkuAgGk2CdMiJSQ156of+G0xUKhCW/1wUYU4h7vy
LsqrreE0CZOy4/8WQ7SESROzCRrZqMg07+snZ03kvURQBuBDQu/m+k7qFBIHkOsdf10Mt/RBddD4
VFBNM8afpCEeZnPGx6Ait34Arg7hODJQxn/cC6+hdTsJDH7OT8rwXW+6kZti/HMbxSQ4tzrfWtg0
JdCjbpWvErC4TTzt27tRIzYY8+Ii9ohbUkosuUvPqdq444HJNkcE2g+dsoLDEw4LLOCM+IicTA5c
AxSIvCDkiIXO5hYCZvrjVVfIuL3j0Axo5ZcD9A1htJ9Xg6JGPhOgfbOObrkbPB1L2n7s5zkZwOaE
RS3tb9gf5+USz6O7fCIbTeokMn1tQ7G1hnbjbVZyiA0Q/Cc3TRAacrfvyqk/HzbGGZje97gigDh2
uJycS4okXuF8IB4myzpG1Q5aI/IpOcb+hY/gxdCfA4WFklrcFNolQGs65NF0acmljUDEYDddKjgt
C5TrwG+kkSFtcexwvR0Nlp6lJO2YDyc20aqxOxZ3hpTtCtCUqIxNWmZq7dvht8fXsOzZVsT3wCWP
dQT4eFsj/S6YPNFKVt8czqedtFE6RtcQOt6PowST4dqP98Lu30SvK8elUHe0dvk5olmklWg+oWPI
2Xk7dcUASfYcckwVy/OfckYiwEwkw8xVFQirn2HJmbUJ85bhwFojjNVpEI6qb+HeWTRilIoaAjY+
vXsMAij8pyxf5ijxFyVw8QO0WVOv9vqMuUwE5S/XQ++lsO/DEjBae7/C/kbvFI6gx3vPar594LdB
bGJnvXhadGDZ4fJx/xb5olAriHBpoFITQXOix19ZmRc/0Zanvq1jFXN23qmtsXAS/U3qsSKyKpOK
lChyUv1N0XzTzbw/lf//2kh7SA4fSfvqfkuX3JIBccvI/0U81rGGoh0GridqrZ6Thcm7JL9j9h4Y
Gy9JICEga+0kWN9yyhhYsEFT/adpVOkLEsj26JTliDFw0sgzCkQz4zGykQW1Je8U38yUfdAxdOvF
n5yee/005wyWbV1PxYOhTSVhtlDBm9bWwchLbvZldz75VNRWuMdDyG1UpNLDoXZHE3sTMuRA8T+F
m+DyBRQcBbZp+0+kksRMEjusRrGPsorp1ox9IAIuj56OIsDAO22OS4X9OqC5h1rXe/bAPDNJ2NjI
K6hrhTIf8y90MMdJTDlpbh6zksNFs0IxOPsh4eh0XdL4lbvnleE57lE11qQ5Sq5zI/8bnuxJo3al
Q2EmGHsRiTe9OJWzHmkDfssiHY7A0a0gEBHteSLSryo/KCK0YsqLAOSUyNfbuBk/QvLrYEdpWgAn
YHj42g+KdAhOOZZBdrm71qP/ChcqCkpL6ns4LHuA7FiutpI42Nv/ft+k3Tk89oKShxz0RMrmNl//
a2+Dt2iUz77Hzm6fbNHqq6kX4HxJcTU/RCZkN1WU9AM4NHtADkVkHY2VWlk/4OLeEPP5ZFdWMjZn
C6GRktoFDCVT1mME6PELrZh3FOXUwXZuJ3mcVvMq6wBfzwSv7n7K0e11w5n6fhrTCEkOFc4Fym23
79wQb1n5sM7q5f6AhJaXYqWMJ3fflBnxUX2b6Pa03dlpmx49z8/I4ZTVHkLniXbFyXTA60Rl0HC+
b0YowcSqvsunAFqWiFqhXFBYLESB6pVoocMCsIpYMuW7tpI+31xK3lpKPy8c42kTpi5TvCkoWbh8
d2t9B+0aYfoIyVppfH/AFsdSSPuP00nb8wDcVE2nlHs8bx/ZITDodgNoYvcYszXQAlQ6ZOzyYnLi
A3kAp2ITmOqyHgAkNCTJ5Ieg887huUbWBIgfwVVU4tElHOl/AM9nDFnjtcgbmPT0ufSaS6nP+iD5
OBxAoSpNqfPGQmFdc3alLYiKBQYAoNAlQ/mj0JVc8d7NJX+san4sESKcYePN9jlOFuPRYFuk5yF2
Xj3H/CTgqvaY1XdTJfZKhXdXws3vGcwVB6X6uXpjqtg0fHRAYbLa8yqvkjobKshiOHUTnbyq8Zid
fSwGLI03akp5QxBKx8uyahGPVwZDGwh6Emd9ES1ASRENFqtCh2+TDB3xlrsRNSLHKI4zMvYfEbpx
VyHzUau3kFeiPTPUgrWEaKXpNy6t1FgRAvlqF7+gRFK5OFj1EjJD7LMnUDIVIFUYCokFhAGEki0v
Y3cPIIkrC0naLn1k9dEAetawVtcjBm2OQUskyFpSjTO37ZXkNLseCnVIWtDhN8Lh9UTXmyP8dzNm
7kXmMrI1rWZczokaJdDDK1mOQEZ2H49cDRwNFixDo+52Gh707FGyBmifxIZvYjYTbYUxh0bXdkXo
/vAfduA4s7e8CnOY3L6I9svUA40bNyuE544fVUJK9dQr/GSoFy59LT6tfuWr5uihn4Vik+KGpsgJ
DW4xNEIP/9fFcEameAc8RXAC2sE3bq1MGrz2yTeharKHXHDcikXsxejPH+RHiDijFM5tThIbP/MS
Sz5hmnLG+LpvVEQIJRy61DfBrY3moJCTB4EGJ8KJsOKfDdrwfG2+EuPib33fokO3gXXv962AuamO
qsMcR289Il8Satw9E2IVqBAdYaYag+VX96yMaA5zOs1f1WgqeZAQUX2KG5yk0+DsDHhPY+ckcm8i
V8KgQFfrjm7Eoye5g7S4z3+ezDn3W783nCf+Nu9DAIAjysBe45KvbdeLqJzZJ3F8MUFtB+bUPPmo
achjkFRtZaMxiA1YD9ie6j0ZnjWRvbrdFmL7yH63qwZ7SKAbqzk6nqJZDJpeHbLnEv3KRYek0YQX
1NOfeVSnXJnyFDQAbzec0e3eqJBSX2rzTLm5GZEO2YRpVP+1B5x8CkMD3npusCQrEIa9Mv3MJdpM
VXhCKevl5nSSo9QjRKsHxHezjOfXHFfimhnH5oQtIYcyJtwACWU2gxzCM57DA3jCCvW538nEooR5
2T3cuf5UoXeUKZ4uL29t2AUwQoV0uB8O68Sg0uHFuB/V682shvUHToaLQs9prcxqoAfkyZ5wRYp7
fA6gDbWLMAJRVJysEVulSOjo6mVAlK06c/JmzX2FUGxG9mYJak7xANVza7xl6XvwhEi/VW56yYkC
lKKTlm37C7jTWM/iPVLyjlmZrNPM4pFxs0hu9U5IIS9zfZHmq5LyEbYtX8XXshkrsnneVl7GHW7o
uk4Jbyl+YW1nthXPzsR1Ru8uTBh3ob6yHahq1EyhVB2cQO5GP2vvoae8KwWyeYT8BdPrrxLrXGmr
JwhZCL9DRUr6BkG38aDLpcyqHjDs8TMrmaIqA+eQ2Ikl0MeEYVGLt+BlJ4F1d1qK3cKhVI5CDot5
LYONZ5AkT+XE29oDHTdADw7ISygZ5oyLIn207fbvGEZUvfurxZSX+q/JQKzGr4PUreIEyl9WYc7Y
Byx5mlbyuT5ueswhbseX62Bn7Tr6fmYFzOmAtILgwLGwf6ccnyBS03Z9+OrSD7RxOGOVHlTblOW/
L8mp9I9ML586mThSwhcBhuhcIbJMu8y/FIMR+C9fDsoUY6oKZRQVX82tXlMOl0HDeBweZ78cSeQ9
KYE4WP+6M/LBlxjqpUR7pDz9/5qOZZycQK61CvqoR154qkzQm9lyex4P9+Q8ckTGLTraVUyY3IWE
rtDFKJPfcOI5EXBbzdn11uDCv0feE4Gc9R1GpwQhuTXaXhoy6AWHrQE4N8ZAeH7KZt4ArHmtm0WU
HSKqkm6dcfxmW+IqhN/UwGMQAoec7iFbE8JGwPYQePFnGVXaI+tzoWiMDNozhTeWpAuXTigkON1W
mHu7jxI1EsdbbHjU5tIAfsN6z5cl0m13lUSORUgB+pcZjRqVN2Jf+WJN9JDxgPZ0pygj99YeAsAF
FzdlFWcVVyPdLmLRg+CqRER52lOUeYyFbeH+yWyBrGXtfP0SCyWVGD+vij0w96fIQVHLr09LA3Cn
BSphIZbGcosJ6M4gMphRvZvchtZFc1+5ngKb+UAx1Hceu4Ktr+tT2XHB4TpPekWZVxEkBv8pl8jj
oLoWpiGdAfzQ4v7fmIC7Z5nsqqxHsYaWX3Ti8IAEoTPqC9ZTRri0fO3emwOec6fMop+LWDwY7mGQ
o6JZ8Rno3NvyeERjeS82E9IgJWikbAZ5ez2j5pY8tJp4z0EqiuYhd2Ot1MrvGtB+I2g0uJ0fXBGP
YEXVgKYohaXfO9uQccnYVEHPHSDlzRDK3Hc2ukqoNpF02xdAUP3ZglOGXf6fPvd/i+OURp0rUXN/
9WZIznAyZ1WYflDI0oqZexo63H1zBVCjCq6lezlOh4X2Gd7GuEFeObjdyUyvZvehXgQ08RHynUh4
vuqOx3fOM/6E3Wpbw6phcGPyYx3ZEopkVGWcJ18yrkIMiZLgvX7E8NtRvyVhsDPfRgqD2Pq1zvrB
ZYoHKP6HW9ukGrXDd4DJyOhMk2nHHPNsx2BNgjxmm0SuaM+wNZ3pk69LQEz73BfqamuPmMAfZ5PY
YhM6aPhqBoYhBhM2jF/JgxAxLTYXp6Fk6W08+xZNJybe3f0FKkiyo8sLRJdhn9ioLzC3s+0hrXVl
BVwKCIhbPm0WDp+NqFIsGlOTeH62Oyw7hJF48X4Z0qruvgHCTA+YJhzvmhhDs22Ft0tRCHhslicM
NncmWh/vVQ9pkQS27KaTtS3mhc+y3Jxbou2jGxv/RKrXN7GS6DaN4RUn+tfG0HzZVW6XaGZmwXt/
Bj6LdaD0R9RIiva2aR+Ae5ecaXKWSfBIB41ZUvxw3f68MJgQKsSH9VmraD9jNyvfHSDBSou4NMlm
/INT2Nfd6zyIOwDs4Xz5Pd/sfqZu10j8CitpaVad5xVj2LqAj9erbXSXM/f5Tlh3pvHP1AAioBAY
dGcOtls6X/tx5sRPudj3dbyWfhVLqlkwM2S0uOCSNWGEoVh6BwROHSCloRG/9Xgz9Q1/PAKuwdug
XW0F8HM1dK7R2idkD4jT90PAf6PQY4O7U0aRVqcgk9paQisyh/Ejqf4LHe+Iu1UPh159yibaU2I5
AGgzdPSd7zjxemtUSLQHzGx6uVaU+YvuKQY2gftPLmKur6ZEA10fpKAgo1G+UQvXTuRDoN0KlfOs
OHT17eHDo0tK9LavozymzARh6jO+SgQT7x1U9JlPkybTJfuzVZONOuzW0tamPm4P5L3kyRpFckVh
N8jJzUHOgmnTabhc37lmu15SivUSewBWNefctmQ1kwxrOndWt+FI6eDHZ5+VZ9rQzMPNAMfdBVTJ
KDfPk2qenjEPiNRmPZATErImH1UIrVdrInoGtwPbiHac1+oF0lF+JXyWOSE+pW8Ry0OvBu+wky3b
/Vo3im0r9UWoaaNrD4oY+aOYVnmIEovxXVgbFGx/xuI2/Fp2sRk++pq1lvR1mEcExvRslsRX0Upn
gkvD29kUzXAVanIGSkdhexsV3ASe3ENRGw/N6apNUCpKMPv+9YRQ4UVVQAzj3XthudF42gJ3CzM3
Kycox1m4K/Lib4DZi/aKVNKXTfeNISGOvoTMn8cMca6jC9jHYu1VzwVidTuRy7PVyD1zeKwwBfeI
bqgrFcqifn0kAE8QJlf3bpIWrqek8xexG6X7v8ver/LNFVaf/jfKw8/n1zBceKEE0tvg6Jd+2bdN
YQNB/bdMIWUB7k6S9cLViBugBEElv314sVdBB1Bx1z0RD+wVb0ZOBnqk2WZi5exSMZZeMmpNY2kL
mw67fdjJ1ZyT6hJ/2pDjDQdeEpRa2vPd6u0Or0HNAhe/X2IeopvR2Q5pIxYYSjsLDc6p81kw4Pa6
8f3jrFK1L852L/VmpjmyBu4E0NQCAJhcs5vPKk11P/WPKUPRi+FliXwnSSw78tLiMu5yD25FUpZ3
sabUGYkHjWjrSgXBjC7jR/X/H7Tn2wEpQW6fnop1DSk1kcuqB9V8sgWqFtoEBP3V5fmfLp6GvG1K
6MvGdCQfaxdEc1W5RSgfu98ULK24Xz+3T6LrEM70BLQ//sC11+RIbONwgJs5Vqx2DZ41bkLBMKRl
/hbsLbNh6b06iC7vIboa4e/lIpo42/ldIMftNampGrf8OWouft370y3Aa2uUvnZ+eY61UrOsJKof
mfljfH8q9aNeU/D9Q6zSfeI3JZGJNfd6MHO63gOHY+GqSFS+Y7gCY1lbhLtyUBQfyJMprhfzAo9C
oSyk1xbdief0hXtuRxUhj3lKa888GCyEJr5ZQl6xsTdAUrN3QIiimb/PZm2nfeowDDTkAmw06cM9
aGcKPrZhkkU8supGVTQI8eErAg8L5Qffo11DEDVnEJdW2C03Iism8sdLhQutDZa5rCrGbWg63GO3
12IXD/vZQkMjDknR0++vrSwCQQou6rtHSmcOhql+DhsU7hVemcm+V7qmEGBmU9yORpxZROz7iTWe
reTkciwrIr4Ut/+FQNQxzLo/5sGRliEU2dBu54w2B+7S6e/zuYpJwfYQhlc/tt2LIvavjURmn3Id
gAQbpMSpmYBTUz/WnP97Id8/vYag7IZ8B9WUANZYsQ8RWlgwU13E5BaphfUyXxHoeAQCB8cJOmKs
XzpPAvyBvXYefxuea63oZaQT88tTKBqer33neGM7aIKfcZIMWmn6nuFr6zuIXhBQb4SIc9QIGiQ3
qW6RABCX7HYjBlxV7UqXBe3vxfldqu2JpWjMclZKNkZUm/pTYXHy3xRpcqhmcfh90jhgEKgHfT1I
ndudQxyF1cRJL/pyqOzMW0UecJ+HskG1Cj3G5waSGn+0XO5R19xSjv6mi38yKxvo4jrsF47iJJaj
fUVl+5lR7SKiVpQWiwgNlPqIwMY2YPi110xGNCaOKPx1LBGu9e+iS1DjBUq8LM7thb0G4yFrCpew
naFkhV07pid92QuG87bu0MJkHQ8fqEjuSns9Srhmh+ZnqnLmaGqPrz9/DAQXms9L3yxRsClbxzWq
qni/3Mqkq62bpfWrv3P6a+nn7+Qq7ZDRsp4n7BtxSlZQoh4kX6o1LWtNXCosPTaWZ0T3WJviJe5L
oI9K8CbFBLJ3S6l+81Gaz6/y4eqhz5rrxGoZl6lv2mQsGUUqYlFIw0r8q+ZGlmmOHplKo+DUeelM
UVzTDjfUSRNBeihGrgmj1BOL3FzBcQR3dd5BUB5P7BbEHmM9Eyj3Q1ack51R9xGr4s+EEcgTceu6
4iYzDZoxHKnE7luqHYFHJ6Rzdc4oMACqLnDJuAaNmx3hXrQbap2ELZjgYIrXuJTrEreeCfrkyqJk
ssHCXlEqRgxnTEf28jGTuFRhhv6k3f5fGZ8tkTT/Yei/o0h1sA01K5olv5RhSsNT3WDbDPagD9T1
W1Z5Bz1twP3ppGI4APIHPiLX1fl+xxLjxUpqxQIOTYgd39Tvba8OfCNTw6uTMm3soRmhJ7AV2WA5
vbcXRf+VuR20ekLVH+kqJeh9fhy1of0qTcLf4a+8f+m/jqZUoXAXEgIeA0bhrRo24uHUm9mg1b1M
/uKqWYydh8DlNu8b1ITgvWOtIs8EgzAEgBeTF6LeIjmCCEGk82xlZn5r87wSWVfDuyhU2Uysjmsx
p9Z4/vRrIwf8Y2m+pATOe6Hjyu1HYPEs+lGWxnJnuneWjPnwB7907pHIp7YZGscY48vFZ+4kK2x9
KFf7kbHt1ysuqeKcHiOBnr9BLyxkkKtWFHy1irYPbyKm48TI0dqOydea5S2Ha62vf5rmARHwCVCx
Zcdo4y68Vjn3LPMns5ByQYQvrv5qMYQ4D8rmwtc3smfqV4+yaVLJYSDQpfCHiQm1VYyrQvrz1F8E
u9EwM8OECc+U8XifIq17ymNtLXgykaJ6uiVvefL3u8PPp0gwqersrLtF7ZPyrfnew29YEv0cSK4/
UjiZfmdzi8BOlBYDC7V5YVHk8XgwdhtGbmbCtESehZCz47SwZA+gGSm9nW7UeZFzrFz0dDGz7+Sm
fg1OOdzZ3vqrl2bBsFaq045H8YIWe4aS55HIVmkAyB9Cg1UUby2MvK3O9rFCXz9jxyIOhtLqHzX5
9Vb/08unNIhFtbYD5PUdsqsS4d7W9jT3kiWocw82GLM6iMKDrluL5gsmEFIsmor8XMhNh1wJ/AMD
Rg/HDvFHiwcPVFqHV2PPmo8nKwKCc8CwKboCypGx/o4+vflqCbzsY7wmgInPmyHb8YWBjxA4N1x0
YBTzXnsEhihP49W2pGI2unKGF5uVkxbBie/NpkZo/Yn6DtDGaTtvcAvx0TbYHQqHLonubcE02kDn
ZfZ4kZWE7IYLeY1j5EpJLtvlRFph95obL6+TUeKrv4/l5YuVPz/UAVUPDi/kk6RYdfGkHsdG/R8g
7bEdYHFPfJU1fx2qBVjpM6vpmJEpRNMsQtPxhFiSP/6l1wsrukJNE0DmFB/NL3wKQhE/p3D/8ZEC
FIhr8igGTUDGEOpexB3M0pjjYD3iMaQ+09hYl3h1113jiY5lybj5dZOF2uQCTZq6TXX14qRPWYEK
1nR6OoY7NWDourA54n3yDJQVPBw7WMmnNAorc/0I1t1hqBaxSLmZoZJ56uF+a7ewVUa5NuFl1NXc
kdBHv8zObkNxunKXmGQFKYq9/F+15j9wcOVJQ6ZH/+hEu7WZybF1ZqypFU9KpIqQPtoDorOQ483n
S+pzDzgD+TJBIyOKjbivtFYgVs0EEOGH8JdYOjn+AA5FGI6RIxZpxcgGEagmjZIgHhiePQTA/fNh
HG2knY/nLUFSeRH+hYpq274BPJdwRuiKUFEouSrrKsb2mzez2AFtxcxOjPuFNRoQrQj4OvsPf/ic
2nnL/NiMvxQmUSRRs0v4oMyuAA5bhtBhQyOdpimD3PsdEg0pdFN7253pWs+1wTFytMg0Kso30TAX
pdeRLfxtadp2Cgm4j3FPMnTaTwcASicgfzQweP8sdiFu9m7+Cj8ArEzn1C8KoRJKVbAGpfpPM6Dd
pBlFKFzq0nTe9euZBD6KIAJtuQA8obM2YNKLoXxq1DWqNx1YaYtKel2Jm2/9p1LrftDVwd10LXUF
xhrrjIvLPUWb9l0r5p0I7Ui+xL8mhDLPJEYQSU7MfnZLI/Tt6bpzcjZAM4iepZuunlSChTYzqotd
LD/i4IzDw47b3Cb04e/MuWEIF0pz+5MuZhwSYX57cH0thIE3xwJY3ELro27OfplgOrlMwLVGHRCd
vLX/1TVZGg3VcWh1dYeaU6v0ivaah2hTtiEJb/CN02XBF8KCQinLz9QGinGzwRiWOTZGP+FOt9Ka
wnDDDcMxp4Hpsn5lHelVtVPdCUefs2iyi+rOzs+3ovSCi63CB7wCkrtKSaxMZ2obLfQueImXGCbD
F4WCorMsciBffx7SsgPS3JwTewR1aOQSetqtb1KcOhXxtK2Jn4hRbpOPnPceUNB9xRB+NvD2ZAjP
B7ccBmEYmDbsV8b3xvEHeT5UTzEdki4jneBVNI6Vn3pkNZEsC0iM+7xE8JAa6OGsYLqIY2Fa4yc+
TVmdxeEvAhqfQmMWH6IMcDH6LDf1HGD7QgCycVUnBd7KDRKdTb5nvc47ycsf3xj8s4UDgkxpbgfX
WeblOtLqNcsI8SbLmnaM6v5nG95qtQbJe0QhCe3euJ1f5EX4tg4LcuScNo5aeD53MXNSeg0bUkwJ
0uOldHQSsEacIh67I8NcxmsJJ7XBjove8zEG/1f2if3EBK4r/UROB9+xZB35IUBomTncZ6iStFy2
dLGLP1uCcmkT0qnJV6fe/8onbF1NToYW/jjs3TBuiOivNtSg9hSAkP4YJcgsiY5pzS/Kj1jnM5wf
FC21L/rg4bTf8BHmHSQ41LFJe+E4BNpW8XXffrpZMASo8U2h0hRTQ36q3GMMTOdPD7VcCmv62gEt
1LoRmbCYY4EAsIjwOxmB1p7VBCHdPpgnLd9l5AkHUv1JCdRah7up0sqOUVqFREfdCtv/4H9usHJT
Q1Wa+6Dlyzl60sDTpxR4dzyVMxkOy8VFPQ8KWyerqDS49Nq2mWmeweNQzkfNaLRS5TSSnXZk6vvK
Vdb8ee6k3wPghjktLaK6kRVxbPu3VQ1OlEz07IjNajHw0fP+BT05I1YnvW3vmZW9hxvu5SZzra1y
hs8D0Tqx8VoWHHevwJfnMErOjaGq/S6II0CXMNhVlkoOtaWLFqmD02n6S4MZEvr2sZRSOIDfZSB1
fupO8bLHCtovk8Ymi3JFFazZ6Pgt9VrqjhGz+Nq8X8rbAngiy329co1YEtr3PvhGdj6r/o2MDcbO
ApYClYF5eIVBrr7cMlQnTVYod2fHBLNBgvOxErbWB/YKTrf0XJ6F6yv+l8pwbVaAf7QwecIvAMoA
v08UXUblGoSnMt1qREoLYz3IWbbd3HHsCpth78ARhAzQTKzmO/YWOIV8Vx5R5qFVPOi0WYQv7zTN
uFW/leooVMbAxAWpqJnuUDd/+275CeWAphcWo7Vt7aYgPt3qE0VNTTkWjRbUjQX6TB7KcQpcyWjw
124iLuQmXa1xEFtYsoqeu2oMR1d4volvRDf6Wbyas1rhj0x6/4RATrWx/cC8f358jRHy1JlQhlUq
d9hcqQZ21DW7Auc6fdxTYK4aZtWBBxYOArv0f0jMTCVjWSUj3XFLwLfeHJAUP4OAqVy6xkHcbs3Q
iqYwM7ZvJh3+VO7zjJZkS3vhXBBmQByuAhsWtXp8ZSV1fe2IyuiFSE4HWUziYCX6YMvfbBwjL4Ij
m1lZzr9YgCse6h8nte0cgSBAHZuMSM21RSMGP3wBbxVvY3+Slz2MLIutXnsEo6U2tZGh2eRCw3Fi
fmiRDIDPMlAnWITi71iYhNWQ7MwWZKrf+/d7S6OZhU7zs40nntcNIGMufxVXbtQsMEEy6PecE6XQ
HGItrFvjqwTW+YP/yzhRcoEtlpGigW8CLqbHVuk6f1Wd5NzrR7DGi9W+HOJdn6L6VyFInpDZCQxb
RLkgJyDPTxM9F3lrizqr0EK9zXKygat+bB7F2pUAQqZY55Y2Sy1IhwSXDW9V93rN5CG91hVYkmDm
hwXbMAOvf+vV01Q+WsqYhxJ20Idc5VEDJkmL4eu33zA5H2uWjts5LmBqTrEhfMfQMdhlt7ja0oU5
GYChQ0yTX6caGdyZIfxwWwJJM3tfWBHnq7igAIgsLbavlHwMTd+4K+DQSnm6rr+Adoz/fpwV/0F3
I9tO51llUGv1gu2YqmUj1GqyUi6SvqNi3eMwnSA+IHn0JHOq04jkzIbxtLFXAZbfmI93NyEdRYRB
YGkF2VtaRVCGeR6yD27qspgzyWqdJpS235agbRDEzcPWWyu/dd3dc6/XI58Q/HZJ+CIUZn10/5dO
QT9WGedyVoy6r59RZzgjaKX41Pnp1zNWVa+g3CaXhQKUfPTHX8CuVJ0Gz1sGkXnXLW/6anFmOamw
XHp6h9IPWhexsjTafS4oxXzU09aa/ry+HS6lWd/38j9eUNm41wATDmoF8cx4aGwzGLuHtQb2oE7y
Eb5lZTDld2xUGfLGlVHBKddQ8A+KyJcD4bfK4MPrN6ezEHqeNjpAlmIcE1gEoctYBWCJLHAFifxf
bWo9yA4mJ8u5vbnQ6bwC/WadwmrMZyCReDL4iJ6f9FHenq/tpTSy8BXKO1kf69VdElkaAPCeIhmF
JCcV7UrzsrE78Pq1/8yJG3pFYknBUguadlmdx31HhLqfsg2b/gQXTjyAACKLGDdB7h3WLlcXCw6Y
A/UH+8Gd1y7S4PsYHGWTCIVmua1ezl0+sh4Dqz0QyWxv3WLwSZHvqWJIT6XUX24NuDyB3qriceaD
WJm375i4DP2Sxli6Twj+BRFQM2WEQH7FngYjGYHlYBNMj42p27Aop2nihfit+tUi+1Hv0Eq80eeN
Prnnoop/qr4/KzVNVqQP1nfl3+r5CgDqX2IcFx8AQuqAouMcg9MzlejMP/vK/M32STtSCcGgPkFq
4h9/THZxk1YIkRvoXLoI3u9kgVkCrK5mcDedp+lJ7s9gTQaB/u+ciWVf/U39cNOq6fbsgYu/o0Ir
P/jq+9PQZUwGP/nynpTHwiSd26Gnfe0Huol95MmamvLl/FlDQMySlHMv5cJ+EBhEVrfvuy0OCtcL
W5rhpr4BmRm0OVNoZQ5B2LTWImg9j8wSlU1ldDRYxkCHPEZTe8ftjHTVLvPSgl5pV+cwY6CMY7Py
X/DinfGzH6QEDBPPwbeexnEEdDUQiMatCJrpLmYki2Q4lkDQZy8Km/MzV0aTgAzhNL1rihjWcsD1
mX3KWnNr/eevmtsz8I/7Wmzi2jAlVIA0+TWuewDH30XRboq3BqZaOT359uoXTpZb7kQhz3zFvutJ
P9gTG5ocJKNPt5Ze+KR4Fke5S9BWGi4wlcRuG9cUjmRgXZ2rVJd6DLOGUwjP+qN7bcifyVEH0CMM
5aRs8dkCpgAZxsdjwOfk5tglamlLDktmGMzfu6C4QPxQIHG6VRuhWGcsJZSsTcecAYaKITPXgT2r
h8ACLQWwAW446kTDDQy3bBaMxU8A4hiqQe9ARqBNgMg8FWJJTKzA4zLQ32rMga4/Z9XnZsWCAXmK
u8ugPNrNtk026Fs8PxivMbFe1wAc4vbQfzNkFgRmU1K+IUD87OlNjXQcx7VOtoq/eTsmj+EqmH0w
Z7LI9b7FZi9SDO0laE0vcIWHIGK6whXipfaPGZR7SFA80HNMUeu2HyKvQI9/JQ932HwNHyHKzB8I
WwpIgh9o4y6ex/Ge1Df6drucLs1AExqJ3jFTVD7Yrby0JsXtCLummZMq/hPYERcjq3DIrLBpnUN4
LxrPzrCLgpnEx7ihr5aw12AWIn8+HTKR6vofL1dKdXgQooFPKtxgQLCcMIa48C+mJIJ1+8v73B5c
cp73H8N1+XLVyZYtSZSX005ydTHzay3lEgZWJ/gt15o6yP088SedtWZAo3Uk9z5KcNQwXPFF3NI7
SbkUPrSRxVNoqEnVZEFoX8VoZz+SPbgLb3IiRQKAJxtsYXJJVRb8PR1OoZoDG6yyOPY0T8rfBGoA
f8uRQExzO/SuA3edVTvJemrV5HbrqPPH74nY4TT7PyoYtO7lWOwYyZaemFtCpSznJxRFXIlJjtsY
h08LTNrx/jfaydK8YuqDz9EsVyjGj5IW0CoGSpi/M6Mg8JWMGJw+zZ9Fnx5IB0AdHDubv5AiRszJ
vHs+hsp8Jg5oEvpk3hnjWFCPyrbcp3ltROMgHj7J/eKcXG0bM70Yo8IuAIgQsb3GfIFsZtxZYqYb
GlwLkOxmC9IN/rqYdsKzLFiBtnE0ubM+92skhFWtb1NAAE9pLgCa36vi9revAND+TE2KpAtf0H33
Cm6RgI8tTZhhx/ShfCDT2NQDIwz3Un7zXeaEdiCNam4I3ykRE7kYQM8goPkC1h+w7CnBNIAwzcX5
plS0vwZMhHh+q+db5Ke46HuRvA2WdeYThyz+hhk3dHMn6QN7p4vx5RRMlGKPdIH3+xNFaMQkerUR
vtqvvfYDrD0HdH9PyZ2Kx5M7hM8LyBRRmC7r76FZDUu4XDlPvpxxnQq+obaofoDEkzpunM+f7qth
kEZyoNBGkwbyvZIBGVqRbuW/1xxFD7gYeQhfF0p4azFAAmhvYq6kfNc85JSUIbiFF5GAl841OGfL
zbYLHr1EH0BXYH0TNac/ro+egaiGkRqhZGLGESomEJyse6vpFoW1NrRCzkfAN82rowGB7m1duyOS
hHPOYsedX3inEVnNsAeqiO1XGF806nFO0hUOKyFNvGIdf6sSoFTZX5VkOpp5ll/CDcJEO/2VvTEq
IE3omuf6XA6cwhQcO3zlCh/sqZqumRgmz1t4iUZsp2vEL6GGpcH5N0HOThyaOahRWDxZL8Ehtf5A
OmssG2a8rVq/GExu+yQbIQPUqXBdVxxlaaKgiiGF6kr6ZtyHa+vJ9m9E+H1DHqQXHNKZCc28rgOV
YAJPN2s2eLddKfpyY0UsSLHNlTH9kGFb3rwvVF9UIgraKdwERMWnqf9tTIfZ6xafqcYgPx/jZ8GF
HCMyaU7RNcHNBjX9Xd0ZS4E8ZlLWOamWTsafKe8dZAWAten4SNKuhDK6S+oZUOtKtgiYREd9AzeK
BzF3zE3OB1dHx+aZychHx/G2SgHLdgNr62EW8QB7Xgzc46/s/9UDkUs7ZqyvoDIuYDbgt+0kggPi
fcP9qT91EWAi1+5CaI2Z2is/F+Oo56WlFJF0qBsJsAAh2jlBlR+1xOSQEm5aOVoV+e7m6ctpxQdg
v+8gxP40Ed0pJbWadK5e520j69lEm+pW30NJMWvM1QYOFSbWlVLwVMUDiSPfGfTjpiUgyPbnG97E
byhUXPPfVqg9BynVqC56WY9rvJK/m1JDWQaOc9NqjW1pXomKvU9wX1adlx9TuP7IJXuYzGL67rmp
4T6NL+V2X2HZlyiRFsT3vWH/4+XK2yQtjApXYAlM8LhZ53uXKu3RqytuJr+kQdiwxX+8vIVnOQhY
qq51mNLk1IYd/Jj+X7P0JCVxObUJtxTJvupyywYk4K4OEr1JoAiF4nHlW7EWLzraacEooWLyZHC5
crtRC0zlaxBb7OJn0TFSXo9/guUmFl90e7O0HtNZQ/sAyb3zY0Xt389MP6HI99nJHDOG+dsLIYas
eI2jkgslyID3cQEcFdT4jSwVbXD2y7amjWHmsGgay4XiI/V2858JGIwBwdKLNmie4sQCNoHDNpbw
hVAQEhAjovL/K6JeTLDyUyYzYA9NgOkpxSYmtJTXBBVqRnI60FEfHwhynVYols8lLnWUY1nIKGv/
OGjqgn7slHXu8N/mvwUj9SOG3Y3Pw3RFlQl/vuG43N8F0XBkXaYbiKIGn3OsCU91SVqGLYepokfi
u3ywHY2JDs6Pr4UJ6M4WfIFbsQxWQjN23pxHagqCWZUgesbb9+bpEJOWgs7O4wK0G7FRevZvHeUz
/SD2xFWuhVDkZQQ4nUXb/8esZdA/64hYkeQXT7TC3M8Ou66BAozoe0ClwoFe52cHkkSGwBm71+Vy
bJOBdS5CAOyw7hYpJvhFsI+lG+oh3yy4Tv5cHRlKrtaUpxGFSjJwaWEg4O+us9SbbHBa6ndcaXO+
rWb7bUPVTYe1+thq9tJ3REBwQtTPJfi3f7aUAjxRXZGV8JzJquYswrOtHIAWROhAOHPEK7Ps1/TK
NKFT4yR8onC4gOTf1vR9WWmdq1RTOuayxYNTGFwQ/4FcT8MKffE41yJwctfV5m0z9E3EQh4I3WFk
RU6ZwbjogaV7CV/z5NYDYajEgTxIoauFnXgll14ubiFRFVFAl7xKs7PEofthDrs5RwwkOoqwufcf
IsnmHrR3OBkAvGJhW/CAwWMazVrpKTFSxydqPIhy+unSI8/WL9NIZzhqg5DFzDozujgFzvZNxSje
hrYSHUW07QCpxJ/XwFiVO7QqtjFuMQ7k4iV0bWMiM8lL4RDHF6Vom5Yif4tx6LTytw4y2ZDMTJX8
JA8LexSfrEjIQoR4YRB5GXWec8OG+/Cqy+9WATFU+qMhsiZaa7EjtUKwyFDMZ/j5W0x+JWnlqJ5S
raTJmMggWoCqqiTVLy1WMXD5DLzp5kOeJ91Cv6zzgBnA3Euk4QDFIOI6HzBuVphXhsrWLGAfoyz6
4qS1+hahQi9dfcHxShzOPuE0C+C/GzurNDdGvrzt3Vtjb04Y8jt9DNiA3f5uc1kPyyAzdcQuL9GF
ifh5IDhRiG9NMIwv3kCx+0Pmv5qxbl78GvhSB0iNzQ4v/rceeU4NbsdKLEWMVEsX7yx/2IVPyxgu
Y5Lvha8V4+jDxw+W/0d6jgFOfu8OnI8pJaeSmWO+hWy4ZLY3EMtjE5dfLqUcWlHOQGgp+p9ZAZqL
rQ5tpKjKFu3Aexwzg12hA73XKNV2XTaHCITBYEiffFqjkykxlLk6vQy1yGW7eojPaLEtjFrbwhNT
vf6AqkmaGSMAx/wrrenhJ6GCnNdkyZqZaJFLx4p4miToeJLMH0quEekxYJXfW4Zsr3fnfT639HpG
haWjUFUfWDLmhmpSTejfhTez06sNGrPw7sMY1z6WWAEEc1i7fuxe2kh4KNVzkhMbQva0jeDEK9rV
D7VVOYrRm7GUNKXdkHxhk3SahQum7aqRTA5roh1PIvhTjm47xJgQHotzpnOOJsiR8H2YWa9+izYw
iVlDJ0B10PgJmvv8w6HOZE2jbO/ezQaikRBz84PMUXtBrfJT7h0c4Q2LSTqTmcD42o2yeNJspHJ+
IFgNcdTm7UqE6CR7Ojh/qs9Nk0QC358tlbq0zTGr1nbHSHD3qmIMrrfkboeX5dnv2nX2utFGQwJT
RsFAbMfGSgbqEdggCdUNayS7GZgx5tBjubZQa8aIw6BNWkdTpl0hGvfFJw7+FHFM6uFARiLr3GcH
SLPZZhwqNDLrAqKpsv+YdtQVJTWZpKWf8YuZkQ8D+oFRk3UvT1Fd0rbG49oLbcQAUCagTsUzJ28M
6N04j39tqTemmKZ6bCbkLv6KIICnwB5+4wWSmINCiZriMNbXB+sB4YnEAQ64KcyR+Agofz0EOm99
b7Slufh0trHG5vBcQrMQSGIyLESa/ri8DDZqp0JoDZJFANXSzmtjrduIngdkRo/BdZ+wBRoKXA+U
76SiZC/rnetEevVPup4zk96wETZF1WCXMG4UzM8MQFV2avn6dW4MNAUxOfDoOZBZaAfdEaXcPERJ
hmfkIUjWGi3ySBYgwyPGB1EYcsUzuk/NjsLX+ZeJzxgubUbl6O+f6WcnOKaJOZ6fo3q9O449nB8g
IkpK1EFwHywb6Q+U2SGYAAOSDXKa/Hz/FM2GhdsZKwNizoENHU/fr5krOJieh8SeKrWZRhHd8mSu
AZtT/muiW2GfNRoPgDDgLMHhChqYh0H9IxF5JZBqDH5iIuXLP4uK4BfMI9FgaNOyCBlUcnS0uRBf
k0xemp18KeClCjh3Y34fhmvZRAM2OQV3l2TDt7zVcf6o5+93yzGASO5Eep2fP275HltJpasH0IaZ
2SD6u+bJKsvuaRoqFPXpG2g5cBojr9Qny9jbNeXaL3RI3Jxcg/SkeAdP+Yk+Q8fQgCEgB45uF7PW
XVe/niItNz3M3QuondnBUUMyrLqKxDxH1Yk2AasOgNh+jX5ivldCidt38FMMn+NjgmgnExfjfqO1
hUFdD0mBJQLOhVESwGOwq3tsWOHXuix2RA4BfZKTQLqG5OnVNxrTXnCgSBrhpFrovvbW1YFIgi/g
BHc87OhzHtYd51lOtjGnPMoYIh4hLC5oYH9KSY8Y3pH3oNKIMoPdrH4XLuFZJPEqPXNs8wMajh+f
tyfUQTUkFvuUQNeuUOkoYkisuqSN+L4TFsjr0nCWI24vWcy6r30paclqMlC4AXZJVsBH/0s7myI7
9WqPFsZ3OOLXe0cPyjK12xRVqIvWZD46THJrwSc2FLooEyTOuOP/8xT3V6/Z88DE6iV220bZGoEm
3i3qWkQCrOvAFqGKXbxkD+CHE8NcpRadPr2BzK0ixB8wZOZdkTMflh9O2pUwKaNB8xH5IUqPf9WW
XNtlkeQGFuO9hEI0waBcAlPLriwF7Jqh0rDh1fvIHPX2Wp7PWlVqtIsXcs/Z3fPBv4aTjN01G8tq
bZBypb9/lmfvX+vpBQj6nff7So7dME8y1ZVnQNBhoELsmPN24SeLkRzPCaRU2kJvSgh8jKoK/MFd
/0Waq/Lm5qR9vQ6Y7AM+PahVjufyPQXkB5zKrk9nTfZleVDmlr33gQZYIoMZ+nbA/8GpHC62qSYC
RLeb3h8cNZ/Bb2MEIYdsdlrbzmUao/itHOT4n+TPfAOwr1jHOYfkdnLAwENovCKk4WWZQTREPkdJ
azgZ1wRvgS4udHIgm8RZe1epLpEVNK3eJMDV+ZBx5E2ZcCu5T2ciSw76w1KeO7uS935tCl33qOOf
bYAVBv3EUybQvJLp3wI+Rq4+at5Ucv8vcsIMEJUS8f646tgl/2vvcRoxg7Ag2WkVcgP4F/0kLboU
iqgE88bikcqGUnp7WWMNkSH548HXe1bDYEfZeFyuOZ0yKxblSZorkBaFPnVsfXXtmaU7bRkmKs4w
iD8oFaY71sug66YfUB1g5F9M/NeH8Cw3DAtldFHOJNmrysAKBOdbi0UJnuI0sH4ZG8b3AIKzJzxE
Qq1IyR4lVdQ7E2UI5HtJkSJGKxhB8uDC1hxeANV3bfWLunBxRp1RCNBXC++ILmMwhxU4epiK3IFp
CrXdoY0bsl0HiSB/Oy0GS/sSlt+JYOrLD9510dUsO81ftT/ZdWTX433Wc0FibgWk+LmcOCORHVTC
wYdcxybvhhNgWPNKK94mTl3sstH++RrcBx8+asYksfNKCu3wKcqC2oEri4VS3hva2anW3Wg4OOCz
fL1OCDrn6qkVYCdKuhgwly9ER7k4mx8wA6ItfrnhBBfJtTmZ4ubT7BD0LpiF0UaSAFNtMCYQnnZQ
Z20ttHCI1OJVqKwXC2zceJyF9lPaWmLIEM+kujzoon/wIEt0CqS6NaxNKoAV8DHCrcTOXWpF3cqN
sLZ+b++WPnV4yTgO1FhCb0d+09bxeg+DGsgpmL+5TklPRIGTTfm0l9BESEIFkUT2JVa/RD/XlCN/
M8vawlpf9X9veggXwC3BEDRvY/DKRTHt1OBoqXhgzWGmDJ79qeyDSBuGxLSOwLHVV/v4zhiRUlWY
U1xv0UxDzHDPvd0pYbIyb5ZQEpE6QZWFFJSBMu0geCgn7UFC2q/QNyZo2X5hXy6DXLJ9auJOJQ20
69CXTkk+/IQi4dZu1PcMUil4sClJH76Cy+0kJ+fJ+RfclCVV5jGJqgVqH5IUkrFhXaV8X7td8dDW
4vx0zGULl30Y/pnOkhUUtWJN3TnCtCVjqwARN63UWFzwBxIwFbh/GMgCSsq9CF4Zr67h1na8lKtS
eZYSFoO2UcsQfAjVd2KswyYwbjkcWAG8BAHABPvIDOlTm/u5npBtNkS8NPhR97uKLeTmPoba5uuI
kW/vXLWxICwTOLjUv0RVZ3B3Gs5F7HtqYH8okFkxz8qxdShRxlG17iPV997UnSnYn5wmfhnr1XvE
eFJTMbIeHdkEknmfSa//gdyohbJjwIUP7tMFlOAqLaEYdui64nOR/SzCou9kSeC5E1Sz5QbSNNe8
+XLafx/sOtaUo7xN+x+K3ylFhwgu2raiK7YKZrRilrj25gzx/f0ZubAZShnrXen51QAohj9RR98t
2rCp0lOBBuYWlpkGI5MizoxSiP/yhEkiGdcva/iAJ/qId2VUT4eF9O0cGwEzSuD0eYzfr0iPOfKD
iDOjf1U9cQ5tBn4y28WehuwgDfBrpDvEMFFKhQFXM3EyENVo1062Nf9ueIl1OBSHFIJGpPlF0PId
syQHY6WZJOPy9kPAhfsb5SQ7Prg+vv/qGPF/63JAeLkcL6FEAImWYwvp8B4TDlJgbX4KBZGretQs
Yqub8uSCt04N/XTHNKNsuzKQiL/yN5LQj6kD+7kqBwNoQz8nf4pasjCBCjOjDiOSdlOq/m/fhXZN
GTsopZo1KHidsQ1ky+xucS2mYESQfiiZgINeMXJKlU8KtT9QNziybJ3HtK2+rSMzf2NKt72cEHas
JB3wwCEWgW2JYH6qKwgXPsPbMhGUoCXUxRN+EllUUJc15EF+XEBKkFhCFML1lebIKkPoy7B/pue7
4R7Vv9piwtrmvke2i5tYK4kAFYoMJV6CA/lWFYC+YQ6gvGLzqfaWvmFkbuGpqoYm+OnWCbZ1czYG
/23gDvqMmHKXIHosi0Y4YZyNVl10axhtRPQWMU0J5knicGv3KojJ9Z4izG7J8ss2XjqY5dY+IPO2
jdOn5juwpOvUIfPHjlFa2It5GWUXr2APPLVfy6EF0/cowXHsG+aeXOf01ie3gJnw1nM87b+sOk7H
8Pr/VhvODi0Y5JNozeWyFD1lvCpc21t3NoaSLQJ94ESDFnv9sWeALTxObPySEFUVYDVdeMXZ1Ghf
XRbrS7/rzXG9CpjxEZy7UaW96jsa8U+Of6lyLIrvKuhHj99QfVh06yigc0E/Oqy8oTgOyL+lVW76
P+brgbGGhplir2fmeP8xMTod7NcEEVmDvn3sm1qMGzyrf9ffEE+UFfDf0GWKGGhT1JFNCcrTf5iX
bFybAQLPRedUoSIz3qJAv1wvV8TKsF7Rz1LGiLCVIYY56wz/NOmhnvPvwUMeDfitYcJeXIwNS7kS
H2IfffNCxtzbkSEViOvYpJ8FbY01LoTqB/r0eSCOI7xhxuUjqRvolNe7Wto3wcDp8jfkYDHkwLtC
5ypsTinXsVtdBXtVlC7lc0jgyR9I/TIP98ZTK0W1ZNPenGfnF0UJ8Ol0krn2e7ZWfHnzcEi2kuRg
6T5KN+G9cYCL5A3TWwRgIOSy44CwLUoTpBjb5NhPR1Lq/1RXEzwB9lYFuHNtDxxaMd51dggzpTEP
81fJPMJhZiiPVCTsDR3uijdxKzz88m10PSI6F/M/jjxx+zTKkMCJ9X+bLunA2k/X1igA39NRRrxg
HU4N2HUPBjjviEdgSQdQ5NYkTV4t66Ec/Mftd+dvqL4Sf0SHBNCquV6SIKyD2hJDaXg2Qb4Uufgd
FHzER95Rw/+Sx/OX81LOA+6NGbHXfiVdpzCNkdO6nOHpepGwMsojRbPvG2/y/CZvJX1IZiTnK0Kc
eplJP2swy1uwRiRzyI38RLGe9bhcABeM2VvpwjTMxGJSKS5F+g4NiEsx5wo5BFcRhk5a4bBJkyf9
xco3saiJbpBFmVqGnftFlbx0dzyziJMQfdHNPZLIti4U2/+frnJ3sxZyj39qVYUF7c4dBRszQlQN
JzSTVrk6t79MRnQ5n/ylYe5jWVWgaNgDehPuef3go1Ur18QKoqZQqiArx4ztvK/zkuGioB72DRF/
ieO5zyFCGaW/zCN+vi+60eQ4xeD0EMKBbpfQNPGxBHnopaZb9bfc8aZ4XbvgNG6ANmRi/CHidzqi
8kFQa/iv/FRwMXOupO/HxwZQ2luuKPeeuIM7H8RlWLegDRIsinbr5cMEDlQS67BN1gY+7+Ixk3nd
pTlMn4JaqYkOxYZxohutjc1WcLAoaQl04Nni/EC0Hc1pc6aZnvRPqeBUZzNAVSjlgL4XcsPq+XUv
VMt+ruAVZN03KojVtpq2Tks3Vt0gXCpM8L0nk3aXhC5m58U/zY9VKcRUuClhJZY0zk+rnh7Hodv5
c68yDRyPA+Q8LzYJh0x8uQu7jDh61zt7ToYPVVoKpUXFIl6TqgStQh4tFQ6wiEJ3eomMnANz7eX5
QVwc+A7OEmFdYopOtBy5vIVQBkX/lZm+JtQi4hLSxuncCHgtyFrKOjDrx3cqRm6esQDVppqUkbdI
peEtGxJ2Kx/hkb8V64VOk2EMDcSrxz4crNPiBWf3Gl3phjGiF5Z+CGphIqGNLaZDy9Rb75DO/Veq
GNGbF8eZCr/yZCZPaZGQLJ08Y7LAuKZW9Co3d97r3VjpPPTZnSP1YHVm2Zdcf9y+5NZ39S0wOX+y
vqdn3NS2HqceHPZLBT3PmsYQ4kXK1C/r0uw5E4D1NXPJ6lA3xeQtmSoeDlqwfB379hCHkIDyu+m7
CgLcofhK6MKVcUmDSm7X5ZMsqcbdzXpC+bRi13IKodJQuKpWXN2dhf3RynxAhGONG1YAuves8qSl
7j2tkjGxi+O37jaLAG6l3Vlz5wJb5saruSpeFIIhMHIq97eYy5TWgUhSwqQ8Hqzq0sOWB+gX6ilq
fNhApUlORrw07pf4LrPywz6yDJ3t6JLLJiS3v4aqHqW8W+Ldc5ykdtdo7DvLky/wN2ywXPyCdI0K
qx83r4CVws+pz+A09cIonDPV+juKnx4teo4nc9c0cTCtb+6szl3gUyjhJ1Nu8vQ7LJVmw1F92Tpf
9ukZLk38P6k8lMgtNSnjm52Qe8tyk1qeKsp5wYgP6n/PrzcXAPs1TvTo8cOzaZw8YIbPtkuM4OEA
wP9RTExfnk9i8MC9WNdI07dvZoT7hK3a2HUNegtk9ItLkbtPdvKq2LbgSODCUWmMWihrGcxnz+G0
XxZG1rqKHbw+zUBQINHUvSP4ODQKwHaEnVrZjbIBfdv0K8v0Oy6aVF4eZmAKcB4RhFIeSZBtLDHD
KmU+PKceLGq36GuJJw71aPuqzSVrFDzdM26UmmFzvxuihPrfTDtoQMwALNq5Zv/McsiMs1rFtXO3
6Qxqq4om8PFFAIgKe7RFpKRRMBYzdDKKwTNEXp2fBwvI8Z6gnASmtRv7VuXl6Kd4V8Ue0FunQmlM
UwsiHslkdTelYqUgrHGWzaYepsV6CXkO3jIn1dGQkhMgC5G292nPTNg1FVx+BM47M9QfJxmuuu1d
HJyWk0XyFqnI9sH9VSAG6OTT2DBiMO6n6TdydRy4KvgsU+TxaheEqKxAEWxVlmsOGuZ97J0Y4evD
lQP8vxLzg3tt8ABWPvojOOXIzWpsAGMqozk2A3ia7abHmAcSR60l3F9OJLNG15HHdGjt4jSvlZ7m
yyGwKQ39iOblLWebJz9iR9N0EiWcbpFnNClK4mWOEObGwlpDJQsF8WtfsDYEHxsXu8SD6U3O1681
1XtO2AbUPU21Rop1xX5wTTRrPQ+Sd8t2R/jXoORXIh6AV9IiCTV80SgQu2SbVj0AGNg+nv7K4v0Y
9DmJxqvCUfgeOhv8/mbkUl6buzBSYTJzJ1CebEDM9RpMPfBo14NFRhBptyTFnCEqROPVw6wRoNS3
dA+BtKzcfybDJmeP2/GOnGSW04gV9o4abGocxT/5OcemTiqXUR/RVYkzd2aZi7yG1LD6MQO8MHOn
qQIFZGeK4EyMhBKKRDDeSPvieOOj/4pJLZumMlg/W4x3BwAa8Id2LmhmhI/CzXSywbsLIW0nFEQI
tx4FNSQpPiq7iivSU+yB4MivLA2SrwFRcEgMFWJIGO+SWznJyRQczTumZjg4153RM+uulnRBv87H
WR8EvD/8EnpKB9oO9orkdKb3oSI5g6P7VQDfwB5EWPfFUi4/xpqoKLy842AH6q5qc2wrAd5W3zvU
13FBwKJWlltGJ1hUs9+HR9gzZU09qD3Gg3hN5iLIvtoRyAmDcNUtjT3qxfnrRkKf2h09/mnUrtFd
hpCtOVpypPRKz8D5RcrMe1207e1VvWyFsWMSQEx92vuylqZ4R7UR7c8Ul/JcKPOynSPIISttjmyX
ku+8DxdjJgzr74/47IXm0ELyutX+yOpJzHySKghsty3Z2f0hNjxYXGzmJktFvAEZJ1lhviZY3hBo
w7BIWWBretpVF48ONkl44I6fzS85VnJz1hFbBAW51eQOt0r4mY3iJRR9f814ysHPkjkY8CjXU+9o
Lsdp8JmMcenClifDr5a0R+M10HS7o2nhkt64YFATHAPuUX65aBJdubcEWwBh3TZuPiIf6wJsDHF7
PdbK0eJU1i1knOjPgcvgHiXy35wUThkH0eu+C7GLk77C6AVYIUEqygl4Tu9JHFjo/P0Bg3lzT7wX
NPqHLIpEqcudnB6iR11bK525FR1KzwQ4vzyqUM0LTXVzUYzt8paupO+IYbZSv2j0YiRm3MMEhEXL
rB4JeyMf83fPwUmujMqqVaQpsK/O9ZWt7ChkgOxsZYgsoeHLRJzioeMLPOR+XsoCMUsNnXIWvcwN
SVzoLSPcKy6K4P5go0oW9HLGdhwvQUjA099EjHDkbyqK3Monhp36g7mGrvbtWUXwcuKejF3boD3w
Njc+/cgwe9iiVjMW2YssS4DVqtACD9SPOmKARlKS8bTEH/YvUsT63bS7d72NWn9bQo9p9i+t5r7L
qNPKFrU8QKxEAoxtDujz8cwcwuPAU2oMj4KCQGjycFfvUpCee69y9XXYisbM03E13pGJNBurBmt+
Lq6NfDC/z6UifwDCzZ7VVYLBYtAC1bneIUsaDvFYKDMGZq20U2ipd/CPfPHPr/xg5COWixxfaE3S
m4QPhvu5llpwUpBQpFtiJCOuhgICaLHkJe99lo0Ibrza8uMWvYBfLkp+r6fPGOFyMjqpv0/ng4r9
oC+A2aoeEeP8mJZk26xgHr+Anz53rqNSBmae27r/akEzvuvz3antP+gw0oKB34cQaPlrGevYzoFg
06lMmHEIPBntudHrLaIJqTgCjl4aKGv8GWHaNHLvPXAIDC38/U9FpZtBEchXMKF9CZInmVoFVM2G
czIkkJBqaPCka5iwOfzTZK6VXckXA+UUtqAgUhvTwoYw9HGWmQw+u/PAbrEa3xBW/0mATLZGDqP3
AZLOpuk3r2rszGG2wPfocwQpRFWFo9SlRr7kVo+3RKn7M4Ozqv5TTCwshoAsAmaBN36reaeYPCtH
k2FhCeFH0LceVFwdIkv2mTAHhMjL03nABR9GUKOrrapZv/5Yr+WzyER2OZBtsziYll4K4B/P0rVe
To46tPB7VcUErOfCHrkQa+Wla9iFbTQ0maK28AIsRqruMuGJJtQmLjcAeNB8n8p1843S3FYlxlwT
ybKZVYVnPHwT0Et8x4ZriI7SYq2x1V9N3Fb28D8GJs3rgxFjnl07YbKye+ldf4rotdDNyXUtD5ve
Sa4E6eN5QlmUiWuDwFQuh1FXnHScgHOheDag3kVPBFI0ymS6izXBWpwmqmIIzNx32IF/ErU3navw
gNwsLYLaW2tKpC556uiNZn7T30woOiPKT0EI31S7ETrWJ3tE2rU9qZcP0hfz+RAaY0DrAQAXI0ax
g2VOGckCIFEb0GFoeKh2hthfLtRya8yG3uHldPi3ckuwbziWnPXWuMY+JV+HTPjMGsnbylG7n6o7
CpiOCgxh1ETz3rWZuqf8STC1bkqOnNglDAwZm0FaV4FyInj+ZkXrOiSZ1FhfnP5aOGhkJE8lAMd1
uehYF271yVU0WfqQRb0fvXLb1Yy8gQFtblZPDJkYA7Nc++HjZMw/iMFWPalrH6J/U2TJmI6VdY/i
s5Dx1z7DX2mIZW555BOagPwxR98khwxfa8+C+NpKgv5sPvsfDsIruwEBFe2pNwJ5MLqcMYwRA/5n
sg47L/LrDd765v//db6w37qfLpzi1BfCB0n1qVo+QriQeSVawpFok2FDblNb46iTE9Xs9q5BZweE
QTaNLGAtrEUnkJh6gU0yvbPZsX25Ut+bB9+4aTetbtKorUi9UMkccaGWPDOus8xLgDkMSPvUfZu3
fzxeGOUM6ybgrWQdbxre9W0vNru3fh57JGmhJ8FX/38cInJ7dR6Dac61XJEVFia0W+lc5AKtqTeR
CV5MKvOYjc/InrHoifNskpf1rOktaJzuXZOC0Gnm8DXdAlzRAdDxqDG2SZLp0blauNKi3e8lqeaL
vi6v8/5dUKaTUb8Q0uYqLyNuBtND6/Kn9c6wDh8H9TgJsYjJd++a2yjQFXqSYhifLQkGSvvFcB2S
anI10VBgIDBVY3NOiQeuByqIC94WdbGlm3aY56PDAgHjhja9F+DMX8iRBUn7SV5buYv7/Ob+0VTe
Yr0Q3mR2dlYfeIz/x6cyFd3fBhbsTicMAgnUfa0sLL5ogyw/55kSYz1hMcEYLiECQPs4njz+s0CU
W75MJbjALY/bIHJUATCiNpivz30KuZ8oxuSm/dvz7LDXSSebfAsH3E6pqvPibW/eSmTj4ZaDV4du
nc2uupuSzzlvhzGUA6fAJKCinAQXpvjAZNZm8i6zNYUEUv+IiACcx1/ZAz+QhfNSCqqrbe6yjMvp
SZsnA+oIIHL+qyVWu9Rby/sIh6Wnrfw4fJTsntaOdiPmLJewwtg1NyXyw+ddhEQtRY6JE8X4a81N
oqAYbmV0CqjNa/MIqn7ZoMW8Hg3IG+cQw4Pmbh8x2PfBn2zC0g+9v9PLn//BjMea4sCoU/KTPJel
Mf+SLIUa+AsmNNwGUYQjocEHxYEAVNziraWq26ofCaHLYqUVtC3TXfz/B0gSwNusJ4Fm5nQgAcMq
9yQfgsKCpk92QCeC/WGiyu4dFSPyeZMLLFh9XGK3Q7x7lUtoJZGoQK1QILsjqxXgfE67JTrI2q4u
LSUeUZ/EVO1hKas+1MJMio359jNtxkmfUL0Q2HAZiYsozt/Rll6fZYtQwhnNRHVJ/VkFFHmxRAV4
CNjVCx0V/pAWNpjKU1Ai4+nkHs/ovHQzXK3nW1J8O6gkSCnxtpTNh1P+G2xrgsvHAHWMQiLzU4K0
FeB5FXu5z9r19BAHHaeLSmG54Kf8qYOavBhj0RdnTiYllQeljuAgJUHoxd6yRpYa4tpT1H0kqL41
wnCBtsGrPWG0ZqNM2qyN2Da80egLsjtzYGKQSZz/n0K7TylwFZ6HoS42eaWwql9hwKigI0iFplAm
+N7CH6rfXKW1qyNvLdCHxByKVsVq+iBvlZjCRKa+/PjDS8YmmOM+qk6jJbLVnouDgop+V7Bh5rVo
O/pRHYN6q+8mPMyykZnLDLCHsDFIgZBsOU/0O4mceKsAaHWw6f/+pm9WcJEU0Q+9Yt8cQqu5m+bu
x/ORg1DHq/km8L+kKA2f+Sn0p9jnqVkQpPy2n7UUuKV4bEUJ2duvypWWFL49JR2iz4ZHOld3Gb4q
yEZoN1GtFoo4LeLgbJBLVm/LjI22s3ssEudscuQHxygE1T6hdcxnepoBoXbcq7y6O3IfZDG2voYm
D0Mrfo7p1zUzXiE/T+Zo3m9XMwWKVt+LuMvaKcjAaFvVgxEEbdG1qDEVexWyfuvG455i3tMFhweF
mTnnN7ToWcHtxTS3adfTRSslMAhb3JeSqQRasLeEvpwmmxkHR2wd9wPHn6F9Vid+2wKafcouyq00
HbQiPP5JO/QD3JCJ7rqHtCqPSxl+W/i9gWuUl3p8K/sOIxdDA0SSDYf4XUxovmkaqiF9q1FNfcMM
/BK5EzN6JR2OeLR51eviwZhpgpY3oUB9B6ra1OXc7YHAU7DKF6fBo4wyKmN/+yJ2jA/wZ79V9Shy
65TKEq+c74AaKB8OjDlcHgkoY4wQPsWYllswdpWVvtFe5HVXG87a2F+rwyRynsC5ssZSbF2PBYyz
zXrVLE8tEe2LgZogIUsgdZyEGvuHLI0eLTtKkCMLHhN45vGWwJjgQlYvLjXapTseMQ63f/DJDZeR
cIf2zpeyxpD+l4vLXiR6KHzFOG0+aVbvG2VE9IIoP45VVlc++0Si3s+zZS5FeK1n8MlYilRuHKm5
lFPjrMEh4PltvTH5zcOF6LwTXitAdi4IIns6/oD51gcvGxEGR5KIAIGeaDcuvVmLQjGUu0VNkczd
kwFGQFyMOJ97WsuOsWg12ufghdjLPTgJO1gO+ji8PeNkJdv+qlNN6TV2wXy02qCEjJ6RwCH5gish
ALYZUPZIPs6uVws/mqqumBzP5aQszVEBBcqSpnO8pKRkB99LFQmnUiDngaT6mHES19tV8cE3Fylt
3mrXljbG+Mt4qIfJPz8MsuQeezIEmpdoGFvY4Yi+pGbKButmey4cst5bQXbGDkpx5GqlSJeKBj30
UDpbwvo5B3nfAq4lE2rqDWCftUk2Bsw/UqSbrFlL0khVsPWTNgVsxAXx7l2YpI31vDXDQ4mlYovW
nNXOTw6QSa70WX6G1gOhmHl4oUHX+MAmwiGhep50mGrYICYC9UZNiWgDVIgA+z1xmVdd74/Oy0gr
l+48ZqIAapqm0YLcBQ2ifNPF7GD3UEfjtcW27tfvU34RpT21e7sR9krfv7XqjSLLsOAZS473JvAM
Tcfp3DJf1CZCAC7eQ+PwqM2lBZ1j5nANEyrAHkPiMY56GcOKWDrDFgk6Q1zO3TsEYMyr+9WCVdG6
yUG1V/txCkWfPjSaFcmXV3EeVMgj/c9wa1WLjBovAJfgIF2Jib1+1IsNwuA77Z77Gye1FCanxAkd
/Q3yDW88pkG/2YtBXbnVVnBqtnqqT14BUC8gwp/aXyJFuVeQ8c5zHZS71ih9yYYblauEaidM4Z40
ftuVCyafvErlmRYQ2eB1AYlRJl2Zxuys87tJ7N0DStoZNzEjzYb5thYCVefRzpJuvO7Jx6l6U758
xYRIjrJzbRZAVYQFJ8lEUjID1Zf8OxONMuMewg1gwV0cxO2dHyy7uL4Oa4y8A/5QMPHvV6wy4Xp0
/C+MGXmnOS5h7vZuZuzvK6N9p54fG+hcOIOJNuxCq3s7RwaxLyVxY1nNIJS/s8ivkt/X7l8UNxX5
ypTsV1BgKLn50a2C6QVyD1QkunOCwVWOC6zB4YWOGTUY9tcQi7GIlmKqTKqHTUO5YvFbiIyhBtdw
nmHInGA/q2o+TGsI/rKeINxrlUGMUHG2mvW8CM99ZlNqcOB9Yht8+TqGv1YAKLn+kOgSBKxpUcv6
ewZIXEB7Ux0YFh/Qq/J+2stXcl2aArx14aL6KQ4+jN1D94cb5YlBCnOzBsMv1Sp3JSVKw7tto0/D
pBbBfXu+HmEryeNessXU9Cyb+y9hgLod7kBoK+ScLfxHtM7H0vH8auR1AD0QMe8MtOwZnzVJ/2y5
apSGBWoAJRhjDmxphOunE0EFl3H9e3GygiLQfTR6kir8xiSgZD0yOXgdIp2BWYUOsLqLhPRYFdW7
3QT2odX+fUtk/J2syTY9Q+lWssABsqZ4i6eZ7LsciFGvzG94Xou+CdTZFjyo9oN0VH3b/ZoWNOsl
C7eJ0knPH5La0nagcHE1lSI61sdiApuB13/umzKwFfX6Q/bLcIvsoSwo6LsTscFba3HdjEfQIiLB
Sv1aLRLEm1S1uWdm3fue+QynJLuX7OQyDqEhZ71dWbMvjPaoYnRcjp++phwJfJtAlH020TGv7bXl
0n0rN6ok/3Gt6H+x29LEBV8RpEKIOPVcheofPa/UbbGrNLqRR5dD87CT5h1WS7lR/5QkwYqacBEs
7cradoRRZqiDcg0BFmOxKn1y68X7P8gShREFhriiy85DisT7ecP8MsGC473GHVSG11HTbChkqSk7
k5kDdpT8YlNHG2fMcHEs1/BYrfH8PYruWqQAfbtVIXLt8UgLk0XZzJD5QxFxKQ/NohcmxJ8qNznF
mN+86IRr3AIs82zXfVqjxSx12ubuRh+sY/uWGym/umg1pPCAm4bI0+b0ycVciVMRZoc9vQYhJb36
Yk5vMMgU5CUaZhiaTeixp8XonICQvXJfUGgFNMucEBvrD/KiuqQdXlbTX2X7dkkjK7umxLLUh7ey
+yCe0QSdx0G87ZJQJnEKAQP9EpyvZFFhj3xxnXiyIVObJhpmAA1MK/XQWLqyqQ9E4Q0prqD8iFww
B3tsKZgFugVLRtI9VrjeNI9wMtabto6fx3qkKkCKkcCn1LSxTcBLTyL4jQoneu+Gjso1Q2IGxvmu
DZNc6lbuQlQd8YX0z/ewv7lbUP8WB31m4ya5xnnr7tbJHVvoXSt1k0dEdrZWc7VCuoMNV3rjYgZq
FQ6CGjWXvX8jDG54XTo5eYDid3hBvW5T2HN5Y40oQ6RghEGwB0diiBMU0w8v2EgnmRJGKfN1zi1r
23p3Hh3FZE+uHxFkXu6RBkosGq4RUwgvqn9xQLkCeVcS6GYAk9x8lgdmpWxFP1kOAAvMVELVC7uj
HsCz+eGpF7Vm0vI6UQxJ0ykwQUDKfJqOIYmy8YOcTShymrY1fbTIDTHh07U37U4aaK0O7GJA/BzG
V/IVRmOvn0Wdf6q6SIbpTABtLg8XEzW9InUlciLWdjncgS483HmS0zuEzosBaPyyJj8p0Z2tbM15
FlLTj/huz2PILZZ2nf5+GH8BbACB7Ddy+izBQknkh/sTJHhsEnyonCjZiEmwCtos5ikh55dqsIPF
mNhw/nOuvDFKjny94gsGAVUpmNeFWVTHrOzmh6AspPx1dn8p5XL9NeWJ/WYp+NJscufXywfrgVKm
SN+eqLB9qKW5IWBJNWCyX2fe9XNKXYGnMoSxDZcHwqy3MMFriH+J7jxNJCYu0/lfiZ5FQoBroQgm
2USumWoCzmyZHjgYTCTO3agNbcmrw9p3TWiowdhoJ5NeXc0MwS0F3O5BmomIVDjkWwMBofdgtn5a
lXV0lzc1RVYffnMsN0IFyrFA2Azm0WdGmesZ+P6YtgcJYOGNopbOOggcZqObGmpQXbAwHVGZ/5rx
gjAaBJojFsCRXnSPTw4H1AJC00mgMzZBaLoQvIrJMkhHoFc22nRy+6dWLOU/BA+bhZDyXW3EUznm
hOW83qsedAVV3q87/DNf+HR5CY9OdhaPzt7AIwkP3TyAM1m/52ylkO/PR5TgizS7w8bhhm7Vt72r
q4J6vz4ClHJvp0pOhRJMYckQEpb6mVwW6YLhR0j5h6sivj8TRCXYZdYPHt/gfdbi+fQbVHHrv8iD
8wbUoKHncVDkm/5b1VNA8/R0kp/DiW3mMh8lt/jAkpxwtsGIexA79H9oEHhofoTrzGNgJCrpPjc1
58k09g4Ej5JNG4RzLvHKq2CQ9eCCNzPZKUk4wC7i78BHgDqpxELNGoFY6WAabU4C5PNaiCcD4I/B
GoyqnrPOG2PoSCp4ULBycy0sJtfDsCpmPSxaRwKHFppIzTkAG130tJNKq+GfezemOQQSOs7/DBPw
Ay6+cMAWIAaJodyV4siKSU63sOJUfGn79uj7dODmY0DFMY1DYM1mKmcfY5ralE7PTnObffjvT1UY
p3qNyLX+O413DajZ2NrvZlTVooIUfXnpbzRWoA8ReptV2zq9121sTEqwU10glNDHkbKRWJ11NeKw
Z3hxy/YNlS0nukMTOduljheqxx83/xFjoJjSJrjc2rrVDlsLnonTcRhXiekzIehfbLFYhAqCgqTx
F9UjMyy50YAvHEEepul9GHmbT3qD3pmEum5swXTs6zLlhHE3vY+6xHIct14FWJHLTjOCTUiZVA3B
32pLqgzom2ZKnnPlj7iu9rmhUHivk3ASNEu9zysjPhmjUzOhh4RefILHoA/JWBDV5mP/npWY9xa+
3k5kP85KDRhHTVmvGt52IdRrS+KNeBwRxD4tw0jmmx0w9ubiapeGduUgzz5NbfzTL4mkR/P0CmMU
lPuBbhSM10sr+C6ul0RP1rhdcsiWUkdgKI58GvuMlf5nufLIIscTi9nQPps5miRCenZmSJtPTKFR
LWYtjJTp2hJVrVYsA6x1hpNfCvC0a0xWCpCa2+gsDnKzNaueRBSuaaWpJ0yvKScx8peQLBHD/Lt6
J7RiOexZQsgbejp/kHbgySdGXWPr+xugHygESLaAJsLUq/bSo2mAA/QlGiUJg9kCi9YF4ofe/JLI
8tNGZAzQ3vWZrHW0pCSqH/Q42XnPd0AHQ/gNrrO6yduoJ0Okrvu6Z5v46IbjF4HRe3igPyw92IRD
DKBOoCG6eJ9fPaKe9x8M41qv7F/gt/s7bZPP3TsP8EvvdsHF+IkUNN+DBZHyj//aJmuiLUr6cyo3
RSUXtdsDAbB9J8J5MaYm7m1ki+Dg+g4Yl6ZsEJMEThVFWbPG9+J9aumWdrix8ZAOrk0vORtjOFTM
Fb5p36d++7dqOYgq5fPrNvB/gdlEro7L3WgadjRboDeQq/7jQzxNclh/Ti62TmYt7WwF1oSLaAJd
W8TCDo6jMc7XyGZk3KKxCl1ysXqjiSxyx+TTKBoas4VzTVGqKcSSBcsRFn4hYICqFwIlpR0IuAHJ
nWJnJA4kzJlAYVz7mQL7RBlqOr0aUXlxEHtH0L5izj+HQC11NYz/mBCo/vJeI293qy/P1R8y6UCZ
armiiGHjd+mpzGJcSkyTEdXMWxI5aIBJ0+C7ekpExaApusC91bChgP2FnXJtPK7zkyekYKqOvjN3
DlvsmRtLIxFxuJFcduiFf+/bt4zKKVb+5IZZjRn/v5c3KzMrDdyemaLgV3EP+arTA2d3PX7hii/t
V7Tj3n6j04/OTR70Ef/89SkxJRoNlj4wHAOnBWdLNcsQut7PzPEHqq58PapJ99iRegHbbzsPgyEO
C/KksTVM7sGsXoGaAqnIRMdrKbJEsidAmyKOKibEVhGM0FTwAMCgTSXMsXgBE+8dHAMVw/CpS/cB
ESi90xncji8TMir6iFhne4JFO+PQNGhouGp3Ny2yq2Zo1CjCiC56vKcnfKshjceXeywEKURT9I3U
JtFFIqqvSm0bkp/4r7Vb5XF5yKUYyLxXerqbiQai+0sKbHD7rgxtZIar+198Lae0mmI5mn4zwuBy
Kgx9QXfkLu5pFk1fGiLP8ihrwHhMUhA94HN+CXyZ4M7IVC9YVFzVMlI8H3TKrh5tP4IO8VXNChag
Q++dqM+1Ahgo2naqwJBywlgTzK4rHfNHGGqyDDM4tSx0TVXnYe48Vbzu+7LqslgCZcuAKl98EfWJ
MWa4ntnLUTtv0mJcXRyDG0DNcxuUB7D7kIs2tvz5BNWWDRIf6dQt966oVxldz4znE95JGqiXzO2C
zoxnNTl2fzRqEfKBoxX77CDaV7N9VVJvHMeVjHN8ErLaKu+/DB4u3qK80vq1dMWYDLbNJElxmvjs
x4S86tWsZ2l9opmeB1QLUJQFLoOSTHUGi9QC2Chi/uelslFGbUrTS7EWkWeXv8Gb7QKU/KUCouDp
hnrQkSEYsiJi9DQZaHy8T3bE91WbcE3M5tmRgHPamHrgPZV4TDSiwIauCP5m5hOUL0rA3yZCcViE
apEscP4Lb82a/3p/uP7PcPWkpjDouCQbDB4bUpu2wTlNzplqSdWk6W65CH0EasJcWlaVQRXZJwco
oi8LOXL5W2n8bBl+vsnMQPR+JXihSneJhfC2EIcluwzpcFm0SFnJTvSFKndvANkqIurWozCimeQa
RcDclJm3MYMj2alNy8stqYVk4B1N+hjEuXxUBVOgbAH2m+iyQhfPBIOgCoLd1LqTrhxoCHxDOj5G
5u+y9RzpGWhbvAnU3qzkXTBimy8LtaIQYFYX8iSF5EgTb6HUQKsOTjqJnXLC258JJIPeDebWlDvR
nR/9sXCEi71quVnXtB/m5yhtPQGNflsZnQeOhQlZqXxC8VwI9SiBm6vNdVQuncYxkbu1oucds0hx
FQzQq6qYMmOHdYvQjsooI8a1dRT8K1DOwtEKydOGd9c3Eum4SZ+9JQIFAhGDIvKFg62k1Spcu2CT
IY9+Abu/sKmJeNHeGXaxTmhaNGqEhmFH6bzlfa+sjI5qh9n9bVBcb6lB4Gs3rlq0OIQESTTOFVgn
/1uhdjwnMpkYjwN3xsb9L1/AAHFJgrcSF9nJxVsGi/HwrQxAW9itVx+aNuGrrbXNFkjRbTdGgMp/
nloRnUCJSYLPj3nDFW90720fGcCdACv7pOJ8MZzWlbzTTtORGl5bMThYKIYjzF1cZkZUR1TeIg7O
XKsT+nMNnuAcMRjMKquVFIdtTigOApGQ9Qz0Rq+iFgfb5z7KwZFv2R8zIbjELbKGIge1iIl6jsdL
b84Iy2YgM+uUui6ua6gTftvnafH2+pj4kdyuJbqYtePaTIZp1qd2FYuVkw6eYgupJRFyxcifLH41
g6TUGcZDYxI7itaRCYXmWipmsMtdthsul0b6F1F2QLSRSetNnmKrIgL8TcY2+CWZoqJMw/K1bmQm
ZgwUqQalKytVX9XO1MWOBiX5ThNX7RLC/KsieGCsu+3bxahJUNMzBbzUFV5SYC8iQH2lyVGjwpds
4chaLDK/kdErkmIvQYYpW4TrqJ3IFPdHXjVkRUZBTK9gqRVGiRnVDCGJ3awEg/SBM1dxhpppgGOz
7x+k8/Ongtkh5RQ5dnsbY3oSk7Za6ZfbyPgDwIRJereaazQNPeK6a7xFjzrCIPVvIj2zT896TBgn
xkkgg9FZ6NBLdIeduXxZILtVCKnBRFKiomsMlRX5zkNGWde+H49qnX4zTXBmuWhlSVeggjpi7mW+
MAoklxamXwbhD00wbFhbmfBBHyCgS5cesGXYxGg2FOORQ4LSkoOyMMg4KsNkK/vTDoW6DQI/EfG/
jt4Opz4DgHtnJR5/tGvD8muq87ykj/0FI8XN673cs83eedFLPcZlJVegtxFXRQBLQnbR6oLNhXPw
v5y6DKm3OO3ykrZlJuJWM5MLsuUPEEbLxZvHMElkHH+x6oR2k9tUoeOYExP6CQ9rRfFfrwH+xgMJ
GEwddVnChAm2XDPdbW4BfHDLxw/Vw9PUKUds0ryQFj0UHTwGJFWQx0f+JHiMj7Kfzb/SxAKfHz/4
Wl8hQMzr6UUYuUwvK12er4kP9uhLG2XJV/TnC23f6pUj5XXBO/CJq1+gyYn1dD4mZ+ypgjhaNjxN
c+peBcaPDte876/IL12n9xMYjYPhr8+Cqlp9gzlQSuAJbJUCjQOG4A7iwIyrdU0n971DJbEn6LQs
xuDZJWVlg+aeNWGNNgzZCVEp5j1xytZpiiqkn2b+WlmzLKzkTN/T+qd38IFz82SPu8ANKSAClAzE
sJm9cBwsthgtOII6UTM52g0K4QJsLFxBIYURPOOaBEZJuljlcSsaojHB9aDW7KrwAjW1k6WYEAhl
owQN6+RckTojVqVDFwJkHnJoopl97mJ8XhBxhkcJE68klyake2GieDIw5KWuBfmT/mHGuF/L4DOL
lvtpqePfvg/yCkLxggeKldQdskopEo1Pbb8lDO4wTxY03kyUCb6jJX+p9KHFTBHLzWn3CupXzE45
Jllv/ASg7U5UHuzpUt3OHcN/KvxAbxXrgGcua1nyjaA6QY/1L9vjItw6viN1feBzJkcVL6G+u4eT
b/6AjYZmWJh7P7m83+ZfnfN1PujwJgzJF7/LXLEQjB1Be90sggSQdq/LZgZhEhu7OuR6ucD2SDo1
fR0WIbuA52j71LXd8++o/fbJX0gL5doFvR4gF+e+jt7ULJX7D5790fsNLzet56V+autlwDG0sNuC
BhTuzUhlcA8kt+CF3LIXGkzHelhrnl8sJIuh9kat6r+Ju+v/F/WL6RURjss+X06POLJgbgbV71BG
TWapnMyuJ1qex/iu+/5AZlEU0M9XSyOWrd4ts4cZ/nD4s6qtaHoVchz+0YvH+Uernaesvs2EdRDo
tXxLsTkvIuUSTJUqM0OZW7gMBpOoRfpHtOAzTrV1/PN/OsDyhF77qbicMsk2CEosOxPjRIBEL774
ruhS+6+HkMLJC497wKGJ5SI3f1nKa/HsBf/+xfHJ2Omj+BVg14GT9VsVph5EconFEz+UfE6FcJuI
wRUQJzfPoWMa6TAcNPUK2eSo9XmC5dx65Zy24anSRvuB64DUiAMdYJ59AfdZ947FHpO4O3Dj2Bly
oVXZpEMQWhfk103GJE+CvrxnHBvp07FM1ao7LRKQsDK5HaMgthuhPn+Omfxr6237XsP6QuVLkwJG
VgKwmf8MR4dnaHi5HoJBAvOckJm89TX32j5YrafW5d24Mkt2ppuYRSRa+CpyVxtUTVtqJVgcv+Lz
dX6bQEHAwh5SISrJ+Qf6A0VFMpGWB01SPhrKUe6pD9Soc9i6PnGm9Eg21jsdOl2kN9auK311553w
cdCvdV5AXJ0oIllnxNWdBCwP4HzNEjV1fNrGQw/or3VXmioO0nbgB4y77GwwTnqG1WZiVnt6Nqgh
WX7OdPrmmwldfuCJjUlwerJBdp8nFQFMtxhTj533KcayjhudCqGO2kU8kZmOfXjXZvkvmCyjzGFC
3ums0a/W8OjD6alzkfGNs3fj/uy0LeP8Ax76Z5Uar0IxMYmTfwif4yI+iCy8cIDWdX+fXc7Z4yJX
lskU5L1EU+Mr3JpidG2tS96v0UyBXLhM5iR/+5dbm8Sn9atuXWu+TbXdxCVwWQSJYWmMAbXb8qrV
CkC9zLbRs+0uUV9ZhCXwzfUGuvnUQCHrJ82GepseGUemRP3Y7iMFDOByLPXRPLYXk7XphPDnFAxe
iN+0V3ljkm4OtzCchytnDRlfT7K7kWe20md/r1z4W3hBS2Fh6hCfbOMurueDxkNiAovCzaH+2qsz
cqpcSyjHRQwV+q8uBTFr9tBSXvsfc7cobNFSS8pyXuGE/AxFyNzc3vRgYaOPzajkqQfmrkKnUv2Q
lU5eRwK9nYAt3YKhSVwovvZ6k6T1XNYE7h2DNxlIWsPUgU56xTwDz7mIkZ733oOZbrZmCex41rJS
kPSKa0TM3zzc2lwbCzXKR766STt8sysoGZJw8bY2RLFcXRqgPn3M7cpBY7ePCPdR0eSwXufpkSFL
G+X75wIoVNpYEa4VMa5mXAlKnuxUYW9WWUtwd9Raa6rFPWHAzvgajlkGQBzdAQre7xfPNdj9dhH5
AGdbksA0YNppcv381ec5I67Y34xK+FiWRLYXaLZkcrARurBHHHUIcPXpV2aUDBk3RopRxTQQNC6b
UC9y80tkVc4teTR+BbLWVy0oJzdpVEsf8COClX/QvSKTp6FexQUarL7LkhRKB89jb2hc+6FL48Z1
vOREHGypTQhHW7o4ztyrpYJ5cbNOAC74YKAx6ZcCIe34ZF/HyfzY3pBulFvVaRVeGRRfrdc1q8g4
Z+0DNpGFAZkO0KdsRchGbyEm1ee8JA3A1CG3ScE+ZokoH8KVp3br6wws0Z4Ne3//oqXVx4VQOCX/
/CwZgqxOxkLwJB7Ds+HZYSi2z+vB8Plj8MN9xMx636NVbO4+EWfDhws4/9fEiuR59JWcestxYHIH
SxiDEGUBk/BoXOgh7+A0US7LGl7ny86VUk6Um7IdCsSPMyG2GvDMt4XG4hCdYxlFNRIctEUN9bD6
1iOpKjaSRFOWs2Eo1BcIR13JQSR94VYqHNa1STnTPuqCPJKh2WE5CY+83zUinliRFbEpwxBy0o3c
6BchgXCCJYNZQTZkDnsXaJe1Tc8J/lxHon41dFqCG8XUpb2H9Wi20TtvPrFTRnpiTg1ws/YJScDj
9ZP42JwgY/nkbxSQOr9DFZnEKlnW4IGjOKLECtwbrMDDtc7jRgINOLTdScBp3jiZYwAaF2E49U6a
ryWCkAY4xFZnmsETCGG4onIR1hPMVvjtcP7PJMm+y/vWDgaBokuZQL3FRAsy7lGMLacTFgufPL7t
nmky6oWYRnpLoSkYCiM/HU7kPecB9h+US9hDk8zu1q2uJlqR0JkSOJMsY4N1oFq0rACQLBWcpLCc
Bo3cZ2dx68sGUz4vh3eRtSlE8dobLaS9Ml/9Lm7rThNPt0IacMS5tYA6/aCT0kZx1ihulxRaUSs6
bGQ5WCDLkoBJXOFz7oGJnH9o8C/U0f2SvdhshQxMNF7oH+PGe05QzqY6VUtl7/RN+rUBF5fz8oTl
r0h27xq2lrNmOGBwXQxL5mBLjv+slLrvha4RvCYsu0v0ZGS2kd/RcpOb7WpTJkAEyt7mC0Menehc
H0mR/ZYtobcjAcknpO/+F68OX6xLyw53gs5DfY5KPpX4TnLjlo2FDMdSRy9ViNV7CY1jFA6FrQCx
msP8FeXLLMW1j+ZrhpCNMlBp2fNEfXfBv0pyMOlH0H1iEEl4an7pPAsA0xx/89DT1Ldn9dY1DO3F
++Lp7nKlmRl9EBkppksqHcNkiHm12mgLLGCE449aAkgE/gnqPesiPf+q1K8reGx0YW97rebIWGvi
z4qfmoc8RTyUi8jJK6z938f5AerXyMdoq0HOe+zeBcPOyTFmwHsX/qS+k7edtMvFmuYzGisMLusa
WyHmlyWD0BEsLxs+J8zuLvwXrUI2AjbASnDq/LGupUtURpc81ArMThBcJh/bggMdbo5M9EpiHGn3
Z6Ut43OWdFs4RJXMGKgIzC13urstEfrmRIjpYxnDvzSqkLe5hK5ZoypLQ9BaVpqJYKYM0qvh5vgQ
lv/zoMQxcTt0vq1eIC66bAvTXSp2gApxzUj01AusqtLE1sO1bTEo84lhhOrtrTs7oDxpskCC8qgi
vuQBMVqtmzUI+zxg7QhnxZ1NGlODLkmNzOeExhXgJGmQrrovvJ7j+Pft1aPmHzdlGsz/S24fMXye
w5JCnra5Ca9QvI53ExUwKRjuMSIS4uMqh6qbXRIxAp9RfpxKs+7PQYf4Bi41QUv/US6AVfUn1mSX
ycDBzgTDkGwOIW/Pk4XJS5JJPN36Qsgyt750Ov7nq2CHtBLHPYiWcQl7L2M0q2wpn+5X5+70WFUN
eTv0EzQT6517gGUVRneOI1PuvUNIlqSu6XNTOgerJTSAr3Z3ok6+7GfK9wTBPC2MfJtsz3BfPvnT
GuBD6NfqQHJZT9ZF5mnf8zhNEEb2ODDWvppe8ALbWNfAzVfAI+NGmp5IRmd+BcxSMBwlUNimDZnz
+ZvrELCHC4nm/RfjWAu4ncJiE4R8vXo56n+8TLXkq7WgYrt0bOHWGFzO9cBVwK98VdZfwZDOJpjY
TG6MFU2YB78kcYFxmIVND5Zt8S+9uFXeodjg2RLdwC+aPwqu4cfNs7ikYIWAhvD92vq5TEnIvgi0
4mvdhbtzJgj0ynH7DwVc5KeapyuM54FX76b+pNiwEduTPI/Rr8U/h76GoWVx4wjmyi64q8lKG07w
M6Pq+8Cl3cc6TdLNk595wjZTZYojOIx3hzftsqMHiQhPyLaimXy4cAMrtUo577011H1feRRCMflm
7RwvxVCyl986F03wPhIxk5KSj+/nPeTgAJKSBVJ8Vx+GhQc+NPWHYPnIXYvJh9HeCETcV0ipEt+K
+tylpE2Vxa0Lz7kYmXRb0D8DqQpzSYd0KAF1BS1H2f8y8RwYNybEDi0aUohiEmXnJyxqOZlgISs8
rfMUZxbZS663t44j3i2RePJzFKYhIBTdr2qN+flR0z1SZH8P51RhdzBCN1MYmRBYPQXVsBhmtaaS
duJk+nhEGcwBfiwg8aD9EMNsxgYOk89yVRl02DQ525HiV5SpmKEuNd+l50eO4MvT+p5OOfqFEopv
sKvDQycf23xu1LeU9uJ1BrrNnYZDQRxPuq6/Vqs29CHXrJpE6H+jPgx8bu4KuBNKdhuMGcdt1Wgg
bZ2uUFTIkmr/5EdLsFG3I5AZupQd61KDLd66KY7Iplmgv+ZGAE3cNHfQRHNkd8UaZ93NJ3sCknP6
NYQ0ymtqCo0SHrmsfkvgVubX6OW+nND24ctAh1UdqKosl3gFkQ1KsTQFWUAQWrNLzy4Sl/RE6QsR
4xnjdUd5SQikrvvIYWZi3CRNTDSTo13ySaMlCQkIibsfQA+h4Na07rptUNCU6L2sHjXZjs++WUDy
/AMk3VRw5a0Ig9Hy4EtzHhJEHNtr6JCGcfj47lzOJR2AIBlnrv5tJA24JGcix8uvlWQShuOmO9ur
kZHsq9eBqmHpMYL+2zZXlaH2eLZbgHgpZmglw2RhLxrSWv/tNPryJLvBE2D/nmRs+s6OZCinSKci
emuJvnqG92MK/4Rivvd/uX8QOIVuZCmLIkFkCBPxexMm18JXafu/rc6vYdRFyFhn0PSzkX9XHhPf
CCUOpSPME4E9D5vPAMCCM791Y/d8St4kua00tD0LMxuYyIBOZaP4JIsCYxMbvwqhqfYEbhf7wo+W
ZMOdXTvQqfAq0b9z05yD8YZc7xspIc65dJASzMC2Ez5UWwxtfvzOK7g4eYwsl75eHRr6dFbpYc/N
n00dVmNFnQOKSzFIa0Hln98SYmJiXWvhkuPEVbVgIh/HfKEsPuTYUIxFHYNC4oxBP7eX8ZVnNp6A
AeEt/XEai/oRycnJOS25Fh+x1w5CEHOFqvgTWS/cB952brnUKkNMcXfrrIJH09d5JxOQO4WQOchy
IOYAuGS516OXGw8DpmWMb1Z4zbfyYqJRfUjoEfE9AIeWR6r3QQFx9qveAxbRyqApU+0LjjkmFpAQ
nSZGdoGi9LOHM+qIqDB3PXF51D4+/Tt2jhCKqzKYoEBcZHVAcRwPpxWQ3SPhWmdYEXNORQUeejD7
omqNCj79Jc3sWhl+svmSEOpuoakk8RBk4AYHmMJGq6hYvbBYRAIffWE1FdKE6kqLlWWPNLLPxaOD
kF4oY6pP47o0VF764lFPMXp90Cle3dvU89Yq/xMAhpIWkmqXRZ7Ty5yXsmdIj69Y/tlGB9GsuWzJ
hdOeBYb2VtuN/h9PjFo94gAXp7k8r+TDilKIp7fEsehJs74/EbIqZCH1JrZllbUjrMztDuEQaOWx
G6/f3rZII+2gUORRBPd3wEP74MGQoGF09doaVosXVFb0V5P3x6xaffv9KtuJkYrwW/uQ9oWYTMdY
M4V9tRktMG5qUhbNk4aOYBrRRsXRVJBkS9fUASmJ8eVQkpPh5ljRifRQmqWS2CHiVv1UpeVdl0F9
ZdQkvhOApj3QBXNv2e0SAc7sxTxLJt/JuhCjJ4vy1HLHSpLkQhZGlqmh/7Fo/NRvImqPYRCCuzmC
K2rY69tlF9rI/vcGIk3pqMb3YJbn4SZoSr6Tb8se3RDYsfj6DywyUF1d9edzXydvLv/7uIKAMkNS
L7m0ZTwInS9F9H6Aq0IUlkQNU0RxRXWH3m187NiI8tB72Vmjqp+tgbx0SpQ6Lw3hDslz1t+daybc
+b4eXTRI/L4ShYEx2PbpFRNkVj9C5TRSEOVHW63A1MUIsDCmMH4MTRMrWETA1ykY9JX0FizOsTQQ
VlFn5ije/t4l2XuMILb8PBWfegREHGJnMByRdj0J87vOUqFnZsYUMhkVsrZRYzbNcxUmszlVGmbx
ZNg3mD7mbxeTAkeC3k105qTatU1jloOTXe3lLCngczwrcMPfxX8U4huI7TQ+KlGSZnqdckMgmtkU
jICxbMcxybqD1s9P5RQYCssJQH2N08gwe8XPGu5lJtBKiD9zP2ATrwkR3515mis1vk8lEWCd2Qyb
LZKZxfuKBbNNohUIMecm9cu/8+GLqdBbMROeDhoN+t2h9UH6sIxftEm99npIDZj43qf41nTCiDWv
8ddVMuw7M/auaeqcBNuV6DIClQmtpJb4Ft1fyd1waH+KIZULdlNwt14UjHgUUvCDsC2WZ0do5udf
fD9lYgg6D7mbE7ILKWAo9kc6hkYdQrGPpAm6temsFIqxe+tvEMlv7OI4QFWili/OqYm0e37VEY5R
C5Z8YEKugbyxOXd6G8HWH88o+s9X/vDAPk4MJib1IOiHqVF6ckaCb8khOMRGgigyGioIdU3gvtXU
fvf/ULZTZkVYguFLWxf5aGNL+cnhsjTp1GI/09wsARHRECh78TLhDjjnEftOWxxlz+JjlD3nEv4Y
EI/yjp63ymQaDe9NSOKh80t1pmPwQ5lKRMXUuMbF/AC4xkt//nQFSkPnAeXJQ7yq3oxa+RFvy1+v
tIqVEG/saOoDR9ah8qJBz0zNVX3PSlifPvVcl/yEGNNqWo5JaCFd5TtHl/WlwJY3x30iQXB4Exxp
TxkGORexTsZX4z/aRWi8tRzUarM/Wl/injkkup0IDsmqlZQWLobia8qaUYeR7wwhXonH+JLVe48x
HmFZnyHJDm7U4dex/wYP1NcrgYUJqIi5UY3VNdqyAOTQmVddOcOCLd9a/zUp/0fV+3z0DQvliUAp
qsWNjMzQEGE+g6jMVOZN0dtZxmsuqyKO6Mc0EN24BCSQGSdspuDsiqPUTpEDtqHk35vTn0aKsTl0
MUpThktJhVt5DH+Ho+8ufPNv3itTmuwdIQgMrXJbeelK/KT9RApXdr+2orVq9wQzE7Bd3k3pThC1
RjfcLKD1xrLlcC4Hc8RXu+t1aFywBb3DB+aXmqL4IlbfE2zuo6x3mnTyyZU5lDQxPIIs6xr/d/Uu
DpJ51XNnSPlPk7U/JhIEwhn9Mukn93Er40kFMtXcrWjOG5hAhoDR0zuSiHstGRCgh23t7UJSO+/n
mzWGnxX0lUhoeHRBaBs6OjWuxRk4AUmBhOOpyfEYMrnYrT7VO3JShAbESeFMfLTFvyeC99ncnqLS
+WF/thoAULfVYCn9lDk6ONq2JQOIkcKeVdz721pY7taQt45WsEDGWh22wlo+jcHkhUI9lRnm43Rg
mbJDDizagxUORXx6ecxxyS6h4ncQXT1Rh6u0Sahoz6u0a7a9hrSGb7XhQzA4r/PRFFVKabQkpkP+
/dJIkkZTprbBWRa2FtXQXD4jnW3lTjkOaxzx1geggKVr+a0F9AQy2R2kacv1WbrXH4wnpd/AEMON
Eb1CJXfc1afowDf6qo9GvtWM/COKj0FZrmvupwpsJY/BTcOJ2ATUwenVCShPQwDjzozIqCLyyw1j
nw3IOoOLcOIi70/BPNTEidN5KSjl023JDVTSZtC0VZ+Jcd4ELcoEJrZ8GZdWXN1Jj3/lAhfpvZAc
BVsmD6QlVVmhc+P2Z2QQSvXx1QhjqGvjzXD8Ht4sVSraDLaVeayE0RSo/W15RYxfXOt7qFXUuELI
sLVaPzve5lajbbX1VhEmTXeFAiCo5E5Ua2twRcPhCDdRB3cwvQIAggQnvXMLQTjj7CJa5xKOS2PG
IeLSPgUWbITNRqb1J1no8dw++QWobjfY8woKvdxb0g0UpfCouzlN8p+dR6e7Rkf8b/WqmxYd2vNl
2llV0VN00cKWJvYX6i6KoWxhICNz96c9jTwqbUpLFR5dWMoVPscksV8zzWXOrKQQ+3Or7fUvSPu0
cAStnldBli6/yIWX61gRk3LGgzqO7Y0JxmZ1tlWaYMIRCxwjwlMsqNclXs2CJzZu4o+/ETRMBOeN
L5PnUj9QvSBEFnrMVXJogzRFq3qa+DWmw6yYxqzWnpdW0vlk1v5Nk9A/0ApjFEOQY/s+zQUjUNaT
48xOBej6M/Qh/bfxhkquFE2DbqJoX6aOa3NntRRxQ7hyrjF9qNqpiT+PJCBYB41V/p0a7Cw1CxDl
j2nsJ8lBsczZP/YBOgQwuUxr9WzBFMKbY3vwfcZ3DbHvKXS0OJ23+HX1yrqxfNa+3c6yNzdolEIS
KfODg9KD5CShVfpHgQxV6sMTZc4ObZqSJLVxeIo27kcpvpSExzPu/OvlbNFKfMrrdZ3fWC07QyVH
0+IoLNUTKF/IBl2eeofSaE5rZCrxVrS+jdn6dbqbZYzV8k94PAuefb7rLG5IPn0jgepTVFM63TCj
LImq+NEbXA0frYs1ZRChTcviF+zahZzLkCvSrVPICHm6eF1T4C8CyWGiukoHhg1Gisr4H9J8id7W
F0ossZI2lb87QcFt6qLyTG9nCjgFmZEPLGxKT1pUVY59zEc6RqmXQmF7IaRytjIPasDW8iUK4m7P
1oi84XOBoQU+KR2L58A8qc08Sou3jVNvrpvFU3L8zOCprCKPz+SwmEeDIpho1lwJCEhNxr/oimbu
y1WVAWcDA1IBqvrcc7EPTAWoHhX0c+/jgoI0lPx/CYep95N8Dtat8x3m3p0aUWPds0jC/yNd8A0I
NfbKWsqqYLrVVtxwLs0LpBe1zdMzxiyK+4L9Dguriz3z+NGJVEcICk2wCZZHUB+iAIEYhk4V/zLR
dy/okD0apusJFLnwuac67Vx3++RZPIVEJhfYTEneRlIyCfEUv2OXh/gkjd40vh9/qR3BGIcSN+5y
FxEORZm0HNUNyuT0GXTN2e1ROkvsdVwiR+/8ZMLYHd1Zz9pnbBu9vxfBaJMbwZta1I1CKXmCKA0D
CSTng1JYlkozzR1k+8lSmIVsA2XbPWnOFiJXN6OmDnHIZjno9C/UL6tWKA8qSr+2SbRBR46mfPdT
6Z4gAsDpf9nA3xPTio6VK/n+TIlGt3tmU0fkwnKclOPpbv8vPTG8XMGSjs7IFet54k48nSHxXmvg
D1cl8mY2T1w/zrVPTvL6Kg8kDDzMVGbyBF5h1HrESA4FraVXV/tqP8VuQcA9dtN0rBGa4h5sSKxt
xswrIillAalga0EqAUKXyrKgq1N1aOhtS6Ify6LLqcueuiZT2x3iMDubfncNMvzIkUI7EuNEXfJY
LK3+sdCMgmJvReqHwPFNolSYYY1a6+R1lNchfEIct5F9/d7CO/LoHoJQyviON3WRJgfnqoptMt4C
FV4lbxkuCUzyh9NbJbxXrTeStQ0V8MWWmKO1DaMFV1M76RQrqVwhWoO8xKOtuglnUsP/6BD66e5a
XxFC6uWTTdwjaci6nnVqgkTV/eN6qridpulv1doNV0SO8MPOlURDIr3Xuv0R3yF49GEU9jDIppOX
P5pajzriUF7bRaPtJxCohp0EiNgTX4Wwlm2PIn/RrdIjMnJhMLxn89M4dCm1elKOHVqB4dRRgM3I
LHBuUxBkaOpd4mibXP8T9FkOQ/AqFMA6Plalv9JX8moA5ycHBr0cAlyNHh77OCP9sZaIZejN/Uoh
FmONhgra6dJfP65Ei/o5dAiWHP7kVrQfT6jXTqv1/eqlaKPi//L4LFk6Nd635uJ2Kz6CLKXbfnvX
YiKrfLMPiIz8JXGuFph/f/Su1ct2gJX0w5i9Fo/xa7Ii9u0BFfqqvAIwaxuP9TiiCdlpJMp5zVJL
4EeVNgYtK5etVDUWt3+UYoV0itvOHgIZORxDBkZ4v2F7S+HQu5V3MQp+0zikI1A0/ptl//3yF+fb
3PT8oKobPrprrX4AP786zpRXDW17KRkdTDCyo6RK2oGPdJ52Mo3Hj2bClwQTeFMvzptEovJWAkwL
YUZh7J4yPyLVTmatvYUQBfIQtl8+1vH+Jd2O8NjrMQ8hx8A8hhDWYqnYGMkfhtkZYTrTlzO7ogUa
ndakDMAS8jHUStgMK6mOIttzR43GwXGPTTUQtrqoMpDMYglZ/cDHyMgdYPOo8FBm56qq3vxKU/NT
SizHjnoRrV25RU9eSSK5fRpmkSoORgc0PYcu8FWxAxmxQGWymahwhWrHFxwBMjlzwUJUaRB3nWts
jbOLHYgHuCkxBstJ0HkPHS/JzQB/+yAn4c9hs59WoX+hOphNku736H0clAr5Icde9XDBGcPsd358
+lDYq18LZW5JQl9Os9Qtu9588Fq9cZqHSsUvYdUxW0fqZ5mbdKB5vU83yC/r/klSuwYE+QRBzGjc
VOSpPXhZzrJYlBbvL+oJact+j4Mxju5xQOti9sON+q20bAlSU5pbWWsxFDn3MFkukS7xRb/uUDPa
gKuANXr0EZRKJxUJZB8lRYsgBzugfyW0tTXc4nhjIEs2kYBqh9HPuWgLrU1sq4D19zaoyMiUuWGY
n7L1dcaUu3u1/f2aTQ+y4xK8nMMLl5qcxr24UNFHQeqOe54e9rsUOn99JS7Kzt3FuT+Fy3CEahCl
PTGVEZzDy7yIn4U83ljFF/UxUwvrqUU6MSd726V8VWza7uUyiQFzBid+kc3VxqeLfX+ehzEK2wTW
rDAf+AFtWKVSF9XlFAEylGBtiTJhLEN7ZgU5gALgzmPTBybkod6ZrNjIAgO5NdKcX3b6riT2hOlX
DZeFQPQ0g2LM+EZIr+Q6G0NZXhJkQDVy5LuNYiuxpTFS+64IexVW4JCsdj0BDMPLQsOSMgBMKxoc
nuepM3htilqjS4HuLymDJ/yXOH/SYhOeHlEyc8Pr4WhDqubkqarUiKooJvHJrDPONQGyBbdsDiRi
Ta/CgKsQSfNaxbLLtIYJ7oBTT9ot/duDWhIoRyEw1uNhP9eYaeSLqcHXKeUhRysOJe/5okmouikQ
pohvvp2ePODhD7m9R7vd4deDz+Mr6m0W37QlFedHtbRWln4+CFjeIRrql4em8wtSYQkTz995mk4W
9I/JZrydWlczEkoXxjPWM/jrvw2ATGf1AF/wxQkNlDugtG44BTX9BhfUVIOMG51nmWFgFACTfBEj
vGEMClomcxX4fu9rFIFHnDsTIDj1V/DT9vQez2bTC1USiJcW7TKOC+5+7hc0gfeaxYeYWDm5Yois
Zv+9aultUWkv48SvKdFxIicNdWpMRIyH383HCIvU7wcNadmFqfILcQO2LRtgCl0dEDU6m0pHg4wr
nYPeh5Rosjo26hZkxmFwy68U6BfQhVfOSZBTAaGee6sKVYVu1N2YZ279ltSzslAD2bk+3Es159ls
Oiq7+lsTIm4XG7/3b+S/OW6o4YypSKUhmBk4Rs+O1K31M7Hj4DUqDv1PAFFEOyCcN308cgJk8EMo
hOaxp6MpgI1FGIAWC3Ub26yEndSpxNQ0vdAnIouGfy3Xc826Et5VA3arJXqfNs/fRoXUP8VU5aNN
y3oQujs8YKtDdqxA3dOp2xoEY8kVYfmQxaLOTucusVC/rQ98q4/JDJh3KubvqvRoBL3YyUbu5k9o
j+67fW17n8NgB6ICxIpsbOSjyAdj7l+1LcUm9YDj4dkbfZSDuXgc5u528tfhCpRZ/Bm1hOV0w3U6
pIdkG+h5Of7rJkfDWEX2jVVBzM4xRAk1LvJhjacP0aLqhzmzX2Xhes/9Xovs6nZChRacw8USbfxe
UEvcJ/NgPpcDh2xTFSkK+KMWcswio/Vh7EuB/MiurZKrcLJQk0HR5Y3XDsv4vu6tDjA4SznOtv4Y
6D4DoK9zp61sQMpEdj17Hdodmv/Twl15QEMOcuSoMd92xk5gDUfkZqotoW0SooNY/rw+Hq4xqKqK
Ubp7fzTadI2VZsaUeCENemQoGvQSI+JmA75W1Sh15E379HfuB+K4pQc4s8s6KyOCrwAutOGrpgrW
gexjdH/efONTPvBh3TnCw2moyWBZIJrhGCTt4y7rpoouI43N6+TfbGv41cac0MSwiNMCGWs4BffA
mx1BxeTeNUngUl+GKSG24DYpZTBL521vBSu2HpHcP4e8/8T94BGm7KtqcW84GOJ2NWzfEclZ1A2K
WPYClZcmiwwF2l0ix1QuABpH0Dpr7Ow/O4hMUCl0ndzBgDsqCUdi22JPJtlcKlw+yWaVpeWPav9C
VCAAGuFnKNwKON+I3N/y7TQM9cWR15A+HUOYMSK4B6TcFiAzffcJPvlml1+sfmmpTKmkuhquiR8D
9lP5hjNw8TNYDgknm/W4uXOipFMOuiMRSxS5TgEeSev+Z9cDBMFsbxv2GWyCUna30PZqsEe4mm7T
rAs42qLw+uvL8Jq0B7LK4eS0HHUMiMs5QsDDedA+VuxpyZAgkaOXK20FD9i6m6COqxzs0L5UrJzs
uLdCbc0DcbIYhSqwpYWic/QfZWakCHDXnlfdJJu9MpB8po9t2dWUm9Gc6fZQfToeQrSh3KNfoA0Q
OAc+p9VeeKXLH4DRTNNzf+lpmEd5n772kWBsgFPftq7Kld196VJfXXoLJ9vu4/YqjRb4nhA54jBN
nBVbakvJC8EYh2q6JVbpCN9qpQppES+xMSRSQPIbDRmrDaqCsZlutN3mtviVrWCQ2JeZ3pQSGjk+
18vvTCEOoZ5bEoMcAEPdN90WrklDFVS21IQFq7tlbW14eZw43xGDEJqKGWfVBotR+isjYreLDM6s
Kr52UzTiZ/jOCqkT0RclBZV+v7eGwthcVrrJDYw5KtnYh5C5N5ScfJG3cEq65kWI/P+pjPfmvh/V
UprQRtCBro2lA5EWeUkiF7bzULREGnJJ6WIU9od/knENJI/LJ+aT4b77jFxM6cK5tVI/HJ+BLXL2
u/i0/0kAsvS6Ut+8rX39qEqcmFpYZwFbJ0DEVdBasJcjPhXpjpmeL0rdUfsr4js/Ip+01zcnjzRU
NF97tAW1vqg8yHeJU0oCUiHVctDfTUVk8+zp5ju55F0Ww2HXK8mXLHGiZIKf2bXcXPeHpVewKaey
MZs0VTlEFbVkxJziprKFUvHDHs2mibjMtLD8Tf+YHrNwXETqGe3biM02JtaJjyXoq6fMfAJDz+33
6RaqY7gfrje+an2LtBNUAdvoFnP9lS3pYh7nOAB+KqLm7sdYMNtauUFUSlqkNCYAvwOVg73y30Q2
+Ov9rmVOX5nhjcDXQCW2+IN2RUUPImY3Pi3M7eVIJXRY6qDVlClvOv6cZBOrdo1L5nJ5ntWAYShO
DCXpbL2ZMLg1nzSLOGbYQr9ZKY+mlgHx4ruRtVfhTSo/kMn5jYllVj1liL6DHW327n9xLK/tEv67
C1sLnRerg7oKsXBkD1Qbir1PS1RomRkd1IH48uIFHo/A7c3jFzfB2PLYXgDMJ/IhjhoNOGesYTiX
ntxNPxZ90GByFLzsDE9kAW+oPe1shJBUruF5Lu1aQD2BBLxz/Sq01n6ddxyXqvgLUGiuHhUHoNx8
v54Z7bFBzZGpH2tl7z831/0vt+tCzuEAszM2K4sTkWJxWO9XYDho48JIv+25WQG7+2pooHieuv7+
kiZ/vlKxkoEpgSrgQJOl/IgyDEVTBw/wCrQ+GqOhA8z4sLpA9oP4vq26/H89BfHqYAlUWBt8bdDd
8NA8omge2Hy0OrsZdEBEXgmat5zSrGunLn+iglMwt5s5F/DPEdbvE17s7Xclxfj7pNvNU4B6nwx7
/1qqgmAqI1/Slb8O2izASgpQALmXOICoS8l3w54XiWxO9QpqzvrCzLcoNcYRrtC7MZaEKO+E9xiu
EVICwS46oaX8Ylqk4DNGgY56F7x4KhYkd4Eslwyn8bRpk9UBYkZbSqGOiq6II7V06GcaHEIee4Px
NbtUdDF0vL0o7+3WJ16Q2DP01PREeRwHmBXaFzNGpW6/FaKRtnYX8Z2FX6pSkLETgUOzP801Fc1h
6FPQQpy64RZv+NVBg/HeuK4K5WjCSldMGISfR5wkYUjW+y3SdsBEEpO2WHyBgtB7NeFeQk8IJl1X
F4eroXN1YbvZ2WTxr4WLRyichsSEJ+qW+EIv0+p1MZTdhO7bZv+qswEQ4XTzk1JGmk55eNv+ZOy6
/HTUn5eSUB69Ztyq+oCae4z7eiMzyVkrEPNDdCNfuw9CgDobCmBuJ8vVKltnqHD1nLyluS/J1Dch
NuU8RGVJZVSuHBO+9UUDQNgB8g47KOlZdPOMEyrBlUxSkyurh9UOzIIC7pnGu8MG3AbBb2OSHFRR
BhIgic5vxhqosyVB/gBacvwfaR2b7zt5qVy0HBaLh4y/L1xPwiqn6O8YPm3GhOexbHUC317Ge4PX
CWi3hJXrTUnzc3M38pZ3YOl9nQxKzM5WyBHVr3liz6Z1tzPOcXF8L/1Uc0yUIk6xP2nWuA08cqT3
DSmO4sdRPmHtc3sjEp3zomiTk6xIDj1ZnNyAr5OogvsxOw0bWw1rQeqKAM7BPWqqjh9CQOES0lWE
DvRG6dy6riyhK1ujEFC1wqhhv5IWhvkHOGNscSoQ2wl2wrzZxl9ChcJou0ZxxERLa8se4n6lWL8g
9xke2w5qGd2ZDOXI+1UsgXLFHERu9J1RgLRDWqP48fiUwM3zHAtZ/eZc9jt+0Km/4mnIDIOLhd6/
gGsgVX7eUxpdUtRIHW+mnnx/OfVTCwBw/l7cKs2FJFgi5cHLBUWm4TUFahsRQ45tUQ0FnqXElJPx
iuR+27zTyYMDAS8lE+n/Wqh9HVJVQNdxCcsRt5OEo+6lPC6nMIxRBroLE9vKp6LLY7aEb8YchXNk
D0CzObJKcTpuUq9R12I6GAV4xuZbCI/a1fNJ1bqpi9rMM+kmCtCqUYDbh/OQGtkAprAotGYelAio
Y42vDdOg/SAiKRKNbGW+zZ6rXUID4xayjNT4DCwkYZtq6kZQKs6zYA3QeLYo3lR9pe4zjCxYwMJr
vZJVLrafS4BZ5PlrazaNPXGoVt7hYWF+hIdcqljlri1MZznHU7vO3hXdXnY6GyW52s2kICqzuGk1
xv58qU069ohqntp4ki4XtJg9Lu0x9wwz3+nkbnku3/+qBQgp4yt8Ke19mR9hPBWZRKqs9V2CUvid
P+2iogG4y85gSr41bmDd4bfxmHj9oQkiOYSHNJCVeKL7t6GfMN7Geh90nFl1q3RA2z3fNA+hZM0p
BG15947OordTfXhEHHsrG/fTTM8jz4DHbC/CRah6h07EwuPY705ChU04I6OMGtokRjTKapt0cKv2
iLTgoErWBuSGJ2ecUrYaPtMzmjfopNGZu/+Ujm+WhPlP7j+2SD+tRJe9rntmQ5XF/oxBRjkwZNoP
z/eXNKXDEjYr3fBt82S+8kFpFf8Uh7JoSJjb08rYNqJ2PwsGf2ZAVvCBqPRqBapT9tbNvLBYWl0T
yhqEU/RFIiL5Z0QQk4yFyTaLz4QSk1sOn1qK09Fvln+UPJAMErYvSqVoGjOBhcNLZl2fdkxoYOIo
Ib4Uzm0QnZ5Ygcn/W2Kb5xYEs+9yhltgEI0j0dFo9tvjlcUvSmJxB6wZp503ZUq5rAqRjx8WlJGo
rzq9Ul1XPggRXvMoQS3fpD3IeLPPy5SIMsnwTZif8L7tJjxHod86T8d8q3ixQ8YFbW8YuxApudH6
M/ubGkV93OJeXl1SqSz7WfhvlxWnTDCyOh76M/69C+Qx0LY6auDwmwAQ14UO2/EZujsXoUMXPaRp
tJ0nXEwWAXEY1Q90aWkGgxsUr0nyOcmraO9nP6Obriwi80jA/5IfmStsUxQw59Dk6FuC2rA309kd
QaiKfvTT6TjWiFEF8zYCbNppSCWiYuWMcTX8551C66burIUbwmANL21ocqSEv9ECkSuzsetsZxeT
+CveKj/Q5WiS2DnYC4PqzoIXCenFD5I4yrPs9bg1ihvyTeZ7LiZUA4UaSzDHGIwEi4pVmuMeepoe
u+7at3YdozJsFY4e9TBXMP7WrUmIDHEgo5BYuoeFqjelIl4jrDn221/8q6IceYRZlziFZehLlZz6
34a/icwDbqVbDyhBUaLYK/uFGJhgK6bzncUHEwxXcx7fQzrSiOQ4sEZty/Q9rRdYpYKqAOybyEBL
lvee/sGVC2J8P9KBqDMKrqEZWWU2k8Xa947ce1Kcwgw+Ac9L7mbiZ0PN6MPhq0mi8djFOs4/4Y/F
XJ5TB9yusSbGXFB6nC6KEgS2+CgjJ/OTLLq+ZQ/Evb1k8KJARavBAZOjUj8akgd4l6nSdgz8xndy
eZWAn9OhxfVbRwt4x8xygu1fEDZBN4MrQcZgRBOTIDGE/9lnXlpBBtnv5L/2B2mUnkmF9mN/n9hJ
ftOMVOkBmdNwhXRY1stUk94KztbTWPcX0XSQS6YUjwBkX3t9Sunitz5rg+7DLeL3rYxlO/QSX51c
62vSV6h+JeDsDhcauzBpmvo4twFGCgo2Al8c7STQSCKuK2eiMQLv4ZufuoUcRT/ZPCMVHP+dIbUx
Y1NJK3dPoEDnetXrXWCcrGjopW/5lq8HdZK90wXZETzGcFGvCIu33QjrfyluOqDccO/Ra94Er4pj
eAvYdQSIVQkRCFsXmDsIxGfPx5W/gtL2vI7eTHXr91pzxIOdK6UTD0kHiS1e52J7Qzol3ZfrS3at
vpm1h+brlL5a5fYfoz6j7ARxXjW+T+5xh0bwLffWF+oiQWTf494Af06O09WStT5BHOD6DuKUKyYm
FPD5CHJzmYqjcrm8XyRTVs5Jvs4yuQ2g927RQ1WJtGxzsdOkkwTn6bJzH2aVGPiioH8jtUM3B6uz
IKOWFP12ZQ5Az25cGKPOsU4Z+3YnmR+x/Of+ZbP8n562PsKub60NDDlHJDhrydBrcCSOgh8oNeSU
feEe5C3z+r9VdCAfuKkXpPgepMAG65mYiYTJK0+lJrq2/IetFP8GA9yl6fOf7H/T/hhZGIBP6P+n
YkKgy7+irJFQbyJilCWFJHrkH4c+S7h1FJRyWyiZUcLWcjAmbvkA15CTJPoTaTfnaLzpBGgGK6JH
Ad+gbxtWDprvksQNCFQDPhiyP8whW3vvIj7j/gzXYqx3ULccjrJQDjxrfGJb2/VuF+b9gAn7Codq
7SkBioWGknK55iZoV4NZqu6BcSFCphwRLuXcmWdFqPWr7g8iSTvTR1gz4L20eUURL35QPzgg56rK
sBUULZ1gl34iqzdjRMK8HPfu+c+6IcF7rkQZHqdcS6xusGsSYhCBLxPcE/rQAL3xIQXuS5q0WFRZ
VaTjBDgnSe6RjdOMS0/d3NcQEBWlU8VUPN9J9r9f1rhKRtmdWPYYKuwujxlDCzSVqNMIB0zqZl26
uwxKdhA49DadmZ3FX+P04Ichu9UB135qjmTBnRrUGxOqr0zjGVwcuvftInUKuJWjD0nIDjgr+u4v
OVAzxQxQLpNp2/+jwM4chq2mYAoUm8+Oj3M4UI2hLRlDq1RbHAwBkOuV2AgVtoa6eWhsw+qwVP7V
uCQUFNaRVdUfajQLHyZf+c/ei6dPJWyDvhgUfInE6Yp+V1FXjMuoo2F4NWvlQmvP/030yRCya0nV
5SGr2FIbcuOztqLUFT0Agdn5gkJiTbFyGLQc89tbojbRTC4qNuGmYWHYI225+apikRfJoCBNIy7Y
GWqvQcGV6NGA/kUjQY0o8waEbl2KLv5spbMA5uqGVNfM0uObG3AnEf+wkekNkUFBnE58Zp3Y42qL
t0XZFSikHG8AvA+gkRGdQ8iPoQXP+7vhH+fpeIDco3A/Hv5d8j9o6GpWpH2ScwV1XAlyeiNspj2h
sWeiwIab3csQ3YWhstOi2ZMjBELzpIItjKLRzjeumsa77F6RfvpyuqPlkJu8SnWRjX+vskminMyN
NFleU2OQJ8NlK/E2VdqK8o/TBiJpi6IcS4/2wbWzenxM+NsZn2Kn1LllIuCYUVFVAtSxFdBxBR+b
U1CYc+7ybQzPRY4a+sGUzplLsQg/F3TfKNP3WNFOIMj0eyoNxTmXrI2LW5XGYW7Vh4IL33KGvJ35
48FOwkVhw6aU7MFJAOQOle2QnIwvzG2Sz7Y+6TsFfNK4yrHpIu/52ZM2XAxF3wrAuRdzPQchJ/8I
9Uc03t18K0pVLEngjVy+Vhp0cs0Tuhf4tNQk5x19uXDp3NRhq/4vhNFI7BlxiCSeVuHLN8Lrohvj
e89tpdX0/W/7aB4PGvV0+ldASmTviP0B3yyUb/FQZg+09nbw3hDs2SQNg60iS+Z2ClBu7c2b9zP7
Is87ukaP1gHYDyAs92QYMmmtRsYj74ofMGBvJgXeNwoLdeiAo3PENb4PEq7L8VRnGunK/cGKZv1t
2UyJWULVx7GneCtx/zmc5UgX86FvG9daMa0aRUkbFI4RG87/2tR98X49L+xfXs+PGlGYrHcMFewK
Y09xe4MTQQE/z5qsKM6R5VAUjVesJrYR9CFf+5bVRKly/4FPrxmpsEAAaxhHnhufHvsAi2WAUlRv
14tFtj6oY/Twbrb5F1L3ABezzoPt1tOioB2IFxkXMfCdbmNVgsWjhIPB7iQGUxpXYKqdw6YK6JTT
FFKreVrT2bSRc/zDN7hlc2yCjL4a6TtRx2F9yC29OhYFlBRjX41G7/DbNtHzYt2fCRX8rvIGd7uq
DTQlqV07yCo0nBu+z1tbep62zXSlWa1ThSr9B2TR1WOH0Q8YJo4oUf9OwQrcMwziC7vdCgo8607k
AeKDfbYmG+yr47ReW6Wxh35Sl7EQqvYnREnTnbiFLIs3tZSJu0fh/BZz7NeRHZ2wZMn9QfXm8CVO
9OHV/pYF6ndMdTcSZlAPvLJLq7p3DEx9t1MUdb6TdynANbXwwOMPa6Tm4bkh03WJ9DqTRVMbdN+3
31vtEw8Zv8CcL/AxTFS8ahH9Ip3CQqsINvQZ44pUB1hBi8ASz73FOI1zODBGLuTBqe9XXY6p8C+U
8ZF+W8G0zvx+2hF+CMsgcfyIYYLl8ke2g6SZjFnp4Zl5mUWUW4m5QU8MjEbwalZBo/he87WflB8R
yq6ups8dGtjFRHUrhSmegrBJE9UrLpZwPIIA+BUC3IN6jZLBxUWfQdRt3HFrnl9AuTzZSGPiedSg
rtAtkXW1MVwNaq54dUXh0jxbgRR5jpyHF0tCTgULi9t0AEgHdayRauJcUfCj++Ifm7brCY5bEc0Q
msyxfKjO24EKs8Jz2fyLzG7vG+5G4lXi5QrTVgFNSQ9eDToXaXFPhdhf4BIaLTz+34RzwlZI4pVt
0TnWN5yniB7ie70nGi648N48OYCAJJx0DE5pE6WYv4DwBPQee01iUhTeGKTcoOB3V4g763dovsos
yEOpBJpEyBS77FuRjtO4TFgGypW0nRvEJNJDr9XpRqoJwco5wnmszrzLF3bFwjbxXJcuPNnktebw
RiGmnNpUuuqqTAN0RMCkuD4RwD6Tk1ys7j1RYSjrd84Ju4nsO2QByqVKg7S5AgkZMKkJc75wHLA9
12DfWL+DIt+d3HJ5pkF2yB6JRJcjHBng9TJ9h3Xtd/WaNCSYYz6/xEXzZ5ti5MegvsdjRuEtPGtr
9sO/ZFZDawf4BTH7F6Z89068PJ23KKlTpA2Z06bimSQaxnYbR6qKgUzHab/aN3Gg2Jq0MFlWWGT2
cL4ZOViqqGOxUzPNJFbCxmW0ce7g07rd/32cTgJvCk9Ll3P9A0b0i7oj2muoURerLAeTzY6xEOpM
ixjeCDJ4uGRJD3UNYub7hDsAwocFyw15hrysz5seS1uby+dIiHaRLjwtpFUgbX04k7K/HeS7aD4X
R8PwcFv/lYZBX+IUuqDx+rSXoxn9j0iIS1NCyvfDqaFS/utZjCZFS63dGoJRBp/NvoiOmawP2CaL
4ZB9DSakbgR1NCiUnHXxtXoEwwam30WOJeSj/Fl6W1dP3lB0CqYxJ8bXczhjkH+ssN7Xha1GRGNL
rOPPI8UMlIbSROQ02WySMVzYKy+UawA0gnqvfoN92bIe25kwlwMgaeXgZlvZPAH4yiKK6zKBRaCP
CqX/ieBW9fr/zAai4Xf9oVR9PBONy6yGPlr6RVj7x4mtauv5X3a/lhNvfpGAdYhX6zGrRkcxee0C
MuQLoSJ4jXdHtJmfkg7du6iXuFa52ismKR3By0WTWoVz1RWmn/4Qy2ydcpXYjdZtiB5cFlApQu/V
4oj2SAXKN0LZHPz4oH4F99IdLPBzp31JllKzHpfcO/5P6Qm+r2e3LirHXzXsdOW+sexS0avkj5TU
YphnkFJ73LB7HwxF35115aCuhX1X9Tvjm1UEbfWz2g4phsw46KssLlbdClQUR/nYTSAMKmuuwT1j
VRydU1mvykLxC2X18JwPxI+5xU8iAxsnJKxkheAyYBpFdtuviUr2fy77X8+gG+vXnOhHugvsLNmy
5fJpx3SsUo0dXL+hNcQ4QO4mFQfiNn41ALWtN6gyDz9tfZPwqvlLZ9qyauUp9KP4jM18kXnYsLFf
8lAeheM+zIKMEVv2HVYordRQP50EctGidMzBLagGDh/alEOFEprNgAuuzSU+QA/aF/R9jtXzz1+I
buBajJqepoRgmCZuItGWkqf6VbOm0oFVQoRTEpx1+pWsIb1JE6CCwi4jcZzl2dRIMT1ONDeZONw2
0QkMZgWsZG7DKDjcoGI+how4IfeCXt/wJ5Y76lu2yrd9PTos5StOqYLCjNhgwGEECdq5uLrKFIfB
Q5vMklFncNFq8kfH6oT5+vksYaTs/CoMzMXH+TfNDuyyIj2WwQFDRl3Nygvh7ge/TzSYXpwojKup
CptV/+eyXqOsCjn574UcQqvH8LaOhGhPnKFAwz7ilj1BfGuWf5SXUL2vUajHtVRWDu2kDGIIDaYr
gWzERmjBpRjR7rTk5UEAbZVxa2DmlNu07sOXtQ7EViP7Bx4bON6XN4GcX0oo7zZyOCVQPhI64ST+
s9mMcpLMTmYJsG6hcUx+/XTKBwEjdQhoBq26t0wXilWQ3aUmHRlaCflOpvc1QDbpUDXsT1NMoAVX
Y6KUc7TG/beKRa9wd9Mb9BqkWFVfPiwIPDmu1zGeRgLiDFcapGqnA/c6ubl772wX9Yja7sN9pYjh
KjbzTBHJBEKBaLb9M27l+65d+xZyPUaDrfQyocw7jbO0hoGorcb3TXhie4+vc8YENpbBC0cw+Ouf
ONXwdBZ0XOaLHWarbiCSffawhLgHm3Pfkvg6dBgO6/ePlBgoCGzvL1r7qxjQnn47MnK4EPHQA+pa
zsKPEpWfD3MiLD0CVdMFgjT7erF8KkOuAh2oEnewBusN7yLnCXK0TqoYZ6YqMaViawvLXp1mWKOE
9otD5PIJkimJ60feyGmWPtgZcG1Ij9FsgoZgpp2EVPCQVLuFTF3vwsowKbYnSnXBa7b/N92CmuPH
y4RjaQotXxr7CKqzTc+PA88VDqf1l6nwNCag9PK89hE9OZBFGbXIs/9iQAXvLP2GZM7PV1TunNo4
gV3FYWQu7Saot1+njLmYXg/yLRDhs/R6iI1o+tL+yc5zvM+MrdttVxcRvQNG7JUy0yqecOI8KAam
qF6bAm6WFLENB5vMu8zcEyjxrlZHDe1rhkV5qpO3Zh+bNC3UzKi8Q7Dh6YuzucAjkhanvX2HnFIv
34+vrMcgv2swqjEWDMffq6405U4roSK/KNgdL4Kib9BbCfBS5QtzGjLzekVAEtJL4xMMJS8mE87i
KqcRnIIOjoGs5nV84iv+tST3ZX0iuXS2YpD+8GLhM1Xx4QbZT8kVIPMNGlX0M6o8d878KxUKuyWh
yDJLxUQdtqHZe/fTzZRGk16k8Oz2nqxz+ovvPNKhzz1dFM1n5ch6oy/91NvjUx5m+3SHqbbJNIP0
d5D//ohpxQajLIUhmnXKlJL0NpMI/M1R4gmXcnxoK7AvkDP6/bnArtsd9X8YfCmkq48Dk00a7DMy
0LflMQu548TYfdPgerYfFFzUa3Cs9QRwmKehVRrdBXDkq2e9Gay0dav6zL7gn3wSIlPbIqSLeO+y
JS5UnHTz6Fo9tkCLTq35U3G+CCv6mGHwh7NrYQcpZZIp4rkXgAEYCnYJIB3Xrgbn+yYjVXqehm9b
GjyEI0avnqreEkga8gTbsh7rB8XUNxL5Ic3Et8t/8mNB5dQzx11Zb4qGNcHQ35SwnQaLuQR3OpBR
BvSEYmRtyrFWfL+cAvEO8OdBQCgH7EvUzY8lnVnTxj4RTd/bBcXDLOnyo1KbXVHKDP46mUlqHbqD
bj84HPcQm2FoljWs1H7Xu6yXNAu2uFh7SV+Yx+fjkk8EH0XscsJpqqy6n1ElJeG2/jfJzz89Hdk8
M38fgEa0MwgNu2Hxb50Nj2fRCw9lYzQfueu/4kYWzHND/229sE9h4ChcQ+8/ora9cd7u8UckA0g8
/oppIBQIr0ftcUFfmTBpMiB7cdZBIywYWvdj6X3wFgSff7ijxyHSjFpfioCOaA205kFtJcwcL63F
Oak3mwB+5UuNpv96e3aq1eG3IazZXM8vJn3Y8wdKosNzdLbrMKYL/0U6SrHxw9Y9AtchES3A7pon
MhLzGqkKqThoo1nM1M9i9pZCGvzQpbuD6xyMLTkg33tOUNjFxwoiG9RQUpJPzA/OInRObcqv3q1R
cGvbW5gwL/N5+nKLVVixkBOGgdW2HBPkbkyu+78Q5ydPouHNCYSFG+NzrxHSx2jAEPA+f3jqqZJi
9hie0RmyRVQzeA3F2Aj3KichqEP2ytvXNNzJJp7LX8sJ40iqeIIGlEoQG6ynnn+W652nFZAL+4JN
cZ5gNXCY1nmhRFBU0F/yoreQRkfR0vkhfby6dSPw1+ojyZcB7mvZSdlevgubVj07kJbZHklCfY41
O0+WtIqDtuLAtHGLCeLW3k9RX9ldy8gWYdU1QTLOPGAUuvvjzS8hEWVw6WCkXWpgqaRjRocXQu4x
qW6NLc67Kn8nzUa/+Md35xvDtbqgXn2RtRVarwEOrk0aKeAfipfaq02rsqoXWgHK1ktG7dK/od/b
V9gwMszlYiHdrJZuLvXc4HWp/Q2p6KDdjecsTJyK+dPPT23Pb9GAM5oVo7e4qP7uv5syhMOlU1wW
FteGzZg2hTEbpAsZLnu+IAPOk6ZeeO+ppLfoaSNcPk4G9tf8GZhhG/Z8WxHl8x8dFWMun3tWwO+O
KnkH7O0YZMLAiUio4jutJTZ27dTHr+5Rdg7Y+6dmpRMJHh08w10kSq3bppmOGc+SqhDsWrENfRBE
7HpS33flgFJ+y0UjsLwxzv4eF8g79kzoIiKUagt3yqi48KV7ATF617Er8M7u+JzcMbgtkamJpukY
Q586RoBVId2LzsucwglNrl90ds/a394kl2K4MlGrVckVWYkDuYbMNNnML3XNQ7RkkIOejWC1BVP9
wPBWrYknk0B5N2mkfm1VFJgNduR6GMQskZ5nT8/EKpCVn0SqU49xs9ehGsD6YFwYIhfixmK0yuLe
Gx/GRScx5Y8HVifASS+NRsaUUY5ktlJIlw5IJFEuStwnpeBBjHHJjrEY498ey76EoZRaPaxHj9e6
ELhX/DO4kCqprWUPTwaeSi8mwRmmd183L0Pv8PLaNipgjjxJSWCRmBaO9dStQsRNKSFXyib9l1xU
E9VELUCYyQbhO/NabM2Rf+kLt3GycIOzK9GFP4o/CM+L/na8iXz9g5EZ4UXIlNn6D4McafOK4bkS
KDnY6T5hDn5NIitIAIQCCuQBJTaPrB7bOI44a+P/yVMJjBFNuDs9qiMThWckZnFMLpCYi78zEy0+
JU1ph9BNHvwtTROKTQYb0Gw1BXml4MhDJ6hG4aGmlWf/9IqtAUfaOUiz90BBtOc2XoOMjTyRxeQU
xrHIchdjgJsK8D7hmv1ERnOMFdfB/dkhRRYvFylS/wTegjK2yxLYKEhdPrkyIXGWhVMHGwCIx+J0
FBPVC5zMyfSW3c+F3QwOEvGqpMtDKWN6acS7/+LdE9VnPWiJtuRsR6LJ94YMZn2JyrLQt45/qJCC
mCQ/VxYe0H1sJkw08VK8do28nXBBhSlKo8izb75bIILOLKcSEXBOZR9gyPwjjehWThDE72MMJQ9e
wO1XxDcRfwTfidJb/xCzx8TecTNFz9AzXkwsYawoljF/vGJ0ff1hdvdOuMSk3jwr9GqizW10+AGD
0t3ETXQRcUllmc95GXIEVoiaQnYzSdulrNlGO4j98D25+M8jE+eu16v6HpwNLczFEz4wxolFtJgW
B1WgOlLWurIrvWGW/zlBUrntVikrpjVHu7qGx7HrvPy+t6/aYO/o3U42f9zadgzC1OqAi0YMRbdn
VAi1rRiw7P1vqHa5qAcMG11l5fiNoKCTez+EXvMbua35ZU+NpO0SAz/yn4c4CQleHcDpTxV2yIFm
/i/ZigxRmpuoDY1IFi8oXlEYcmo2GW+sG5VlprFUYoiqcvGbJk/7FkysXTT162odFWVZPe3AEpan
tBkn2GcY90419WJVNsfxyO+9OPWg7dvZ2aoiku+kCp1PMe87CeUdc58Mhz8x//5BwdQP6FxLuvT1
2xxYOanzc5txtK51VbRJc0TkYMoPUIy6qm1z+wJuUlz1mZCpLhYzrcnzPEToQcVqUyW+AzakfFhz
s6o6ZCOUWviUapJf3smWUaTEfy/IkdiSQqoPgH/eO0rqakBn78yATVlnjMJlMhyxHEHo2HM45fip
0kUJPJuQHjZjeXrkHL1llvkkYuWch/hGBfj3yOz7KQ7plhAoqyfm6ibeZY1S6Cfr4h2NytpUDtXz
vu6UTK+QyQiZ3xAbmkrEXZgQcRgZ4oTokebwThrwJCNVEQcbFFrxQS5IuXEsEAuQxvZ2e3SJXo2E
6Z/4KjW5JBigpVieNFBCzkBZOij7O47B1IszOpJoZe8rHt0dAchBfo4xSzwHCIoSA1fbsz0PmMpw
o/M1bct4QutTWfC8Czog6gOysFtQT1mZ0Fbkk1D9haF1cr0I8IUmZ8JTxoq+gUKYA/0aDp9XXKGn
uCY4bTfub5iuEyRs2VuabB8YWCl38Tn86iGljPsI+Iiwtq+zIHs/b2UlgXjNvKftUbxjQ7UxjUSY
EVv25A9bYPznxmtgkBkZ1toXOjlFvjzM1TsFeXO17CVoGw91ToJI1eZlip2YHCRQ0YGK7AUTr3Vo
1zEwWW/drqIZ6rUlHLRiQDX2gkbIn3IQgLolZObDeMarQYJxjxdqGxGhIvLFBkc7N+k3JqFeh7Qj
86j2NY8bPYnUO3b8BfYZ/asXrULgb0GvZQ6f9zO5ozQY7u9cTjUtMygY0Q6HWQXHJal7GN+Kb4sX
NXTmzBLJAZZQ0kqXZ+15e9xGUDB/wY4QhLeVm+q6Mmr8BkYRda89OZRVMpcrz+GotnAjcCoDj1B+
B5cp0YQC9b63xzvmxAQ6y9UOR67n9oLG9zSDwv62eiuGtKi622ksSWZ5Dw2ItVdYX7jmVH+PSLH/
owWW/U8YHzn9LYfPTmBm9VnJWnpAhfNVbkZS8POVCVfQakO8t8vqDpzcoJs5/WTY36UXVpHJvK9p
PuHJNBG8Mn6aI5tQiQQ6QuFv8FoFP8p/lf17vUmokyi2QYaHPROCaweiX3DmO7VDgPx9taJEfsR0
JVsMAqGzmYofoWIzwTkVeXhDvaCQ3TyCRV7jFfZ8df3gs3LIjLHH3z24lmfZHTc5Wsx8zHrMhryB
87o3xoP4S2afXujMMhElI5o4WQbrXVrJluoxuRMyoXkKpRtd8qT2NS6fl8aHZ/srnj/Ay37PeGXL
Gch3iEZ/7zAk5whqql6i1UOiv/nFinCpS1vzmVEnqZMTV4A1rXOPCAmOqOjfLJchpWyJIJsxRysL
gEORiwIVjtCijYw3iOt9//DMW6lDvfj/0GFkcQihrjR7rhPoiVOLAZpjUkM78ULwVWqNLryxcUA1
RcirYfKmftbgHwcuURO9GxuX04i3RWkcp5FNxj0zoY9329KaIhjE0NNaHPP29z7u2HJ8lAtlAQVi
44E7QvEEuBnxEJJCaH4CJQbf036U7mnXt8Xn/PPkgi2d9pmVQZM323AESxh4CoNd/OcRxV1zyuyy
pCiefsM6KYy1760fLN8sHachGmhs0azBqMeNIOuDyfWj5yfS4x1m4GNdKOVPetLrHb2KrW3yr5Xd
1CBolMzZXn9pDTtRkptKrL/ytLu75BaqQlP1oBxD9iJ311T4V9oqVwWvGJ34EF6tc8hdbtpJ4JN+
j1+fgFXGmUHu7pU+/BjL3t4nDm7qVxRxS70UljsEwhhZPMTFZafIawr1U5L6k1qZUtFdGThYRGEC
D5yZLHVf6jHx/qig+XxC7wcANKosCcM8w1JCjIIfImllOXyHB5kXQ+USoH6PbW5cWCpv8e5aGVOr
8wkjEqiufBvIkf6aI5RV/9AySbMR9b39egrW3MLzJ00RWObKExKl/FO7aMNKo/qTCMnxGj67ZuD+
XTFRFJh2nC46bQa0NTv9vSPZdlVFM2nkvMk0FRkKfhh28AsaQ+5njZ1tc51lBYxS+tW7hF2Cs+Il
3vkWwIJ403I8Mck0MkATkIUGZ/CE7Ma9aUI+Durnyfv9YD71UxwBDxQwaCSOXOfqUsR/h2B/kV9M
tnywPRALITvx5mukAhc8CAyoEs1VW0qHkTcxOQJ3HTkuO0NUfKR63QIu2gup9nXsRFA6EibETJJG
hkryWDPKJd+Hmbq41I//ZTZyGg1ZHHaCODrVqlIMHdLO0LeFYrtfSJgfT3yIm4NgFE0z4BEFDJQP
QRYqR9KE4wizhHPZD71ddhnkTPQd5+EhSFXZPiV3qgZizwXzI+w03hI+GfDDEnmC0yrBYCOpST+z
UnDU4NOWIHmkkFNkcWsOoxLXpP0hjmELQl1TwfzF9ksS65sRiHV8S5tbU9AVtLUx3CNzVmr4UtFN
nYuQemtY6Rsmj7XGRiYlX0g4DKuRXkEwkWFY+TLqNGuVvkFR5rRGT2mpHCA32cY7RKTElkSBmkX+
HOfh1yz5i4Qjh7ixAVjUvT1l6PsMKTVLaWaekWs25jXvU8UhEiNZUoYuIzq3pjZ8/f24lzv4qXB3
vE/6bAFZq91O14blB46yttywLHSkginZUdc5fMs6SjcnkUIozQb34PkrSB8NfKNUjpH4XfxociBa
fS/aATvdlSDsYCsY4H/iImZVGDTiNk8xD8tT62t+1K9BohVcGInQF5SPDuPEk1M8au8XNaXhJsm4
XQH0/0otyAY0+OCQXXecKGWYb8OyoFUYO/4OA3xZPRr1hL5YRBMJQPd3qAGyYOPLIFCnHskpRh2V
q7uyRneoFcmEUbiWoM3uR+aicSezwl6ppnEZGlVZOYp+QcYyzuWs/3HhllEs2NVkM3cGyhEXG6k7
e+QPk9XY1Pp1C6ZjIiXOm2QByyxuCccLqJjZfEqcEdZMZg4aoHmph+Axf6KxKLmXkaKNEWUyi43Q
A4TV6GUi4/DYODbhL2L+3ss9OXF6GLQhO4pDxS7yKpwvFsE9LGtF6yfWHhIkE1zP3heB4EQ2VTId
H2YZzNK26V1jJKgYCLls0PXjcLTixihiqCxFFQkD9v+thHtoiBmT9xQBQWe2po3WMKIZS/+nOBBY
omFfs/X14SnQ7AqC7k1dhlIU1bV1mb9wYaZEBDbuUTyYx1GqCN1+CsYB/pS2CYepT8wW8wfGBJks
W0LKPpZ6x3KdwnSrRN8J5i4Qeha7opAx+FVCxkJVeruwGum/823beTDP3mFvxbe9Do4cNraX8KmV
o4oi70sDb75x/kb8hIehOOLT3RDprnCQSYY28KvYEvUW9qrWkZPEJnHK2r+Wu3xLxXZEzK90+lvY
MGiQ/q4m4Ua6EMY3+/r6/vOlgpWfsBs5aoyfF8TDUPGHrkMhbewa0V1tQOrcq1yhiwWRrZj8L9v2
gBaLNKm/24+7yri3omMJRVWjhdwozB+g2AwwyJJwQmQ7CGlqsTtjl7vImiPfOhPYpfiRownC/cTT
PlqvaqHAtiVmyVzYS0XnrbeV+kmsKHAe9J/b5nt+LaAbv64QD0GgObmZgxuDpfhm9ZE461hAuK1y
svXOS1dBJDMX5q6lHb1pBctIkDtH0Jdq2eGqmwvjPYHhM424CvCscxabn0bZ/C2YNZnhT6Uzd8E3
ZyzCU75vaRrU299MnfDbtK3uDpwWdfUG8BEMB95kdCfniKurVQpvLKHhpV6TSivM2m9Iy9rW3wq6
pGd+DUftA9eP+Ih63DZtUszTqDbShqzcwKM1l3G478bpQhxQAe1q7nNTSSDZU4wUngVRJecGDB9q
Vn2FbpthRxAWIpAh2GUcqqqiA6gbuuWzVivTmbz2hpTz3Bgjr7ucQSID4fZ8dTxYY2o0dr9OuGGB
cZq+GrFz52Mm/bDOCMWln7yrWoeIZFdaM/OUYGJLG+z8u84WMtrSPZAKk9YA1EQnwT7Fo04xrgrq
TExFRfbH58D0wyO7I2vAMI9999UrCgZHcszbZ0GahdpOTzlipiQExTOfHr+1bLpnMW8hP2PWi7Qz
GXik+N3tS/JzCwKi4D7viNlnkNeF8IkLkU8MkgmnSQESWGAFoXLazE60IumihrSH5GxfKzWxFnf9
6rZcqpbcdVv2m6sPMJ5t1/VAZSmBpShmXA2OzXxEi4o+Udq1RqnLrnmEQnWs85s2RN2Am1hxg4mv
ocNu3Vcj6aWVNNix9N2nhC6ZSg3744BHLwgU9ONFlfufXJU4tb5PqnM56Z2asNO7ffqATv4pStJk
Dad9yDfhnl2xHBvNLfmDFdIiK3kradnHjKwzF6ZXJN9FXz+/k2XE5fWuSg3Akg2pkT/ll7+46xNG
wNtW2XLW4wpsnVNPzJkO7TaPurEEDMY8ABO9VrZakIkaFznSkQHATkpcTXCahdohTsVSCjdMzU9U
ylhjoivaciL7GK8Mtxo74r+kWqNiCU9h2wSsfJZ03kYiEEBTnv9nAeQdmm7oYklpLq157cTwBPSU
lbaiLShmHKVW8Q61KzR/zhmocF6Na9PPSsT2PJERGNox8kOIIppZratiunh9kHaom1a7aKbIpuJ6
jte+N2Gd9BnLiIe7cYvjxIgs7E45ZjLGJ+MF2XmLuEEA3OIeJ3yUk5RNldMNoTVEmcssy1uH1zMf
/o8DEq2Kns9huZGuP4z3klFVoGpFS0hfbE1e+67gjxJGsl0ldg/W+z6za12CJRD5Mu4iOBSqrDpq
7v0NRsg0pf/JekWa9h18tD8SM5rRWa8/xONHJ0GuOr04yXuQbUd6kG3qPlvggw+gE5p7Jcc8UQWf
eXEL/oVDvSG4IFdg4mIrQ8xXhWdsMMdh5Av3d9GN0ds8yCQW/7U0B7M4V1Y5PN5CwhcjD8ijPIcF
ngBPm6KpkXrGCoI34aEi8KvcY60Ib9N0UZ0ngMVsLxrjCW8OZ/Cjd87S+7YbmzB4T26n/u/0OfU+
eg303tGkW/fJG+tjPDT0PICJhkpvgAp1LkpwYMDDXeZ8W10BD/88Jz8RHniphZuM0ZX2+rnh6k1W
4vwgsaw0Ix/c+oBrAQFeI3aslh0Hzc8WsbQKYuVxg0+zF5sR81zV80NF/gabOupxldWboiWWshPG
ZGL+SPECbCs5jEd8fJ3s70JL8ppEnS8nj1m46sABIcG0Nxy1Hj44SVuHP3uJE2K2OkP+M1lw3lRL
YLIIoRJB7Pp+68r6fezn6s+LgFftTGRgfJPDMhV6RhFk6/u+rMTZtc1J3chOGO2pZxsOzbxRFGMZ
QqOETeqv5xsubND7GAugzrpSWtkVkTfqHbxn70er9LxhRTodLlcPZshBdEYyg8co1QJRcnXmoY0Q
tDNIGMtRnJfbEXFeslAfMLjiOxtF7vKmHEWM8ZiAn0HBL05X2Ju3Snv5a/i6mo4QRz++FIJZcP2P
Acw2/p5Gy6lIGLONF64YiRY2f89PsObEKPmc3h1dUnLUVCe93/qQazu2ToXlbqMFPwiLbjnb5fk3
L2A5ZqH5lJmA4nqWWyTNIwW2SJE8RpspMJ9ukZaUtd9gfqhCERNpI3hvIU6XNGFpYH168LolOU4t
VQwrpwyw2TspGG1+cS45E5IFvKwtlx79T+KqM+/H5PzKc681c5r8YyaEIIU8Jw+yXuZ9jZ8rUzB+
F+9yRZmHAAIaPl+FjpaaMTrKlbB6iysC/K+jWSJ4CHl3Vm12pMajyTh/1dHa1Koc7LEYtIZonoqQ
saTet22T2q97qqJL/pOZ3IfGGVRQFMzf8dQKIlTSu+c5RcSTocN+BAkuSd1PmJQ6qRcG5AyFiymE
Umer+1xDXS4/td1wgI50IwLFbHekyWQKgcSqs2KtaeEEdRMQhiTkm3SIzYcqiOPJJhbJQMIrhqqB
EHRliVeUicM8N0LSzkW0V/GlgXKFPf7J7difRViiMFwt8kClL85QUVDobp13cX41/9RgKTDkOMD1
zWLIKKyfOF+kjE4ioOvB/HKQTzjRIZaKbQMRqvTk/5PbtjlSnvSbj4D6d2KTCvVPRWIxwaBZyJuY
ItvlP1tg0kvCLm+DXB8eXqL3lbrCAhXWFlpLy0Hp5NTA/nK5CqL+hyZnt1ks1SbbCqpDE4KLlqd4
rs2U0InTTSwjTydOg7fOfsuWc+XbDCPRWMIz97punIPBTvKB9xtQ1kJl0JaZrezTOAK9L9T9qgXJ
bR3SucNpMKrmBUt7H1eXSGlBjwRjF2f4phSvWvnMz/pRzRT7ievl3pGdHjB484dlQvyHUGKXbOj1
G6jIcuGNtBBQDjsOhcyTjbQFOgwgH/WBukv7EH5rvkbgkrR0Nccz0GlysEm/dYo9OI+lHrpN7wae
AfkCF3BbXb1j4y8zVU/BX+R623Fs1CVMYzhoYYNUg+lpcG4aZRH/DReKR8g9+9SvX8Am8b5eCjP+
nRmxdhavujVke/yIS5iCskTp/b3GgxGVOXdF4OqC9bqroMkCGQZ5FOxcIlEuXrDWBqCALyAjcRT/
40yKonRJScuoeaoO1Ox4z+vtU7r3CRg2j33BIidfHQU4eV0pJ644Nqnp9UDldO+Cl26sJd8olZIi
JVEhevhq5SsOIsdEJkRE8jiTHOK02JXVktLxcaAirijEOhSTTNimzVe7OxqE59/W7gbMBXilvGFB
7si/Be753o2fC8d7SzjVhX1/71XhFewonphSTJNq3jB7ri8dsvQGg2AA0sppYhe4UQbEGozuW/Sx
L2yG8CrgbMLSfZ9fYuxU+S8NDsz52Kai8wFXDPHvE+mSDsuKb9W23AWlPVEbUgvqmZIZ7dUtZ+u7
K0ljAa2JFdVeY0c1Obhs+UpgXjqViKBrsEWy88UBBIsxNBDYiZXBGAdRwNBeAmDVnWxEw1359Hdh
KPY4N9qpEG3kEuG7iPHin3jRgTihuQeUJK/twyBwCLrl+bMlWQTxjkbBSeaAPZ7l8cPklTCnZV0M
WjLgfC8iLEqCInxH9PcFoeOG8dw2FPHzgyWzFM2bllYaeNx2QP5o3+iIOBJQEKgMD4SBObDZLiK3
0boiNmB+3VbrU4FxHaEAwmSp81Ik54q/D9m2fJToousEDyyf3JZNPCXLbU7u25lcy3+fsfz2cc9p
LRJpzM3CDa8AnNXSDVrEhQRuoYcTR/gMyT30KFWlSu9tfVWtJsFVlNN2xng1/YaVy/7fNTe1aZD7
mIHC6oyEpw2qMGz7bs6946zM8NPF+H4J7+geH2vYVRac1FVd0Pu5uE0U12683Dcu7phul852eABg
FpZhz25EpTRQ1oC8In6oZXZExmsouYhbVYv4yri/HPPpa6LodztwOGtzifMJUo3tc2TTKMa6fqj1
0WUMM23j4qoamFSIOeJX9U/FOLtMTlzIxqWjqBTJgkzTnbBIXXUTgLacmgSMuWqx/iJrIoLuJ6SC
26xpScnxnyUob+bRte356C1Ju33/7GJvCOQDynZdOy6t4vJvvX1kOeiZAXslaRfHrVpJ/kM5cgcs
jsvFbU8DUuLYypItiH0iAbvBwwa2OXifGRypr+hBsXZ70rFAOcDH+LA6NaWmyXK0pMniiFOfsO7H
crU4SkBP6UWp1nYQK98IMneBtrsernaHS0Sv5nKngZhuvKbcLYFuoVpgEiWRTTbxslbm1gwNTUje
Z0qt5xfN4fb4Dmh1sxtw/Grk81XtvxNtbhjYlIAXmH5+DNjDNO9kqe7L94qxKmmLpFtrAqAP7ujQ
yiHp3goi0w2SCNUZQJLb8bZdePhtGVJXEaZc7L5Latwy3ZLck/8QQPxKIN2agaxrTr0UcSWYL8WX
Q6ZWbV5BPyMgXP0o0AsQ79aewvAZ7MS5qsz4ol9pslfYDlReviILAkgsuJTt8jwDlI7lEbQnNifI
fheOl66DOek+TaxnAm5IngAQrVBYgo8D+4FhZ3DBcCIVid05G+LhRBp/DDimGrTem2XUCrfiqlnM
e8sJCmxF13YhNmx5tasyBBil1pfvssrLyYZdMsU04iazFayVulNtHuiqzenDN1fVcnY7ggt7pFu7
BP5JiZBigBYsmrn9n4jjIqROVbfbUYkNWGK01n64ld6OabF2iGJRDpjkT56UhEuA89nCvPMK3aqw
NGyKA0VAX42YvvhI1aNNcvOnU4JPvG7rXMVlHTX1OrlgvUgjzaGt3Nlt9PqFlnmSaILSmEAjxVo9
RSDQTuQ+Fu4LdYalUrPPMkPIL6WrZq5TePbU+epNthPqbg9HCqBHFunjBu11c8oguz5tnVNd7NbN
oJkLeIph3CqrDHoYS/MjtSn+fFGFmRUqpXoavz5Wej+8KcFDHTeZ3rykJGMpeGjPTl8rH/J5P9VK
qVa4oCrzQnmYsikoc5TCwWS3plxH6+KaqeHqpq3dlfWi784tkEkdMsgK3x3njQfOgF5MAd+zpQa+
oW0zYMo6m6TmNlvzQI6dShr9gGVx5lMBuyDBtz9BmblyVb3bzwsT0r5CAS5ehwXwv5RCXGkoL84t
TY0zSQ3cVcE8Qq5jXZAjzau7jgmoAk+O2yYsMOBkagMJQv+1C21fkP9CAr+pLYbfwEi8ymQ4XQjY
arGn/shduplS6w9gxlk7Y7IcVTY8y49WqMvR/3opYWEZKpKKdNYsZjXn+p13yAGuBNcZ1HkG+9Th
UU7v0FUBE8nFrFwo0Xcno706bj/XnWRDNYKm15ZojazPAk7Yk8cN/uhFhdC5UayeKukExqja3faY
La+Lrm406046xk823NszeAU/YjXnfmfv+CVGuJ20LKOFBakhdYs5gdFSwWO+fuLSXmeITjDOWEBa
duJ2BMx1WJsaaIZgWLafrdwNQZCWObQGjoWaLagEAk250bSKzEILSnyy38x1d+QGLxY7SlbxoRd9
op8pcMEO8wt78GrmH15besIwObWcvmb8t7H86I026VzUkj5IkQboLhCrWKeS9fE1ikn0BEl3bUxF
CjrqDKrGDhhRyS5tdNPNo4oWCLby2yy+q4S+VYveWZSSGUWHxQGlImwULDJKW5q29lUd8Ucvza95
8KPFuvDeIZID5UkZgZa4LxmkqltUqq3IP5bo6mYbNBqtmohmfB1Gsc1/a8476ir6aFJazEA4sAuJ
OFpGtwWQ8zWUJidYXSIgCaVssYhJjCAC2lUGpgbUr4OLBvZ/47aMbko/m/HV45E5iGLKvj+BVp9C
Cf/lglHU653JzMEaViIwwkyfYL2n7cYwnp9Ml3gInx2SLr6ishUUVJJUlVUw2ThECOM9vOuZKmFD
bCLkzxb6+tR2f9wllHMJbsd86cWYbE8wUv/LL+e4nT0UXky5GRFy6pE/RQ93I10/eB2GRObeKOkP
LgMgUvAcPtfo33rF7ONrEcC+QB2xRFg/iLYWUcZgJRlsIOAb3Pn0zWxSEtzxGdXYgqU4WkXGJ2AF
x//nm7pjMt5FPNFHOyoGWp9y7QcoiO2iTVJ5aBPRl0RV2Qd5/IRyAGHgLZzvf2E9MFwwsM8wGu27
kB2aW6yiwiR/TiShC+OK1sG1wwDaNH/TJjlmy5+ia5986lELjzxYhtL3rlgEftgeSVR426i2OVMj
u1qFiml6+DR75GsCP9+O00Qdju7GxAiAs0HHzd0jh1ePnM/L0xrovmYKTIHmUaxb7e0Kmjo4p4mj
rWEZI6H/mLyZ+WBw7lYeGxH0PyYFpCRhDhOmGJNGSpNjF6uSZ8uWZVGvkmhKdW61hI62LsBSoUBl
cPVGe0bjKVIy6bF0TYTg1a1ICSp/jq2+TtbHM5D7vlAxT+PSFK3RaFxX/siL8Pq5Y+XI85rGMkO3
hgjWU4aVmvnSe/JqZ6VSS+A0k9sL/cLaSBHEFvCmbIXNUG1jWKK9sE/lOmdbsFanqHGyAPcirYPX
5UFqlmlyaOD+OVCO/8JF96E1c5djcBWkrLjNNo2WCJaQr5PK3ZhssfBou2huagPj6kqfj4npUr2Y
yoceppyFnymOmQxyKg42VkalMD5u8S9+3ZCB5pcLqYny9JzcajQ7IAgpUN/G9YOJdxGJPzy8qKZ0
Jx9xgFgGoAW54JhAR1xHmuelBLcnSUy4uRi4om6pNy+ioIwD+wQAD81Weymjv1eovQgKW5KqTdCm
mRa4xRRGqkj0f1teVXM/LDPeSCqKt/l0Bu1KDmEMdUUusPPANTRTzWuproIPM4jI3L4xqKllQqUx
HeGGuDHqshJRi+O0E4d5QUv8YyQ1/IGtyoOe9hfcthwKx0KmhE0tARrL2f8xCAQVFobNk5F5U04C
w1Y/CzE2kcBlIOE4tvpDmM0HXFo03ehfZDBp75syaU1RwrLo1zCWmeoFtncVa3sp1gVRO0RJSsCB
0sb40e6Zu7y0t3NdVx9mwY7X8Puh+pva711ldsORcG8slDRFzXnIislbl5Mna5WoLEW866uz5fET
SEuXCPmZoEd2hoNZSyBkhNcM/XX+c0M9DhQq8lfs7MYniBTd4jqkg0/ipWK0RWqz7t47jwVh0Vdp
1vS8eyvsSzK//XWFf8wpr0QKBnavFgWxifwzc0AUcHb9lzFYjE2wc1foSdjc7pit3TQEe6z9jNUv
H7KLCS9V1+j/fIfNOISz1l64/GVC6xEqiGQ/N4BGFaCHKyduSdLzNTRvU3kMaXAMmbpe1YUFTZtf
vZWDJXCHBuChmgZD0zjcVk2h0y8yOEmPOH/5mBv/+gf1UqHw2FOPQN+f9d9M/bUB8mCoZl+ggZRn
lV/UkWV7T/+rj6tpuHJXJqHm2JxwYeoknuuSMOwbmp7U6i6m0of3XnQXdjMgx97CRiD8rR0FpjdB
hePhoKkZdDpZo9Zc+CLyTB18BtYwzF93/Jz0TL3ZnWB44Ur3lNZkhLY1ORKISnDJmhXIMFjQYYaL
sC5oFCMCLHVy4fUn7nvwWOo2ZzozMCCKKvAXgh0Epfst+CV3A4G29SjtcjTNkMmvF/Y9C6VhaOmN
A9jHod37dSWOz+vGYHSp3rmp5Kj6Y2YtUv9YSIWt8NqQ5feWZS5DF7LgR8Ycv5gQFbHW4RbvJNRL
tXIwnhSQQQ27fREWLNANB+vLwnjxISJghUB+B5v49RciuRhgNLl7Wc7BQvDoeGo+diIRQnrXH1pg
qBQBq+jZSzQQk3qay6Xlpltf7eBE1GQISMcoYredIlGQiW/KVKxlWV8mKKTRFovY1QGoXvdeS3U2
ay+QMVMwcFtM65sBJoQIejVwkPXBIhekE+nQkSgdCM2llNqna5xuWVt6MdMc+2zLUQ7Dqwdu69fZ
r80PlS7k2bouaDKlzAZBH3G7BN0QkY1DAcT6iD2DwZYUsT33Mgjm6KC2kh4HCtpCbf0gOpq1lU/A
3CGzESQYgh47wDN/oR9q+9mYIt2VjHrCSFYg8nA/CK9UZU4iPcvf7fXVnO/M8bZlKos8zii4dOj5
bBIl9tp1nbf8YLNHprI8Vc8pNjKOv3H+j96/lZ93Vh8AyRvXicPH+ReDare/TNG2YGnrkFXiR3Ox
n/gLsy6zjT2izeLkZAaqQ6sOdjAwmEhNeidq3L09TBK2AFoxb2ki7k390dJXufIgGfKounUT/hfY
wqHcbGvjBx/V0wb9nJG1P4/VnQXj9NyUgO0ONHjR7yaJSkYF5CIap4WrZz25MnUAC5RR5zzeF/lJ
kOSnzZsu1FF7MoRpYWgiURNnBwfG1dXjJDYWFr73hbpITVe90oDMS3IMIaoLECFO5zwxkw7l74nW
fZ+LFHxejaOfChPK1MlXyJCZQ7NhgmGFtusDWKtLzLNCgh1xIjLuOX0eIH9z/JriOdZ7mlMKCS2p
/a+hcvGEh5i20mftWUd/UEj9NfM8eWxYEaxC3oFD0P+lvypu79BpVwmyL6zsUgdHRxNrYSvPPDVE
sPdtSFn2C4TvfXMS/QGYsYVYo74NkF1rOYuwOaP2np+XiWtznYk8qZnfO/jE/+G46gEPLPh/gLPT
jwIZSxe8FU51uncle4UY31zCAkfVxu7cn07ER4n2iWd7FzSNGGhJyNrccdvajZ0WmjtaOu1EBuBf
BYdlayDbyDBHHtElvh4jozLkdgqS/ssVPtsnclHlUjIMEk/jC7pYDZ6Hh5z3sbFVCKpsxFRBTESp
QxMXA/AbaWMVqrMj76hIKHnGo8qDyD5ZKZPDrD1MQ9M2729MZl+KtSeMK8EsnBWNQDTTrVSE3dVs
/5TwqKWOJPrrrb1twpbeCrj+5kD1ymO9t5orRYLoF8so5/FZAHPZACoBA6A/iBES1aOJ2AqZu1Yq
9ZZrEuvT7tPEDiKXq7/kldCgTZgPbUhYwYAghttp8WG5VkUO39K45N7ngxG1uFKygOg53bym/90z
OJXW7ovmRsRZdsYBXjFbdfvHMwIX5zCvzceDInK5lhlrHrXhu0BnWrmHhegoerOPnlqOGgaKRRh3
obt8o2i4hMV94yzKIrekghMMOYHxlVOH3w9d8CDazH/DLbZOoomve3pLLH/wNFmY1DwrRT601APq
ABlILftP0oIu+3z+7pcJxjSiqkWXh4a+DLTe6t4rpEzXM9tNAM2hmAirrXw2QMuE3iVj+iN0Z7ty
lC/EvZkFm131DSap3Fs0L3XKyJzXsl83BR1OGrlxHn5v6saj7Cauv8mMlMbDDT/s8URW3paJDDqv
+Rhv90tvFX4GhyvHAU2BZES/WNrby7YyI3Jh9Qe0+kZEML3yAd6NkR0bcXPAx8eDbTXxQI8kgCKs
uH8t+7gQmDwYB2oy25i2gvd/plNtxhEAcK+sDEUx8/Plp7Zrujj2AEdLKiPVwNGlniTuCJfO/UDS
iMUhcLwpuoa4TP3UNENynI96kW9ca1UKCMDickrsoJFXs2HdsZTsP8YfGcq4laTZwlmukU3cH3og
mzgN0BQGwykcqZD86DlN3/hU2PtSjAXvb121cMz/CGUrvSVz7nLynYTyKhr7QJK6nioANPgK3Hno
J3pRLn1Qw0qNU8hNfTqJWbZotaXJk72VtP80WOyLL7lIzGa3jkBGUnujNgbooJ43/C6mpE26xY3l
A1fkG5wFmZlTnT+GBSkNSKri/gnDjHH48NTrhyD6SoG3Ye3osi4ycMgRSjfpoAdYCy0AjQkr5hX4
IGh2elK3/Tz0oTcQg6mhP5wzhxXBD22praLzuYJs2pspUt4ZSAbWTvFqhRUpN300HI4XpPPmfmOu
Hupe14c9DCQk84IVhPzFn42l12/L/OR5HgB7FmzbnL2mTx5dLBjfDG3d4G+/3P+Ytl3er0IXYHQp
qrVVTQx280tfuHWaWATJyWHX51CImMzZ50A9WH+3kDipFcp+q1pkFVNn5w0W3vcY/P8yDCuLo/BD
B9tbUuRPv+dV2W08vi7zz6E3s3+Lnehne4RoFVjDlyi80/jkXEG110rhVocPiN1FbelJSqxRc103
3jzfe2ihIPNiliobKiqFLe5yAMc9c07Z2wpF401uybQ6LIIxzA+v7Q917KYThhf7jWRp/l3SYhzr
Twzd/348DEMngM4Syjpdws//W1xCgv0iJlRMJMgf3qiJAyaJ7DFuJUIi7WLzp5WWLuG3AxRF0zIx
bo3fAMu82A4MNTLIhEhcrru5bBMdyd7hx+F3ZxPxOC5kSU1/GRSrHodt1HZIBxQ2JK9MpEkTaLql
uacoTF8Ii6f56OjfqTwq0/vIqESwgxmS8VBcv0yRpfdirsVv7l4CHr3OhAv7/EFKe0q1S0a+x4Q2
GKK+R75fBBuchvctWX84NGI5EezwyLCuMd7mcdDdypdONOzHMQ2o9ok0FZQicKvNTceEa3IYo3l1
L30ACKXN95Xx4MGgmIwq8sVtYE/yTAIP3dZ4A99PS6Epa1ja2ehAyczK6yy8dbehxEitGPRCrvH1
QwfDMvtdkpJugboubA+zFDEvWPZ0EIlX68NemcW8sYjPWYsHSMmIDK+hnf+ph5al69nUugTPJMBN
mqt8hkKYnQzq/OF1fTEIDFlxovlC2S9n9Z81+Y2zVwpn+0i8xN8K4WjlYYd3eaAPRxNLAiEO2ncD
Dk6Zqq6RNPVs6V04uTkcYdAqezeeZureeqG4AgZapca7nOUsaeu2JxOiyw9mi/PrgaoGykD7AUhD
TTqMji3nxPvh23vCsi9oNlwKOrAncoBNR9Kb/d3k/KABMWONuGwQyKJtwflKz0mOBbmyt6ukXbAr
YVmXYEaECmIqGcGSJTZT7l7d30rkExs2urvFmzNzKjfVPR/dFqJw5R1jtWKy7nM0bKk2naTjd4gG
TJigKGYlkObZlXnxxhEqiidZsGQQcXrpUWAPnIYkyPkSWF5LP2GmyTlLz/UuSzB+MdcdvHD18j0m
UkHIjgrTK19v5i+0vXrjVn/4gQn5jQ8kmfK21WFrnSO+BDNepqxrsYQv+tryEiiM6/x5XyW1KYRE
nSq8xLnVwdu+Y5EcIGWxmKH9rWDXCUF3mUtlyXawSfC65Gv3PouRmXLfNOit1tIaBaptsXtfOjer
8mQptl+NmFHfGF3kOCxrwkqsjgpfOSC/AaBbEAhVk1Q03L5cNQqRet7+LHO4/vLuFvXwvltW8tF2
oXnnFDh0n2vusLfU7yXc66D9uMkmBb0doXHGibVHrQ4w1sxdimLA3QBE+MZOypQgDl4PKwRsdrOs
NRZi7T054dTQZihVgkwpuaoEIuQx08gInifI1ArXG2uuA5vAZc4laDXpIaWFrj1eerIKJjsl+VLe
aPqwxKl+WIn2OrV/0gL3KRqByUpYHsYZrYsU/c2v1mf5q0+U5JOFFpy65E2eUPz2oz90xUw4fJSv
gHcQ6i43BScfA1WMgPQa6T+grHotyyABZPQbUmQVE7TCW1F/+8w6/nDWwKzepid1BvN8WXBKoFJC
KMbsmbG2ZPqgDuFVnCyHefyJOyJI3wMxKEw7wXsK4OAzeeZWl497ehV0HuDhKuF8+Pay9yDkiFsT
BqOdGtYnG5mYNbrbvypwpsA7GRuY4al+stgq3p2AkSvJl1CcDuZOjDDKN4D2T5g80Kg6L1Y+I/HN
knVlQ7O6fJf0g4OX1u/XdKPS0BPrh+0bddXR9gdpHdmTKy8791q4DTUsQKarFpw7ymWelv2mx9Gs
09z9kLlpYagO4+4OGKlBL9qi0ourxHKlShC3iw1np1kWhV9h/iq7K5W7GLJjtWQtQLIK5hw9AbXR
VkII375++WCyLnMp0A8ql/u5DaiGWTtrtPdi86LOg5f8ANSkkGnazs1cmzzd28fuMKEVRdD16mQZ
D7iX9vZB/POHQDiSNQ8mDNs1c9NLw2BCtmYhhzwjTN8Q4mcr0IznzWogxn6J5QWgKCKysoMGMUIH
4YMB5gIXLeTqXlXNeW9bCLncBGCUvFi67RLAFxaiZDHsm1Jzkbg6WgMPRpj7INpoqY0sOExIRjTg
OduIvsff2InkCV3veEiL+a8uWMA7Q4VNGytMrmWuFObxLT6VhxehuG/Y/gYbSbUJ11vThTdvwb3h
fmXMLedgUhJnNGE/TqSHa5L20+VRZWqRUC6C48ugTVRxXXI3Br1ppjXM05A+gyH8rpukuIpccUaT
HZ/zcAY4vH7h0IeiLdcZCdwBXO3oTvuZcM2Mmm/dSxt7edcpHRAdVO4EkAmqzKBySW9olXsy8+Oj
C4YHNRU6le6Bt31lsVcGwJp2r4tBaklm3xiU/d9HnuxUoDlYedfcelYpqBVI9WPmB3pLzD2i34Gb
dBcNdGSO3t9bTOm2l4VDKjk+bdW76jhqb/F266Llru1Pi89OXjdfXWsV52a3/8oqhO7UjQV7Uyjl
FOfNRAu92YkfDBQ2j78hLp5nozJnKH5C/55zq0nnjuVPuVgZJ2qXLwMxRP5KmYjlJkCocGcmn+qV
FBUExLr8BY6jSHNeTl3dEqjJCYt2bySwDgv19P9636zXtn5OOsoXmt92wRmazRY4CAswSmVjD6Yo
wVHr2kP1f/6khCVLD5konsLXyS2S6NbTynsRSfbogTTCAbMm1nv06hZg0FuhWuAnwnnFow9tGaVG
8VQxpkFbgnOZZcr1kROl01mlNiNjxk7/i7QGjFC8wR5xrlsQ4z9Zb5cgjMpmtiXn5KPySTUoAd7x
+4dBWo2UHa+MoP6iIKXdwoPe1YI848yt2LaqPFMt/uxpvsILmktyZGr6KXgAj08vlCZkDmam++tn
PgMmrauTulrDWpATYgOelzCK95LVUPFZjheGCk0pl0heC4VWGrFZFKbGrl4sOu8zKIbPG32zYJ3X
QVfs4pe8rah21ifzeRoRaVZmc+fUWhrovLxCL4A7CwUBxyHRvjINsa45P0nQ9yoGFZFuGQqZ5/Bn
Etrv+bIWhOb6rWdm/1VRavK8WOi+tb8+1EzWgUIgUHwEWHJhTQHgul8EJCjHkdeo9xjD4ICi+QKg
tT0pV6BgN7KGgJ3XjuRc56fv36rDx+ukjlv32cHmTOSFfxrbdb5lYnOBN4sB+6mYOe5jJkHD7zK9
GuRwK4txYYQP6xPd/C/3BqaO8FgUfvrdhMER+dSJUvL1D3jOrLCx2AeOBj+nHBhoq9Ow+3N4CxnU
j8/SY0ltlPVHOjwrgnAXqRnBlfJoRd/zc1GrbaQjs38g4tcO86h6vafNnWlcJtDfe+nIJhd5T+9Y
4/XZozCkw8D1Ga3fNxRHoRdU0VbMtmYdsZPQEg1qWjpoiTy9OPPDQ1hF59EPsp2369vvNmFRHlf5
h88hrYG/rJqqhzP5ff1SfN0GtL/zT98hJtbZsrnIPNOoeW4HWbw+CtZyApul/UZ6k2fIGo7jH+Oc
kOZ8OlcH/vW8f7va6VXTMXrHatG1+d//HOZvu3OpvF0UPgN9jRiCidVbjlv1jQB+Qza7LBlEaCI8
tlrZ8xPHcS1cjluqiVL2LhtyFCUt5nfsEr1Lx9TCyGEoGB4FhZeetkIq9ZaBOdGKmOT2SL9MdbN2
B09HvY3kK56sAnY9IHR3Uyn2OVXPyI7Jua4jTTVOUVVhOmKi68AN00v9fk+IryS6cwz6d+nzB3Ch
UY18Lx2d7dOBSpQf+HU+nSNgF4GsFvLATHhH2sAfP0I6y1AoJgu1QJGa+LH73qH3Lo0mc089aYDe
8xaM9fjq6h9CGQsO0Uhkc6vUgFUCVPSIMREllT8T+To7jal/CoK9RqixubaJON9KY0qufM9h11rw
GEl0M14TR/LsWTSMsBvcxZrPDNfj1dwxJ6KDGxtHzBEG62OW0olWK0kJJl1JSWx8Y3tHt27cD6pG
13bT8jvB5dhsUt10aAnxAUpj6qBKmkVetXzqmAFoGOKt1BAJYOVkECgABsLkGU8T0Xtt36aJx8lq
CNzLX3SntZ09+TXUGaE2VII1dvU6LCV6+5ODsleSySj7f8kZz3gIPbDnlKyUjpUQ528NfCH8nY3X
TfZwz63s0X9rquku2whu+m8MNUeuy7yVwSUg+mDes4ByBA1mw0Nl0zwe/e3BSxhSmKew7JIUvB6k
M3W26s7L3Xw62iQqZR2m3yeUSSUiC8+vbhNA2sdq3EYt6NpUhLhh2k4VqjxN5qZx/SJALSsjLGL9
pxFSatvXp4NHbqm1YV1sbaA0VShqPr+4XbCqjQk6KD1e3MjFgWyhN/gbcXe6d1f5pLxPgx7vElNu
OOxjiHyIClYd1Zlv4dRkzFIWKOqXiEzklTBc7NfIBNM2LQwl4w7C7j02aDw4cPxNFLJAbZXAV1Nv
0L7ouRbxeemW9Eg0j5D8RGqnr0VHQ7MufUfxraPRMfQxWyuS4ggZ7FSDlKQROGnVflcmST5KFjBM
ZatWE+l00xm4XLHvVG/ckG/kK5+LNcqAZIo0gcXPVLkumPOBJaH4NYAQ9LJav9Oj7XriYmUEVGlL
KcE6NTiz7/tYrhv+IHvznM2bu+91h0VLWpjTw686kLvziKYqelL7S+os99D3wQG7WIh9TfF9qZpF
+0X03Oe35PnbBhj4STMB+tPJTQuBfJii104ppAduofqoi9ynNfVF70gap4Ui+nPxBoH/kyVEHHYX
tvwW1uYD2k0lh0rS5MTIqFv801yabq+1KrLkjt2SxMkZ9cZuCY4NwdthE2oaLAvHsHbXoeP8zGd+
yE+QzEqjqLozSr0J+wL8vO7tmhQoWPZJKnFZPNGfGhd6Qi8NTe4MW/KP7UWq/a6iVcn4oP16G+q4
Qk+xnoc3/k05jiKMGx0XHUwBIQ/EpR7EIWVsLXeb+RYf9DgyWdqbn2jsMNOvgiX+K6o0zpi72W8T
5NGkbcXMacQa8gIhnWMAkSSKnQi6W/1KtR6lub8TDQ9B4Zy6JhX0MzpMfxuyymUuLQadr6H5z+6l
CNPDCXfFx6kdjiFGlbB1dFfADjVxccSyegeMgiLgQOfh0ePil1a8Ya45EeQ0SRfVawVUM0uQ3ks7
ytpuzOq3Jfci2wCaT8M6ASlPElbc9al2EF/HT48OAuTrz3Zgw96HzPpw9wGHjqMzNf5rRpy6Ud1K
XP1s9NyHwkh6sk12UXp3NwitwbmzqUJkVwX07I7dDHx53Bx7kqTVtlmpPG56i1hAwd/qmGNp5Ucq
ckQV7N2C/8ISKS78JLHw3oa8xRnn5MeenZpbZtGtKqZSxq0cCsXunsqIQLRc1fM3qtqgfqiEAyOx
GR44oapiY49Un+VgP6ZM+TQWovXtilFhzTKiHvV41Xud8nOP24zH1Ho1bR7pC8k4oU5k0TdBC+0S
5DTQmGctnL0ldpRWH37FFwvi8r94jsp7awbBPUo8dgsZ5aD69pS6romizTVxr+NjSaNC79ce47mp
ussuDAs3NutwnWkWNMt6gSENWvY6BriVISiKaM4nfq3C17RDxq72i4X53wdcjyULy4N4KZ66XLVP
FJbZNwAywYhJgfb5kxTFcy9DYH2sONMy/aPhnDq7v3q+tbYRUVwHFoto57JI0MFgxvuTOO4mepGC
+DnCuqmGnCRdDFXBRyRetuuu4UWZFm5F0RlOLc2PMVWNfXBw1Qk686TWO0vxTC4Lam80HBvOK6IZ
0Vke5h+5Wj3KNMLtOeK3P3afMpusXtX2dZVuTEH3/vNB191G7w5hUDLkLioyADd34hjQ/jiUsKRn
QsBgXJC6ansyFH64pmkgw/n48ek/pFtSjxQsEvLXdrMDn0tDGc9fQmT29Pnvblg3KJQp+HgY0XZi
sF2u4Z1RAPcu+qFkrd60r+MSTmCfrNsY+mz2sBoA+ieq6t5yTCpGHvk5HONNXwN6IMQiHUIsoFjb
3eT8F6bhYVlftJl6j6nTXTXXj/uSyLA11Uqk8Bc1Gst7KUf8NPos3lu8TgZt4SBza95/ImjicVg3
TDPnwPJWZyHzy2m45TY55Lvj70HJMYVGTZp9b7haooNgD015Sfhn93Q61mUM/tyXcEik0wgJbW1w
040dFIGBPR+WKJXdBZRN9nLBTnLubPys/5Ck8Jj/qlCeln5nyYSVr/L5suI5dsT5P/dPc9RQI+d/
FmuD50CNPerFHIHUuo+rRJQ11nBIIIgDCFbi1Iwk0Be52XxzwCmaZcgrBbFGSs7FitXe69vj+Lf4
HsM4Qyvp0TzP6182zwxZMIJvd0mccLUXMfgYWbnYJAGD+nW20Sni0qCFwJaX6cg2wnlpsqh5irBg
Goay7GSYLre+qmJ5AGJ6oRlDCb0xlvlHdZgejb66oVpOJ/eIwVHHTqbTKtKusvuMAHHru3XH2Yks
jgK9rGnFkXdXHayP9nAMZYjjedMlOxVQLoO6VCVlVsK2wM2/5hBliZc42OPuKH3vxH2z37FF60xD
OYXKEF1hGfpBqmaMx/UJGOuG6c/TD7iWla9m1ENb/6oi74dCRBkoGZu8IkzquirmDQU2qcYPZHR4
ldiqnRvO0F2Gs6MzGm81ZRnKRyXnoOlYa0hGHqPh97Qxi9XlMnxt1GtuAsKM0A7ulz4YZ+bhdnvS
ZRp70VdfR4xvDKdPqP67kqjWLwbC2qmPB/eBm/VGHsN9AkW4pfr/U8WyF2s929y5ik27Jr021pi9
R13r8A6oG+BjAl7ZBHuspC5es9wgkMKgW+1GpvAisN8anjk/9pxIbSaDLaJDO4tPP9Ma5VDY2crW
nEJ4vsjWIh9S+og3QSJZm3R4q6YV0eI0CnCgX5OpIWJuO3+Ci1TKpVnvc3ws59wjMUE08tKmawkc
yISJy3yGKKltYMeAkJ5GNO9KAHgEhO1X2hUXBDVjKuMlHKVG9rBkaXZfX5ewjRc6zPV8X6ZTMyBh
LifAfkv8Ic+x1TVMK/tWBiP2/VFRn4aKnabVXxKQWr86LDWzh7YnOiRqKUr2nv9u2Hjb+l7C2QAs
BINXFZkpBOm1CkCW3Yl27FIv0waGAX5RZ6HsjXlRKZ/ET/a9Uj2fC+U6GsBKNOE8WnYIXbPU2NqZ
E213L5DOCr43Fuzac0KiLw04HwKEi2Fd3pnWkuKGpgp2PThfm87mNw4x0NnnvGJTajJrsypUZdWZ
9bXndI5c10IjdAVbK1ULthoQTm/+RPZM0xFt63qC6JE51X+nXK40F/h92aY+P/0cOcsOY4Xmlaq1
XVthzUkJZ5JZTxzFslXMJbDs3hGXiq0+XOuYz+g9Pd1BhHiDpqlg0faYzZHiHUkM0EAySa7+vstO
EYj4O7oTMCTSD05VVfGl5I5WvMKaALCQci7hN6ved1E8EXZRALuUtw/SXvs1nSD3hYL6ttnKdk8C
Prk1LoWfh5qMUKnoZUr60/Oxjr1Xu4fxMC4u2+QiJjo1eANAhDWVPW6dp0AZxLklj53CE3Y4qVQS
pVcBc1p/onJG4WMfUw2hNSfoAFJ3X9utQugxRGRUkdgnGuIouFJlX5aWdqvb1hB5at0fGzU/wcm2
gFvMLbHvsIRdtQ4wEQ+fST5DMT2SK3Xyw2wjFcT5bCfHi2mUOI/qSRqr4Jp7uSm0DzBlnSD6i7wi
onpu+VggPwGsoVhTrHcW0YD+J635G0ZjpTWtFFaT5nPEDJLQZPy662hzwyBZAJN/7l7ZZteG1Agi
DdKeLIRcpe6/+napXLSNd7x8QNQVjMlo2V0Us2LMKVCx8yv2ZYsw/Tuqd46Rq+emUOTDCiO9RiH/
ag3gXNaLY7mmIvJIFd69jq0Os0g3AGhTZ839KOcNczoJCUG6niJ0qpjJATOe4a6lE+G/+SqBto29
6HB2iHJp2wpFSuoTC7akyyHK4S2Aql3rMEJaVr3s3Y1kOXpaLwNW2/zp46Ic8DfPGyyBIAC6wJOA
WffkVFQC0ScFuoWQmNniRZkN6X8Yb/sQmoFarFqp7oCLLsZK3QveNhUVjqRkqdvq+lPR9A7kA9Id
02Hv7oEhc1r1db4Am1u3FdBPiY2yfmIdaAauararX0qqQFDnzBenFnSKD+zcDy1NZ8wklw4fT5EH
9nwdaJD1E4c2rDxUJpPyTJEqiPzG8P+WfzpU2rABDC0G2cDcDe+fHRywt5DIzH/ICyI5nXcplJLC
Tiv0BhXfWkrewHqLOIdkHETltwhOkXmR9A1rhV5GVrhrJJ91AvWrGraCE8nITYSW04lcknj1li9m
V1oxb9SZLILj073GkQa5bj/iad6C8gVqDpAm0gixsih1GBGZthE9ANPlWks9BqhmGoiKbWRRNBVn
+Kn7siPSsBbdb7HdZyuePE1hRv7nczHk0qjLTNPCq8e38h9AsxHbOMcEKv++/dJr00FdbtObXMYr
0j3FsYF5lBTWIWC3Z9dgWCvlzYdMjlDz8otrFdup40jkeBOic3apxKyvO8rysCfiVIFw4yAcdPtQ
r582heQYxzrfSO19RDziUO9KYVdMete9nT0B0BEs8Zl1YmvU+5biwX1qi3iP5eUWWlv6DCVxjbmB
pe4B6iE/B9vlpyZzCK1iMpaFpWzngNdfUCrYyDmUT1OeuzKAkkyK94o8HjsAomm3kCYRKaU/UCtQ
0qVwY1/RIu2LqGlcXjqeByqeGvvtj1f0PZgpt+Rhx8tucxJ6G3bb4ZxTEzlgpdPYYpR+99v5lf5x
BhU5dbHTY1lgOVRinWZdlUwnwpnYsrL038J0pJkO/u44gWyqpKTGxFbzGlRB/lseQQTBliU39asC
WM3LTcMA61i+5xLeseFd4sFVSOkoKHhznlaLcXyWMYv+u4Z2iAdkqgimig/WDak4KpNuK0CpfqF8
eicDHd7tUHsVa9/DQ5krp7wvbx5zjK7/eRbzFptGxClTBPcGwQAHaG0L1B1r6DY6dpJGzIfheRYk
Kcc6aIl1HFC63k8NvTgeoingL/5+iwb3OltD0DF77KNYNblKwr3pQtJ+wj3EBH+LjgPXQs0vLMFZ
HI57yZ1Xq0kHcejxfTEhsZ73M3r44GokIfeLnuH3uPnR4dU8g5ou42p/yGpOOv4706kWy9EOlkzZ
EMn3p44Rktyq3LSzTQGHl7jbHlyKouL5YUeMt7macFUUC17JMioM0Gt9PxYwajZwWb7NSMM//Ji+
nEui7rodJ2W7WMQhz2hgQtNv3oYxin0V4op7lylgikVk2o4wfgouX6OZvOlOiGhM7+8LmeKrKAXh
KIKLVaO9R5eYut+np78h922A25nXayAJePn6KLgoRBxHjQYhsWeDa64y93Dxyqqt+gXrLd9J4k7P
OHP8HPVmp7OWYbvLGOvevPqnt22PfATehybD6yJWOGve4iGdPx76INm0eKr+9y8ax1lkeq82ZGSz
w+0dg63YyvLxsEn44gYwMRwAwjKT5e7G+cOiVOrLT69sUW9SDstJeP3qu+/6XSsjid5kfkFgTmv6
7CrIYRWt/GrIaImOiMFW8xNbup5iZfaoWynv7MJjWaHzvGVFWDi11W1Jwtp7uitv8P2QAhnUS0px
6O+udLxePZI9VOOVLNVmXXXcT4WfGexX9H62rMCIsOIyEPjeS3zZk0GoNF43keX46npG36Cz3eFh
X3PeM0OcTjuNvn5m85T8Fsfmn2/lDHUf2XTKPYv3Gql5X8xJsJC8rqamyFBu6YHT9WBH2yTTh0Is
aUhgE/ArrH3xhcoU5qV72kMwRQTakC24Mm5ZDV6O7U3J6ZK7nrbHmGM98D2LQbBypq/+KAs+fhuH
lFnE6GHCvZ8vcT6e2qgXzqZCgcDxFjex8wqL5b9RS2UI79EfVL2ewZlysww8it6gQ+Eh4binsx+p
VatIHZu8SZXMTkCk60olaBBLzMCC1lIkAozhuDO7MJtR7roVX6SiW2roqqpWW4QfNVL8Og4cQqzu
SStgEwJKTXtBNMkWHozqEays8Jj2d8xxir3/ys0a1XKJGC8lpYwOwm7yhakoMzZFreS8sX5GWTJA
tUWJA0WakUQtwWWqGXr6FDiYkuHRMVwxM34oQkfaj6OyKzo1LD4kFVJVNtnlOrWgb/yBSX9TA4T8
x/SP3xpuFV8kvYCFmLz2n2v4t5pPKKT4ceDS/ryexLJVAY+2ML96o8hIyqIdBwoh3hoxX05MLZAR
euaYU+kL+nXQNMnT/R6oSyYOZpjOyiWmE4XoejSsXaeifBgkN8BiMqufYVwyizEgLgAyRgnjfKEK
0FoU0crmefI6v6KaOE8xCuMxEkn53KIGvbhEENlxTrPX7t1bV/qe10dF6218C8OEtATOUIZG7wb9
AxaoR12OSzRaksn0x8yhhv2VgNzyAZ2RsWQ6Z8TekX5bTt252b+cPZKw0DogkeFZD669+dVSawqL
7TSfD/pEye5kEPIwJMammXha7SvbgLo7OulwdHPjvT/8oIncu59I22evOvqrulGunXjHR0yBybWK
YQe4b2YsY0M2qN8msGH9AqLpWn/IKHuWpVXI5Zn2qwAuZBY+nS/S9ZQe62W0BsH0kI3ruB+qvbMp
ltPuCFGP0hiOJz1+10iau0QtP+/Su9zrVtG9hTjSW7aCFgC5UYAy/7s1uIaekac/IVdabG+GVVA+
LVjDTWv+kutEwTKnh8wZAZKj07BdGMTZfvPSufv0ndwJoXzTOWRsQGTsv848oG/i7wF4fwuyZkWD
BVSJV6tQoP7JQ+LNMiZrcl3mRotX2KG2/ciJZkHlawlL+qFPhC+PfTLrIf6hMeIAfoVmhXtKWKqA
sxFj3hmXlESddND4rq7v9Y9Z40KqmGSmFx6tGh6twAXcRDI3dodmA3zHNNQdhlh0PU+taVCho7Uw
sLndJe5hIyiDcN3W7CNQyJEktBTow/+mnwsr6l0yOWMd9vZS5V9x2TVi6auxQaU49YTNZCmq4sIb
s3T5M0CkghyXjltB1T+xdtdCwmW22FZmoi+iJgGF+wRNMTjuHDyEo7zijXJFE9nJmUDUK11nepQ1
jlXWOQsf4VOASPLvQOgJyY9swP9fibh32crbKlXpqBLg6J+yxFBzfyFNOGRO8Zpc8DThxDjJ5CzU
766Wu/8Lf82rfWFueM1JGsvmJVfEDMSbBGBF9qmkTF0LZ/W1AVbM6cQN+dOex++BrD9toOBpUH5M
HrkdfgdsIMcXCDbeD9o5pFa44BLhntcDHdhgRXFeS6dHdKLdgq3LNnijzIcbaUxr/5eUdFQoHdNI
YKSubfNVY60hvvu8aEn0g7g8IFhPeDB/cpBrgAOPmeEPWW19QYI0FQFYvRRgYOEQ6lggSmT+WFmt
aID5z5YD5uVdmy8kAJZ//7x0++fEWTO68dcIh5Y4sPTu5Z2BfZPOCwe55ffv7s0+4nHT3f2OxSYU
fm/Loa3RMGhIxqVt678/4ioDW456WuF1NKyPJqw7VEuao9rOch6FuvMliX4Bz/jGjF0tnz8TtwK8
toa2qY7A0P6qmx0a7PbfqJBEAA9Xjn1eJfZgv6m+IiYyM4IW42WrZzfGdksCF4DP7g1vJvJCv3Gs
CGRkMSHxlzXWkSmwy3on1iRwRo8oKde4gzws1t7HBXWVBiUMx3D5xdKbQcy5yYnore28Itt5I80f
JhoJ9hU9m1viHFoF8Sidz/A5IE3JpUePyaG4/Oqgjlx3tp3/+mHZM1A2Fn91fs9XyT4gGY/xAHsR
YE4TuXF+1dn99KZwJLASvR2BObXSFVUsti+v3A+Nx5JzQuPXKVuBWHJnx/dpjQU31wj6KD8jDEoL
RZpTiiZEAFgjIenRqijWLY88A406m893f1nArDmTBytUAQ0G1CJvxRuPS4x5+H/ATr/t1KNpGHEL
jNja8sZoRNdG955L8jWSlq/HDMPAL4M2+VqR38jeLA1YQaNbvzSyNYbCMrnzr24QcasJvzYsBfEI
2K2lqfeEdef7WRqMQB/lh4vhQVSnAZ8d30gNixLNPpOnDhWm3Ba3YETbwXhoMK73wIOLu+TKxT7r
Mopw2sOnS5Di0d4kKpHJOA9FH15FQwf4fSiYGDs8gnKkzUn9NjubX+nvS6hO2s1JmwoWmMU2M6Vi
RCYP43o01zihHi5rVeCprGU/+kAKKALGiX8oAVvnmLTwFeMPYcLVbRLLyH0UsDu4VpEbbS5BPb2R
25wQ9MDxRObEb+gP4k3B6/21BaLxp2DUDzPBLEE7JmLClDvvcryL6mQuNgHXURl0QgCkOjGyFLaM
52eSXI4oa86R0L+0kQd3P9h5tQmJ4fhwiyewi1hXWHOmWNpT2kVz4L1uBe9Cc9kH8tgwdq3xLBj0
mDHPmbOYLBV3nzdgrqSmJeITp1JnoTLz5WgL0uWL4sa8TedNt6RlPUkNd/k1Jk25LPOopKHbwrW/
VwmppHNQo9GxbPBUcOPzzf88h9P7VP2fsEmPo1Dy2cBVkntC9at+ZnY/6VLoXsK7PBSUk+H8pItU
rbZW9nck7vzAnzpguojMO8lW9he/MEPkQ7Ka9WWJQ86iOKDl/8RcP7D4q47neeMTrw26UqrWIjhs
9I5mfsETkCaNoZ29soLYVBs7+/UoeVh01Sn3vOzwzoyo6/kvrAEcNlAI41ot0YHBYrKOSGrYK1uh
vcxZvN/l8+Ii6btEoI8NQ1cDDeiAs7uPFZBV3+WXa93TA3eUC7nYzLioDO6EhcQJOZ2NeyQJmO+C
r+i8UEbMlef43XXHYiRHg0YbfhaRz7D9MMs3pSafNiQyuSnTlMtiK0ZplfmSKwNUd700RFBy9YoA
tcsdXJeiZEOEbDH9PTEuwWmn6s2DzEOVhPhxbHyi+xNzC5usXqfUmW6A4fo+u7xiArUxPQDqCXn4
r17a2j9zC7r1DAclj/1KzsL8134g9rR9RVnA/10V6XOmbmOO6Y+oL4VGH+rpxV81NU7jDrAauVNE
lDTkYtcZlcqnOBquYWbRmsp3wV5uIryhCClxPRcM4MRzrm4FZ1KJa3FM4MFE1bOEKhfMQ0V33Hoc
rQ282VxiugI4P1UKlGZ1vnlULQfy16rx27VM97jEeMUwh/PwsgRcs1kayMjkFNiMZ83UwermpNEt
iPvARVSbXDER9ZdbO7eQrNHvZRj3pE1VKboAfjU+7zg7JMIsAL73KXmUKFdFJPD5gvs/rBxB5kiL
bi9okWyYHmPw8ugLNL4QJOKkCTCbTa+gfIWG3l/AuAcSwPGBtI6AnlzhpPYES03WZEq5mkMBUSNb
u0HIJTB1Q8e38MunhCjV0eNMiIAOI3cl0zN3hF3Ja93AFnbuPZ+HoHKtnrhghYzldSq02Kpz+Mf0
tFrrExOL+vEBsPWnn0eCemZPzKozsU/6PCXU0JXj9sL7ZJbZpHlrhx7S+M6j4bAgWHYMm7hHCnyd
vxk4J+DyOm2hvDLRmI8SeLnWkBOO1DJNfFpG7DX3D2em0HCbrMKsU46l+dEwAJJenKqSgQUDgN+z
S7GaLujG/F+22Amhj/LbzpLEg63mIRQI6+EUh85NOxOtIdvqmUPJc8/vKeEEz+qZqbhyQcYDpIFh
+JHoe2VOP8v4bJzlRwMljijYH0ajY5ZMVlMsj3lrOicx5alokgQft1qRdi9ktiEJC3NVktfudRry
D5DvjFhOGKw99h4kY4EJD4L7n8Aj7Rk5ZUMs4mI9GAVZUR0i6GGaVCvIdKibomfkIM57pgrS+cNe
Er5etsyqLJ8Gy4WttyW+sQu+znBXbLAiXffobdMUVdLXnBwJgo4zTQCBFOG9Weqx4easCpLTxC8I
SpL2smHyDOZrRrKvFSTZKWDNz6SF6QUpiflyejJ8dpMVOUpzzUqqcmcWCKmXJOwR6bbV61bxUHj1
JVDmRGbQMiBQbScXP6kaCKCwmqCv+Ff2v/wai7kh5vd8wvthabDv9cKVgHHqVzr4U19xFzXH5W1c
Akkxms37Qpgxx7Wkhzfq7Ham/tNq0l4VPM/AxLobJHUSWbL0tOtPp5kJUWtr/EqGJp0nBkQAgV0u
b0nf3nyFsjWal6ewRLqFizUtDWCnCW8zg58Y2+bZETMXT7XPZkWz5h5yowssPD8EZTx9xcBNBgBb
f96QZFpaJdHzpnUWnJ1YEEcB5Whbxrd73tJKD2sX56olR4Nv66DSYV0M2Y2DNipWgFDuS9S0rZ98
zQAWwnC+ZBg8qPMMucrQZADhbveUFWhHR7e5LqoaELz95eHdeKkchfFT8peSINCfkIf7Qqcu1PCw
3rR97OP6KayQMdz+6VNDifIGoYwBZElBqcjNNdUbQWPK6AwVR+ic34TVrgBQmysFW+ijHVofurMf
goX0kuRotw+zS65egIF1IwqCJqbqPPgmIvQnoDIbWJE6UyoEC2644nEoICi8BM0mlRPvYes0PsF2
pkWapsdOY2b0Lhbs0f5PTDQpZtfNvn5cffv62vyMKXTKsuR9bFtynqAKD6ZtjfNhJ43+vXiK+DLZ
SUVsgNMeBv1jUPiSWKn/tH3nUDlk10AKeQRu7GSCZktwRODsUWG9X0ABTKr2OzcGP/oRj0dbNraq
cs+zFxjQoOCqunMOZMxuM1OjCoORAV/9+CiS0zLxNk+toYfsgJs7Ry4ynscNDZbaU1gp8cKQTqdj
G7MsT03m0guFp5LXYhxtRPvG5fv+HeDTPynUzxDjQ67rcQxrqRhh1kVgJsbEiXtF0Byc5w8/aa8Y
ylV4F5QiTAbRqVq/cHjfMsmb4uW8tS9qSBlSBZMhFkOAN5wA8igRRxCaRYr/xxkQsO3Ws4MZlWxo
ED75Z68i4c9zVQZaz2VyJz28Bt1XFMwQ+kcK2KZ5Hz3R+fNGLV0BszwJRbbjxgRRdmeU6MXEURaS
4pfLzkiiAuCgYLVLycq7JJO3oFIed9h8nSK7PP9jA3197yN7P+npjFI5IqSMdAqy4t6vd0v9t7Jp
7vsiscBrSTWbH4vlPo5KokX8RtXhR6tc/SKdvLsyMSpFSxKBZ3fubYhxcVqwYQSSTlH0fG6lYhIe
69TgTsMQzmNlTv34Gc9wVJUEtkqKGfMY53V4Me418a5YMMdapG0fvWN6ry12ommraM3ilnv04a1e
QoS+At2O/hAnI6jEZz6qaW3Xh35d1PrUFuolAbodT0ih4jxja5nnc22CGEDikYwklMMI8YKwiN0X
K4oi2me3LpWyJimkcBsaybqpqC3JVvy8OGnSl2OMfIO8AAE6/VgJxY7cVvADifI7XjQJ94S+50HC
pl1stldhzohQZ+jO2rCteqFYxt3C57TeJHA3FP/ac0R77MMzJpFMj64+JHHcBMxcf1sPsT78uwLR
SIR9C1aheXnozx2UDCibwPilvo8zgxcOQUjFkpo+pVV2nOZvIr6Thk+uk9H6WhP574qN0VP6MQ1r
u7dlkbTtEoDBF4UUlpl+gppMXCX44x6ZKtUCoQo3Ki8Ep4/BDqbcwtV4ZPUsesQnER+lGtsjPGhr
H71V6XQaN7xJ/gsKTTGOPG4qu8kLGOQZ71HVzb/0/LU+2EgmsFTb11BMmAOLArstjXZOqZPsY+rw
LnUkBt4aq3RcjpINTsha+l/4OvP27DkE9PhlCtgNqFbqiNU0S/91NFXc6z47YYwKon2HooItAtBR
AWr5LojjbSdf5aCmdJ8Pt1yArZJ8HMglZdwk42P4Cxekh4e/UjOEbJbE4Aaxlf0P3LI2NoMsSCBD
oHQi+4am33qHPsE5nE/p9K6Hbbis73KslbuzuLLni3j1me6oLkE/tTICJwsK0Jkg1WawrsQOR47u
V/2hlmyLSqsrTP96w6FK6fyVrG6cD7+8gI9UdBrpD58lUqwxRNGAv35F7GtjhS0y8/k+Mui+nhju
tOKmBEOpMsVWOajgHl6ceULp8OjVmSNKrG0iOdzp/O4PQlDeV282aJl1ivG6REA7uf8cEQt3KaCb
51s44kM0bCP0lLa+ZtMyZiAC9h8hmPzbY1BowNCaial6XkEi8pQqcXEdf5CIbs+EGEHiFdH+4tmK
YhayqR9SRUsmi+66sDMWZkrJJLIQbP10c7yPo0cdyybPEK4taOnldNdyr/Tx/yiywX4ztCEMYhEH
rRkUn6AKxbQ/tGndiXVi8uvDtVJ2p/4fszhlg2gnlHp7quwME5F0+DXqD/mPxgXxmm7MabpzakZr
opNOXwkZ67a+M1ezCauRYbblWHOTCCeasVqKxZOl4mCkgPhu0LqkaOvg74Bgaq3hNI0ky8OMthi8
8ljEoW/1oboz4/nZDWinEaHwOILOTYW6OS8M2CRj9PAo4pfXQKd9vlbOTmNtgYHWFH0MoBKZDq50
UjoGKiz/TEEah52jy4k5NPVsdW/Uw7zZglPaJgMP4rxfBvzpWytdfagd7Nw6RQ3KNSQPyM79Vhe3
HdHbX91HddHpdEeZuGzqPIkBsp4ZjUXKEIbTgVx/ND2bAWGVj3M6qXbSeO2eBLfSvxPrbmaRAEju
jOowJ8rFshvEDWcT9lnWbba0/qZuuiyDM6su1YeJxhM6x8t1vjM1J7DvCvAGyG8xCOY0FERUC4pX
m86/+PkV4eV+y33y6t8yz/1roh9O0Ng6enA1NMuC6q1EQRkuT5/bItwLzVPOonko6jBBxTxoXQK+
jKKO5TQAdtoecYff+iSlqLFd5wkk7m0aNidFDouqn28rSjhSoDBAXp0OvG74hNim283l9aNgvz0O
48pk0PmhtvRLj1+1GsvLWlC42bFLY9WrdxuGltshCbvo4qle6gtSQwg0aZb1xYON0860ARG96fKp
DYAHk3tsxPiTs7vUQbbsv2V3nHsk5NA2y51LEmKNUM5gzxRSShiQhO7NRj3zPI3rtcFYf+xR+UCK
iTfN39sgnNWeGzArbK0HPJ4mW1N9QO1YqESgtfSm+qXskkFZTyW352GjjsC9ao2HtoqaAU00v+5s
2J/MRyQSbQN1g8cEljXH4BPAvHaQlXrfQ9D0aeG2NoZRV6915Ld5wNUgFj6Szzr5iER1y/sbunBj
IuSTaObxxn1xiLkh3MQ72dQqKbNjcHKUMqKtUDSHhOTyysmIMPbdCJnXmuk9zYr6f1HS0I7RTEaj
fX9OdtJ1dVsHRo+Ewuj4bT3PGK1hqZTV5hwz2R0nSt9iCSLPFGJeyTcDySaB9/DsV+yQzW4TRwuQ
0FmFDey04M06gMMzs7mH2az4FatZadZuJTbhZPP3knTST3VsjtpNg3meTaJdreVvo8M8OMqr54fL
LBtPcRjz7kWtvbaJ5lTmjCvd6ERFsSphsLiMlDtYALFm7WavAgctf5X5utg/dd4f2gkxVYEkET1u
AdS8/38bibzUvhoVGodF5o8EJD0Edf6qnwxgEz4y6dWvPaFwuF/omVwFcjxQcX/QDp92u1L4RIdJ
L3aJDQ9ys9NggdLKI93/KwvuekF7uCpV9fMFjtuLGdrpBcsBEg7knaKO7+NFuk7VcNmwKJhsFn+m
eAEgX9s1nd0wtLn4DHv4X1FMOSFjC+NUy811OQam4tcPJIuy1anpwQfPVk99yt+v6fUgpWIcCRP/
kabYK3yB+lpaz5yztYGtrn2XhO0g3u+Cxez83nDk9p4siejD+YkvT8iuKqX9qrFndqJVErYp0KJA
J4CirqjYNARCgoZFsFWTQeVSGqbuHMa7pLNm8e4Nbtqw5RdsjHng3SpnLHfk0bOizKCm9+B4eA2b
FIFoT6Iw0sBOPjHMCZ4mNUyf5pco0L6OBJsenTzsU3WfdzC2zdb8c29FTEUi3oV9rKJg8wbFGyfe
4EqEeMbkoEeBwFpz3NtLM/o+xN0N1a5yq8W8RFseRecOHdVDKl93/fO8KJPxtGXrNyaqtp4oHI5G
yLr7u3zZnBXWiChyQpiX3EBp5+hB7Ce91Bm4/flCzr3syabykar6E1oKAvHFkRmtQJQeTXPAcp8x
2xrJo+S+LTIjMAN3G1PYG2/7uRZ86ZuDfiu+Vt+yp47Ag9hsP25lmLKW1kseWwUwn7jFf1yhl/i8
sF4B03FNRUBc7EuBV0wz+8cLjKXdhOMx8uQ9jdRriy35oayGSw7HrTea+S9tqdlHNfhSqFVzkyC6
h0WdwBQgTNaGRlUPwzV/IKUBgt3xFew076F8c+CLqWGHBglKwwq1ffoRwcTUhvq1MTrEnNtr6vJ7
Q/nY09+VfhB1sxYW+CbDBTWHsHClphr/yCw2bHwbs9OZPvRNog7mk/56QnpFOGs3tEb7EQ37aNa8
VUP9Ynpts4WHqAXv7Vs1tQ9OoUOnO4RuT2NqSgIQukestK8fpHzFXnwxCMlS2rnfA8SfmgSkWx0M
R79U+/LDYgfxkosDnwcAL5tcCnjQ40svazSEFPksgDpiGdmbtBBA+nIH2OJR96p5aAEiBNcCy/NG
Y0bWeB4wS7QMrqm2IoK3OnRgjUgzo06YNZP4pA6JAQwUZ/ISRqq8z5dmu/acAsrAv2bD4ZaLCaNF
XW8hM4q/qKHzSMUP7X9mpgVHL3AbJsG9PeD5OwscmYBllGAfctZ023ZzEdYSF/5bmIzHY5Vv0rdf
t0r1Zhy4R27Ua6B0oTF2Qyc1jIy3IyD2vEsrk2Dh/ZyT11TQBHPsvy1Dx33WWIORTd/kUj3WgBD6
C0IzsSlHqnS9bZgsGagxZ0D6D2s0Io/2h445JaoCfkFe8oYGy8k4T5axH1iw8MR3FPbuWAACm1UF
ZGK8T4uiuYUdQh6K8PedeF/vkvscREitQJmbwF+c0X1VwTNOBadSZUH0mgu/EE9n3F3N6L6ukWW6
sUMYMc/KjtWsqoYX/Yjd0K3sVADSOPr+Nvzx9PdMfAAgM2+79oflgpxzoR8OXaV8Mf4I2Z+XdS7q
zZBctw8JiELrHHAbTp7O6Pl3ulIq7L9QxjjCWbpn3vLviqZduf5h7fWmQDinM+KndF+45PFHbj4V
WssYcBR/oTHmQ7lZALIUcfrhPcJjhVXNG/4IpoJYcKaErvo4KgE1DUTTiSSsZw1+Y+FdHNbRVWI6
F0xrSNPoRDbD3JodTl4crCr+B4F1jANsU5p9v3yWAVoyR5DNyV9z5q1ZarjABo13wQEH6PF+Auhr
RLgmO52KWOeGVDcc/NJpwNlD7Nwp9eBQJ25uuMYaJUg87FC8mRpQ3cUaDVTmNoI75NlHTCj/RUaI
88+KOOfy5I73OlAWAXDH7+lMpAsx1coEX/3kvGgNsND24K98rGvUlaWQbj7zTtA/r9b7Xh13ekEc
k5oBHsJ9DnC6Hrk9cy/zJnuVngQbPLweE8vVfpI7C3qH7TZ3y8wceQ6eRwkF30N8H0P7xTohddvc
LI4x7OBFIONUnyd2NgR7FVwzP4ThSd2QGcT3uwvPmOefAe8rAmlZXqPwt9s+7g/eHA7iVfLz5YrN
04iJ0PSbSX1j5Q7efZABE6+efwiKEr7cJb7Owb0e9GR4mze8pQnryhnRi1c+6o4TagxCRRwwm+IC
5ze6PfEJgaBHF7Mc13nmZDZX5XL4nf7WsS+loDB8YZTGERDypMG9Yuy6awbTtdNT3QQx0yNPLNJ/
lnFv86wfIJE5DZNVC7oMGcuFbzIHgZy1v/bmZn3G871LSap4XOaAPGJ58xBpX7yG5uOIAnxFxopg
5KdFAiIN+H+8HSOx8M/XBYUWqnW9SA8ZdbaHXC3QWE+jQLRArVWX/vFg+W165xEZ0cuK3xMevqWv
FfUR25ZUlOE7TDozGae4scHjpAeazOl1XUnapc5hVzHg+EJ5jivqzu/0hS8uIysiuaZcxSgfRk4D
SQDdKFIqU6AC8ZAGJLgwYHrN+bepbfC422FQI0+RuFMuY5uf2hfq5ysFWy6Ex8bi0Ne6JahGf2Mf
9dG1zxd8+4bbp2Z6n6R7hpqU7911BYLi27U31xKWm5Vm2zJP4+7G15qO/FxkmRGTOPyxC5jX4XFs
Kod9MwrFWckBFyxt1FPpUBgAlKtB1uGW/qsju9A7Y6rD1QSpdYnLO7DEY/Uxrvw0Ng1XGYA6AVzg
ftyiq1Lkl3daP/3FT6QPZIKvOEgzvIyNykAZCgWtGgQTCMqK92FhlKgm4RyTTvRSVXIekMWIPEwc
7yvYyK9nJKkQ62BqU+H1MafzkpMQaEonSkydcURcivyzJ97apOeXo3PBWHNqQ8UdlspDvty6anrN
KsNDlX403dptte0K86iNJrvbFPfUPfL0Hi8sW0Jae4d/uQn7i8/djVe1z95/nL43/TKccRzv7/EO
k1+NDWg4QA6JJTT/TMKL/phhkFmSVU82ZK97wUY9uGiLgCDLTlecUgN9MOe0oD8EyUIhkQQA26hn
zuRZoTUHgMu8EjrxzZFriPkSyzh7D8qAY7Oc3KBdJq7nsuC/Q0olErwhfwm36gJ/N40BCPZ/ai+5
nLG53TWA2vf/+jgjLbjcqHS9C7hqgaVXZ2VRXD8QicZfCriF+YMR6v/PlLms0F52AJbrimEarvSb
k7vjxdi7AX54WVyVoMIsHPnUUxpFwx9QbJxmG7u5s7Ki0UAlc8PVdRhGI+wlhhrVdfF1QcxJDt+n
xOkAqLIuOpGnD9SrF2lrqdiS0YcrTASjMwOiuV6efc/0zmzGx1+2k2GQRRTnkEcD5wu8uh38S6L+
6B12fcjpNztQdobAFWBWFzwd7KCQ4aCgru1Ax29K2fT8wrz9Fp6SZJGaIdc4qLmDDxq5ADV7p0br
LoLpE3Rme2yAhAzHry+SVvSToKwNuDq8G69j9Re+xluquCWnTkkEMx5V8fK3U1EiY4ZY2Rp7fN5d
Ftb+jrvW75PhIAb4fjwDOCWHYGl/Hlz2jDxGYrSHZXbc2sLQRGEWowEuuf/av2v2PmexddbtO6yE
KZaKGuCUZqC3WRF8u+hQxc6of26zFPhHTINWW1MNPD/xVTrC0tZGYS+UQORyGAODhG+qDnboh6xu
zK1q6NybKJqC7gnkxR7M50/8F/16NFWAiEfp4t0dKSJ/+evDAvPIle5WjSxGHN/NzEksZOno0tms
eY9M9fctN61kEBxBvy/AgjCHIFSOIS3CzU1rK02C9zFzrvb7jlYHjnUwCbhmNenwQECw+SYSxWjL
yX3L/wraHnkwjiv1cJZyrg5amiXDWxDuMFS5MNIxEBRzdWuJDGIvKlIA2AKtZhHQYC/vRlfVkTnI
uBI2E11nvCH5Deu/e/pTSm2Y/e0QgjO4BTfyOcj8t/f6KsniH4uTyBNjsvqqvfdvFpqWUg8vdSEE
NzIkBGif3Q3BVGXadJIVeQ9bR0ybZR5aExoXtMPOP7EVYJbBxYriaM1CPoA/9B3im1mwCGjBU70X
xGmojXIaEx6V/aOeYyr17tSUkM522cXEGn1qA8C5+q2j3DWecKl80bjYCjSR/JU8KK1eGODCqN3t
LkdP3qTurIAP4WFoaSH+EcQNpxZ61AZ/uLw8T5i465GPQ1dqMjh6SnKGw8HcVZHnMr8d/1lW4Ea7
bjxJKj6Dl0r/+b4qaJCvXUf5TNY7p0D8pzm2HUJvgRqMbhdqLYjiQSYFjzJlmpFntzDefdi3349E
uCFHBlqhjP4DLEQOaNApn7m3znipfXMYsYO2RW9n+iNiXTHaSF4ztx92UTMSqZHmNPZTcw+TfD/q
wOWcjlPPWgKePWAUfPVpsEXsm6bXEwSILAMqOPcGHN/BR4OzBdpj6kSmW4aMThr6LKf7qeUGX+xQ
f+uFFO3sPS+yogm7T4OiYez/s6fztCTSAdniqhfRx0NgwS1Jxf+uTFTS8YEmMpyi1/lTZ8ZC1QjS
qrJD9METQCnnVjgZyB6sHPafoI4TvsNq4bZ4x1RydT5vhHKlm/IGQFr//09ttSe7LP8WUyl94cbl
lI2Dhm1CixnaWyXbxUddAUyNhuywv1RQtyC6LhNjX5X6+T/x0V6OVYzE6rNUXtgEf6nemMXQOJ8a
JKyOFLFZGXCGdo3lJUhsKMcf3nP3LbemhE3mJ/+YSM0dnEjco1bCdkdqctFHn9vgqU9TEtDLG8gb
Rf8QknWI14pN4ntKnFfY+Mv1o+7o340ivohAFGQnmhxeh2IlntqCjVKSFW96o1iymj1tIs9eUr+N
XZEc/yQN/MDqDagmneGHFDIQqX9enQFxfJreY8uv2iBP1OHaK1sfvMpveHY/baqHXNcl6VghJpoM
WxUjvX79xOPeBHiRa/fiDxBcdHuH8BENu3wOaAcVTouPKe6/JH0E2MoUD8NDQW2YolXzERSh+XUS
yPZ61I5LtaFqvFwv6UeWPanuL+Yhzz19e4SwjryZrwZZrk4/YxCHScUeiotgjbkJiMdpmVOw9Gtz
/8FaskqrL9IcsCqTgCR2QxZgwF2Mtu100yAqXYvS7j3uczR7I3Gg1gLn6av42qv2Rmx5JOWyeLap
0sDKPYcLnOOzNp5DL0fl2WnefMDV1RZzmTIZ/t9OQXkstKDVs1OR5/jVzbSCmxpdqQJFNlFVJq3P
uqik7b2iguY/zgphceuiZK+Iz4omkhNdju4rm5wlcW/oPBvVgle3lcBfdDC6CgZlhY7UylqSYKRB
UJHkZH05lhKHHEngbpGRML5je/lPgBjgGfd7/twCtGwI0EvlLInnMnuomTJLDjkw8Ft+AyeLS1Ku
V9u64vCSkQ8A9bXEJIsah/JFLIGLsAQ/n5P6xKKtIEI4KIY/nb9PRhZe08VDOLzUmxBhi2jkqrkI
dkaYys03WmHiw/w86znAclx1VR9jkqbHbYmCXd2u8yA4mtCYzJc5BYJHepsx+8jntGTPvEneF6sQ
0sILoqDUCq0kVtn7pcOZ6+OLR88HmDI8EDXLGfVDjudikqh2tdIqwN0o6p/9k/mgW1wGQbJI215p
2rrcrfH3nwtCs1Ma8/HHZkAQOcYmKFpOPo/U4ehJl9wGmVF+uTgGMUw0AFzCa5dR4whULxMRj1tc
jb9gVaTyalVGICBHROQiIpPfvduE0AuG7WvGY+IR9MotaXjk7ankiPNnwEmYa9iota5YG3cBKcKH
aJHG24OmKRAIPMxQTLs5OumnX0efkmbqTB35QNOSs7r08g2wiVc+/Lwvhkw/rK2by1pbtcis4gG/
HE3lsQWqjWt8BJtxekbbtVgFldIIqfhGWJiIswXRE2xZzI1EMsHBb+MpXoN1U5w5RkK/xyBRzzbZ
xLr3i+6xeiwB+T+08XDPpflSwLdIRCed7o+ds0OZgQLZ1ZyD5bDDLC65kiVjalm2M82io2WPVHD+
GOqidtyea+92Pdk0l9TDTXcn9StwBL4o0lsZ2THz9lHoA1zIQ5EU0P4f7LK+83heUUcSFsq2lajQ
OgkDAgVmm8EWyycsUU89VfX8ry+zquLzZRNtKD9LPrgHdndxS5M4WF0tdGuEZzMt6T3/K8rcDcxI
smEwCD9vwdGGHzn+J3LZIAEtJn1QmdcvvS+rW+qNld8mDz+ElQWyyAcrIDWynZwyMFCvKbvSDRQw
yhcoWgp0qojNWKeZ4WpZQhbf9jXk4y5y/dcEC1rV2FdQukBo6jScfkYSVeFIJgq3Xx6bgr0Wfb+R
RTwPm+OP8YDd3SafSK5FC9Sl25TG8u3oogJ5qygcirCPDlk4bXuelbt1gUvjTPt38+0DS/H4hgvQ
04SyT7+RRskrNAUBUyE5i+Cybjn0fLYaV3HzWzTTtQc1sPbFGG1tqQN7vpTSf5O+RmWHRUtt+jtO
qBQL5y62xoUkFBzeRUwird5juoYA7NLTKcuQNkSKetz33k2V6T55YaD1nrSM+6wI3vpdaQmZhhaL
7et5OiIWm7O8Gy6JC63DKcL9xu5UCr8xlaf9AVimO6QVGwq6Jn5ZvwlpB8r/pWU9Iz2NXn3DamPU
r1QpB+fwHdKiCROJnpWF/2F5QXwO6yck8tVWfPgb1Wy8nI2AJBt4IH6T3ImsY8eKpzXU/cHSRKr6
FmR1iCTMR6IETL9Yui1KbjzWIk32p6kpH3i+AKCcU39t4+5ob/tjTB1zCwtPhSCnvCOaa6/o0QIl
aahViveyiO4Z4sAbj+KQOh7NFHPyynLTVS623RqlD1VI+mSqUqhQNPlgxMI2qd7EiuuWV0sj9rzY
dRv9nYymWl879omp7jEDWRlUPENsFSLQsLh5BYrJgPBpYC4K8kj+ebwcjl9sjZtMecWYHeLbDHmW
e4tsm10X72DeUZLG5HcruMDHYoABVyIA16LLi9zGS+9Xy/6PFWZOEbJ6EDQgTqBSLi2DZ+wwmTww
hkfWFELBOBKhHXsKkNiHcBBz55pp22QPw4BL0Iu+L33Asy0YQZT13RX5GVcCjHoQ7vBuSQiXT1Qd
iYUGJkbYxVbOrl9QDhCXQvY+GBs7oUiOLCcPHMcJKGNHBnLE5R3/91au0XAaGNOtaqqiZ4Fr+w/J
mKvzUU8tsUKGhmiMhnPwKVTkVYCDI5/7szyc3UW2B2bKIOhu1v1FGCWB78+COdo4B6GoMgJGXh4W
0mFTU/F9VIlMLxwN3H/ZPy3/SVjnsKQ1DYvmhBZDkhyg+i/9rmzq+h9jmvUnfvnULMXOiLNtVGM0
lkhJQDgx06dUQPUgM/KjGiqqd/46va9mQdJt19RbUUtRi4bFgIw/fnC28yrxTZQgf4zVXC9946Zs
w/KG4guKSzeFF8POJHBl+AR3kpuUDedZdsmq4Sy6q935YSDjUj5mrbRKZmXL2yOzZkjUndbFB4yN
USqsQzyHIpyT1YEMy8gNVP3I1I0EWbtt1Z9WPkAAJXo14Lo3FFp4YRpOduFct0prctjfaayIbvwL
CVSF5+vqMd+joeMHFbW6yDuXG/9squoGRYaxIXxUIP2i9UpEsVWyXufBaIDiLr0IrknnMAk/lGQ/
lVg+IbE0Uc0xPY2aJodeb/EuBiYctHoIlqz1zBY/qmv0eqIydARxeSZeHBDKKjO0/5og8ZezCc4x
7CxjguUW/SDh4pzK93yy6KRtIoX83blil83tqaj6pQwR9zcAiD8JOeLkc9kqpFOnvow0nnKbfAcb
e2WlYE5e7IXh9zi5cbeS6iAROFagnYnQsj73wOz9cEr3Oi7XtLsh86H9sCBJAHkNHAXxR+f2NXg9
3NQ/cXgGXM2VpzCDjALAJ3MdbBTmShwGtZthOFFWQWJJ/hpP6Z40vY0TEgLPuhN+iDU+8doovvjQ
ahGlTPhPa9J2vaNL/una3CYkcrdsZo11BKk2zR1yV93MM1/hAv/1+vTvFQ1lQ04wiY7DkbXAu6yg
vbpJX1rgzrQaObAy+LmUJfy3o/frc0qlUmj4/G1tpCppE53DmdrT/vckrspaM7G17v1/zoz4Gr+T
KkDu4E681FC4UW7mr6w6UBrI4IL0E6uYlkBQjx8YHeqORNGmVei5F5AY2+bBdsRvYod6ki25Wnxd
OkjZY1gpgzi+XZwAAjJf3M6Whq0efhsPyCclNwyf7T/jvjucpeTSLJ+Q5wXtNgJIvwa2NsSC8RDD
NLrm3FYlQ9LHI79u/kDtTss2h5bPhbffl6PMc/jZAi6NzZLJlC1YtmXgkZry7ztBTizu7KD5vjlI
tnDuobFhya9LHaDagso8F/Jp61zybmFFNjDaWzR1QCGuA6tumPdrXwfzKPIzi2yv7WAiOVWlSVmm
VRPl8JYvJICtup6pXnpTSCVLo/V3bGvo2tQhF9exlGN2tuoVws0gWNvp27TND2iCiAb5DRmEkJji
vhZK0KLmIJMgEayGhtoIIVOlf/ZCAbslJeS0dGRc7lMCsyIu9KlDDhlVZ3uz5z7OMbL6hyp9ccZT
iUY8H35oWqfhkqu70QTgEazGUK5uLjT8lx68JGrVw9ebjQXDdls/2NVBoRBQRDySAOdtcRkOMYav
sD7sW/nbXJkl+YnjvzMSiHGbSfE/ZeZkWOBSVl7ZCwRmbvvmC0GmH9M30aJLYBmCDnu+t/hzdTCp
azpD66/JxhTaO2BSOkZfrN16fsceJbJ4lazeui9dnh2fpJUp0PIgx/PTGbHRbbBnANFOabMVoS6W
3pzNulVxaSXkG4ig4qOxOyLQVU4KAQ8O9F64HL4xy2nX7XNneClSH5SrWwiTfn8FwPoE/1IA4D8N
9P7cK62mdTlyVFcJOt89EwHFS4kkgTFqhzu629BcUjGBB5nfYpIsndYo9ky5JvSX0PCbpm3s02a2
/9aBYW+obNPWAzjWaA8EB/hqOzY6axnDj0d7E+axhkrAQ74n3AeuSOrr1wuoI+Lll3VGKZUI5RPX
G28p/CBQ0MFh7oOrpL2XVG/w+sCy2GicqDp1j/ubQYcPJfH4Ebi9YU39xOBA/vDBZ2oa5GtVnzC3
Ew9wBd2lPa37bcct/apDofC6JCChy2Rqscrr1TanE4noes0Iy8VsTrmvyZgcySW52Ixcd8rvyrG8
aZtyos6BS2cfKMskl2OCSbhHqRfbdkZDcVxCHciQWXujqHgmXlQs5Txc9VEMXslKRE7wJJf/onF9
uOv/SoMa08h1CMExnanb5wBr/J86FX+XV7jaYyOr7lOyrTjOFW6sur3VT7lMnORTPhLMI1dJTkoa
LoXsitECBN2rGm/N8KDe5z2ksQZ+71MGe5J3qoXbI1RyffkAImJzWJYXNUn2jigxFhLWPZ/74M4k
cwgknx4hYhQMNjkRE6SW7EUJ74R4bKOD6M8RdZ1mRtNkMvCGxEATfMIPIX2Xnux/73qhoU8Lw7SM
cWQ8w4e3FaZc7aEKSvkVDZXGjLBG4MgImZ3hg4QSm9iQd2H1PQNiVVdm9DZcIUBL6JLsVXeePubq
1NavPqp0y0KC9kpZ78C7uy3+RGLVLmHLwu1O2J/ItTp6Ar7Kfnb4tw3ryJadoM0nH1WjyaZVhl9P
8dnpIcMqI4FSszuxLKpIea/s4jzZNdM55J5ZA39iiD1yJB34Dm+5FPHJUObyA1BdosoPOFoAHJTH
O1wmdAq/5owMHRPB/2wAHFhR2EbVkh4MG4cB+bHsEX3JuwUe9ch9lmp9lxvRkBBD7abk+o9zbeEx
pUs+m1wnyVJWkVa2mDO2N+Gkqr7g5DI8o0UED+wR8+sVV8jxrJ13OZvM0uNhrnQvADgSYusj/UBl
RmQJ8OuQaR4oKJQU0N6ft90SdkTs4fEGpeEskYTry38jjPwzclDjLdRVDFyMaJ63/BIGIu1LHS/Q
PZswqKa6HN305/5rTEZcfxDvwT1wwesJh48gmTa5tIfFlR659KhwnkPUqo30XyPaRAoWyytqmecf
rzqwYzeK79VbTLdYQsaXWrVuOvpi3hlqeUPALZjWSP8PUMEhosluhXhqk0lU2v0t1vtuhuzAqXX6
OzbZMLWyzxQQ4vIJ6JcGGfCNIbxFc2wc9/+HF8GyQSVlzvqOXR902U3oQh3n0aUaBnqHY5l/fXRn
41V9gDNBhFh8d8ONdC9mi1RuV9kMxrBCX7SIuRO24cngKjnslMPHBNnfem4zhAdoMhByfNVtk3lz
1SVZG2GRAme1In+EQZmNS1sgRuSW74CS69JA9GltJ8mMFUhI/oawsFgbnk7a1lrS0wuUCx0Q9elp
VcAF5dCCg0qtuBlwlFeY9LD66jYsItQmiWafxb6FddXQgyCau9+i7i+qpQwjxLHcG+K76VO133fj
xfbEybDhIiiaX4FRTsekLKTDGenc7gnC151Y99de+8FXPkCIpKmNytKkp7U8iHsTyJZfJtehlL/0
MLaQxm233pssM6vwpsP3KkzcKZGMf/ew0SDia35XJHs85ki5oeyNBrgVtND0v6vhw0Thw33ZFxtg
8uCpNaeQK5arX8jBB6lRPYiTGrvnbsLd+DHn3yCbPufQ2t7Xv8Yi3+gHvqseweCjx2swkNpfi0+h
6z7m7P8JsS8pZaFtYJF6eT8fclzT+k5ZWrhTb98ZS45veWkQ0TMLDSYYfa63jE3DERi4Ec+Cj4AS
gimCXG4AUyUUqXVi+CFwFlIo7H6fQYsyIU4udIf+0+i7qirdIBwVgnNnfbpOFY3JvLPs6rhths1K
LXSn/u+nkiaUmDVkNTdSfpbchSpdF346dmWtKaiX4h5ChwCoyVKkf8BUgfG5ZRTSPKGy5Qm5t+ov
Lxjm+SNlEZjGTH1fBzMHJ97LjFZt+Cq5IXCFmvQF10p21bsTNp08Q5/Y99MkdQuW5Q7mBUXm65Jh
9Zi20fJG2BGqg8BunSXi/URXMXULGqQCKOH85BePv7EDKHPlu4iax4dim92txVTA1HNEiqIXKWoN
OZHhQB0RMMST3nIgomXhNchVUXsMjSROYi/QEyTkH1vwNFsLu3ThN78P+MUmPCwGoateWo1UoOet
2yL8bnkZVXNYIPSqUZPlp7QpBk100Ho0oEs2I44qIgOl971uonmigT7KvSEhpPZ0JnsrSlYZNTH9
fDZcZlCZtfs908x0Q3myOQrNbIRE+1ZUUNEhMRTSJxdeGEcIhtKSJZJv9fF/T+qA7ag2ZW9rbSeM
Z4PSo4bT+6HyzLcaJU8AIR9j5ICc9eWAn1KnxIfKeabqNRZ/Dh8D4lBCDWVTArP2sB26zyXvs9zz
9tTX1LtKnoezkww6+MVAbepqARyMnraUO6C0410um5C2EPMrwguUnytkajz2Jxnd9MmS6qntikJJ
5Txeq1RIGyF8bseZDqhn373UD6zFtRnrhaIJvw11tG9dQL1fhzXVrb4v2ohPYEAVHrGV+7FceB37
bedOaMmDRTyhH9G/R+AnVgdR7EyHwSHqQODslitTpdA524sUa+aODC16+hSBi2sibzkru65XgpPf
FlrmO4qvr3xk+Kc+gI6p1ZfcA9lwbCpqYJbLoPRuN2M54AnxZKE7iAOVxvgnw/OYctO5eyX/t/i0
rd6uLTlcJ9qkCPqIfyVU0+xznf6jzQkEpq9PuNl3ZlDgVp173ZnJ7xpPeJhFrMiXJeqFGc56OpAh
6ZBPUejrIP+IrElcZgRKgZuvs+bR2lKuGsFLWYvWH9sdbwlox7aMgsVYGS4IJPwSsxkIlxmNRBvY
ioIrWQa5Z9ryMM5E2s+hw8X7PdntvaBkyhqT5+x8Ueh2Xqp3JNDRlPSV11S7Jvg5WRYeYx1SPJek
4sQuX2Ti3V9dY7CJ35l4H2bZ74ZaHdcJXKi1fih0C3m3Bg04/7ORuPiQV5ue3wgzMIg3TzgVHpQn
qA4NzHRoEfnKxzgACpHEAv6XcEF+McPnSEdouDSnPd0rOx65lFy2BXydazczB2P70ushrvSvNdpv
FOGkO/dFCYB/Poi6xdjwhWHTpySLZ5HG39L4IE36BG7p/ZaTjSGbaFBDUCpoNsTTCOplgW6n+AsR
zqtOF863vEzypc/BcPS2RIY5BWcXfQj8gnj1uLgFJTJ1U9zFIL0bMb0fqidhS6btngEzh9cdogeO
WvCYzHM1mOixlki3IWgYkxLg8EEG524wZ5uPb/f2Kh8d52dF50dsBSPuoqQhJudAARBkdcoE1Ela
dJgxORC3alCJXdscD/ba1g3bXno9V2OvsTFEUZ96AiTzsi8tUvkM7ACtopccK1Mvf6FQpWafTIDM
K/qwsfA3W5BuyvSAcxoce44oqKoTVyOaSkxijXmEeG5ETUDtHdXVyq9rfv3uxyMgTOnxyzsIo7Ux
pYuH4HZTZ7sxAsCTdJU7acJDeFhTGoGc9zyrYwNaClyHp4IiQF1TM80yPhykfeF2YNlVwE1aRAEJ
91hwd4agTyC3RBo5snRU5MjERZO3IJ0ogCJaIZNypzqKlZ57NNZ0gAwHL9I27iRgbhNjOn7rihjm
VArk73J3BDskZ26WM0CmE7QD/k+P/kb3UNbs6Xg+eya26gmbZc1mPT0M7esyvSP1TWFp9mX+3G7i
ZCdgYSIGfHVPEzsXremn+auwkegZhgB+XMMDsFdS1KHJnUvZJz4DZR8unfZs1+nVzxvkYZuJI3gx
Cv5mINeNfn4lQ2yOWXWkJMwQ9Bb061Bh4b+ETejktImEAS//Vu9pQk6R59Cjqnork0NRrKjCM7Oj
7wjM9F2tTZjWvGylftNSjeUMFgGr0+hYyMILm32r5wf51xD5cf2YFrCrNdbEUXDPRCtRKpWuyfOa
4V5IaxIZbzE3yNvTkZ2cmW3K7RtAEc4PYVDhuomeLyoZQVE/5QCWa238B4LhJsrk+GJyR5/iLhl7
c0erutqjDNYT1yn/0+MxxlHGE4zJ/ts1HKaHOo13qfMUwre26twx3qs46bfaqVh4etkfex8CGWaK
nXNSNb8RZRHC94UwLOSuo0IcePIOYQo0RQEhbNxwTHUk0W9VEDhtuG8WMC8Y4+Tr9qEEdQeAmgv0
hR9F4pfVIOQ3UmOt8w2cpLHh2teefyKtO5fD6D5WzFBm0RqMHX8cUvA0BaMxlyQzskZjLjGgA6nE
tVb+E4kzdttrHWKdDkbVzJzaqjPZNGLGoXKKl/EOOnh1WDSU/DEXBeEf7Tv85aVNYxbMgXuA34GP
ATyZzSQtEhwnzqdzP+f51OwTLMQ2CmUa0qp6twYZTFz1DAE0VVgRHF4BLmqBMlWFZriihU6W+R2f
hhUDmeu8M2DPaHrKfW83arSduGeGqegy3eoWYtNOiuu2cjCLWA13c+wHRjdpjhuGr2DuDlMoM5C+
GMLLvyLXDUN3Bgc47dJpIpR6UPxSdk1m/UxdNbqq6VYqUKcQSGnJDJgChDAMEIVCeKz2Q4qHga2w
R8m08xf/R2cM5rB1hlz4L8x7ENar/LxH86d1MlDPI66UExQJnG7lYhdW/7O525S4uJmbOeJCQhuI
pfq3WYCxRzquD/e2mkkrGRc8VIR+ojJiaMcrlgm8bIGnXgI2uw92vfzKjFW5q7eGX1rxiXh3gkLt
V6ar3jiYYj0qJEMQILD4sScR6J9jkLzBSd0udz9X/K2Fq8z2HqDLnkpN2rX+xcvqFGJhWTg+1hID
AybntgI+btQf2JCvOraFW4URsKIWtc+ZOBIrIRi1RuR0+VgChDSvvM5xJmHA9sxk0Bm8F6D4G+tm
geY6q/W1N8hkbvV9PKesfhdpOVdpvS7LnhGVJ5xM9noBxL5guUllIdrm4XxBtEW2lPicZuI2w4gU
fJRslB2Soljc+pManltSP/IXWCiAH6cs8a7avcxC52Q3v+qNzqasGbWBl7HLlhE0wU2z5Jhzorxf
bbSXKSRysAADqEwDrKgK9dMWTWs4lYdxWySiOo7HBMXa9uI7f7ffbhTqHSmVt0m6ceoMYTLQcvln
GUbmlZfej8CtoX7qiJ3YPnWnHAta46e8nGnGCrh+q5tQRgGjNGQb2m4LKktwBs6IFTqYUIxtt944
uNSOInN2HcAEqpaqfj9fDaIuNdQcXl+WSLPpq96M99YEVYkZG/wvcBT6qBEANRLvkxpC/MaEaSAp
UUGqW8do6i0MHAWhRlhKmbXemyH4JU1i37JYuG8UJtHTGepY/nvplgNj0uG2PIf+wCfdnnq81Eez
Z7A+eTKbBQf8g2/fE5i5V/prD7h0PP5VlPfzAYtGWYrZe6BAcbHyvsSR38oBqvSHJ5UAc0yqPwMI
g2/GeS16A9LO3X/74bgEa0KyMUjApeGZH4WN2HJnTVYbUpYHva/fWxK6WrDUqqnVMOtuxNVjUFid
GdfYr8MRji0CAOSm1nYT5To4Z+o739vpKJWFiPGctTbKVfQ1ZGAw100tvFEspCf0pp8S1nkiy5y5
cWpEyDtqc4PVKJDjpuusqC2gsDw8VtHUGOb3sb75L0hk3qPs7JnEmfj9MTYaDL39quTytrI7+o45
mUGCOg0EUjOEf48M9pUNsX69ccAwQ6RJ1BL9CUzp2yr6/KZkFJyFuZbDQ9lFVzph49YeSF4NvXR3
hJUZLkERSH3cyp99hdwy7Pq0wKQPuTgiI1qxaXJmqIiAsYCFt247qUsZzOnNzZGx/ZjZDcO7gyzO
7YTaapcESnDcvTw0gnoVZ5lEej+SjbyMSv1BD4f6ZXVIgsAz+U2YM/Gd9C5isouuGN/IYjfT/8s7
1VmLtB6W8gavoUJAZOYduubmj2/eO+RiZt8npQesRQ3z9+QBPNXc4zBsuJ0UqtwqAqWaVWYx9z00
t4xCUMAmKtmABA9cOpnlQW9Ov1xQm8oxhl9G0ZXKd/733vWSfWngitbpNPC0JewetD7NCrzr12Qt
KdcBAV4Fx6e31b68LR5Hu8vZrHxmF5HOM806jsHpo9YRopv7GY8pR2RCJ/LMxUfWLTRfhny8io1b
ZLHzJX9v9UaSmFVrptshsLZxeEcc05wYJE5/z3HSnJIsPilDVSloNdYWo9CIiZHvEcAjwgv8/OgR
Xe8Rwo3iUfndpEAGVOr1BOnb8qnlfGVJvax0l3YxOj+2ix2J7/RMA02wBLmmKNZLqgsJ8rdr6jG1
KRt8xy2JWgLYiyNCTPJC19lgBpxzXXjWyD6vIYXV1ZMgk835NluB/WIq0pmydznnYmBdSb+kWzgN
OBlNfc5bVMFpFmkZDVoK6VC81zauinZXrMTYMhGre037mx3+g6rPUJxqw9HDupuh23nRfPTwAQqG
f73ojxzpsf8EPbCds86JM5kXrkKEX2KgIYUXYmGKXQv9P0dUjOCioq/g8rpVgLX/iDNWkmLKF+oz
Y7AIlFxP12aMu53G2tZpV9AujI/2YK8TKuGNLcuDbc2U90zTK8lnDfAjCojSG+XtBRIESXHEtTYg
bzdXPJ0K7AG7ywvJ00owaB5b/qN58hSQKxr/XYW+hydZrTnIt+BamT65gjtW4qiu3u2B9uD0Q9a+
r4hrV0nogWF0QVngnk/ewB3QPXhfGL1bekL+sHjqEol1i11hyS3FzGFuy9lLY3nqcAyJhSff9SUQ
dMXj5NtVZaa1zD51Mo6MRQASvjd+qlz6xEOFOSdln9V9AYv8WsU6aP2ObSY93RtPOHTlBjPuBlHq
+Rr09webFQnAihHqnYjLy0zMMa6j4eXw47BfAVj0CNx4kLVrsy6+ishKmWOPAi8Db2ao6CNo3j2x
VGFCn0KBB8YeFPxuzcKZkIQLICTMA33mAYVKwKNzzpQYjrXOhO/wdJbH92re5Bem61UodmtHRMdF
JznIKD4+3rhIn7KO2Vt4M/vJGN85/Pj4i4NqK7LgrECFFYvQFmgaBewVyDysou+M2Ra8O4zbKF2k
XzMLXbWJ0DdjZeoJPKHAagSLrgxql1Gzdq1XWDdQtln/klJJVC8GoYZD6ExdbCRh1OxItBRIM3Et
qYgP1UcXn6xzBbLs2v25u20A2pUz/sF+CfQuCovWL6xizoztea4+o+8frUxJQ1xIgwgC/kgsd/wr
C/gbiwtEka2X1rxzNKk3a1pQzao/GmMPB/n3iw5CTb5cUDa16GryBl/cr6eoNYEdIwRRZmECCgcf
N7J5v1y6qafM7xsg26t26Fcr80ZEN76d9GXnxSqt80SR938lbSwGtEE/Vmx+aCLLKcENu35qJi5C
6xxTZoosKEMN8M8U/PtSgHxc7zQGcJd4Eg98PaOLoutjLX3vA9Okl9L+D1rED3+HBB8qgCg6B7/X
nRDLINVj/1ExNxd+y0332ZH4eOXtgjmUTLrRuontOqet7qgamck9Txl+2ef1zRa044NULBwYkCw2
hFszR41uckQF0azhet57v5lSiOJ11QHz5M9W6RH7bD+Wh5d8hAuYP2WoyJz0OI8nXQxcX/GX3H7y
Mb2oLRPsFJKVSraloj1YmA/mB1BvrmSzwaSZQa2OP1RFo/GGkNiKdPcgKLQ9SXKMdyjY9tMC4ewv
YyLbZNyLWpl5pxmqkHzUNS98xS/t8wWGWMm2IM0k6Zt3Ka8SW6M3x7buNAuwxIhV4w3N3JSejlJe
9sfLdEzFx2ja6xsvugUS5JRpeTCXyaRF4WYRvxigQJnZTyzFfzeV70OqLOjB/WLH8s7D11WF3em2
hZPzimn3OQe6lVz7t7HppJoBVJeZE7461t3XKryYj/TCLfxI66F6mByv0NTpeS1yPtnrxsuh6i3R
0FnNawCqPbjbEQdgaxu2Px13j9UWTNGzkkdjETgsfMKJazbGmlh5Vec3uZBVHUbyB1atJDBPpXLa
cut4UDn5MYlxqkYaggQJajazDRlWGoJ9erzL+KDS3UEIZw0ecdfLgidagPVUjvNUREQOHOZlIoDN
RwYqWFknwS+Oj7oA3XeKuLh9rLmotcWiGgYI61qN+bT+nqHr866Rjc8sfI0ExTinZIKepYpYqVCv
f5DBxh3+KBc3vEJSkJpYMDQ+N7Mw2np6g8LAnnNeUFd0L9dLmhEy55gRDyoPB60YCra/yu5kCcyO
b5vyk/nvgjoQWKWhQUTQkc/A94grvKlxjCAmDZm4Ff4jjWc9Vb/9PlW4JiS7Zc9wAePwQIEGOhDL
9Ztr7bSDKUNorRtaJ+TCH1fsjIQK5g8W5dbIJZPKa+wemGBD5udVao5S4DHtXg5kB43ytJ6A8Inr
m/9R19uui5qZpMtILWQfQZHMQesfONO1rAo2blNmxUC2IbxejCFa3yAA4Z9Z2j+mCNZhp1O4bqN+
HKOs9IHa1dMh84UrKP+zQf5YKLzVzzB/hI1HvXepJVAy2t3zSMBeeaRe0vZ0tgehli1tIF+6lyK2
C3I9qnEJVtXik1ZaxJeqbQ+JvvLCI8iWw2wDNWNktkqnXBC8SP3SG3dQLaSLrm3WTdvi9prDOeQ8
cvgKQv6RcWcUihZWD9vrMoWoQGd+/QUah63JRD2f8hiLvuZOtD9Y6cQEQ93kbev8dRHYmoUHstm7
Q+bXpKAiFMvZ2DRPYbGduvFhu13mnbbhdB808OBqtDf2sEvgVS8VIHFD02t7UjeZhszgiYfXCbnU
xu4dynfLjj6aHFPcBIr031CPg3SrzXvTQuHAtswFDdBGOX+6Yl1t4Y91ET9Qh2bH96CAgep67dJ1
O5aXfx/t8NeF8+1noa9Po2+OL/33xa+ke+RDq9Vm+IKewPoCpYYCzAoyX1KkjdeEPVIj0zyBTGEx
okk3R+6EX60KHA6Yca+ze0PechMMAUsgA2RztdUeMVrbL+xvzBobizvn0bj7pzeAM4hzyVwS9LKw
BaNfxta/a79APPro8i/+s7fOrecUkpUsEI3aSfIwEfhwYPXIdyWnjKPQLcLRkkm4zfjLXHYe6bh3
BXPIfelhO1WlSEL8q0Au8faczrtwuRvvzLKPesppgS0wbmpyDOrcxMsWhEiie+nTnQxDFGJwRRJG
N2CITB96gNOCf/Xo5Bftg6fZXtdPvtyap/+gSJ6ytUl/m1Vu7NeJ6T+VlkHnv/32lLFdvm3r4eYT
CyTxQ1zVsuLw0t6UjmO+khkwQ3UY5nqlx/dYEJwnKTdQoof9MAkkK1RdfEJEsEvpDwWkyJP8ndEA
KaedMdTa94j4IBEIHeGv96ikwNpGTNVXGmG/xj10lbZ/XpZEFW6pkZGFFL4/kWy4mLMPyL6KuYEd
i9AZ//mdoFYbTGIac852SMmy7ClKu5wA7SvBRlPuzrsu2Y5hxy6/1j5gBYGd+D46mgEfS9HftDEJ
ZMmUrE9sz7V7u9nb6Y9PPhz7oDR18pOk7hG0IgBk8/cwwBEvPwEfWx1m3DcW0x9P2PqOhnHCAJ46
ydIKTTFpnsDpssUPtPjjb1YHcdLcnhI0ys6zi+Q8idLoNwlEVR6TdjAqjR6TpTwJ2XmSMQDhJ0oo
MaLngkSrlLCXTrhH+X9KSt4AirzD0XDC9wYsAk1tBk2s6rCkEMETKylKnU8I2WLX2s0fmrkXJRGq
9w0OilwwVcgossUmGIiN33va2nBVwbCqTaGHOEeiwsEnmdTayATzGXSZSY+Bt7F5ErsskfUVfP4o
d7skoEuXI/Yu21tnBO+3s6Tkf2PZ3JZK2LsRGjBZFDRGYVmWUpP9skbLHLEbRHA5LnQ8NXOIxe2T
jA4Z9WmwgvKcx+zw7Pxi0BpgL6uowpH5auzcmX36B1WNjL8CliSgbRG4wcgExARhSaJLCaWUxaq3
ux78+ESZzHnFV1S3DUAa8VZJmQPv7MUPI2ZkC4N/WRrg0aY++CCwHts5eYvmOOrt4wA5B+OBP66/
wlkWnjGM5+uyR48NXkWOlcoUTbV6c3yyiawd4DukfVKGgMkvGZfsuSgHaeAylylLEP8JspdVsVDq
rIOuJLhnj+3TTeJz45JQaBpaJLBG9h2sWfA1RECcwvLtKtrzaUAfo9c9Yhg2Dtvz3DWqnWGaai3X
EGQMIOz54BJ8F8t8I0Sv2Vq8jV+JHlKcBfyf2QnFinbpgxJ2agOpKy/GTJRYZFijoDUib1PK4PAe
yovU4r0pRzyYjya3OnaRpbBn6o4z/DfzivafAkSkZ6ooG+i1byTxfoPIdXRmK96/kWPkzr3ZeqWh
hAkyUqIM+6YlZhN8xFs+wjH6AzvJvRhQQDQDj3l3n0ov9dPK0lDGk1NeIz5EzVwbGv6lubdcDQ95
qcMw22H72U2JkM6CEfLRLGa5Z+R+3OJMY9XKElg/WhIDMHtzYSj5TWwOZKgk8QO4aEgp+OLuMQtX
8Kv0J1w4ga5r+Zv5pUxYeeNHnql9eyefSYQNKXPRuQCtrgtTUReA+44IxZXRA0FXhtC4OqjAeWov
tYpqaq9Smaad/gzNlqD4/8clqm7tr3ipE7RaLPKmrKjq4olXhzM/2UmhUnl4zd0GF55dLWW5ufj3
jdiM7/vYJefdbVmxEEV1DBemBHzJzdwM0dLU/2jJHa6AWoJJpiCUB41GMSPCwK/cwTGeqej66xS7
HK2Qu6E/yM8rF3xuZwR5OXZPJwduF8+SMF5GkY/AkyIZFe9uf1G4C+3qsjWqoA17SqLN5LClZpXB
1UxLv838Y2TRpe5gmFL0ykq6zvcoTcOR/3prPG6vNSD7m+udo4tE7AVjrRy7Bys0+JthtYilsiFw
XP8nsHwdC6i9gmH045YNTc8gKLjpiwgXmePybVL9zfIYW9s/O1cK/FqPkxk47pKrGsHccQe7EZv5
3wdn7aAdx4fZruMO8r1F417s4uMD9hsHbJTP7SIW7z9bX0aYrlk74267brd/1KXMnncZE+XUf+5Z
5hKEG/QZ7ltiBppIFZ9VlFjLwxA7hBwNoMUiYO3gbcRz8EloAcjv5lccelbNRTO76c102bcbvfcm
NDoAqge1CRZ6UNJXZ9TeOUCty4NlYe/zs2b8E/T3Yfzm8ukgn+p6pQTVHo4u4pac5Qf1DW3dud72
A4Pp/J2SP4FSXYeF3AjqxrD7rx8ZVUxYAqZh0B66HIJ2I2kAsAbCpJvQA90L23Anogyz5mX2sxbW
UVbX5R4hSJj3epeqUKvXmf+WUD5CjB+/sw5zMP3jb2sXcSZymGwyzTqKcRV1kIR9jeiC4D7b24fX
noGwd5nS9aDca4aHBKoNdhSoT82S3YPmt9l2sJIfjI1iqLopNof1hPuyBD6UTWl+B89grAxJWO2Z
VvJ1i2PJqJOs+v4TyM8zcUyRH9XWx2ite/vpnagkrZ57pQseuHIvrxy6M5aIA4ooIdAikS8Jmm+5
c764k0zBZI5ihDMKkWjQbEjB4s2YomhGdRyHFiGNcuKH5dsKdGkckVf6VPh67maeCagatiMpt8Ax
/goLr8faoMh3LlnIBDMtlCZAM7h9dbfBsKR7UvMCkiKDNl3j0jPFHv1lw94G/dcTRG6V5vkPhc0b
fzsQP0p3us+Iey2jJ+lRyugERIZHrC20Bm6poUbOL/jzAR3I9BIm9fgBwvSRJ8YdqS1McXT6e50W
wBhfLtOq8LLSz7/NjXOfexn9JhTrAK9LXL0cTfFVrqm2PFgOX3aG0eRzK/+l/NKOC5A87OV/54Sy
H6jILODXaO0GDjuWbxLSUwgJAqpWGtHicHVSqF9U8GO1WzqCIJeTLDBopKImo8Tz9RGI8rcIH3PD
BO3660Hr7Fq2MVGyDeIMjXjG5QhlVVNuhQoRx3otAgPnbh2koDjwqKxBwZluNcFPxnYqZvaVW8M4
dxODIKiDWYSzDf+VJGphHahypSoKWpvZJNDxujyKuvv5F7gnHxiIgZu2qGQbURGuVUuGOQ6scMmh
fI209Pv1IW79aqmra8viY/Fl3S+XPKGZFfwZLIBkYXqC/Rzf1D5hLV7klJ2Q+Ju8sKj4YNgxMksu
FPvylxrSHnmohLeHZQziRRgqi20jiS9w5uZCaQd9qSZH+EZY9P4Fdqytv8ZNwe6iuEbZ8wHbdwHH
TmSB7+0X4yTz3la1oa5WNWQbHtpyBGUC7SXwuuZm1krgkzBMkkEvsawT7HN5wR8575jYSZnLaKR+
8pL8keaLHKYhYho3cXSc3HpK5dKxH7QBelFZPbQj50HSZBl9aORt2z510jpsO1j8uD2U6bmpCdXI
uzpvuem7zWN17l1224aS5fFZMDaMdvv1v3plL244j7aMvzRmDRlgUIiMFIu0Sa51sQr2ibpNb4Ae
wJKG2Fw0pUilNH8dm4je0fkB8m1yRXUYRSvYfi/rgn0PK0f532tdT7SOAdioVLva7hXPgGlnNDlJ
caGU8eHhSYsqMJK+4FfnHKoh9xWHBN+oa+GfwAfjWL454sGBNJrgQlSb5jpn5VbUbLMTT/Ug3SKh
EBrTICKKMeHYPFQkPbEj7IpnBOBfUESzTna/+CDFfNreItWRj7q6zjA6lXMz8dylzQ+OmNcSkmg8
ORYB0RoFQDozsbjjSPP89Sg08iUSHdRnIc5zGMjkJeLRF/vl89bpg5s26R06wZV8iuWIjf73z/eQ
YeFVdWqRJWOSSCkkBxkmnsEn7FSUOXWUgT0ti9XCErvPBvuBolQLFDkjKbYHedyfIuGsQjwfN3Qk
sUh+G/94wAI/vbBi0Glx3IBUpqZMIm6nMLHWoq8uk0qXzWIWxbgrpvkKpyJzb39wbhE1V6YrKNfx
kB/5Fag23MFfgeQ9/FnwoIdTEM9MBjeRGot7n0nmvxtO4Zv6NZLc0MWqz/5oDFvWeWzU5eoO2nSP
j/ZxKCB5LrM+4muF3kB4ByMA/s8mtDCM7Lgr3z3gcsXYjEJ8Oz9axkOEV6DZp7gFXvvNxlmKVK7o
ARB+jBMUGGSv7MnRrsYkhnjroBLXUQDfuQmWQ3XynPSAoMA/AJMcZ9cvq7CblQng997ZpHwORh+d
VdcfRjC6059snPYRhgB+MauMRNIUjUvJMKxLM1dsx/SyjGiAufaIDCl/yrDOhjkrBOVSRpw4XbCW
Yc2ulp3pH2DYKPfXxHKcuh1aLXpugavIo95K6ChYuFVMvhASr3XGlguWhmtgBTw/Iq9cZ6InU/WP
OJWRhhLrxLeGMfQKOf5mAEiqqrtDZTNMpDzWp/HkmR1jH0ctGmD6BHCBnZVQCmbvd1xev97d0sYv
XVFaU+4ErB9n6hxuRTsW2dU15IoWWG88+UgA6tGiCcrRkpKyuQaP6WNbnarr7GVCXSk6g8pCQEZB
Jx4HBlYy5uwl84LA20S0Pw4Y61LiLN5jFqwLFC2X8EmezH7fXKaxYAs4OrWIEOF56o8a1em2BN9E
n5iZ3y7kI8IcN2ztym6jQUUl+bmVwws7g0Mx496h+N7qdRVeEWTJMuRCuQge76nybkJs1nQIBE5g
0tk1UeSXyAS9iO2tvoW7vjWaH34qHDAnFzOJz2krmmDTSG7/MVGfkwtjFAb2AVjcGEIoMjS655PZ
NF3jTXHy1JWAwoP22+I7KDfW7sULJZtrW6EsObukHIctYNX84TI39OsXznMYZzmWGYIG0TKSw/Jy
66qWaA2+eq3J9eftqh7oeX4ITi9zNIXUw+6qCaOidM4KTQoBYHQbE4xJkH9FYeTabwK7sYH2OAng
gogzwDQsHMTRik+KoNnlW60Zrg6dAeP+XORtWhtGi+n3TNObj6x1hl33eC+RbrVqDQv2RqGCywl3
dau1xGnCDqhjcxBJijGjZ90GQ59yIDJFW/pKsteESOpE/WwZSeMkhI4rnPgqgQvOnrTSYDi6D6xx
m25YmPc2l5ciccROlbME5up3ribaVIPr3CK7efoi498XY3JcKIu1bepRTCea4KmuL0/cWg+LkvAL
LI/YrmjWlBf1k4eXVeByaOKmT4ADrJcyghb7tKW18wVjA6c223jygCUb2NTH8LHwk7HBDaXjmWec
HNUJ1xW7v+6qeAwvZ5LZL5NM3rUycpCTd37JW8CMCyroQyRIQ9W3uit1oPhm+0XOuGsZ6OgFYZEh
d6lrH7ZG6AcYkmJTZQlXIZQUz3DNBYGdK1i2lKmqI/rLByzFbe8LJSFirfi+ckCLuoa+vL4aBLPt
uv7AW7h7uXVApvHK0aJY2DJPNT6GzxM4CJDua3uSc8cd9WYZu4dRTitST14Cjw6T6m+4J/NzX20S
Eyan2QQeTGWp0hx7dHh74eSgqOry7ptE35kwEJZubUxkEWEZB+KOLQwJwrYRExdriBfiViGqFsVo
1/rehPV5mthPW5h49Tepw312p19ApGnhKVO1Jx+v8foz8pMxXgFPbE5lK2SwyOKeh2RPxKNmloch
LoRHLCiF8NOUy9GnhAqMuVl6Mj+5GVP0LSwh6kPYOH6M8uTkdt7yy06qCVkvxtFiN6vcswbhcWTe
XeUQiQ5wZ5RUI+FbnQUuCYXHgnhF0dUewTAQWlOsI9GTjlbqYDWg8eYNfl+mXSDdsx9JwEMlTFwy
Jb70cBjy5oGK9CIfaA17Q+hVRlNeQYT+0CxIQoC7ZGE9OQPzwGKtlhGOaS0OQv1kr0bwXqM6TARy
qTOLAYj5VIAF3zkW7gD0TRbDLho/eXRKSn0rH5VnRATj4fdTjoUPU1ynV3o0gvgqi7O8IzhZjFVX
TJsyOfdGPUui7WQGBeZxka1UvyR8p4PRDRdWK5s3DkrZxNO6JT69gWqTi2J20rjTXi/0biZyOdrj
dR64zCQt8aIenoYckqXUBepH2TygGzZyCK071x3H3OhczMFklrOCwRBMdi1ZTkYdWS5XS2ynZoGl
SCGKi2pz/nJVRReinCONTVbiCj1AQbVN565JMFayCfA7msbzdxJ9Ry5GcB77pffMydMUhU0RB2pi
rfAAeoHyjSvXEvr9HQ0c2BpSxiYh6k9IR6PbvsSN4vff4TwItVlJl6gvY0v7fKGdDjR8Rk0ubjiz
taGtSXce2JSSNpB3TV8CX0jkgYDJYS9iFzKwc8JrqcmLP4qYwQXJY1Ivd+IcEHqWa2vtA+MLW7OI
+5YlyyyDxqwyo1m1TwTM25d1AiZ+V7YnAeG+xzsuzHFU6l91JdT+ECrrSwsX6uCdZCWwqleeITIU
27xIGBgV4LPdK5awbYBvNQvRxHpNi3IoIehmlTnXv+63GA3GzfpoLvc85sLNDp+6Ihf2BjY5xH6C
kmNEFB70cVaz1ZZTa/4EAHOVU6E7O3pTErv3Q+NAjqBTqDCZ4mHqEKXs68o9xHJzwCaHnGcBtbvX
W+uqhi2IY+T1CIuOJLvFZY1ueC6sSvKxslQrCx/6sjoJnwfS1KIxYOunbpgNc+HuceK7XUn3d80T
Rk45hBBJXjoqw2+QdveL7qgh+EcINsWrnRWjHrD0ohn552pnzZdNAPvIRXavC5VrN95TJXY19DA5
+7/xAH6Ubnyun//hWpGQs65S4IhpsoOR0QxyAqeS8ib4+94TLaT9E+74ImEunwSvtxdQxp5Og+DF
Qz4EKLdZS9AsHR430GesGnbbueQI/jh7EFRzW4p7HHOf4GBZ+RwIuwvFtXK1wc7qSGASs8JOP5AK
LMRfuOQS1dxCAHN3DlKUX2LCKtz5kLifPOHKMvdnVdZjd9gYMNBl2pfLBz+G4YuIP+eeXrkXmOXm
kqNB8499vJUVzI6023LRaTiGeVZruwF+rP6PjOtfZE+28j8rTy6DgDi2dlwT3WhviWKm744HC+yr
ZJ29fF6hNSdLP6Hnv0vl7WKlnvDvYzJNZWY02EiWCpyscdDZX5iNLxgmtRyFYB1BU48+/SMSjB01
T4FuZ2q5jGBuKf+OvbVQ8zhDlXGnrzwXQf4BmiUqmVam2bOVaFdFQWoVAn9UdUJAyVSKSYA5dFwq
7CM2VW6ucLd/trGKn8buej40cI3kTYDJM5v/gu3UVKpvk2Q3RqnCjhOMrSf/3cKkZJQEOjAy7q5r
aBx+MlIHlSugpcB0lSTdh8gi1YvPxRodiyEHXl64SrVjQCThpROtfUiWorjJMQ5asSBYWVhTEBDI
gXqmF/g0MHkwCVnvB4hA06IzG6Q5cberGHPUIb4T/vIaujKLZz1UT+mXp6hYPWZDgRlStJFHWq9f
QlRlrd6xbvW6xn173HMQ83e4rPeMna4gkpq6XnZH7IG2yzPdEwf2lKxuZmApKkxAncnIo04V7CF5
NEC+65ItVmfeqQVUndTTuZz4XmmUZxNvgVqQJXMkOe1MLaMkVOf2YncnYf/EqMjpKZtp657PMwC7
8ZqALrHwA/fmSqH0cvRT56z4rV+gwT8RPKzQjwlcrHqzEG9FbuBTU33ucr6+FWzYkTcUQIBjToh3
F6u3DolYgQnJUGKAF/bJxnP7UHjV5A5jwjQ49rHGxAe50YfycZSgoHB5qwMDbu8iMYreTHwTP++2
qr/Mxl81eMzFfB1D8D7eifQKwiQ6hSfxPH3PeUhmNfkUnP+pNOvnbcwroGvusKP+3GUGNjyL92dD
K3XFf0vuIyKEH5VwOOzkRWtXiK1T6u3oXdpQ4pUra4k7jthrcq1g8tfatByHnawx8aim0NbABFd7
cCxVJvccGg+h8Zh49E1CmxvLBICLkIdLEO/I4KLB95ffjrVos9PN7ttTCGnTkLbl7IHzzm473ynh
YZTcR9Nuf9gHZhjyTY+9bfYS6gApyAWCMfk3EvblUftvF2Hbsh29XwgAVChIQkEn44cKUrpjz0YY
hfAOUwOyliFqUN0+nJt9u9ceSpgtYQx1HDJcbWUCHjjyxRBszBVd9tjng7u1FpFmoEoirwp+kOSf
ZR3OgLBTpCCvZ+lb8x1cxJhs/vjtHKMd7SvwuP6yCXoaCXPvB3cyMc52MzNWztZ2gfDMb5HUVyOY
LExisTPBG6ZvkXMhvIz2dDO05z5b+ngC9/d2v0Nxz0Ujvnsuq2w2+RDQDW5oZSOpODRo5s2TycZd
mBAmx+YNIsMJQw4BpDaD5TKyEGBAL6tOcICQi9juBYT4+3rVRkDvpegRpp/TKr4nvOojHcoR8RxU
ILpT0zOiKQBdJq4HucDU+f85XjgfBu1iBcvHAQRKqwQ/YFavp3k3gRXopBg2mfgUa2i3kyPdnX5c
H1ij59ZiwPDxDTN0g3EYjcxfa3xuS6alqiMXvG5aoJOHSZ5skZW6IxfJbhDEcKX6FtxCHD5b4d6n
C8xzUoIVAGgyjHTxy3154X0XxtAVir1/jtx2Ydez64Hqaq9nLYri73wjM29HQncJxpywaIFnRPxC
bWsT8GnM8atoWjqRTulN2SER5opowXsQJrHWb5RY+QccUlZuCV6zOe8zwca/gj3SXiNqYhdnw+t3
ukT/jnwvMKvvQ7toNw/+6CZs/wliKAFIoptHCJ5JvRgu6ysajOiionZOV4l45Sg6vgALNDH19iWo
nnaajSdYE0HiZL308tKL6r9E/U3mBfhOEj/5eDpkyAS1AhC6wzr2JxB/8U32o855sXSbMkiskUlg
wPcADrLwr8h+ulVhgATPYwQh1T/IQrLDJdqxBJgUJ7duIHsr/O0nGRkGnk7RJdRkk3RDBU5J17Cx
W8w/iSr2/79rG4RHwnoPtk41FGWD205CYe4cbi+XEGhSbnMITW5cBROHtczXG7JXkgMvb1GM67Xx
7IzYu4G0WdwKBYYqziBSSO1pr0lCdQPwORQ5/nQEnvif/oCiS9M2ZeFvsmQ8Yfju0DRujI3e+1CI
nGVkriWJq7lojhL1e668d8dv/cNGyWz6U+L0iqkA8W/cpf+gVawCCoYs+ix8BiPLhY6B3iMub+hV
Xe1DMOgMWS116740x5UuBbgWYY2dQZg9+ENyxbCsVLmZWQBrp3XbsceoZFIZ6TBRUdQGhN6RgCm7
5KDFG6oKp/LAZ7splwetLuEbwl25qExMba099GEwv/lBLCC+e9VL0yKT1GDrX1H+NheA8fmnD9ez
Ww1fhTpoLi7kN4wA+Xid48xDhbnNRQQZHdHKH5blDo6wcMaNXXl5gT443H3hzBEzICMJmc6mxNPJ
E0XToL5JkJS/jpG3FSJQv+Bc24IpF+or5x9bWE+KBh1L810X6kd+ISLFNrKM0xzngxLBfEZhdylK
dtTJX376i5cGDZVe+T7BzcWLIOdKh1D5c0q1Jq9c8UOqZif5tUthsprSYfWBW+juizx/hq257QFo
GJ5Mdwd9iFvfYNAiXK9TfwDmcHOhfxG9WOVaZiXCZR8YOFzV3C8DSaykBnWL0InDTzmnAzFhKecG
DtzwJTaF0Xj+nCl8hx71oZjxHAdZ+H4jh2V1barQMIzauMpwLjF5JpfJ7dN18l6jUbo6T76agxAN
48je6xLJjVqkP4GUs9G9Ot/WfeSNC5sc6yb0n6P65MLhMyzi9invXTkz2N2RZNXAfhM152EnsxFz
ZUX/JDVFR8fiivpJ3PvhxSCcdb6OlbH/0vf69BpSwdQTqq4AVVKio24dJuoD76F545YxrGnkcQU+
FQ3mq8ZVquD6FOGlpKfXRWfXUHh6ce7rEIibEGTiJzk00ZKTSqjz7mYxvEKi0moaaTmbWuUvfM+x
ZueO/vvqTxZZ1p3Hpi12Fi8S4HevPucnXb6Or7zUmYPufoSPqAZxDVRq13/yRwUXq058tGvfo7nE
0WnfiEM4h/nadADmniFsmuzoIWT+dhs3K+0oicq6n/scvCVEIx1d+hSw742ByQjh3R8c/eNDRAC3
0I7AbD+wzUHGVtrWiSTKS0unUzzzQ9tx1DPp7h+bOd8IBzhfHXwoSXrzp8fRkj2NKooNs/DiKTfk
Jozvp6WbdFkLV02HOnJupAOPO2UEgxzqIGQj1GTYDysDPXTdFxByvZbQhvBs4H+pI6KD5Q1nRbOv
KtYihIzUDMyP3NFaUW3mU+y9990rPQwtm5cYGNfVym8sX5k0nySbkmjG6rSXhPfWRjoMDIf8cz19
Fg9Kl0J36jU/snQ3tuItzXUDRCgENdZLFO0FIwmmNEMjbATIrqlzjNe4g6nTZ/02uKzxf/S1oreM
SjsSbLeyM5Sn3WeEZRiGLQpbmdi5VErweju2zc5k0GxmLa3JHMuWf6Jm7CdpbhJBKoCX3qwYOaOq
5ntpO6EwnUW6ocqVDwwFNUbUZm+gRzDKNEEDF0UqvueakuCcczHWC70nAL2h641OBiG9CUAf5qj4
WbTr+8KqJU96AH5n8FEZjw5Zw/uBM/zEVdB5HqJXY6pjhcPnB+mSarpD6XZZsc8sCnMfB//BC4/L
zeSjOI/ah7qrxVYt1iBbj/ZUzjECAL/ODau3fK4bK7sam7C8d2odeLvOFti6WLLHn8ANVsBpzqq9
U1qvZQ04qnp7gQ0ZYEhlntOxnPxkla8LPb2fv4wY1D9jTuMeUlybsyvwK1BvpP0DoIph3X22yW68
aucYW+nY6DOrtnW5yOqsEkS1inMNtj6XsQO9QAz9XTHA+6je8xT97JtEE1Tb5nZFZVFzU5n9x9Jv
sAAgnAhvuJJ368sGa39sWiffV0y4ev0pjGbGDZr3EmdQdP+CPoDLGBqEjNGs7zXq8WSktA28dxi/
4Fzeh/d1uCSaA7YEPi1ftilAQfSvhTSwRGpPFtAvlcX7VHjyZALl2g8Z/HwHRdvGXrFqYrOLinXF
7pEpitcdETNPfRvMLL6+QkZ4128/Ao0lsVFi6bCgmqPpguZ7h1dn/Wnva717u74usdEnBimpkJE2
dgzyq1/T6WZLvQgNgMF+Jk5C0IVSqlNkFyVnQHsdcRy5G7I49sHEZ6RSlX5ONR0QZAMqdsDHT0Q0
ULNnsR1scxnV91kSNTr+gEQlkknOlL5umkRbWeyD+3r4011stgabqZAVs+s8F/QMKPl2DZ2MY/V2
xQSN3U3IX0yKNI2fZ3TyF9ROZC4YWOa2riG0K8/8QAyI3ylBJgFTi7DQfiO4EgjdLtBbempo7YUr
69oiwsktmJH3r5tgnbUOBbMMvHJfPebUbQZNgOj/cz3wVmtVRIuXdHuxXe0d6GeZd95AEPrun40M
vcLZkwPXUPB6NVpitApojGqw8jPxYEBaYy0aTlgZgDaz9Oy3c2ZNvKvr9fDB1oIunLiY8iY6wSEz
zwJbOVLYE6hx8UZpB6It7aULYitmpgfH1XVPhzwJHTxux4hCz1GliDpzaJ+7k1UILwnViXBN2oYe
YIDToB4BCWhYniongfAVqewDGS6Xe+taq89j1NzY+mrd9DKG9iPv3y/dIX64aUCIkd+ZDOms5aMe
j+uN2IZqsA26Ms7AlJo+xJ6ZHwNRjTVPZTVraxcAczNcCkE4A4772vrGAoPozsnXsxnFPqFHcUAM
ApjfHTh58mALFBzbwQvLtBqaIM9AIAwXKhmJAtD29diz5Uzz1ceDDiQOY90vslH9VbpPdFJUDbb7
lfVV/X6JO0ySOHXL7514Vp4H8/oQFuf5nxtwUBVakMzrln5YcY2i5BYE+ZugqB/jqYs/XqousMv3
Wt82e1Q3Iu0RO5Skf45uWwVbGyHbXv7Av1SyXemJlEJfZvBnWhrzhJY/obRtK7JbVuzdHIpRPr+h
IYsXptRAUNyVfdjwKyu8DQBOzzGJdprcyq6jyKHDFUorLCxrYMzgRR6HpaSmwRRMGKCMwEbe5c9e
9PdRO+wivoP9qCFcNPGiB7IYPl5f53cEaXzMK5tmbP+XTZBq8+9yomt/GELLrs0tLMyMd5YNX2E0
gcucTBf+h/c7KWw9BxkXKciaSkAo2D31Rrag4lYHsLxWuP+V38KAe0DDuViP8KCp5Z+OEEA7kdyM
AkxVVcvBRqt8TaiPVhvQdnSP7nloJTvdEkHPsa1wkNr2aBOJFoXsYzRxL+JjQ8IVIyMwOJSzVvDk
W96IzkKQ4Qzw/dFuLUMIzfzReNeKK0A6D9wm3RzJfIalMPwIpoh6W6SnU7GwTZpNX3aO4Ig22OCX
MMu0ZH2lBHBKvFIkXsVx9Qm+VJ6A07WX968+07f93+E1gijn/BVnGIOn9YDrqDZ2XWEEVWZWU89z
H1RnTvlwVkb5GdZbPBRxc3KWuYTFszLr54V1Ln8VEqGG3H66OdKLJ4OU4uvQHgyGqA62CIVye3fg
Nmre7Q1X7cV1TKJUcU71wq5qRs0Wisc0V4EttJMq158Trk7Vl29Ykl5horl+5SwXaX/aFfV66Zj4
a8BurBuJqHnQJE0BAawED7qQsNoz6bUOMYLbKCJL0LbdE5JJhsPNBpEbvM0m9m2P8mcWQ3b2Fosf
t/a80nnM4Hw3f3ru1IfHKw702a0J0eO3B9KISyhR+moSQ10kySzqYRGukDr90fPe/fUThFpVN2Nq
/M0WVHaNWeeH9vGIOxbPylSuPs/qrBYIvMh/EOsBZup/dqQJiT/zbwf8Tmdvl3L8405WTH8qnlEL
wRiyEUXRh3mMsZWH26EHRISWN+TY8dwAaWQMbBhmJeLwEH8B+kQK1PiGYetM02D6PCznUt7q73vv
RxcBj6fFPCOVpy1v4W/qTbKq5XruevLBdpoM/rqLlqo/kzFQxbCrrBCiBrYdKdTcSBUSK09zl5d0
qpmenOPivI6FyEzctmoGdJGLua4mit/o+MJV8dZamr13FbQfVFBT4LZXwgXkJa/VoJYkdkiRyTtB
nHNUdH94ab70Ben3tfevNSjEomw5JifGqiaCDptMaTJFhwuIkxWiFGZpRfRcum8IYk8Qs/HX5AbR
FT/66EQepwkQnVs8q0XlWiyWII5YOcBy4eZSzeGbMeobT59POI/ayQetcy1hqoWKI8P4CZ1+XVI8
ONuQ6WnGwzavGcyFOexmBvbYnj1RQYbJcEjoT6uoMqMDKMeaqC3DwT3/ZclL62zlqSWTGEvs6pIk
TUI1N0+yiL+dIZCDFiRk4FktKD0HaVwvEvlKdieF2qAnNpwK1KVvV6DrlcDuGdFdKMZNAgAW2ahR
8+VQyGIpH9mfuM3PVmD0IewC/i0mDuBTOasxawZpk+p8cvLcHdf8C2lGSJtmzxoraAdmpZSzYo85
KwCv6gsARRj+/AlKbTq5e/uYgFJ0PPYvVYeimyQp6ahrI8V50WTOJ8CNS6KHOZUtQ8tqjbrzqY26
6FhQI+7QHMUo8Vm/2QrgJtkmv2ZaLg1MGqapbCd7IHQTl6AG5Zn8nuBDlHnqKrygX6+osVgYSGxD
lMI3pqqmr0+kCCcXi0ULQFH8l3LVBymGSkMMV0lTDxZs/dF/8+gK/vwKbIqadzKVnvPhjLaJMb6w
Tcg2c8sfnJ8zpKW27D6Xu0nlpYqQsNNi5kSimAC4TN4MFQQKNrp8PyrDA7rTRmuA+ntRvdTWYz9e
DJoI7eteKiDJWj+gRMrH0/cs+KLZhgz3hxnfRs5tqrjKc6wSiu1809h0+ThfrVe2EFjp0GQ2WJ5X
ow0qP3Kng45vnHBQMYN5uGoXXJHoLZYiYuwPmzmjHQpAMuEOnGtbFgQgTf0fj38sAIqMmzeUyDPe
ukVNKStTDl+UZHQ82q7XawIdNhlKgBnaIldSHzzUitCyUtV0QPLR+f7Rhxgcljhxb+8WRRbORZwi
wZyJEtMZbItmRFO5L8ojJF0+q7mFCoyLNvSClXb8GL2ly7HwtVj24DXtzEwK5ruN1cTpy3QwNXq3
BYHb7Twa3CSLSsp6hs+l4jsxzDlhLoK9dnhgn2gJbp5FKXqCf7Ba+Sg2u/6kC2Sx/zY5X5fhcAwJ
BWKFmME/AJLXWNUn14vSiMPe3CFqRey/erNpSuJxYt2ypCqGSG2KiJLMM0t+TS391VI5jWlzsb+e
hI6wt7eZ6Zo4IeID7g3ol2AgpNAS0DqYx1rxPYnGYl2COBhnB2cyZbs6+pY/Ahbaawu+bGyb3OGY
rTBMz6kw0zk7oiUagyB33YdzT9Szoe6TweyzPf5VlmjtTeFjCdEVVvpPcqrqNZwA/as5GFyvmU8w
xu2Pp2gdIJ78ONQbDpykBbxrNBA5YrXZVcL3MvOSblPpqPbtir0C/CfdGGltbzjgXQXDbkadar8A
9xVMBMbYqV7mFNxxkBYt53vnOLuxbbTTJPWiJzmyMKegfIRyVYJ4IEXdIWwXxutmnJPafDI/RWuS
q9M2cOv2UD2YjW1YXvWxuib2bR3iSNuDFLm8fM3xKEh/+OVv+6nG0fsslgXMxzUwoFQLpfhVnIw1
lcXUR2KfYNdMgFjklynpxE2GjMI64Pjz9tsHFfS9b+GCWjflaBUOjFDHTyIj/xomXEi7DRHzlcBH
tYk/krvFCRTRBVptQV9DeoKX6hj8hEWiIT4faiNlGxnPbgtc4CXjTDnDOW2WsSxjbhgqV9D0xj6G
T7kpNK9jyw2i1UST+ahbCm+uYkgSr69wEWlUtynn8ImcwY2vNsr7UdPGEbEY4TGwNOcRgRL4DbLy
IsY0o6GnmBvuxdIysiNP1ts0WlBnnCmN1KPRmvocBrK0SH/o0t5bL0OUAsGIecUKK8hMP4vlEVLG
l/05+I1CbLvRwxiNWW1E/mgvx8HlFbvHz8vKriWbHZ/tTgmF9r8v3VQLaCdBdHovzgdI+HrfbLPQ
gTELS0PtBgMOyTcLEN5tyERnEosVysF7Gc58e4RJMxrlb2kc9dOrspYB7Y/zF1pjkALok6Olrwio
dJ5ltmqRo3dWJ+8Ngfa3p98vImOji8IPaXDArZCRIAOB7733FLxX/ZM5T/1lc9HX2/1ySPAdUmRo
dZHuriKKRwks89EIsZ9OtJuN6KNzipJERElQY0ZZkWtK+ZOgee5hRvr1eFWVftF+nXkeNuutRrer
ZklMAT3av3OaB7wcn6ydrHGHqDrtEvzICp0ZFHTYjBp5zhKnz/CCN/9tFg4Vv+wqBdzFemswsF7/
HoCnh7HG6nZSsnmZ1nQFDTsjQK4pzvj8JadKJf2HKnRh49Q+YCMCRp8V2WTNNVWhGU1BjK1WrQfg
7opyqdrD9S5yfb+avdfHb/1d6MF7dAc+aRlLEmWtmlTk2M0TjSNOWpcPWY1Zwb2J3/9lIzyr9zLy
1Pc3XQFhCPHvi3g9RLX1BoKrkF1IeV/zSIJ/Qczn2W5FopyNvP8jYWC6z/LQzgVeMiZQII2DFNf4
eMe37aulHjZdQYNLe3ZCKPnipNvFHxuxETy9BpHX1BEGgaPHnw3IfljyyvyiD67D9d4eevzg52Lg
1EsNTbGoqiaBN9iFzr4Y3lPu7zLIvlKbHuVYVexfbVcK/qHJBuJdu3/PPYXkMx+EswA5IS+geMNz
BRY2U5/mXzMu/UVwi3IfsKjfa8x5xMngvz2A4a0BO9aIXEN/9VKQhc7hAx87lV35POjNrH9uFfG7
3ea/0S8AdSah3Vxcm7EXmrEGhL3s5TG+EX9qBxVoJWDQeVZ43tQQId9GjnDlXpbiK/TahWcVeBFQ
N09I5nDUxp+sJn8uLEmH4UzODfr0L4O2oQCVOP4Wawa5rj4zF6E+A3APkE7VNVhkA3TjHmBaVSh3
XuvvkgCm/nKhL3qx3k4tOtjsTJKcqu6vubZCy+myMas6xPIYhh+fdqSSS/ZyHXAv5qFcV0o18oxv
ngJQDU1JIELIUdeWgc9OG+g+k4vWJ1SwsNg6Ml0EDFhpNj5pY5o+qb7YvwQFSRZsZx/qwKx3wZSg
0z/0xHkAdr0zF2gQwpD46FqQueuljCfaUgi7gZFEXZBUnaNmc5S6t6DNnboeabnNPnuM+uVKeDhu
Jes5LQeY3E7yRQxHB8MaLIEm9vgv5iIgF1/xVsHIA52uTCuQBvBINGdCLcePBUJ01ZmjjxwC6iSa
p3wycB6PfxFXGS1b5dYPtdauKPkCatdg3Dq5dtaZKlaa7WgZ0h9321VWywMJJ2SO4JoDFXA99PKL
ymIIZX6ItDapmO3UWLbl6e7gcOAZjEx5alPhbjVBH56dBDbigUin/3wEQYgOL+XzaD4Q/tJF5zPs
bXRNAqCneR6E9y9L5N6A5qpt1uK8zPRCy2OF5W36fg9kuZjIz/0VdOCDM+KMBL7tveAWSGI1briS
uwklRW4zjypl4cUlOVuDL+rOgzsPQxHqhD+aeN2kz7VgLnZOLoK3coTFk+zeSovsxXAgpDczBsRg
dBDX6mTS6ctQgVARSNKgt90BaoMscD709btC9TkkBt3qBUUBVDmRRw/U4tK4dWxQ5xb22ZJOi2at
m9o4v+YXtH9SfvwZiMinoYirha8lr5OaNmU3l8Yy3WvYRMAMDMgf8g7WuZvLMWs5j+GlAMXLtvov
oR3JfADbpCLhNs/fxSpDnLq9sO0WLGgQY6OZdy/rnzGhihUCrd7QnDqArraTn1pPI+fekcZH5Ehp
28n+p1orP5Mm4gJaRtPHo2pMXrWW1aeIuOI0pfMyx9fLJjDYRYiV9cj1Jw9o6h3OorP9LGoWaiXv
hbB9e8vSftQ0bYFNyGS6lCqwiKGYylxREcHHuNyovy6ZblonCZsDaBbxHIQAKvLw+W6AfIxNhwRP
VPZ12IyrzTRsfm0GVuUria3bAshGDUCPvFdjeWH+inkdkLwXx5s8OOUx7qiiP5g95EdZwslCe58N
MlE5q6JQEkNj2KWAmGm/7ZAREQz7FflcV3Zek0j8e2vrfvjD5zWctd5hhePZhAIxmvMyck+P2TV2
y+znWxzpYljQSDtFVuPbirKn3f6hzn4CZoe6d+ssqY8gReZ7AGpyLWP0C8ecrTL2C0Yl3zuIp4Tv
Kn+uJohKWUknHC4V3MS6wuB9QYqEa6zhoaZXdrW45uC9BSyCSX5OMnIJQUEc3YrZUHZBzxho1azt
USrLpWAMIZl6giARXS62lb7XNQc9XmqFMG+9s00aObWvFjH7tetF5bxTygS1JE5prZ81FfPTnBQf
lH8T6NmfU/subOyhupSZa2IHdRgQ85hDgS5MEXfq6fgWtEzfcBYhJUv68KTefOcxdVX3argJveA=
`pragma protect end_protected
