
// Top definitions

// UART protocol

// RO COUNTS
`define START_RO                           32'b0000_0000_0000_0000_0000_0000_0000_0001





