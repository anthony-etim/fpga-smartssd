//
//  Family definitions
//

`define FAMILY_KINTEXU            "kintexu"
`define FAMILY_KINTEXUPLUS        "kintexuplus"
`define FAMILY_VIRTEXU            "virtexu"
`define FAMILY_VIRTEXUPLUS        "virtexuplus"
`define FAMILY_VIRTEXUPLUSHBM     "virtexuplusHBM"
`define FAMILY_ZYNQUPLUS          "zynquplus"
`define FAMILY_KINTEX7            "kintex7"
